`protect begin_protected
`protect version=1
`protect encrypt_agent="FMSH Encrypt Tool"
`protect encrypt_agent_info="FMSH Encrypt Version 1.0"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2017_05", key_method="rsa"
`protect key_block
EyYGQkd2q3jAoavrA1E6hYYBzojRLOEgprBLcNCBoHBeqkYJ7iZtYsUgkK3I4J7EqileHCyRdCH1
KHQ+jpUvAWIE3tV8nkdTEZQz4SZKcCE+iceCO8C2e+Knu7/4skVM2klTYclaehdcm3Ee9cLh7oSC
OB7YRaKxH61i4PX6CmeKCBPBXjgkNhl46xmrsfyPeJbenDYwwZGy0kgLPFUtoMgbz+8LWU4acz8C
mWMSG7WEAS1R5KQfHpvf8prEzoPQFH6JQFG/3IdbxpNNrGm/1HV/3WPjQotfK/5H69XpmSDo/rKF
9Tn4m3567UbrMXsqF++xcupaaxXSKJuQRq2FTg==

`protect data_method="aes256-cbc"
`protect encoding=(enctype="base64", line_length=76, bytes=20128)
`protect data_block
/z1QFLd3S04/Md5PQ+AYzi2Eu/saIJD3jk+5z+WcpzH6/D7fgpVaNCsCRK5FKEflqFMnWJUZMvkj
6+xx5i75I6IGlxmtvk+A3JX0ffCD6GC98FGlu6vwWEx/zdoihi0jRBdH9pEZYdcWmTZX0MsuHV5R
asBoj9g4rzqo/tVUj+rrX8BxwXnp0haNW3SNTuGeld4g2BDUlwwmAFEF5B4ywbkKZwaGbfpHrhxE
IZ9ym4c518bEnMWpJN1jjHKhAWIE1rWMmddoZz3x/YSgCO2MMFKZNipn1EI3IXQmFKah8Cs+iQ75
QJBqmxcaRGYNYLiN/bNwx9S4V0YhmZg9FS9FdrWfZs4VFPkdCyoGQPCm3lI0bbkECkGJkEWZDAIX
d/Ha1skDtx1Sz3A9KjAtF/rDjFLam/zud3dQ9GKKaQq+L5ARI75a9Z3a9YaG2dtCeLhTUEklApSw
rkTJgLpfDY5tZpJ2pzYD9PQ41LLXTlf58JHhmS8YnYj/mluc2y8jpQug2Ten47hXierwKkq81aU3
khz7BRhJogCNsAmhw6lkG2xDgozIK43ZA5DhIMwzjRPKbgqSExVGMDJr2d/V95ZeG+MSYFcW2PaP
O4WZwwLubngt9VlHk6PpK158b7Emj5kkpLqARFqhcqRTqPUwkLjfFoxJBRzMmSPYXlJzMZcyija6
n9vN2AV8PVo+WkCDnQNsYKWp3+7jvP7iyGJhdAWyKtq5T/1zAeCT1/CvlKs7XIcypPWNnbekHHiM
JANqgblLCPrl5TVwHxkT1ea89SJqFeBKw269xAZ6HO51GxI2l7SmAIWO45QaeDp4Y0N5fnvVbTRg
ixdBt4tA+zTZyrVsFyCe8Y7rzYYVgL9kGrIGpwZE/RZnOi0FGZZHnZns/JaSj+kDgGvNVztm/emE
P8aTFTHX1ZC9OMvTCPmeDu4MKYVI6iqN/erMyvJvhlcDuDTY+qkrR5877nBkD84bBhG9+FiYOzsm
XB+WXre0fBZbdaSQTwkW11XI24YvUrsWkyJm205z8P6HDA0oMJrMaJ1X5jWGIcPzABAc7770N1+Z
fd8wtOmH4XOVzUWrEd9vpRVutSMQxEt0a8d8rQwmtfwpmi5ULPcB9eYCep8KaeZOWpa1ki2DSUcu
tfPoqfQwXQn0mGk+Me32yrUr8tmvYPC4gs32ppzAviOXaHNRA8A4u07rwyil0R90SbPMLYAOToVc
jI7CqK3T95px14xRKqSU//pzleCpgPEsgSTzXBxgODwlzljcvzqK3M3mlhZ/fMcRd8LO5eQhMYBE
rPg+ApED6ij3edEcyIbvP9b+MtxSxluAM1hDKLGprmY1HAhize2QVOiTmazWetVP4HHe4Z+mCfjc
3mKGLaEQmxq8sJmg27s1uzr4PRAbD7U7HqaghIM/udwyE+IvfIQcX0Lg5qZl1WxtEx6TTIkm24Re
z/hS1NynGtdJdFT/BruBbFgUrD/UycRNxBymGCtt8tvlUW1gI0l1RS1xUuadZlRQz+3XFl7G/sf5
vAfav04ukki1slIbwzIamS3QK3azZavwUdDoIPi3gaPvs8F/5MZBSC+Q+TsQTxyuHT3eKVsABuFz
irZHPM10nXAaP2tWJwF4QozPTmDa+qZWAH3fPDAOQ6BC3jeoyR5iQLCkzbYGApGPv3vC1++14Khk
HnBwUDcmpuWa2G59R/xxyIdsNV3eWwVMYpqpwdG68lwsUefRqY12uHo2ivtZiZbNOc8Yl+C/lZXc
9Yh4ZrPpSrxQG6zukJyMB5AlCjMtj5tk9fBDUo+r/CyxxyemeThjyRg2GXvjOkQhezGEZgncisF6
F3kLwsmZcMUrOkgpLcncHnACC6Tqs5C7df3zgxXFOLXJmVp3JIIPCs7/1u2fbYoBfVPlftrmTW5o
TXU4mBBp9EDsHupRX8OPdVI0RY41SWgPLzdTN5aDDux3Cbdw05EjSh+6OvhsASe1ZoD8WOqr5IA3
GuGgUlNDbagm9DS7qWh7CQEN9FjcadrZJ69dHh0okaGdUClYlE09kRAzw7CRcUMCjD3D9Yxbd421
SiHlOpGIde/ooRn6Z+yHk14JO+0LENd8VqaWG8j+VxUuM/Qfw2gSos5VxVLej3KAuDWKVF9zknQS
lsiHktokeAyTRrD04yfwZVUzK/R2esgjhGHfPIxuAduUziOxafIq9gCBw3xV/uYBPD005gJ17Ttf
ABUoL/D7cB619REjlp36Py6tyCCVuSe4ng63HP2oVdhoGMqYnGPi/Ot0vCRNXZDchWNzn28QiVVZ
xCxskh4bKcVJ9hZFbHxFNqIXBwA802/SVTQrxzc6RBrRJr+Ei8K9QEf8f5n0OLD4P0b+VO5FUdh2
X8E0u8o3dqzhUgYGWxEvQZgefPtv2ZZFHY9s+q8U0INeFDG1scBAHm1Y7zishLCyTeKugOaRK8Jt
dl7Hvc3jHw8gp77SNGuL7bdqQ+Kh7vgtxfp00dxmc/DKcyxB7WcgjWPviGJkOplNiIq6ALVUd3dQ
aKKVt8GPplwgrKL39UAXkfjZD5qkVDWry+pdz59hZ4fuvmX6EdJJO9ELjjYVzlB0iAjHDU42vGCj
pLhaIpWlpHRNmxqdDi32hUvYyeIY4khpqh56H/UcCwF9XDDNmt9aoy9GN1AiCX2uGjyO/vXF0GEu
wSHoE/Vma1up7kTJZiRsWCP5/rIYLD5d4wZ4OZO9DHQJFgQ27JsUhjrx8hHrEktHSd8WhMZEha4V
TzgY3tKKvz8Z/s0zupT/AhSda2OYdfDUpkfUAdbq5amB4E3ecPwXK3MgF3C1WunVYH6k0pmYLx3D
Iin323NzZIBi4lgt1b1nMbpBFcevAv4n5DF5DP7c3fcYo9w7KWQwyCsKOJDo1PdhF3VKlcOVpN1F
4o88mvk4CSRS+DJfyIcttFdyOVZbh2SisvvGnH8jNWu5fTl5HZM9evSrqsTPCoxJR43XSEd8+njF
bZBC0TICXbvUcLbqyg4ioffxCz7VCNGG0zXstKTIt7yZbPf4Nna196n3rrWN33FlbTwPTM5k834b
Dj99Ct8sS4JQicXCHW0WBiulCS12xVRmaHHp0oLcSRQlRFMageHQatrWUAIxOyxR3Aix3PATLx70
axFNFODnCuhSdwucbFs50RqOQQ3XO1Ca0X4ujw6LRWyth8JDyZlUg6+HADC2JF/hKAoqEyuTwuoK
6Y2l4lqBaNi6h/+4Qhh1kmkcBuiMT5PwSVkLMyI5lGLPpAoR0S45HhMUsOdsg6U2ZsDkUbl2n0RV
XnDVi0v7EqG/nB/+TKNI5hgNVke7DJwkeWnFBPtKQPXGXcgsR4+hm8DBXHUNM3BDc4ihq7oMc/D7
YkhrnDrH3aD/WL3dPJ8r4SXWBjHVy0lVdLXwrPx82tKQU9VTXjaEtZ/hKcyxJGM/rS974Nq5w/E1
VQoeGNlSrG6XZfznQoZabSyLG9h6JGKqnGer3rPhlaQ7Ynk2GQ7M8jm6lmMAkbW9lozycv15tRXq
NzLUNXEqZwTTRwm+ui7DbmPylCxpp3hTyiwU3Vz9mQ0jnVd0hImJMTIoFRspnIbpvgPKOW6Y2Nek
VFmwpWW53Yh8ArC0EB+TlrboFPufhjNMwYK97y2pQLYWNLI2YlDEJGZAJqmx9fuXdhGil1V65s8E
O3hFqZhfBpSs67+LIQDbzPrY8T8bdJvze9/w5tPKKzN9zmFsit+6J4tQhEComoan1nv5sK/PW5Cq
/VrqOCE8KtHssaDCX6fHA1HuoBzBmb/HP5iNITpnzd2uiiTCGlRTbnAUYMnMyG3JHI/3KTGGQ8gJ
Tm6VluS0oYTc2T0FkJdEKOz+I7hI3hXlISHJiB066ZZdgXgC5WPSGF8C7rinzSr9dyb+heG1RpW6
L+0ZpU10wx2NA3QK70MW9U361UJ20PuzOWRB1vR7ipSpdfmBSTmYs4pNfr9mxZIS6SqQBPHaxE06
Rf1/A1CC7YTI/BqvK1wfCoXVeFtvMWzjxp5lcNIpAf4TPzdYBHumSqBQIiLFsiKAWRhv4FJjht1i
/f4E/MEsrJPNB4x8b9Tf3NlIWxWWSCBM+A8ABOF9yC/N2gQ5WasGzjipKhQKEio0ZpHYxbrBI6V7
S56xCQ1TfVVjVKnKFr7bPip3OwvctKnTsx9S9BAbypkPFtg7lTMdg1HtvFsldzKKF1Q5bQ3R7SNc
shE8Wa4POv4IufM6Pp3gCs7CiB88Fv/QK1Fp8ufVIZ0WxHtNbFTlEz2/XFIGKOklHJYh28h2gmAk
6HaaefNpQHtOS5W92UYotKT0tASTyK2Cbe9mbEP9k47SQFJUsIlgeL8Pu3//pz4DaAoO5nhpsTdB
xvsjmqHnNVXqpy6YklrkWwTDVgeuFlMzJfYET5ATH8iWnNvVW2paMC6ac2xdY6wuPyk/0NJ3Sc5W
XCATykxpWCYpPCxG2eF08tdeZSuRJ7L3r0/Ep2wNfDcmO4tYFZLecdesDRTx0wAh106PzFGnRJk+
FB1x8QU5PiuNUYQvELUfHIg0BMCM7lPqOKnyVHF8NYGQZ5STVYWTyS9shhGD7BNJ3L9+AQSBCftv
HW0CLyBSts/WbvMJZjgaPIbLvJIb14dRQFUwKrhdMPpP17G55wSoZMtZ2B3Z5baoEnFA6cX1ku+x
GCrzqQUUTjN3wrN4gLUKDLikuVBJBXfzEqAXDpKV7i1lZMn7NW9avdENz3IngwiuWBgnMCOW+eO2
ehXzZal11mKdTUTjvBZhwGxB+NRM7L+O/FX8YSyzw8q+7OAAb7V0au3UBrS04ch9SYkNbJ6bK9LV
5dYnizvAG/HnCunlUcrh/tIqQjYTSu96zfhzg738c7ci9925Jytbe9a0gif2Q5IaH/e7XNRIjM3s
4hZKAkQ4Tq+4Z9gv8NcckEN8z6NI8j8BV3wkeu0tXk1rziJJVGsR9wUJ78rHLWLbl367bCOhWjjC
XvEIf5gCAjZnVHfm7IqA9ucjd9OWgg1eT1qed1ZmQIl4a2b0lFJwqBDj7z0JL4DTM8i0SRvZTd92
aBtn+eZ+8UDZmmBa5IDqM61KIP8oBxQVa4I5I6524BavbCsM1uykcnQ9wO4z/xu15j3E++fo7q5j
3Cv2r+hwPAwOr3tHH5y2s3gKfn0T8HLHSn3gcNybYJVe2CCJC9MnMRWkq81QmMeOfIAwG/zUQdyY
TAhqaKvMvyuEXmjk0J9ODYZac0oMx6axcV9yfyOCZU5nnbA2MmlTusZmsYmAxY4PWsGSgjBG5vCS
OAtUYtiCrgW1ZyUvCQE2q0/bBvn6u5QyaB1xjjlil0Ch60cqmRknKikkZNckiN0qQkC/AAV89mt3
Q2GWNRZ3tTz4MegXq7DUWG2ECl3698Mo0AG/YAmlnls4w2R3en2eZwat1UpAukscolNNkqQ8fnOW
lagifmIujvUsjkXySrWpuuhrfpabWBH/AvMZdJahPvc3LJieHOXhGjlhhn/1YDvF0TcRu4sKoQI/
eEz4zvcphv+SYqnES4U83QBvKdk/VWU4wN1kBoWMqAPHK/P+NW3dtBOttIPpmfmeNo/2Zemov1sO
EYlsScOCAeHVKycstZ1NCJB3Ws524F/q6K9nT3bnqKHtR4akp52FalrAYC5dnAZKUHplp/y99ka2
RABVnAyql8AGv5aEMDU6G8LuUgI5VKlFms2L556aMvhC5fHjO94oiWVV8/hU3HVclWEoYj/PIpdK
PHqepmTmOmUvvgvUALzhTS4zHufkDfd/8NswKVyf9z96q0b8RxMmT0kAQ576lfwTfur4PCg9j+4/
TvMfdV6dtEU/pjvRVy19Gg+vSPzL53bUtiMVlHHLtKGPi6RVdS8foiythkkhJrbv5xZ6QPUc/EOo
FvqoFw0wo7go1f/DKzQDn7APFOL/EZLkmwptFXU97Tv89p8oGb940M0pFGttpUMRM1VPct4uQb/V
rl+sOn6JVjBX3QLl4VprjvQYxnyTVPitmXDSv1qhRhdsApELLrmFqh/E0u6PPKzP6veqBVHvNr/u
NI9LUa0wrbPqyxyEG3K33jAgLGP85bHspsj6n/b3drNZLOQiQF0QVCCkvbRR4u5lxnM/t27Ie7XW
AhiheLVSsWt63sN1Y5ROB2k3jG4HUMboOfCNKhfZPkRaRIIPSLjGxrjzmSNSHrt6qt+FjXga+JUh
We8X2VBynIiPMYLnHTU1ZXq7rkwFzfU/PKPPxkjgpb7d9mPpYrpBvyGAq74W1cDY9ZRTO+w0STRb
ep3+mtWOlSkgDI9tTJxuKNYNz8nOw0bI2q1bgmWTqCRXhAI2sqAyIa7wEcjnKMGf5JZb+kXyAv4O
Z7KIKKrTSEqdHV9qPzFsztyWymjjhMpJ+xQfZDKuUMLls/jT0E0wM0SegvHkQY5tRO9PhW0jIUiU
xPkB1ec9+Pt6Ye8oFHFdIht47PB1FBPzre6C8EhtzgpUC0cPXoBzmljJ/nR5LRj9yh773yL/AiXv
8bhsjit72Yoo5MQeCO+1WiiJU/MjePXHiDE2o0/2tcgmaAwNFkqsrk9uHAuQzbT+iZJMPcUFrfjD
5v5H1GTm/1/rVmFkspZ3QdMmZy1wquYEjkeZgfTGdNEHVDVfDwtrdLLptWQtvcS7E6h/r/rRnYmG
NCYV0M/C+2+SPmnONcBJETD6jUC5S/PLlILXy/7Bjz4r8fBAGEEiu/XtsuDzWV0GKyADSY86wh2Z
8e2N4stM2uSmpnFczRbLEkz258t6i+/h+Ax91/uss+rzjuMWRATATONTvlqOAC283ctotRtqM23r
bmlTSPCqZ8jHsYv+eeetqoPpbXeARDmJ6nb4+kw/0wTeV6i5xs7vbvXoysG1Aee/tzMTOewtzr47
BFEyA6BrJmTS/Fk+Rimifx0r8e3phivQOx8/SAtTk6HJaQcZrzK8FWXK9qSJIQakAHv6IIeqj46/
ZX8KynsXGXRyT5MvbDjHhW3Kda18AiaYSRPp7EcTAPbdSfkETJFE0NXs2zu3hAEQ+d5NdDRpt702
cPPooE/mkkGeIDFl+MnD87XYEuSSTYi7mQofd8ay9fvlgv+BysAYlGuPQbhxZByFVasq3At18WvP
OuPW5sVs0FdtGrz9Omot1D/7GSZzAaPk+yz4dDjdEZ9oYl6YMUsOTvZlPuPxqG8JUUe4zEqcAnMx
dg14XI/SZLXn2I3lwRV9+0jLjePxM1znYY9XK8YdJ1yMIHGEbd4kkB+AR04q0GOAHZ/oD5fqWJSF
XnFq74jiGDJ9judZz1GRanBFQ1gkJQYXCPvO6324ad9r7AU/uDQKjTe1tgxq8pyqyhRbeY15EC70
4vUkH7EQ2lbM701Z6i30mPN6SvWrzm+b2rtqsmc27LhEM2iLXhKgxquTStNOKTbggzyxhiUNhey8
49IwLtKfILN3/8V6VgcGPFiXKEfENb8iv/dlBbxEVpskzKT2EkAj0G/X1vG1OgM/ZtZwN856BmIy
mRstH2ZcAtkvEJL3rGA0LQ2S0guhCHQkG5t8Bx39wvT5eSnuR7kpL6eIAco3ghGSof2B6fWd96An
RC0lBbcA84FHsSrNlWy67EDdDGJh5USPDTu1fYcpgMhHvyfY2rmJoz0AyzXTf3gCcqlZWbkBbRpC
xQUhUWevlNXG/5T2uRT4yvIUAjbBatDH6Fr6skpTsEk1CA5GEwAw1ikn9PDmb3lhqCe5bbC4Jc7p
h5Sam0xgGF/lBiPzNAqwsE99hLTml73x9yDkaos7lCUftaEPP0XgTFNJ+FsPzZhwZMm+/YF6fX7W
3EzoUUGr5jyjmY79WJR+eQ9RlDedTpYhN+Us4+oUyVp77wl7tABR+25sYzppYyMrW+Hfhyid9W4x
mBaVDVi03dhZDDoupM393jHYpS0Gcf07yJ9s0QeXCbxi+Y5g0Nv4NYTV/O6jbWrwON3MqNwsJbD2
C0hj+0otY1HXk7COy6S79Qm2hYBdWRU2wAAkJdlck9eUiguqilO9lNJYx+AkwSRM21Cpzc4fhIlf
MlAM5CBMUIvHdUWeC8RRrMgsp0VZJY2iNhXvFpLzNv0im+TacvtCTIMefp4s/5uq3WWiXEPSEbyk
cjvYVvE0IVEx/bhbP2g1NjWZpbkHRFb/PORUSC25lnE0cdfGYRV7yRu5qkwaMQk18AYgpdER4/dh
5ZN3ITX7URwdlDHQhwTHToo0tHWcBhjuxfTK+hOqo4OodwBpcWfXXZFbGLLwgHpxVGQUQI5Y0tiT
pD7ei33LDFUqFaHs2YxhmokErtR51QtzO3xxdNDQ4J1IGlqNkITCeMxk8O0Z3VKk2FL53pf2KSjy
B2NdcUYUdmO5oIqP9oUfxD+znhWD7ABVXob4cYbS4fnE21CfzbSBcMRa6kEZSu4aHo+UpWQ7arXX
wGflE7/bfQgDKkZ7X/3wXG4aAiILfFHiP/hGoN4NJCrDABdlTRErL42HuwZ/57l7OcYzEGtUZYV4
L28/uoBN34cmoi02NHWW6A4/RvTkN8W8sz9VQLWktL5dDgZVmA9HkubWJSD5qEk/0gOf0JZOxebG
cGrLVpPmmJECJ7y19TlFdd0X2oo4QyDgyoV6Br2hFJJ1OJTVZuhuSG1T0qGL+8KfcZyD4gsoQwFK
Nub4UW/1mAePYuLnLcB9Vv6oO2XdXN/a1mk/wQ35RfcPal/ZXQsONEttvrhPic/+venhU2W51VFx
2xEETzeuAMM//KGoDPnJUk3Jzi5SRmKQZYQdZtEbWZeJhzMNUR243nuPJtErcUM3QtdpBKZzlWmm
RxS1R9TMi9WZeLoKf1YLYiXFX5TK2M2loYDHajhYn3x3e6CVUET7sysjx01EYVZDnkRdaO3VECBs
Hxu6gRHxUoRCXRB8uYeGvjSucas2JHz98srzuuq1y2IPVqSuCYj3tT3KwOHe4lQb/TNCyJP3zFEI
DBauciHGYecQLPKj0WzeOZj2eVauzQhTP4ux93E1I8VtuZDJNj0FNm0QDQEWKTjQpTzNMENxKqc+
KKjyoJyu6TludaJPG/SQhc0Ckpf/mDF9I3iJMqwIU0qw6E4CGg/BFEj6BZczqmrYhR6A14kmvKfW
bL66LWW8HpPus3Ge0Bkep1tSPDVg1WkUoGAHOFIR3mArWloqYdjMMeggiTxkaliag7LZT/y1bLzc
rHPljfdVRzdDc3uYPBV/KNp57Ec3h4mxO33iN81cKsz6VlQkzquFjdZPOPm6JbHZwyADFwAYRoJE
GfoKU84/S3kdOlI9MQwyj/PvgyBsthnbzlQ1VKvu4bcmd0CJFvEDnWQdBK0HiaVAV/O3rkmZB4mn
nD74VmkXJOYabIL64/1a9wq8k5hNs+HZ3Hk0LV80WpNoOUPIgjfHyp84ObBS8cXaRTgt3yi1lrl4
lUE+38PcLDevJYaqncxNzZfhG+CLzeCgRjEASqxvdOOxmfFHSIgEZURHMU3+zKgzob1MIt7c980Q
CtaVh4OIOH13/oabHQmR/FNxfQndPECFKcCCVUhSeJLkt3pvyoH6tX6bh623bUoYiy+7pEITmQWx
C33g9JmxRyYtabyE0F+nLVC8qd7GNeBGWskprkYvhZx1mNFN1rwp6w3FY9dLuJjuE2z/iYvckyTH
zYuYiZuuva39T+9+p6L+FEZZsj3DxMxQecm5UPnnoQAIT35rwj9e2JAdJU1yJIxKVIOFHIX5cXZC
zMNCWGcfbGXvinKAJ4/OToHwBwfzzfb70F667dGIDy1hRlS7RBuDy45e3TZo4M3mc5NO2pJP9nWA
mpyeVdhPIKDoQ0t+h9vLtXO8oVH4pvurg/BZZa90JAJYRf/P5UXkCarSJj4o4X7qbwvB+VzM2Azd
GO781wKCFTm0aKbirJesQF2Ic8/JYFKdNNwvaCge2iiIOWl9uiAye8basT6rCtCPKLqE+0O3zRS2
NII4M4isXBKfbuGdjfdla7vP4i4wTOF5nViwNmV8yM9CsQ/f1CgVJPYydUJJXrE0NEXMRkBW8jJZ
vxtqzxkapLvqo68fmJZN89FV6/lduhXtO/znAwUOZQYMx37oC+//BdZjxqJBHE2pOsssBXYvnqCC
ICz9davP9MStwarPLJ3tEOuUGMAibcHBAeS/Q9lSSj8JtSuRsGFVqaqpGl51jhTTZPrV91Hp3F+e
5F5eBn6n/DSUGfs2e8ZvVT3I4MY4a8g6BuwR1C+5fn0+X8LBp5oYdgvfIiT7cM86GfHXwAul8XZ8
IddHQ8y9lwLp0qBgjxz+0vvVmyjcKzNIhKNtmUVKX83hQf3nHSEyqjLSTb2+vHsMtp3tg2Nyz6Vo
LlXdsG6N/xilfDVkOziTL0nVXNqT2KG3KbSzOB0XonfQzJJF6JRZg09QJvO7I2vfiPJpkSAnVwQ9
mz21G7PMXd+bvfF981EawRLfGmW6qKxEL1oMl5Oqlumx2ta6JHnpwx0QNBlWhoJVVodAQ+/kG5BS
7vIvyzO6aRh78dAgIwhjskCEVF3wLXId0oxbH3lpSbyTUACzprZE6zSfosoFzS51tnaWtIFqc50h
FXgB5Q8g2ZE5mcNAjLWvfEmdlj60Sww7gIHpBiJO4ocfDM1VPYvY0C41VGXBEVI39tedRtVaZnjL
9aG60LioLCekFxbfXCZv3d5IY0GkWdThhWfGaItcZ2Ka9ncyB0jOKznqpZyG78R9XqqhIfqLBAzK
GVULdH+Gy4krBN9BKyBt0ofNMNivlRjvQeh6rA0acivOsrBSxspmNVi4N9a2vxQxKqVIQTNpodbq
JqanNLjoKmuCe0zeP0eIMAAt7FUH1c6qRrMo7evQcI7mS8nEaAnG9rlOVKdTMN+u7s1IvRhC5LN0
vs2usG761rpZIpLGksAWKjAokZ6jdbxBt2oCEBcS4ulpNGir5FLVy3SXQaZJ0o2kyd7v2tRx5ynf
XYjkpaQxoKwgIL+QEd8nNbbsFcHeLsf7VASA/QrBxQPQnSmwFDtwCv2V+gS2F9jYZ4yj92qWka9i
vO/zIt8o1FH4GPHRilNTl2lFU8k1pJXP7JDPauJ5B3PXp8T+/H344e4x8v0bWC7fH2SF2WekYheA
HsD2/U4ZAXKHUsNIAQCXe19m444uYOfaIIj0Oks3YPh0PUpQSbQu/Xu5gqayTHcM1/kFrD9OyF3o
02hiYD0toET7GHJOHoG8CqJkVYkOjxSnNAVs9hX43oM30MVEt+Q1ROaPMB3AzjXT/3I1tMtONrEV
f2gbleI6nkVqg4owiBwvUNV/MBGzUcazF8XgRYjd4LLaiaA0+obWYC3W8H7/1u5N+CFeAuIG+YxD
CLoP0SCTiRzt2IQxShktrnOcXde1gs22AMKYf5EPkJiRY01kTaE9ABjbLf44JqF7mcjyQn3T2gBE
YHp6nWUzh6DEQIEk/FKADpnC97aPBTLYRcb0Vysjs1/v1MbzcjX0F66x6u8Swx7i2CADITng31De
q3ndEoJPyxY190Il/nmrFx9xh7NwgLGFSHL2q50Q+N00oMgnFWbOmlT04YRfiVRgJuzOjJhRQIil
sUxeiLFKLqTHzaOpYPDUBV1hsDEmosRIAumMf7dY5aQCmZQF0ts9TCxtYuyaGrXtuNRXpGc5YvQm
bq7wczLdXQpie4nyrWigLY2h39YdXpmaYqmA0n26Pkomzq93dhC47xV4ImI3fVxHrItGnsJA3yzM
y+65ZuhErACCyg1r8PIB3+2uTVIFPaVCzHK/8qvozn2jjmapvFfxO+yjCFY1tia6zXMn4tb/6Bin
FliwWTfWsxEC537+ZmzVB1hq7kIZwPTCTC7/2JwlD9YmHEhTtRtP5slFP7rvMkDujFuFTmO4TkpC
tcs0UH7BUUqLTR03fIQ61HpQeHJtDHpxhmPTf4WiA2Jx3A5Xqj0HkjIf+542fkHF4zxYzNIBftO3
bhWpjVH/WhXTQPIspUQzCmHkAkSmLXCGQPiGYSdz2GQFqgdv1ZFJUNlT0Ue6dvmh0aTp4hjHhRXW
DNRHScLuxfh0EUKUFDDRO8xqSp6gjj5+I5ckpt5Iit7Vs+A19MVaxXHPGo6ZNbBYudWnIotJPNli
+YES9aaXS84r28/1u1PtDFMn5V35bC7JjjcZSAbCtsrNjWTa4ToQVhgdPnTKoZyNA3DxMRcXZu67
Q0TAbXKhzTg58CWvh8HUdR88q3maDRG9uBQdSXft/YFmydm8lGgweUQro+wo6UOs4Dauo30M0jWP
yx9NdQjP0k4y4V6OrUNioOhH5CCs7H4Anm1IrqpSFd6Y5YLQi2icI1NAWlGH344Xvk6rrUccys+Z
zehAKR3dNUFAaG4Na0bHc0fUc+N9iU/U/00oClkLgVt80gis71DGRnQngURG7Ei65Vs1a0O0D/hl
M4XqCXI17YUcT3M28QqQFvLJCRISuUIyIXqQDYagqikVHbYZ1dCtq/qz0KmUs37KKWGTL5oEFunY
UywgifGp9dMEOCGWZYqhqrY7aSLUKm0In7A9KWwu933XKCWpABj2V9ZfemBIhmi+VHlJI2WlV1Yt
7SRiPRVcIeBvJ68bCSMwVBezQwHlCjjTlwIWKtoHgLDgeo9Dxtf3xQySyaETvWx8XHVDzWWGpO0l
bNDCZkcCwwAvvbMjfm3H5oAK1RdF4GWCRT7NfRITbElndDjCxbuD6bTJmhvGdmnwn1pGC1I5+s2e
N7SUuTLZ5uPpOawtvfHNI0fx71mjwn+STPmn0in+LbdSkvqBeE7v/eIVjDDaCGX7sTm15g4pNuQo
kIhWxQY3nGhWtSTXnVmvWWkDNwvwsVAjJ3TNhyapViXb2KiuPNKzPKQlm1+JD7MMZo39w2rRRFyd
U57arIQdUyezR99Rr9iSCU3oV+E1+G5LLD6P0TX9CPIe20pHhC99kBBp5mNEPNJnJJhQwdMSjzLe
g24+lncKmzC7HiYt45GrCLeAoazpzzDca3yR+KvP+KnlpSl2KTX/VHaJvpJtJ1oyA6+j4sXrZU6B
z+LKaFPNSwK53MyF53ILt0krNUak7eqXqZSVx+JYzLHpn3gRViaNrvUXet9bx8OzfiJaUV76v0At
rFQzosxIYxTa55fkWx/n/Dz8kRExV8ApcLMzHSE1/0el248o21RjYLyqaBoAHkII20/6ZFfLv3+o
404etaGXi9eF0QHgB6YZLQDj+Op67IFKYQgoZicQa2jOABCmlO3kautpvQie1Yet50AeCWEM+0/J
1kfryxlAUMkvnzX792QCKVcLEgUhLMa7zsZ0TUpR6dUEKz5ppoyvXU2eDGFoASi7EFpE+X/tZBDo
hfd3zLD73dLDeMcxHsjDZRmFU1uukZF0HfOoo+fitloBi93k/mqC5ZwpQDa+MRBudnMjBNGtr6Gv
/v+uJc8DFLzuTkxjmAogmD5iyvVC5KY2JCVVnSJ1WoxFLRGJrUfEK7OlCdTkCm3KQcYOeto1lkHI
I4mXvonvIEZsojmzLCHB6oyPrlnDA7LSKUPitXfoxFqQldgPVB0KR3zKgw4bi/wNXn5JjrJ+39Wu
vM5Gg3Gw++YbelqaMP7PL9SMLKl9ktLAJB7vwGU0gFZdeH86EazGSL4EZgTZEglXVBD0ZfMEx3YC
nRQTEVY7jJHyrVy9OzKcNpphooy8qz3Bx66XI3zwlVaLI7bPfTCdiYh8E+MoBFSHpnM/8oWd+IKF
tQfCH1WSXLV64EK9WsGKIIAEG7mTycYzeurX1Ev1IxVg2xXnxcSE4/kAZcBwjRN8+eNsGLOTnVsB
L022BLaED/YIpyFh3NwBaf+lQm+xvA3689xe/DWGJIUOFUxLDsPbq7k2Mja0V7VMzTArj7w2av12
CLBNzvwt+6szfQt+fVskuBaCRmRX1vewD8lvPFn8Kz8QhbYDeey7JLv6sdfMu0L/y31K1JcWmwyB
OtBclNnhhk99Z0LIHLPP8fw6ol9LAB1aPkPtKlZKXmlM1Fc4KKl6/sVg9d/O9ULC+HwzTEBhctpX
vvTtvzvN0LmPu/qk5Rmz8/BLyYEftwmFk/I5Ta0HSYzk8i0FfJUnXC99oTmnE6mO/NUAN7jvXmBK
1g7Y3BecmlIos5H7xSfiTSAgJmoCmA9PbCwuQZoLenz6COijSbwlVu7g//1FjQXb1zMAMp3E2wQg
RI2myfAOoxMIPLGNckZHxtzAdl0sZGVDS+1kOcsLraoFcFMcupaitcXDPt7NdHkn5adSfOyWORf1
sAP+YhseAcrgKNNIOwi2/MD64mF5F/8+VxMryhHPAqceFu+/yNlN5+Sygq26nkzEWV5gedhRakLI
gGLW/HTolARK3CRVCo/XLCfQ0nMxrD5NzFu91kfr1mmu+tHjvZwnxDOnvTKP82QMzihYcHDm9Uj1
1wR2SRR61hqSPLJImPmby0c9jqqxFUb+iBPYikXthrE411iGbP9dm1FwTL4xKSO/QC3aNMIKAxOq
Li8OLTSU2WAssL4+GcnvtejKE0pB9QpPnbw6ZKzt2pwTCPn1uD+IYhv4o8uvi/WJAuTm39JkpC7J
M1Ot04jrHdKyiqDfjURyEeq3sB9dMIKC4Pf5kY6vD1nc6XCwZSNlhj2wkLvoNTwM4dI2jBUdtkm+
B6k8mR0tvfXRLDJV/XdSOBhhGu7YdbJfc8WxumEeVAfiGgMcQl5tXdq5+aJUaARMRphWh0nFwXNr
fkJEvMNxgHjY64ZjTbxBm/r4SpMAzWZSi/dLfFUAnhvkBtj17q7xYqyZP+EuX9T3wnewoPS66YZz
lwNoelicyDJBmG02vJHYzgxNrDqbAjNrAQfS76Fzm2esQ7MmA85xNSL/S0JSMCEkmJMFgcyVtzim
7u6uQ93zeO0iBVkfvug16Jup1HcC/dGViMQfl7fiBK25yg6YNZUx891xf22bqYiN2ZZYhEKx3rLj
c0yaDSnnLX8tFkK7dqc4yvsHZrrg2ataXsJYY9y15CtJyt34R39IpzqggY1DUjyfc75hWTbyKAkw
F7bJCLvyqoIGxXbI2MO00rkNPQfg1POLzhU0c5KK81L3MRlgeEm17pUyCF/oNTKAWuYRLf/N+Kny
eaOPOSqqKlhre+0V86xwx3ozE9vDpsijaexsoQP1QTPNU1BKY9W373iR7FDQVy2AoAsj7az08CyL
S5PobyBbx4NURMms0bDw9MhH4JUvCnK7hiDfDr31CjRkRRRTCd3NRQ1D7Zf8Qf85kk3ftCUh5FXl
fXN46ifP9sqVCkBzPcMHiVs7KlW+bSUK6lmSQPuYvh266kS5O3MAIZxJ4HpuPIe85vGN5fLKCIlB
UeGJ83cmz1SVO/SpB9a/+EfHZMqLhWK3IvAorialJc1TGSbZPMW2YBrgPLC6a/wmKRFHyJJbLlep
8jw/RDFFfIlgIUm9QZXTUK99djx5SoIFOQFWDxy3v6I8+C1Zcq+oRqu8nkH7yCQ9DrMHkOQFbmWg
HUzLIYy++frRtaK8fAtYRgKlIBZiPRdLE/dRZdhFUHiTExLssDekVYOHTO0euC1tiPOFyU1/S+lr
HLdxhNxvhzoLDC2UP7XIwKz7ESAMRiGkd0iRoa5SHtkVd9JfYa2dKTqJScNgflHkB9O+7XOCgYDA
68g6dSUtT8CMeR21eSUStZPDsDaFCFyOQVtVgD0FeV7tYEsh02JkFHOS4wPj8UtdCRsJTOa7Fy6m
8wbjMdB/1AVnUvfbYhuuTsSeFX7my5mReXwCW4ESzSkrMtzrwIcSpmjsFeO/CqrqTW1VhcKzKMZO
N/thWW0Lhy3X6TAmLLWRNHTXpjnv7Tk2fsI89dV6FcqurXo+KreRgYdx+SkG1J8dIJOHDjeN7EYg
rdKP0xVPzznpKwqULB4XfsHnnGZqz4bqWDSMwcppCklvZQeYnCbZpzySxmOKjBlMAzQNf7fXGT05
TQvtEwJx/YRslB62XXWU74hL3iAnv11wlVq2bM+iwuKpl99BUgwIdFEPiIa8S32GalwI9Q8VNqVW
R02YMuOOqhltw9UJ66Q2MJMW/9q9TcVvitkg6KiMZLHqY08Kndp0cNoZ0IkuIDSyjaXFeIpSGo93
cLz/dtphhoti886vV6oW4xeWTCA9jcous9p3EWi4c5F7dOxzV6X3nNwFy7ZrHLT/uHGa7CB3BxOD
oVSsgCvduLi6lM2fQpgNg3Kd6RzUYS14CVdpFdjzghdhxH7r+g8N9e5Ne9pNJk2ujaQHI0u6hNaI
LsFn7zQ3JdxSXhN0z15Q0A3zdsXLDHKv/jJqt2kZkeShHbl8nxkQryzYrVx3msVEv9b9Sh2p3kal
+RMn8VJc5GfpN9bK6AXlR5DRprKH3jeR3P4h1KeV/W647aUku1qrOZ9cj3uUGf4AVuUVSQBlyTIa
Y9rxvoSZ3dS8pgsw+CCZzzEjuASfKRBPwNQfc/BNWhAddAhwAHsW43X33Eb274AUS5m1Nt/MtFYr
LY8/hzR8TcsIb99DEQtaX1jf/kUVc/3B+eKfVFwrUNVJ68FChsbpEdg6tsnZMZPywb+a0VCm7CcP
d5Tca/r8p7TgLoHm/UDOrX+otvoaJP+KrffywFcRUNWhZTqVEkKgFIhlsE7Lz0B6oQCeOaK/lse7
AHSlEEUm5oR2sJ28YOCn7AJ6u6s+kHCI9FVNxqkgXm9/+9ggO3smb80qam7VTltyr+GiV73AzxIv
i1V2JZ1NfiQP5C6UM1vqv9Ke5yhPRog3rRce+VaHftuyw1/68Pc8WI64ME2U4tE2C1MwcvMTxQJo
JgKMmJepaF5XCXsXOnn+ANDLjbp0wi9+Rx/NAw5Sj9k1vdkmSj4M8s2Sy4Ix6di6jW2WQtfEqJ0C
lZHndMI+c7NRA9Cp3LrzrH7PpmiAV5tG4OgigRMMlhmdV58f11sCwGGRr55BtfGVauJUOQYa8+Qy
QWCx3pnlchMS08s2XvGPou3LkRfWvYIdn+/8tiJWJs5vmgH8TxIFA7XkGJZUevLgfqHRhwivVKoA
Wl/GPVnLvAPG3E7/cRajNsPGOnxI7HG2r+Mt5Mm1DFU/sqtsA9tuFb/M/9xBBmZgn8Lade7fj1CM
ksDYC1s+JjUBn9DOPACo7sIcS1PL1+ecXl7JN1wdF0KU4SLrQMfP8AePol+veQdQb0ezywYBmJk7
A4dIzYBbqbmDuaU2nLSv9v81bgR/8/g24oJ41zmUOZkEGVuaPSHSGdwxLxV37iOVRx+hfFVM/tY4
QM5iEm9D+j6iTkI4rewtWrLdV4wV0Z8onjo5A2jReYn9ZrjGRMR0MapuyowiRF9I28HEcsBzhV0t
YouJKVRdxHEE5P6q3SPbCEWx1pcQ6rFZoRKsvV6KAmLlgChl0St0bEKqqOIgojDGaJduAluce0UC
AXAwxbfTy27zhKli4XRWCj4ii1u/hJwVlIE73NjRnNSRTv8QqBHkKnoVN1Flzfqtv70Py/9CnVFz
gTXi47+R0JgWPIFZJgzOehgy4JI6prDTYyEkoKtd4Jn/lfdbm7eVifd190/je8rIxEzTJ4FUkFjY
3+fO3Zfkr2J+nWFURrDBIL6647p0TUBs3M5zaXIWiLIH0GHjd5t/T5FkDlRidgsrNFH8b/UBhXJ3
qrkY+rs2IqYpJlUpght8EzyujFAs40CBFje2JQv9QXCNiVi2CiCXlHFbiWvypWBSnJGSRmD8BX+R
Rjh8lhgL8/CzwqlzakFZ5rLwmOILFPPtKieZsNfycQIxirZOQLmoqUSQ3RN05VrqKTnUSGVkJncC
wk7tVf0buYO9CxLvADqHms2JotGLveTLYcOPn4Aw8miaB4IkyAtz+ijSrqdUDKFb19aBTiAGSYXp
n5PwZr+CrIzCQQLgWiBQJCQEJLanQq1deX+Cq1NukxgsU4aHnk7AS6gPDkUk/TMx9ngJL+o7PAMi
vzsRc6uFrLaOT9sjBDXd39/RqYDLdOdKZhOWNEUP8/XoeM18H/gT+ZeV2yihEX41q02DS0Uffe8g
+ZHCZuKfQvFTVe1XczVFzXhdgdYT4QEGYaJCM/8QTf7jVkEGf1z1Am6tDxKez8cYkOu7fzPC/JA1
uN8wpAA9sBFpjMlNdR7r1uF2oUwU9yqFPNtgeNluhVppM3CVnbRwxz/VVcWpa0CuE+EkACaLud6q
bN7LcSyA2kF5fq4/h9Ue2p8J+uhI0IBz3x+7AdU53Wvn28qZRdlSqAr5k39+VT2j7pB+1jB1aaT9
0qOaAVfR7TlFc/o9hu7wJJDRSE0B0+qJqQiPhsjIHJEF85eFfaQuV96p6dX/aCzC2WJP2p76uL7X
NUNBM2NUPj9erjPaVCSgyjdmk+++VywBVO84/tJnqaIR0qhzIne7pwSOfWygU/+KUxl/akerJfr5
e1hs7DkbxEKNu9vo1qGI5iUYcwFeQjJVE14z3Cz7JGbh7xx7HkIvzvwKUFDtMiI0of3wNM/SNC0o
YzThsNbofwCsDYiNx1umJhvLqkxESnBGU9nhK9Qu21FXqIvNndVOSRDxNsr6o8X7vf9fWZbuGyua
tKITTGzQcNrIGIvAtsCseO+rbC3qzQgErmQ8lKJC6/sjZRWrkU47dCLNJOhy0R63mniyc0oW9lVE
uF/L8PIx8Yp0TanMeSEZHBfkjwyscyKnTHtitr1H28TuJmJS3ZxU8oH4Z1hg7cn7mC1OBIf5yZLX
BNRoESEtnnpZux74DaId+0n3uETcbqnswYitsORaOyi/luCWYR41NEp/uzF0zfRFVOvGLSX4WH0H
Tm+04uolIe80+fHuRd9tfi4aN/77M2FTecHYavhQciBcZwYJ95JBRSKq1I4p9ANqtgwrgJrG3g9a
YYluzM1I05PwDzAMZDYROPnX2VUlp7jur90Ttlk2wtOVu4XvjCrZ02NnQqyHUqt1R5DGLIA2iSGj
1XUyGxM3lBDcUTY2qtP67Qw8FWKk3YQtqnjX8seTYDUdU4Y5qpo/Pnkz+vj3WSK5a0o/jxUZwm2N
wOgLr8BVDMTj5eCBArl7In1eOlHyP2d3qcrRD3g9ah4nEjGMmmU0Sti18UnbMoNAEwodIhtRFt7p
KhLrFIWNKVOph69zGAx4idtj3cqHJ/ku2Bgze7/98I1yLM9LO7FObFz9MGAFJEF3XEHVlZ1Dr37v
G59FBTVloynbD5OWZrQmcl9XZnRvFNOVBW3Cy7Q5rIerHvQGcZXpanRtv0Y1cmSrdl5C55vBMjAy
wqEOY5CquXLWIsqQsm9hoWKj9+r9wUFiUcEZCGB9Nv34+GfnOLlls+c+A9DGG/r+BK0VnxQ0Okwh
8w6WEd5AvkgP3Mn3K66Fbt/bQfhCns0vNQk+fP2+5LIlV79hiakioIdwdo5UtWQlSQmhJstxvjoV
P88Wic0tTQ9pXVPlsLvBra2OpnaK5G2/XR/kQu8l/uuflaPyHsH2BOGcEjJvT30orcVIMBjbUy7y
AcSBT7NLhyi+9hdSFeEs/OqcUd/potbqulUWSMq7UTVvoozSdCYYIHWJJ2pjXywPI8IgNPtBF0BJ
OZMWJ6eRRyjBVaF5K0BvnDMyd5g3C7jk48Ei/P+ZJ9q4mPLFcALFhefwJOGApeXYPrXbnIWYFYTN
iL2yOV2t2LEYh/i4x7lEoytH1CYn40nshzKYtVmDgOetdL4LjJNNdUBbG+Ofc1mLTs8lBT0bYYXY
Nptkn4eq21mEU2U7sWpu3a19gskcVhcuvExeeiXhQk6q2zwWBz7R+lZvbpUrOI3sn7Ld9t7yWUy3
D12804M8xSR/DcyzxK5v8SQtkDjg9PxQUEnQjM3iDcwD9sLshSja8Jl39R/J76GLrxMudvTVwoJB
ZUHgfSx24yK/vdUdPWf6GlXVIR0bImFwM5U63QhKhm0N60do71BjbBMo99Lu83wbpfR13A4Crk15
11qYtVVibP3WvtaL4PPene/jWBfGrrqzxrZPKp7An0g439VWJ64t1u5gQk/ShHYAUUz4s9yUyl5f
O7w3uqvgl19C12+6l/T2KSYpPq2rYAbBvEOJ9sK0FqyHdjdkCTFwstrxQhQzrXeJLqYB8LqG8weB
uN4Ahq1Law+BLTTJQzMq6qYWgf6sB5dIWypemMQW4J6xImuLI5hc6Q/bDLHlQACROvYnEUHUI5I/
267xCVVy05MR1E3ZrA/zm9Zz+uZIPcBoDf/H8XnTRYqoaxkH5pbHeqaRi8jMOn64mcYXi0kaiJsu
soONkkW71nWi1mYjn3TNke5jBLqlf6fG4UZsZgNiemBrXhZ7n5zF94/or1lYeXDPbsNvgJWTFgWr
ySMcuFl0ICAT301WwqoKwJ9nFeN+wC4ymdSjrDPuH786aipGkPqV4ZAAX/ttQZO6tQ34IVGfoP7V
tZJE0Ed7I3uUtk1x7lz4vxA2Lginu+mQFhuoEuNAal3JEn/S0+VQoFp/NCQrfpka+Jet057Tfy/s
o8wrRiAPLfKwpXFbMIVGycIr0he244xsEgyv13XyoozFiOK5sl3E0Q46meIaNtCMQfIRvjPF2RLv
KFMtR/D/7ewO8GR/5Z+F39rucTGOxKN9aqfHt73RGPDgtAgETFVfZGJfoqPcP68hv/t5IB+3949g
O0vSr6Rh37HvQzL3kd3xKdHUv/RHDmWdLGjlZW3C2Nn//RK/SGRuVL1GrcmhA8QMCLS1dJ49hqUo
stMn323KnQ0QU/1YpK1X9iI9ihMKE/2d+QQwy+J3eTInxkdkCDdIdgcCmkgtgcuiWPsrMTvim4Qz
kajSblojKUfTbmHn9msP9GkKL5M95fBBvu6e79oyF53wZnY9tZVOIO1JpPJG1BTZE0yKz5taf4/3
ROPorBV7uH89/uBQVXG1OyVyDC8Jl+TDgrDr10Aq8N2qOoKH7YOuP6kqpFEHpEerwSHWY6+aGgbu
MyPqwnfSwPROXABHXAnYmBsGVd7mXyfjDa/oHQpUaFVXbbXUVEz2KU9NdeMyUxf1VEF6//GSLXOW
u1Ob9SmFRpHlf1s5QG7Q5KxE6kCbM3vlb2oyU8LjU7FEU/5nf/PFPhYzFDp7ABWvNFYAzMossM0d
GIv64ymUHUtMZ2HEQ71vY6bQtV0d1CGSDCaySrdg9CGUKPwJLv8QjQJdcOL6M/OjkXhPLfUbT2mT
WJJHS94b9DSKudyWHmQ2Xkmym7CB/p96NwolD7x68K42C0+PWjc26kqPIpa9XczgF5MSVlmCW3M5
eBe/BXOsvuz6gEehs/p/LL5NsUZ+qFKcWtccPshwsBVk7xlUutU1TXwp/qdnAiaZ9Y3+1u9xeUIV
nK1xv2LyIdWiQm8isBm53POCr09h7IKSwSSpoGGtdib5enYZPTe846Kfw5BmFEEEsaLKeJYMAZM6
PjjNhnjznC4zM+P+1geiVFtT480DR/O6YWfcwxbXun7At3D8kfOgcHF8L2LGSExJuCMqyOdYZdmk
4Z/5QG4mqJ3O1B0pkwDkbBLe32HSPmQVyDgCjim+bF25PT10LcE0kWPaRYZetwDjoKLQbxO2Mxk5
5mgyp7SLP+OEDfR4WDGzN2/NrKLA7rSHdO70tlMfp4LnNa+K/8h8rASfgju+/3l6Z6hMITeD282S
AkxarjMcDIG3OViJd1j0P0Btk/6jwV5Pp/4u5tiNPzEsJDsEYlZ7FtW/7Z+Ry38WTUNg4bJFGdtS
A+NP+feM/OXukclM54PKL141UlHNctQ54zgOia1vLSUqnLcyHwNU8SW0EcdPgnbOgTNC/KbKXI9C
nXudQzkfI/y43UZFjT55ZFbkAAeiRUllyK6Q0FUmlq3+WG19yS4Hi2ud0bJPy2hi5poGB/+Z2REP
gRlgV8nTbq7DO8m6hzqS2I/W+v6KkhVzsD1IQp4rD8Lc9F32RdRU2L+e9tWnyaZDZo5Gz8zyZxCy
V90JCJz1lmlfJNLebYOyCK8mFdGh2lhoJdSya2N4vhbfdG9zK8pKxB1TXkAt+vTjjYmKHSwbr5pP
07Ln7j73j3m4qqtOqiMFr27zIkxwmUK7teISLzWRzChJ1F8cfGiuHRhQ10bdFd3ugjDg9QLz5mS6
s+no6OwxVXftIx7XB30wc5U7MqCggCezBJBO0El9BSzO9WyycZrkmsucAVHOg89iVllyyGKs/9CZ
0+OoS4kDJZNF+HTQAXPB1oMm6sATG/x36XEFKDX70y3Q7JssX6hTtQBiFIBtr4ZhJD/wYdTNrOPl
U7FEZCjyZrrAiARQ0zhdNZOajn3zr1OfM0PMr6lkHf7BGljtYviLJKO8ylLCG8HCIGEnMt8cESFL
QgOqIlCSqp3olkPjIelaeOZpZlo7vOBWCrUoncPuXoyOti+lFZ/g6sajHa7mX4fqw+wilECerTQP
51ZEcIq0ulaZPb0ZJxwMMtAmfrONd3wNWr2cXyWbbX/j+t/KveVqI1OMYazVghkp3bTHU35lBlR/
oDzEgMEP0wxN1XYg1g7f59rom0y4+L12TQCjmeyeeSf8mUj0jTD3xvq+rkYVVzILLGAlxj+sRgPZ
cOMUR5pMAhzUT/yTjisNKzUbpvtwtbrFBLXmCUDbSS83Eow3z20f1oIT/6de/4WYW2NDekQL7fWd
rXCXI9edaeY1ti7f+t9a8NUfw3RJDqRSsGlcBz0ZwzVLp9cIV1yGqqRRs/HZoYye+MAvOP45GtHq
+5ZRgJAC9uapQoewNbScsKED4yudbHuhBGb9VxfZea3SZFidbExx7wi9tO5vyX06FBJyMngpeQxG
RXu5xvhmF9fowDssRBLCepZLtaDPhJdGnsm00/PEf/1UU8K1MRLn//7sTE8Dj6ECJDAT++2gPt/8
U5pRqhHaf2p/I6+uxgzUMDorfSTDW3OUTVWr+KRT9hAMpcdBe5zaqs9nodV+8YJ94qadKatl7Tfb
vIRYhhgXkWmlyu3PO68jehhAeAnwIE+vgsDv/rk7fPIZzZuqDKU2fBfUDdbvzKTLLS4vT9xG+7Zr
Tb4r+guK5TeCF0ODJ1L4N364u+7+M5YXAcgxurNqZ1haqLgWJqk3zP6oFhou/9K9+cRpHmkml9gW
s+vaNBVsMdoTDIIFpwoM2MjWII5j/jrFxlmWJpgNdeDBK+8Lq5pIlNPqXB8cqpIusopHvVnk0cmJ
mEAntvVcIzB0vs4039lHYP+WmJ+HLYSIXvmUIKd2RjdhPyrCvsMJsuN56dagH21HfVe5SDT77QXL
sumMkt8O6HztcYGzcgzqaqsfgWsA/bjPw7SGiDthd31Qe18JKg3b5YUMBHWiI9vRa8Ew6GknfqpD
ms7kdABxJdIKY6dFxeqHVqWGd/alq9PA9Pn586rVasFxN9bFuWdlgwASzmvreaDHM3lJhbDWLlF7
HtftnZXL23JPztubncXENk+/Dre8GIlBX0xF3cYA6BFm5OH+tVdwiUrDI/9W1eNLvuvn8PwWXs9D
OdeHJJKGVyFs4XXx4a/h4DOsvZtsWZY9DdTdAN29k8mZyD0vlNvHvbjG0c5xWrMw/kf6htIJnrGA
240Hr1C1sLkhEBfqeeiaGhayo2QvPcElW6Bv48MDSa80Kc030gBQMveSuUtdSz3s4wujgeNOR1lu
bb1BJ0klgObLuKx1sYkLcuAK7AgGVYJCqoadRZVYNqtbx6m7kvS4eanIz1MdhouMe5V767KYOoT2
hGDrPZG3Km3s4irqJEBEKaXoqv67OsH3fqc8hWDCbzJWvXHdIn9W9gO1UQhgb8yx03A8UjlXASJD
f1x4rYD7L6SfQo1gQOz7MrcmPMV/tccD22cjHTDvkyQxeDWYMIGJ9394lhegTzTVDmOWNk9EZB7S
ioIrN4AUJwCg3lYwtlA4BNjIMvbGnEYFmhLKqH9jqaq6VEcsg1A9iW3tX4b8yOHjd8RPJu7nOpmB
TyW/j+YjORrsYBL4QTJ5gt/Jsh7bnQOfRZgpOhKLoWYauKbe2do4em3THVucPEXWA7BZ7HzXgooi
mPyHwMZEI3IYGBghU7NoEL6SvqDbzUO+Yj4qq5kJxGj8sRTdOlZjy77dvjRhoeG5vaA84hhrfA6L
Lxyl1zqdxx4zfFerS/SVP3QlTdoqjS4t/qISk1GBW+thbqAXDdNpzmjwN+3ODOMuPsA+EE+2SVxU
HGb9lIrOsAM7QeNAFTCUBXIFFp2gG1OZ7L3b38/gzmg4IXupo4HBssuEGEArPwUros6PLYc33HiG
OWis4MKfbu1Hp/n5rgYQ63wtT9cVx+AbtC1WxYAM7G18lObN/sVpbU2gUT2n26xmwUdUvVftAby3
eGGamz1Zg73+/uCEcFg8hWCDUP07TbzE3PBCUGx5MGkrTt+7A4N6UqKZtaXfcufQ8aSk2VO0YypN
mdEuTYKmOhNsD3kyc9Sn+boaZR7nzffZjadGoNBmt8xv4Z+JJMnsnERytXdSlaL0iUEq3llfW15g
lQSM0dGeicVkmM+GijzX4Q4rPVnligtZKpYTeeHa5rX2KgDhQ6oCLPT+JEgJ1Xu9qXTecCgtn+Bu
IFPn7jPsLU+Oba9mxY5sEXk3ZbFnk95YnfkYvUhX8W5UfwRASd56FvHKuEE1kAvS+vIbWjoUYqom
wuFXVTWt+ISlgc1IwDOKlMadaDTNBNVJHQzQDOX9GjScWw+uEY2mZSm9fYWnl2w38LgG8V+oyTQG
OlajI54JifnhNnO26IJnkgnEl2n0AfZ52TY40qwaWx2G/zqzGFd6Ygv/sDerq4/pawdQKBjy6bEu
pkgd6B75NHQl9uxBX0A0+pFrVA43Xslh2fOzYcgdfLcg7ENyvsOU9lSR9HH3NqGKI5AQ0FgrLzoM
NiHLklv0ln3OXwhbG36rFNJSa/+AT3w8/gwIp1wRw9AMdQRg6YIUJpJPHIFq2tXdqL7cpB+eTD0o
Qc6zo8IHwrdYvzYIPiMK+9g2hFCm72EVDK9XsL3bjcFCI3p+nV50Tt/pUQQ80Zu4X8QAirUeHcrb
zgEmbNUwhLvSsFAPNEUobvwttlmBtLmCyx7Vn7o2gK25wmm52aBvhrtYzgGGF9dHQOPoXF4A1ZWn
64Jl0GwZMHb1ZDD4zSMUkcA6c2bmISjSkeMJ+Ipj+coWIXkVsxC8Vov2sLeOFvYQjaYAGMdlV4Dk
Hi6ssn5FSIt2CM9qDr6bUe/Qb+tTAhGASFwIpMJxk16/igOUE6Tc0kK8s2jFIkzrqf5Dlz9PooHR
knkkK7zfFXG7oO6UBcEHPB+5hFnZP/h01ogyjbrzWfDNjFKt4/WpjIp1vHl7SXMGiaz59vEw4dA0
8vc7+HLM7oXP4b0bLeSFBRISilzQ0n6ZLTJjuKJm9uRO8/1V6AgePp+7KdMNFIbUqx58rV48A85D
V80YY+Aqmr2f1t2j5RFVqlapm+zWG0SkPmZfaGEXV8ZvtphI1G6LIZMdXrXBnrbRqc3y3CoSr02L
xWpnxbjD/BVAALRh0ucZ/Azn7szKqwWN/NwYD91aAWQ33TSls15dodBwzq83f6tUzZtQXfW7OcoW
5z8RTM1yh/aVFUGAUCBK/DMu+Mt59BwPCvXe2x+nbxU2ywlg2VYE9l5Vho8FIm/pWg0KqNFATE7p
ylUZ/yPk6JmP4CtDwZgNYag42wnB48z6IYPrbz/Ax98gK8buo3IE3x581Tpi10I+9vz89nDVg72o
PaR+SoDi1RK9bLFqAZllj226tYXnAtJ+ta2AWfyDFLdfm2XxZosJGxuQQK9FurTPtmNaBMq2rA6H
8StikUBLzr2PA3TFTAqC7WIy27/sifSvFYPk2aMYQZ5AREpmf1L8/cMxWmznTX94cJ8FL7wI+UHG
+mvv/AVZP3WDfjjf9Lu705tz9Y+BR+WIBTh2xM9IwqSIl52AKFqyYeLlNjn0efqyJSxg3vviBY4l
2kcpbbjqqVhsGK/lr5ASm6kIJls4x1S5u9egm4y+6PpY+UAhxO9vPGQiOUqislKaFHr1guZJrYfA
F/Mms21iPnl24TpyhVfhgX+xokPIGbJUcSVx9aZGNYVYN0Fya2RMmQ+6Nau2D/M5MTA0h+xCMA/j
dSlWvvMCi8FK6zqyJHOL2TLpUJMI+L3X94NsM6axwaC3sAUAXKAfYVC5uJdPfvGVn6CUdD4sKi+9
ZL27aJbMHR/OAr8iCIuuV24F/JBcVM7pgOXi8LkPGQ5s4HJFaeDWBhdvyTikqQOWJr5ao6mufg/0
s+3QRMlV/ICsUY3y/JgG69uycbweP8Q8DkmQstfhk6q7ZiDHpDfMx3Wp+ySw/FLyXT4TxGo8I9L6
A4+ucWuC+e46z7IldxEZqGM2NEJBgVyGG3H9BVGDKGesFMa7tyNzYHKpvHrBg4yvD9bDbf1EefUr
qYuc7ZgdbofbjwxTZtSa8beJh7+Xp2aMcfSheVZtIxbxrM2i04QRH7Oj5EXwMDEdxs5TvE/a4OQL
tJG6jG6DSDafkSbwx1FLojP0RYZOvmhc9Oaiym8la7KfaECzswL7mL2s0HvR387z8dx9+QegZeBv
my+9sCxVY/1xrj7SVl2SX0D0Bz6cIV1qn5xg4zp/34+SzsqcPO185GFiHiPM/zCbgVJTPWOfDxSc
wfWDcgYhsuhGzwGrGlN5ItWl8jC/IA9Xz5UyTe5ssbfIotyplGksnE2KNh2NgpkOz9Cw/bG9cRRz
G/4vkA1qTTylr3o1zDAYYRTvpKl/lTnPwVFGHtkCTdMh5wWL829oiXAv7vih39Eo7doLXAxDRXjC
PWuVnDeyA7KenC5x2ri56uJ//uMkqTU67J26ZZMdbuRXQFVyMDJVir4yQJxBinVQtWKL5o+KhcUR
jmWlBC7+4rhXvWrOzxOIwfYZzmBqLbcXB16DFGtNR/swxE8RP8I2RMkC7GH8W/n+JdniQ47E5UOp
IVq7UiU5jMW7V08OHhr0sQ3nmvO+zSU3in0EfyvR4H2kn8IrIPTUbKPRB+6nWW7NLcdHAmeT09c/
qzNuDqw0NI6k0vjNhMOtl5dD/odOzdUctU2Mx9ws9RPAkEyYUZOp3PrvY1rvOQeZ2o3M3GQ/LaDM
j1vmt4A9NA==

`protect end_protected
