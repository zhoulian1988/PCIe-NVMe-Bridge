`protect begin_protected
`protect version=1
`protect encrypt_agent="FMSH Encrypt Tool"
`protect encrypt_agent_info="FMSH Encrypt Version 1.0"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2017_05", key_method="rsa"
`protect key_block
g2jBXS7FWsoQPpRnxelwhzhjXHrNpcvmqFo/3TXSj1mUvdQbOSprN2XrfBlg0hbhGUjivM3UhwFT
+NNSI2EET5yEcaXnPU+p228rlY2w75G2EMnC+ET1eUdEVZOB3a5FcKqsFYlwPljC10AKxseZku6r
6Wtu734g1Eaag0F3iMxEHqfR1xDbSyb8PDjTo7X8ezrmFkqc2c6pRXnr68QxTqjozlIdLpknBoRT
Xtkd+6Yd9H9FBcGHc5++QJT8d2TrvYzS2fddun5WOh9tsgfihx+en4lsECgjuRbcZNLByHMVf4P6
5Svwptajjc17BJQOiUHVD/2IvayJuIzYrHDAmw==

`protect data_method="aes256-cbc"
`protect encoding=(enctype="base64", line_length=76, bytes=133280)
`protect data_block
fisjjlgaeDUieazJWRGAJcuU6lSrB1C6/CzEZu/3VbKxCAVN78PMmnmoZ5Ng0eI4JJtlK1Y2Hayz
POzPCAvsh8m2vvbQffCjviaKa1P+UErImlVKpMsq38z2JfcqLKlxmtcAjfET0XEFXcq+GSbb8vc2
rs4By+/bgpAlBW4IhEuW1qAqyVROQsXg1X9KPyqxzFO+xBZmMZXvdcufP0mxo+bzl9Vxo4H3Qb52
OExcf/xNlHEPB5wnlVep7EGpgicE9YFd64YyPUpwmEtIaVtz04h+7fl2qQscK+oTPIywLZ1wyLwD
yivy7uCOXKTJU8kR1XGSiKSIzuJWdML6bA/OBCUFtHJC3+ivmmAEXqtipOS4ytYcVK4dhtLBgwUF
KEo2O/AEw3HRrc8tvhHLSE75zesWxHPkek4EaWh2KbRoNrMXeDxepX/HKXI3++cCplhbK7C6ZnUY
yWb+mak/RPdKWm0h/fQWdW8HOsEbZhTEz0SXqmPPStgkBLiqxDzJ74QW7QgGDOfpGC2xRwRDBvYA
oq1PPvrAJTZlnEMx12CXl2DPq4bmTDvs7SMN70zJtzhpU1p0gm6e3Yev1k9bf6hreKm5V2SvSPXt
eAOC4lC8kWRXyx0TjyIHOICtTjtYQ3WIXFXZgcpYzHNQ6ltA1gqlvMmKULx7hmrfnAEfSijTLuB+
ZLGRhGokPgjFWESEJSs0dDlXTZhR4VJVuXGDHUfrPz68Z7VJ0YiKflKam+kMepnIm5QfozZj0b1n
9g6hi7KsbdGIoZAvEbFxPosITkf62sdV6DdANIa1dkXIplneoF0ANJweE2YL6v7ViG1MQ8nJPC7C
a5+jlJxxxQ3IR6hBp+cf02c4k5F8H+vOwcfXBs2/fyel1EEkKkBxuQGW6dIpFt9DZ2k8/DE0rBmt
lhCIYQok/enclJnZwF3zEFVHzgYenpgTiDxiKFoCfuGLdgXxKoysNgVav5A+Ds5wceeLUuil7c9y
OeK9rvSZF/58DA7r+xIR/s/Flz2eG9E4pBCsJqbNcIJg3PLizqM8q6MjT6nI9eKYa4Ii7aSm5gIv
KRwb4JOzQQy/9dVJLk8dxy2mCDKGSYK1VlBwf1WliKT4f0V1FigSqooM76snusOJ5+j0GZ+73UeZ
43VyJ8yJOEwgEAftMlfyQB0ZzYZz1QQKXbILXpjcpahALdRWM+eNMqyoPtteGhZwe2A7bFGHrTAw
tvwWF1H8QaG5m60NAIIySMbNeTCtcL8L2XF0jHJG4eEKwKYEo7cCJ9PEvFa6CzNe8IeIzf4Wey/d
/+GEOxqaWL3xF1UilPb162pgpIKa8evWtMsb+yMSAs1VfH9g9BC8FWutIqdOYLaEtJpj9qG5HGkg
dAaf/I4EsuWY2gDeElzDmS2qCNwfYqKI9JdYU6MDj7agNQd5nay4FIRuIWZqXvuAIWhsuuaaIaCB
bhbt2KfdYGQRxdXnUgFjYqnx1fWMjVnDio4GJmF5YdcEqOIErMXzkOaZox8CKnDCslFMl21shAmt
oveKNnF8RBkUYDebNCoAeiS5FUayGt9Rs50zM189muxe4ycVq3NnXQuZwuMPJMIO0ZWz2JjXFU6Y
uxN7zEQwgi7/y3Jh3DsGSWt25hdv7YoSjI6PxBaN69Q55cu7OB3ZYbdg90TEJDeNmrZW4AgwG29I
CdgcgYRxcPxMxzP281LzLKV7ESz1SomrfyPqtJ9g/jbP9HDSS6FL2i0CEFZABhBSZ8TCDOVUVlxg
NCULqaPxfBGTfC43V5/8DzWnT2LU4bZctd6QrE/LFNZrXWarTTli0I9Qy03J7xnLzsrr+YHgdfks
zGcM2+qFPExu0QcF5i2oR7h1KvS0hR18OFON9Vg+7p/3nPxBnKFMioq//QqEdei5jwp50OtNYjZz
S7VvfonXtSX/tdWb6hFVAgdlup4/ApoOeN1pYTkwksqYGOdoIQGBFB90vaB1DPreS5AmrCNnKsMM
sOEjPgumnp/8vYdtzK26lsTwLfXqqukl0Oh6SmWZqs2A06rrkO7jupFigGErP2dpN4mpP2oyb4lM
mYBH7MOCKCmm/wiqt/pIxhBJ0qIUM2CnFl2aZOpwkXBlbIFGqUfHr4yWVcMXUEqE2nFMvxRMQkJV
VG/vFviiCQWBStsnVjTdfCm3pcMlHW1mn3J7CE9tXrIb2RfW2yrD5b7YrL/T1wmplFHoR2A0pwy1
IJ88Rt/BZuRpyknq7K+7ZrkOXFgfppeBK9UWK2JTTzxWmluipQpEYZ4qwsOewj7OeA8tKhKaUwif
u2EubjwG7ncsWx+4lUjV9v2sY65DFKwD7z54jw1WbuDv6vjRXGjaxMXIFXMBXT66U+kSeT4yQkts
YhN5bbJ3jPzoOFc+gPMMIkQhur9yBTw/wDjXn53vyVLlJPuZGF9Q7Y4Vxve8P1K/Ih8cVLNXbNnN
lYv0gf3LJ2nDEmpZneHV67TtImyNbB5bPVzb5t6E8BFAg/pTwnXuDD9Xrkbl5okZ3Fm2jgcQcE8J
GckkZdoXsxjOsF1kHosEnjmOhgVark60YvipYapnUWJfoDCc1DcZcxqGxgpF19AE2QhhOm0WP6Gd
2IzSVTS/i3Gsf4kU/raLXQqilgQen3lpGyfIeP6u1VRvrDXvDH1JjkvaOS2+LMwS9m+XSqXatfgq
STdPZWjhvaxkSttoFbu1p5zrW6yJu0l6xeI5edafPLUyfpzZlcT3NQ9Sp8dWcIhbn2emI9f4h7Lh
sdCNINU/gXLmqNJcekA3UeVq7Tl3v266XFnEGJbQ74Bl1FiXXvGBqiYGuza3oSJT90N2JxczJmNg
NqtIrcLqKPOqne+GVaQ4/WO8C4qqE4s70o2qWDnXH43KCzQOmv132W4TWBCyXC4Srzjq10sbuQqO
qUH01sK0P0HdEdaiQYYG7qemuIZn6gzsshoi/nqx3MkHWl2aYOFolrnkSKC5/x30ThTfbwu1HF8f
fDNRA7BX62oDQ5/yGvhUH3Y6KXxfCumTljKxx1zsjg7td8Xx8sAfDEpi2J/8r9od7NlF875Y/mG8
d13Sk1jAha8F882A2zYz8SLooVQ0fa22c0Aj0ZKKMa05R1YHVnEGL6J1H5RYYrvMlFchjqe1OOS+
1Oi7X+62mK7VCtJ9ibnoMaRqVxJExJj2xso3+fEyrzDUFYE0be+mZ1sBPWD3yU89WtbeqHQYyuO2
HoFoZETNcqehM8+3Snr0EYKoA9iC6nnP/xz8eIeumIu2x8Rwo0Rk940uopvrEapwbmS3V5uDzCPa
0G5ZyHmNCOUsKREjTc/i4qO+xE2V6QZLmduoi0DSfDyvXITctrQ7efp8GxuSU0OLqzsbi7p+Sohr
TLUelLE4b89bHqkDieJkCtlmCvjzGgrIJrXEX2RTpvQuoAtAd0rpoi1qg8eYw8S9LOdczxBJ8R3n
IdlrVvV5DtWTeObMT3uxQa6e3ZsDTU39O0WfaFFcWWmFqnMfyrKdSIRY4plRAUpuhkYC1wR+woMC
HZEh6ra6NLqgxXYCoWDGT1iMDpBm/ybO+n7qB361w6uop0EgGx6bkIzjXRtOBUarkFR250+581XM
k0J8eFX3WS2Z3oXqYWv+JUi+43L6kaAWrf+bfyskZuI8yE9Uvj9v3ygvrT193spbjsWhWa50bC9W
Wjy9yQem6TM4ffkpvZq/a/SYpMOkBPFCrz3rMZUmpAzxa5oer8yGSTySHFqXzpNzqkIwnvL7eJHu
7KDvmEjCAZhiadI49d4FHbapCYPtjzq/oJRhyfaf5bm97aZGTgA6DQxDSV+pKax2DhtzF4yni/4x
xkOJc5Y/UtMpexZ/rLQVwuH7qRxDTon1bcqhl0i2HuSPit6VX+DTNMVRWmxL+dVgBdMBOU8W8Plc
75ytl0mr6hkYEEX2OjgqCvuniG0jLSBI5Y66Hux82YvPRBpCglHpIg84GspD68yz8grJ1WRDPlsI
EzPSllRznKyoYSEaudnwAAJA1ooO7euzBytWzs3tbvxxkgf+HmiLKM8IJmypDouYmZolzQKf4s/K
c/Ss2kIs8rXaTbHIghni+yhAyZzrDEQ3Xb9I9ErL7jl07H4G6pwpueeS6dzALreIuUMlquDxo9sL
4jG2kNzYHV4FgM/QY+TnIoFGs7bTyQyHpbf03Gctk0hSf/IEmq5wfk4ZLVCtDdRa8GBHUZVjWvvE
wGynO6x4KyPZMML86ufiaCwIth0moiel1/H8O7l+LxgOmnzdcLF1XB0Wgkzkgxb1uqpsYsBDtKf6
EpccbD88bYNsldgTZC5TH60h5QaVCKw3UH7RzBvtdZDRo8CzS2/hIWul9qXXCyMlYgcEnQAuiRVs
KFZ5LtAM0YciLP/KtYZ8VXMRlsfT+NP/TAVXnvlmY5sv7kEBgB6oRJXDrg8eHBMi1lx0hspOuyvK
a1X6wI15HZS5EVGb+xGULfL6We9qQriifTM6NPtWdREuQzvyDCXVI6+d8b/aoeIGfFaSeAuvYFwH
z6mzdf52QHcOXK4rj5DwaC/ud4DCwfWqU7A6HcFfZQc192+pswFmJpwsMmpkJNHtQmq+ZprlDQId
mGl/S+kBO5rOhKzBeObof8jYvlBFQy10ogGkAPDOVCM2TtOjwEOBl8skj0cDV8k09HSdiJ52NAB8
9BrN/RMabTis4+H7VTlrV6qot5dSnnnQWuOaOiBuybxzINzqpp3pw8KgWU8RhB2TKVEwD/07Dhe7
AFIXAn6AhwheBwWs15g/mqEl6L31vlI5CFiPv8HGk9jfUQqwfbKwlsgXxWxdw0ZgswvOolVF0wHI
oTFrJyI8fATweRmCd/iORLvd5gu97iAdG5W9fgZKRCWjbtXpQx9Wl7xy/NW2ZLOfMwcbCNM8XAdJ
fvmMZhSRUckO/RQhFgLPe9/AW9t9ULhg13Kh2oI7D+jvLcQkTbN3eUiBEweiEBaAO6Nb3tB72tX5
LwFGhEcKz03J6FlnXWE3GH3QqzdTic/oPaEo3emQb0WhevvwZn+PGY1O8Og1j0lazKDRap7WoayL
MJVIc3hPS+iri0PyRKM27vO+RnILMwgk9NSl5YzTdsKt+xYSCruY/9oXtlINc5LJ1oU/Yolmp047
vxK+5LsWeIiJ2TuU2EJz5nITj12WL1AKNQF0rkM46Xjr5zOv01J80dIm81i4fQRHw5JCQ01Qv7Y+
kND69XdchFyuWqUcKV/edGzVl+9PjHY0LoHQENcK4LasNOqQhclplI4F9u905aHKPRhCppU52njJ
IPZlDu1BPRHK8zhj/WB42gMIjuLsAxKx/9Dl+LadZ2lG3YBKoLZxCctGsumnpLXUsTgCreAiR242
0SgdacJUqUgYb7HK4eAXXN9zlLVT45n9VF4I0Gxf/PgqAcdkDqpUwd8e6+LrV41+BpTZD6KsdDXI
qjR8D04HUC2V8+71hn/r5HXK3gsRjJ+D4PkD2uxTk8pwea6pymm0jkyrwKuoF53YszU4AAXSllp+
QW1H99Ckj5I2tiMmwMM0DJrHXkshCjAh9Jtta2u17S+1gOqgB5K8Tw8gx/+Khoc/JlSspgCs69su
uBVJDOUbv3eLMXl1W1/6zvZ04+nX1/YwJzbcKJ+AqP5SqpW/x3d3JFDKwVNrfRAe/aka6VbyXFq6
gMWLMijR0MRiKek38UH+j8iEPYYvBzuhVSWeQKvTDKhp2J6PKDvh4ZQa04L9sD5y/tnFMPVral9Y
D3PKX0yIBmiA7PvvkRALCyGIJH/3jk796Fi5SX9xJHAWTSgYC3PD90FlJn57spgiCH6EdL6DUwll
jI+3AAvFa5WCAs7oJV8ILjZTY8AjxvsRVtW1yYU/qir5x1i1yvGPJHHg9lFTCxQeyTu2Ym7pD6xO
XzYqCJD0ZRHWoR5io3E/4kMaTQbpNlExxgVVEj85bNxtapvP2C+sxPMpHePHrz+GPVNyqerW1VnF
9X2obVSafbBZU529oKg/m4KWPB6CpbdP2dklApARBa3bgSfr5+mAKrJLKkqAjPz3KvfIOIN/hGUD
TkcVAXt0F9ojttDVIjB+G8RypOTJgmpi+QPKrqSbx1t6U9+90dLmSmItPZI7wINswDlq1XpVP8wl
BMuG+4p1sqzQFDnBSMI+fhOH8nSo4DbGKpgxG7tfnOxudLyYK3Kkp/xhLF3Is4rfdcWEynr0dqCx
ODeHVC7C3fLJOSuwVAEtNk1p15WJ4az9cL4juSDpqEP9bNT2pwWd2UtpaUeYqVSvYaaskfAmNfYQ
5NkCvY6WDcO8do7GR+k5cjJxyCurbjNgV8NSJF3fTzusqmnWtDsuMrz2CpEQTNt3OmXG4hPP0kfz
0CL61oIFmmWAK3EUG15vmaVcvEqXa2OF8toc+dxUnV+5/1Dw40Q87bm8PRBoTmAb/MVEB8oYFKja
/Lp2A0u/+VlkwGW1j+VqpaWvd0l+mDHxriYbQ6g8H+ouxQtQhOCzxwmh/OD6IqZhnxPWhiPTz4jN
mR7EOhlMg8x6JWaB9/Fn8R7im3h8goG3NUO50LPTq92kCEI1w5afSJZZr5HUakKuefkjijippB67
X2wllj+NBmiLAp81sOA5xySgcJzBDR7M8OAVspAE+8Hg5ZKiyCeVP5flERREEhNUtPH5/FQobaVW
OE6sCfR9NEw904ohqLEqMrWecApKV8kC5/5eUk+l8BIWyJzolR5nq6woQNFxmudFsJJcvXCxWMlI
BVKX3+7ns4mahDm5+Z9En79OJ3SjXgWbS0SiNNERqt6Dj0KP6RrNkgKQzsNObfx3IKFxACB3ijgA
jX2dYGCG8JlNO9N4AeBpn7GF55TGxYVU+l1KL+0Y8J3A/CawlY5D2sjY4ZkUAi2a3EQ7MvaQP4RT
iSFSgXFtCSjsXXBK/qmP3C7MERFhSqER/8FiE39rNOva0fkoXlYgumINaSk4/vokLFCuMJQX/3E7
KcAiak1mUyPjS81qsNO3Te5tyVcXsnTrWBVqaCgl2ikKfZHULSL/5EQN8U/LlOFx0ey3l+j+oBgT
I3KLPtZZvx3M9S4+LKMyhc/Ecn/P4IY6c6Y2RzXE7JJCbWfwBC5JdpdKczOrkUsSzCtbBC02jK4z
2XBKvCSlVr0Zw/E2orOhI1BPrulb73qSfh4VMbAWgfaJ/EmNe8py/mB1eQdgLALbKFap4pdMl7HV
DOvCGNlwLGNPfZC28RcH1wuNIjFlGvXmMckaG8C4GagXMwmLw8BkjjBItNvncBb8+p4lnB6lUtzD
7e4oIyXecFSfFYs0DWbCEIaIUOgr+kxtHZgwpqyX5hZUj+amrXSjQCG5mDMvqmpvgxGxKfoBNjDe
d6gJb6EEXe5jivYxEestn9LC7YQKlMqiifjuvYGR2dbwlId3ePk1DI3hXCB7R7xLwCsdlaykXvry
W4bj0ehsd4nRrnx+D4TJYxFP2WtTsbB8T+ElGQijQFEXxyWYHttwx0TtnjFTkOrBjZnPbLVb0J1g
WV4zYBSmXWeUy/YcnrhhFkCY7F/qwPrfxinh9/TOhI833nWki2hq2X8f7wQakmIGWdYPWylcqnDp
gL1CpDH6oFcS+58EjrftM5YhKOG/ZgPuzwkryHfB9J0dCvDT5f1jLr6yjiIK6ogd5WW3pyYZofGr
2U1J02lHuZdCUs+95MC6EAFH2WXWpRXdZ4q8iev6SbRG/33REQEzsVAcIhJ0E9xrZUMr5/ZSTa/A
kCKaKAQmIzq03rOEvfiQkTx0m5F6e9P8pp2a9JspZ4vO6vvjXNDV2Euacl7lvsIQW8/W+hl4oaoA
RA4tQCX9VL08biGwe0lu+9yRv8OFlsIvdLuKMgwOLyzhUC3nxkEmrxs1fmo3xKpK5hXGdXy0pe5O
0jsoIpPu+4zLl0lO9CMVfPrnQKAFObC1/piu1DSHtMLbnNhBR5zoSuBjewEbeK82/pi6M6k5lRyC
QO3sdayo7JsAN/uahsFK4nGhfgD44sMrWwAaSVGMq8u4RaBTdyNRQG7M2eRTJRc408bUpwba0oGY
bxC2T6lklFNz50K+uJ9ekOSgS4A/9oWSNtj9Dnzkmuf6vCpWKdpB9EaoC2hW1xHRr2matiJGeFxX
oa+96JO2YXHJBlEo1Xi9JKTIh5wLKJMV/kyi1S9TpZ2J3qDhlUBzOfnDg9Zo1V8oeO/fy+Jhm5Ew
J6cAwdqDptaU9hyGCKQe7eM2Lyp+TV8+bk/D08aAi+kOC663F4pxPXqaMpP1xyUUeElmM7YdMDwN
ADlnyrUeTSLqKM+iPBbgVoTGZ2w83i5NRKCpnCmex1AyuJItTK2ejzSUiQUgY1AcONIjMuVcoomr
KljfN20g5iZyIF74zgt2vU7OapeWlfg8yvnUGOHCTrs0TZysMYwOYxgVHqeC4VbQrfkxw2tvROHK
cxTOM/35wmajZED5XxaYrVa0T54L6HZYUmKb6VR9P94UQ+oE9LBKlmk983Kfq4YZE7oyPwcAqJof
Di9vR+PYCuTbwhdWwRfwhTU4m5YL2ObXjrpaDG83lUB6Mf0n8z0NCKrtYJs+7Kqh+k7bpfILxFcD
hf4c9PeLIglSHdWvaIXAJe4fIPjiMVuB/tRRyZoP3WZKbNrQscC2cLCO5yOk2RgnAW0NwIrFiktG
1khDHwIq6SwVdIJgDIZqrXVw7c74rmfy1c958RO0ZADoAQzyzlhdG39Ull4AgOlL54C1fd+VgYdT
un6Utr50Wc5sHiFnll2a1x5g3Y9mGMWcKZlRpl+1yjTH/KbzT7MwQwnR+ppELKjKtZbaA37RVSeg
pQvgOw6/cQdeLrJN17vheWvUsNs4vtaQEQixBjaIBjCpPHz4tiYrIklxM8SrjfZ/FHuCKdhMnjv6
5fb2H9C29OemdJd7DWAvE6jLC7V0oT/iBgBjqD9JsjAioMKYiu4w93jQQ6rmqcChAxTtZX7wA7TI
ZjDvX6pVMhlvVjLH8uLWyj9Q6eMOeYpeY+VqRf0T84CskjOwmMSaRVNWIgxrEYPZzFHFHPUYqRXM
83z3DchfP9J9K9JoD+4XhxY5zAeGFsdYVacfFajxKvplvdMHbgm5QLXAflyR/nir6eVRH954+V6v
J3QCgu7TOSpRyhFS8PzfiSAhm8TiHkCXIF6ECDCTJssPXWQKG4uSHuhMPry+UY731FWNT5CXITox
yTaWZ68J5ZPXp7Zi9tozpOHt7XY8cR9kL62ElXCO22ypDNLO+OmDNqbafyb4QzIQgkdHPjYLNa3u
LKwOmcFS6Az8iHxNDEhgjqmfX3SO2WAF0hNXdwIlnqO0Nrs2dB0Y0/cnjMp3uPxxgx6m/T8DnoEw
R/u6Bj1wVLCmfqvyILoDPLHgPnSXckaGK2dP3oqsUTFk21Ryrro025BasGszk8sND9RDmybvIHC6
yo/26ABJAqCTS2W4b8tnLu+ZvNXNxvPtkImJWFiaddiwoTwniE3xk3F5YLyAN3B6zA37GiP09WGq
MiHT5NT7wgwXZ+IHByZAuKnH8/YgEE6sojuGhVhEhDnFBU2l6/wiTCvlL6XD4wk9eV92+Hr/yl9D
iap3x9uZJ0k5KZG+sBA++RVj9+hIPm71MdRIjCnKprj/TQwnsepv+0cLGZkfNHGupTk8WTJdV9bg
dW9UIGT+TVQVLMRwBn8FvIVxB3s9BiTREh5a+xmilgOsxLFAOWVx1SePwS/WE6UUYdEvrI3ND0Qf
QyBsW4ZD18w8eOVgqThMp2GWWcI8m2bS6iXX0TgmsJNqbU7xFc5PopPSqkWubhYuXpjd6YJMwJSe
wLsBiGRCbTcmb08Vqy31/J+Xen0WO+EBTW8b/6E3aTrqoAZzhQZuoZzaizCYmmxGXqrw42uhtfQn
pRmuKVEG/pkuf6xSwq8sYL/pwsVXVIQxJ1jqhv272CcnIG8UfIwuY6/7oLezGi+2KHkwhxp8H7O0
KXwzwkyfY5L0YTl50NNO5JIvAArZ7WBm6OWUhmVcunSWSurBqSnsDczpkt/h48cUeHTh7VZj9JSw
rVYdX9InoqDxEK9jCpJrR9A3uphJEFcmlNj4COUDv4J1+iydEcteSxb6TCt/tjgMvlMi+knssO2l
PN+G5QcbxTZR06tQc8VX7M33gT+NlhaHkdmgNAv1h67gkm/kQIqWxW5X2xHZUI3ztCMpEgt4Wwwa
QD2prUvz29ythvJiSAQOt1dunTjNHDgzDtanI006qrslw8R3TY6/cJFmiSbaQBkGB++CLWp266CS
s13iFv84mMBJn5qM1fe+O/KNmoEa8IwNwEubEj3tF8evitilHEXAMelTuXS8VmTVmgDabl4mQKWD
EJjBzXumwoq1OHaRxW6iBvkITqCJhCKikgyMFamXOfslAHYA75YauID24E8o7k6UG+1tDzuElD/g
mQi3fi87lZbbtlq4Vbztc1C7R5UkOhS0F9xSLiiGMVN4Bki9b5IqPA/pBMUCoDx1NwchlyOWGRDt
An+qMGMsAJ6IZUJsaLjGUxa6WV2pjRr0YuEOn+wlFztxxn4lHAlyFneu5LKxFexjyTK31XC3YzBK
jX5W4jfto9g6XXImmDqsxNhJiIfaz/S522w99VwVoa3aCbrnCtn9+xzL2gOnZWLFPOFJwxFeQOVF
dFpeTDQaR9MirLSWeXud3Shwf2AlKJ7wBvkX53Eh75eEW0MqZflZ/7KXcWuKMd5EGkgzphS4ra1t
6OE7LNEEse2NFuDpr+J2xAEFvdfb72Y/YGh2MXt1vDpWEk1g0w6onWP8LKZyoDYdTRxiTq50M3WU
iO726pY8wGOlk39PuGvOTWS55nGopDLg1FJ+NiLGMi1CzlvUnKCCP6NwMTkJ8AVSoZGzPbkcDILQ
B3bfJ/nzkjG7UHly7KlSap3qhNJclEJZsiQiMjCCa/M/8TyuJ68hOaV2vEVHfFJpKxBIYfhwlOTo
OPFKOZUQ3REZCMPKeQ/jXV9EG5mS3z06XsHg7ddM2uwPa/1sYfHpy6PrpaLrAXv9M5CjoZeAHnog
qAwHM2t8h3jMnwJotyGUATb3AvcOhTtyRgyLw29Gqov8knXCrdSogFPuuN6/CdcVOg5E6L/SHXgX
8bmu/cIFC5+fr0CS7N6SryEIPcY548z7EQUe4RlQhXLXnu/zUq6lHiVx08LaR1hIZDjoWnyr5HG3
BeJ+w1lyyGJaT5rjzTCnwN27milkea0V5uX5dsK4vIbrGsg451+PElsLwfHKfB17Y4XVVYSDs+Z6
zDBYw69cKdZoXwjBPps1QoQ/baWKcZYdow9Nk04IjP7uw7KPyEcmHHAwsdSOElym3qNF4TSxVfol
Z+Vxr5Xed7bh21uA9m1exMP+wdiU7b4REUGyM4ueLKtHgYN7EjGsrsTUnGOczZ8ceSy4h0tkxHdf
hvyQqFxd2COdWo/bvqlXKphPrXHIkWAwmL+uJboLMrOcsq5xU8MF3mM/bK3i/Jz4H5cVItOk30c1
4cqnAKGNrCe0DBLksu0kHRIfcgXNf0drV4Q6AAvECEU1T3H8XEi4gL+WJAwADQANE2FeyrehqOpP
eZ2VlWJ5R/AH8YeXgTt49ouhLjHuSmeb7inZTcxborIznc2sqYEKVdy0z98GA2VBBNHFToijlMMl
rAmOjrLDa1wSabZ3DDFV1SNzB2ITmRuPfCHebeiEJwozuKBAF6twYUwCUbk8rMNrin7xhBv0qWjg
23KN5pyfDziLti84th+JULQmklYkgZwi39/WvmYU3dBhBqksChmrLUrky48MkpTwUyqoFyuniicW
E7FnaQe5NvxpkeSA+FnuFy5znTNbrjPX/5+sO5jkMuVTvufhDiIh/u9Pi7iSHKk54vxRs3dUCdhy
luQ5x+B/2nxZ4kqWVi8D7WzxlUEZMxfdre7QWlHj6LQKtJTop622Y39WSK9Zp1D02XwR8gl+24Gh
A1Oyn/Ny1g8Cw48a4ilXQu1cMC7sNO+oQsiB3jCTX8h5Zk/mNzKUr/Lir60+3hu4s7zUtYtRlLbb
BcwM50GaRYrXgZxKPtdudm9uhehmSnK+yTVzLOD9gIY0STru7flJYPaW6ZNLkw7BwVB/VLNKd0UL
p6cAQTFaWvx3cG0naS/XfNV7eatwTp1zGkBOaoLHhDCWqIuJRqWpQhKrpGJRHV/SnShsd6eHspP7
aRe3bG5v2Dv4UxcIFCLFA/UbjJjylClI5esG6bp4ampjQqujfQiwd0ug8L5jWn/QnzxVl3LsgRe7
UkdlnIIJfULD3Bidf70xyLFGkTxVAYOnUDusII4KkLBb9/LX84nJ1hL9qNl1qbQRz6glcXEKn/ia
PRiiYc2ac+uPfefN3Z32b3F+5r+MCp2kpvGed4wpljdf7xkcLPqyttglSd3Yxfp0qR1la41tspa/
liarCIkBZse4irBZ3/zDSWmlUA9YyLT84FdOViYQdcNZW5jli6fjC/rcPtDYGEsbeHa7XU9hTlYW
P6uRQdOzn0qwSXptWm94sEZuH5bfbHtXA971gYLtvhccx3XdQZUwA+C57mmIkv8RQEfz3SWTJ+Ua
FuQnxqgNwtbAgStyUF663ZxK5Mumi0G2yXjnepvvyqFntqfQIh/bAWGW6GPFmqEZUQuTHYNhObTd
BNoSgbxTe0zp9EUGvdSLd6mlKoczuxW6jgrkzZGR1pR/MIVCxeDg1mzi1TGbawEm8V3jc+Gp9uCb
S/HrnNEKojaTgHMSTKhBrlJ+Yp9expLVwfhPVD+spn+zLtzs99RlQKXPywDFFpZzSkJCUtFH5dRz
AiNqKk696UNo5iHKOqmEbaJAu5b7GkFxK+6ghaYySVfbAxx/vtpjP88zjLodDtQ1XgMkCKBOMrRH
WuNrqJElOHYsPJwxgCv4pDDlD1eqwyef3si0bxX3sTnf0LipiPpQGB2Htrx5V96Z0bZA4L0D0mvK
fAA53J7WlGPFfJ4SLwDUjqIJr96CzjI2uagYz9chQtaBjpyXevnL79QJ2Op85L8g8SzwkvO+Triz
GkqbrXzhEfnJnHWkcHTGLd7oCUQniQx+ceWlRYLeIG1eB3T9p7UZO9+wiy+ShDWGIxpUANZm5vR5
hr8PHSQcQLBp1jPBrr2KZQFzqw3OaSR5dA+GsofM+x1/arUAQvWGkJCnp7DgtwMEoKDZ+1aWveCo
B0QQUhisXQ3WwuElmiyP2I3DRngJDtFCZwGvHbYZXSbs/ayGAYSis7qCI+ni/Bhz+TbN9VpC0t9Z
HWQJjzll0blAipWYgfmR9iXCDvOy7/oBfOJ0kBD+q2oBgIaDFlZOVKMRgWn2J1xk6VoX7TuO3CvY
mk+UF/Ph8LcqBTJSH64izi+ziDNG8J0E8dfCEPXi6OhxKUgtuQFvoGWPmIE9NcpzsP8NqJt+D4PB
qMH0UDl5xIe+blxlAWh+EesE2Lu8DIbbupMIYyScsQ0iEn+LkahWHed5cWMcL8S9hzw3+0o0Y9IZ
rBGmJYU4Zmx9r/+QTb/vzPLJOwI/eqHp/T0/puHZuadfmlrA2KF0+JX7otrj3hVrHDvPJFv/Z6Vx
XWeIJIsci7sZKH43lmojIB8A+zdFchckm7DdQAx7YWYuPL0ZY/S3UJJ1xUf4bv6qJ5hJ+3zYJdKw
4Gvk3lxRTRU2RGFBfer4rGqoTglH+mxJRpvIeLCabzLZ56vCkqFVFKu0B2WWc9+o7vBS4PiykYA/
l2Hu9TfieVAQKsv+gi7JHruI4/foecjxEWiR78qwsdzBQ+IwZz6AS0zyZbfU9U9k6/aKNdo6tuhV
zk/ZCv/phzszdToJU6RwT8L8G1Wp5UjYyYNg+8zjde9IPVAmtGuYX3IEXHZeLnezfp9xlRT9RYxn
kiciEO/pdp2aV8VpgCfcZ2xz++f+SKPQC5xPnwS2G0yl2VxSBDtRFHFSgZ1HKjiMi9r6/HHQgTnO
dlp1/eInrfjOdNOcUOLEJqsqJugX8MZKe25umJBO4G4IqVQQ0tgHWgzENBRinqfVfOYAHpvMOcmi
oAd5N9vkjtdQZgL5PT13+vzHIidK0x2j/x7WdY6lxU62jE1XywTbFFfXVRbKvZlTlIIWWpJzuiC+
aLJ42cJGM6bqwDHmXDwAsOB4msL2gaLjBypV5sFViR+6zSAnQ4YSdST/uIPpwsYNuIIJoNLhSmWK
io9DxL4jkPboYcdJggBGmyelSEoFQEAyvL7iDzl4GtcL+KyJBR9ixl6NtfqWhi/XZWJJzyUvYetG
1+OALdUJO7RI33K957Qfu/hUzfJTlqiSNPLLcZF5TPH0t6tU0h/o6ktnJBqY545mFb9OvQXdnHNE
VKyKaz4zjFpD/g37Xb6CyVm/BCCnRIHcaTl860BbFg1n8wbGyRD3qpC0Xh/IkxxqneYmmsZpaikU
t+SgddZHDxOu9/hNFgQDjiGcH6btIXHFwz+8dgY6Cz39zgo3XCarHYHpejqMXJ/vCibzsNGspSZY
0onv8+Fjbqa1NyYcwHUMhAYVB2oufkyToxwgr+WgmR0xe1IBD4LlK+y6XaB/qF+XJDSx+nU/odwN
qzqjkErD3eniSvwvrV36NWINVvtwE8DgJYP7lIw5Rh6nRNnwwe4bS7PMTzE1YqquCaLZP99bOwL6
8b90bfhX3l4YZM8qzF6FU7CrsgRm0VDy7VGQ6TWunQh1gx8DQ/71+KPLkA85SxTtzLzhFNOJoVSU
LCKqY9OhsSzxGu82kv7jRgIRkXRlWzM9YW7s/ofBd0Vc6CCd291IYGvjZK9Z9pCL3ycVxRDEXV4u
YemaITrG4Rk+K412aqWoGiz3Bz2bbt5kuHta2/zbF0PQWmo/kaOCWkUgCrCJEVNwTRwQW6umuunT
BJo7K08jaUi4neTlG8Aq5eOlvqlSAVfjgj6uPu4u6tkrT8d6nXM6Lfpf1fItN+kJ5AMtD6InpWCG
d9GU2qOuWiN8fowHJHED4MA/F/8sjaIGD2GaMrilVBx/efNT3a31I2TcMe8HFs5Ch0oRGkd1TuCk
RWOv4ofOq05UumqzP4RBR8rt0lxtrTkIXUZTJia0dxlXeHWvJO3VlhwkF0DYgbvZRRzMgv/dr4SS
8Hear+rVdTC1jcxmaH7ryvCJAN6oQyRyNvjTyFECQ0muzIiBO14TERhykdT6HzG7yQUDqEWWwATu
q4xh4bgWxLOqn6qJz5BK2BR1HpvebVdO3dGnEfXPfBtKyIBFmEfmYIC3ai9AdLHjOjdUrEonU1/q
ckU1bhwBt1A08RzS/chNq7I1vof0vdGmY03Z8ZajB0M0COX2YOiEyo+3IakSCwLgr9ASkvIHWRj1
pj1R8VtJk4kayNigzDSnCHYmNAngWGKlnu8IzMWAE1LvAGIMvZ92sm/gzGlxYBwxm2UAzAu/ItsZ
tYtqt3N2u8Fih9d9v0hETglaVh91JqJf0McUaZzr23BP963GoS+gJ9fBpEU9VdNmA//EeRByVrWC
+WgtKcEv8c2dQDJL4CuyYaO3+Zo5vVOepFwSxKn/Dg//ByQy1SnHI9UJDUNjmVdi/cn47bng3+UC
o5+slF11Nhz00pagid8ZJbmLtKSnhcxic35XAXWCgBd6+LhsuV28D42Cm8KeWzmLj/n62sMXHd2K
fpA5belYOCN2wEmG/Jdg2ADAUMYIgH9ehXv5aPOQzS1TyT9QfBmp0m2S/POrHT8giYP7D+AiJeMl
cYOwc01VoAigGH+/6XmoSooxW2+YWelQMHyTHi79HakikBdBwFuSQmyCTb4B1tz59RVgTG8uWi84
ciP1YG+PJIOnPhW3zM8Cb3UkSAJbte6NqiZUZAKzKPWeoS2rygoOOs7WchIfUxJX3Aq7W0qmWJfv
mOV6R46Fr/lZ1QrT8Xyyi+cH0nHgiSNQzdn3UTPNWV4uazScrsRtxo6DwZ/amHiD4vVFlKmizjlg
b3s/nZ1mJ7j+zvxsW1xFUk2F+1W1jnpwMkE5qfNfmzv+ItLEeIOcrmslfzf9RBBwzgHZI/CiM3F8
gmbbJ/px65XnoY9twn/pNEhPFzYxQ4sElYO3pQp0C+wfFElccDc8jUCg9J1MUEkrF/iVduz2xYsQ
ixgABnjj2xWHMfDZe727qml2PXgN078RFcpJwmVkhoI1XPPp6t5bKF3kCDXitw2yc0lzr02ApBaQ
5hBdvPBLeZnUoYvNbAjAK0JslglzQuWkhf34p4x7Csl4ynUent3YdjlaZxoQKv1cfbNXXLSa/5wO
qhXJH588IB0sKYh92qMwI/RMULHdqBGhbYCOYfmcCo3z5wC81X+Tz6Fadnfvg8IdKZeLretjntGQ
2Xs53DZFBhdL8bwrAxpvCw1nDSQ/R5lo9U5+ZAgMlevu9SjSYIAtR/a8Vb6DNaUl3PBAqj6ImKw/
nlBTU6HMCnry6umAuuho9aKfw2xRO9sV139DfB0JO9pIhOGFjexc85/JVKbWIEUIy36WWkmgxBKD
HR+NKMSIARTKboc+wtS0D4+q7ibfxiNsIofzY+sElhcMd5hzccgIXmOKq30wu3YPNxCbYODR3iOK
qocSCNwz997odOP/0rCRzrt3sfGlonFw6SDK2ZPgsCh7yTXGrKQ1Dh0al/2D8iwf49jt2TFjgceY
kiNkMlNizHReMIw1ZlWRXvXMhhG3ERp7h0gTrM78FjimV156guo2x1knlkeLnHl1mZhsk06G0dsQ
kNvXLu7bQTkLReh1pqqSmyyVsBQdeHDRahNwFv0G0JGjEeFcExra78LsJMYF8rTHsN3rok24uMAv
2XjYUXMvkUyp3nzaod6VhI1G2UEOuPnWinGkr7z0Bzmmij+3O4ekjr8bG1tJeDpfUIuge2rTpKkq
JwmYvr/pCJVWNmiqN9xLVudvazVFK1MPP3/yMex6z3klIqRCpOFf8YlS2wXjyn6rVxlm5ualP3BW
1ACD5G30v0Ln8OSoJ6EtVisvCn/pCaZ2fSYp/gw8akgrl48g0Md9qIkF0VIoeE74Yc9ziY0pYBXt
uriY7N9WmrB9Kle0x8ub6Er7peRd+BJNv6T2MeaOeBqjyKqu7M0b3qQzv+MaJtbOG2ae9DHdRVBK
+K4kO2aMMARDCuyd+p84GHc4KSqKGVSNEqoeUqhLLO/01OCIBtCKax4qItavz1XecHs+5BsxyWIk
7JOdvp0uHPB1mIaMnirQd1hDjsG+cBXRjJZJVtTD8vghJZDfu5owm2MTmI9o2DAPMkB42erzieBy
55vQS9gtw7QAkWIakJCeAwuUzlZFy/XjzY0MH4aYU3D1Dw+ggrx4bwvixpme6oYb47FDJkG5gRHp
n1SayCEKZElJc9/tT0mwh2gA4+c/DB76oNsXkZ2wq5slET4oMJ/Z1iis833AKRN17LNjPUZhnoTa
8peJzfQzDRfdrUyedCj9hWuuA4uZTpMF47cxa/SXHib+LTe9mHIzxrYm6YOrm5W4REt56nfxxZR7
KywZrcRx8tUKl9B8jB9jSGsxm3qct8STSjp+1G7i0bLfD3Jax4s/rsc008fSt+8dG2bLZk3Tsp5V
0Q158W6NBNBtajTq06ds1mqLO8fj75Tp29WeJJGrTPJPf5AvmQ4tIvkpjQ/QNg1Hi7Hl6YJxcFcx
n0mJvjpOu43d1mc5YPaVsITfvZgSUTFPQREieHnzV2XcsHJbzxInwhRE5Y1IHUnfVWF04Gcy0s90
msXt4Y923Am+icxzyiGvIuKT4QAWPDrWasUAvMQWTS9pZ8F32n9nF7qJWVg6/iQ7JIhBm2y55KT0
f1zXIjSNLbD6kwx+6X+g3eVJs2Th8TClbhZn/eYKeAhX2Y8twgQ/Au4Z/3xibMbZi1ioWG6K68E/
5WMpyh1V1i1oOvNVcgb98/wMT0hIX4yx7QtsF6ZI55zh396M47f/kFJoAzg8/D7YG1yu5dE3OGvn
7LNiIVZx5jt3yQJcTIZCSsV/+mGN6S7PH2ezY62sds8E+9LXphlOxgOCOIxJ7KADV58J2HQ+wIBs
/S7n1LBpxRhYLsj3THruL+UxEdtFSHZVdFzTEYx/cq/nsJQLcpnKFsht2R7WEuU94wZ17v+5Zlrz
NNUXa3k4OsLNKWV0CAVgY5pM98VDmNEXNtVv+O4I0ikWt6uRD9fEle/+lXAJxJxwFXal9cGjr6vc
lLJ8m45kzdspaWB8vkNxjzJnoJTerEx1mmB4L43e8RvKKQotsqJPy2O1kiW0sEktLnvkM5qpXzX9
idccvo9erGqroLfZfTc5CCk8oSNV8wW3JInoOAujo7NYsGCOtSzooZw8rMPuEm9SbXzajWwHjGhJ
R0CGNCseVvzQe2xIoZUZX9AZATDy9fo2he0U52uIr6dZdq+O7j4scFsL2wuHIuDJxzU2vvBuiW/2
MXdEVRPq2ZkcNOYOQza8+CJTZdY/aCUS+RWeTbEkyVlXR9CP2lYkRNGhBjTdrhgSOHG5F7m6y9r3
/1MR/EZdiaY0soISRnzFrfWqoU0UpY31liM/F9ti0uET+/FiD2fhVfW7SVvtymO+1qK4LaqoV4/2
c5JFGddjI0yzdvKd9Yjq5lhvmr6dMW8nsJFyuMN4PUSKALJIVEcIlhJKRkDVd8rsd3IfwfXmcjAy
cIzsbciJzPZNmqe4fCEoXFvacG0GLJtKHPygp/dPFXI4pYWrKPtE+rwnqZ3lop0pE+5TklQVuZKD
YI2hXmKzDkfxPQJ/ssSjjFtV64W4rJOol8Y4rD4THtkBDzjJQS6tdTYHpyf76yM/vByDWeW69NcC
7VA6VeaSSUVgkQOH3ySaOAu9QumJJdrxYWvpnf+MGFr9mHJP5AGhBOMBo961PXMDCqLN++Y1azK7
Ld31cqnmmpYQY7uzXoxPFAltVdnCcKkPGhxnsu9ZRqEh0i/8/5LUEXGIaP+D1we8Hvi0VMmhyYaJ
z0aIlE/3ultyrp+19ffdUhRfilY7SDYR0l7iF4n6KNMSOz2BzjbvD5mD9uf3IaV/tyQyjh7gguii
7Apzmmx88F3Kbpzj178JSjZ+l9Io/J9Js3F/M6YvTZtGA7sVFwOAnofmZ6aEuN/Ne+XhMA/bufhm
TTAYXNZMS0myzIJ8wk6ajRG4Wden4MCp9p3wIRgKcZc+AU3UyQ8tHSR9Vitim+3ToEvRI0HkoJ/i
KQi4Z1OLK9MkNZWrkhwakzGsjDuwdhZvBuaedOh5fFidRuAT2rXVfZIR3RtDmlEmc4cPZGkhjrIr
V2fxdxpT2lY0LKgcXa8yoM7CXPPg3SPJpaOxJcntiyY08IUcL5MurcTdkwpvOjdD9FUyskDgQVo5
UrEOEiBt6ljYnobRPUaF27rlHD6IASYN6Q5imqEUIE756i2PMBCgKowwjA2+Pj+E6a5hvp5w04t/
c1w5uo1GDHemMzKuowwiARub1T9kBS3HCjWOj1WoTc5f2LM99DnLMg791P1/MtSRJ+OWtPLJf3Wr
cD584iykQMLd98ywORaHJ6U/qbWWukcrzVuUAXmIpVdXxbhbDZVEtC4Dw0uh43TpASFg7kqWc193
1SLfjxh4RwlFSBSvx9y4kvrnIf9AhAaOyXjIlKH1uGH5pdwYfeMXvj0f1Ay19307FfxzjtNkptqz
SBEUHd6QUZTCozx9qIfqm0vZzcgrp9rbt2YTwp+5D/lKEwN7iqH8mBeXKqoy+axdPwkq1IPPD4Ua
wev+Il9yKA/etvLLoyKViSMSsR5NW8kEwIXWa852voYwc1K/ZrGhvzWEb7B2esGCyUz//owY0/zI
+0o+R0vzHig/nh4dis+x7m9rPvo6GUVH8Jc5u1BhVccwkkwlDtpjBXLJYO9iAVdUWpca4JVRARMC
6i31G/f4gxXedT2qzOF4+rRJwMYSIvcr580KeGGfrPV8LJE4y7PfwcowKiwc/dHqm2JiGH5lbtcV
9HZo2zKKOrLlmPpo3ZqBzqoQXeyv38LHnlF8cM3GwiB0npbGJSbFI60LMobEr/BQmgxatLLxe3zQ
8xESjw0ml6cwGILorXSeyNURwWrEmxSEd1rVjt33iCiyTawS1rJBXgJh42LIWt57HrdUXRU7+4Xe
gWmwTJQRM8fwN+ctARghi5Q/SOq/hLSxEEwvREImI21Czz0evB1UMmFio5wxMsv1Y4+FM4z3eUgp
QlPtOgcz+/goUHeBRQmKdesV4o71RTH6+J2JiZPP/g+OG0fITRRD9g05NWd9zBBVfRJIKqgxLkS7
atyA9BvkYffjwScBpNKjJrj97FOaf2gaojy8sxDOl2hkg+F55Z+dGZ9/MCYpI5S/wXPWV+XqXK1v
eqLRytJC5foDfuFji+g/i4USouHuvr4Dwt8lzCKHrd1q9qIiBWlwNLssm0Ze+I2W8J+vsy11uDE4
iLc1DF2qkOmwriJgrV5vAMoDNpehb4mf+ZlvYG+mlI1zFMgiUjx1H0GyCGEwLhgUUv9EeISl6boV
1sfloeCNSMHpM7obmONta9sl1U3MTkxy2S/MMRmgNuRBD/XPOHGii30ekThSyQ/n9UWpO0OG7wcw
5rBlgbBP8eglcBOpI/Nji/RnVPNscg7LLCInvx0s7PQAowOQTq+EHvQZm6GYlfFfPJq88lj0tP59
z33cWZFyf0NUDUa0tXWNexCkpftJz8Htsp4wdA608LmJY6Zf1kW0G8t4cj6o/UKp9P7MasBpf9DC
gzlFC58z2FPoNOpMXp0G1FQLyx+couNZCLYSmYS/daMtNKa8Zmw0TNrPiFI+zuezy0PxO/NhrC9X
kidEoVKDztWhJDf6EUdqzJ6WWX3l66N6YcJ5QewcXBGwMPRA0VYEcNib35V5wnSsNHNPJ16UDZMa
7EDLlO/pZJD/g6VqL8ICqB8BDGRa0LelPuk0cnmdAta2jFRAfjxZrRNvj5sNpfbY1gEOTz4+PRf3
Rm72YCVgha6ZdYUewNIZVjC35Ll3X4z7ixiUyti37hEeG0K9RZMGxKNnxFR9dqRGNIAgD7Lycbis
zxfI6OAYyjnxnl3kq7izoBB0eZ79AiuV46UH0BH6rvHNRdi3mk3H20xxQzL1L3KsDHalqRDjFsqM
Wd0aEGnFDhoy2fflz69lTb2q18VcekHo21HdNn2QNSZXMpHCaa7pUFoZs2/RaYGkImu9bMBju7Nx
bkWLJN04eqQ4N1iZw8mtdhgkRJVsVqw6aIhocrUUZFjQK3ZrccYYnDcMeB52GV8guNOwpsU7GXxu
HyHBe0LwhIES/DpDIHcbUp+3Qh4uR/IcCO4vtOZiK04t5YeL6FUEUjAMn9jAFXcm3GEuX9IKx6xC
Pl44/QZSq4k+pDioWHFH1G9yNoUofC/KZ+u5QMEcXnDxSppXiTe5f6YfLv0usn2K7GQ2Vrze3R06
CbifDeakXDLgp1M7JbsSSvefTJFl7sq/T7yfar/c2qDhIEQ88P9bydHbgp9zxZ18BClyVSGwnT/B
QHXCTyjohMh306QRZT+h3E3x0+u2N5KFEE2QeeeqKOXvlqGZ+ZOGVNMAvy4onZQtk/zHI5YOjHfo
KrNm0i2Ypy7L6czmHROSUlqlX4pn2IxuZmQHWWQSI2cjSMx9PHxvt+K+U0qy5Z/uUGD+GSQBdU3o
Idd0XFElqI+2j7dLZl80nim27a4EDtO+YiVoim4h3DQY2sXm5zAj10jr0pkrQtXnDlgULRFtWnap
dvhH2xNXduKxcAVWgbObovDCs7y/LrRwzJ/CWyZctvQky2D6/pljRB3oy9iiSZzfTwheksb3XFBp
6P6z5n1CEOuoz2Ece6aJJSzetkGBF1XHcM8KS78hou5K3bsWppRNTcJM3TsZsC44mURxkSWAJNCx
asnmMnjP2wwO+5/zIIwOzfMNDCDuZHst8hEUiV4F2q7rCdyo/bUokoY1nCTTMbjx/qdhl2U4z1w1
PUHUEXwe8DpukEH+dMCpIOPY5qTw2oo4vAE9nNwzf9zPegTYzzz0F8hIFchUjkTI+KbBp+HrxcA7
jJygxLLf38MnjwA+71Zd4x9OKhYGlKQ+x4S8LMfgs8m2g1o/EZ79qscnCuCFmtZ/46g9kMDYc9wz
ObnKRnlfgnSSGr+wqsBDAGvXBGpAy5vwC2PyXaP6Z5kxTBTi2gfR+RvbA3QWQ734Y+wyztmbaivQ
AbVOpxXP0cfVo3aU9Amsv0QKX5OzXXWlqDei9fpEo89wIBSjMrn4UFdQLdhmVHrUv86nDLwdO/hF
teCxwYJtdhIO45/LyZnkaQG/Gu9IrXI1dWWLON8/pTREAAKPmN82n26jW4dIrQrRPr/YqsA+FRZf
ipKCtWGgKn7vtH4AU7B48IkpjeruNmxM9RA9vpIBfcxHnZE6LampY8HubhnYC0KqdvTPbHFqS9Yp
bX4pJHO1UnCoBI4ZcSeBpKs0qGf79j2kH7VzSXhKH1VTcmE6fKm2OxWbVGmySnOIP1uyY7fC4Mhi
srT8m+cWcrNHQn/QCbpb75YI6pBGuwQA0Iaf+8c1g0zq/wEfZI8eEpGdlZLstXqcOp3RGZgqkCIV
YzAvsS7A0KWSaxmeQxBnym+GIvlQIBzvEENvmtV59rSpsFQ4smPPwCzs/zbh3LYy0HNngDDvQUt0
nlvbhuMYYqbWBK0cZpBi7fWELT3Dr6xLknf3bwmMOqcGW6/H9Vlk4BuD4zT4Ju88aj1aJmoKwzp2
VR7k/3hFATbaJ3Scuz+Pc8g17qMreAQNnzuKCVuMLFekIcJDO0GiXoYeStLpo4Rt4FfsZ0JbNMLp
tFSf8RV6gA8Ig9lWmPJUdBw3nBZ7z6xlkDllAy9EFhjV8xmAoBsAeBPrpu6IX9fVXhwxdNDOjduG
zY2gzubRpKi5gYvl7B7F5g+bx5Yw3BzyQkfR/gRdm3HVvn9CekjxfdpGrA7MbyiDB82d9QHa4/KT
t0eKyjvA9GroPJ2zqdrS/UbiCyRQwNsLa4rnzsIPHBBvNlo6zzvrgt6KHBEqzJKegnv31pWOQ5UM
MYYqQECczV8ysA6fioH/TOLRk23uYOnR2yaC8GWlXtIXP/Z/d08GhH0nUNmAdXY/bLnowJUVDrKm
eABLgtu+8fGJr3RgcMWn8IcewjU27DG2VA2NOfM8s4f407+V3CewGX9nOKzJwOfWYHirFtQEy4cf
0i+d0aanNIHZh4RNRYIH2EfhqTzKvjjnJ4X5JozPXQ09a0/AGOl4zYI+3zVCaDKDfpfRUAtY97Xw
uRzoVAK0ZXlYHPeVzQBO6qWcSMdtrnqjprDnKWVWkviiV+Z9r7J+PlSDyzMre2AeOlr4K5iS8Azd
tMwHMVSx/d9z8C00vtWNDL4FTUttqqWphEl+UV2mw1pVvdO6JxM4cf/a9ARDBcVG6HmnC/wIAwPx
32kOhGzmRZZNK09ZXLlh2EWvcgXt23KOWGupAzH8tFpqOZVkhmTA6ztafSaA1/Dy4dc43TGiDSlC
gMrrVy9uIiUuF1d//SXvzGlNg4ZYygwDhyw3lmUDx5uVNctyBbvCipk+vhq5cap13+DlZYN3gllj
I8hVL5JbHiAJptWywrO910G64A5Aoq22yrk/3xmHLox4LJ5RjefU0H7yWb/hdQtYqwmASdAt02MX
7xp4nvWnhv5+JrpbTNns1dCOWEODO3+xyvD9DPBeP7mMoBbMF2wxDL692lXcIeXLM+JxtDqHknH7
d8XMTEBAVtMLC6/ToRN1BwSeig9fIvRa2GxvLSxF0k/it9EdumCbGfHHetTOraDNmROVDXWIOQ5I
cnftrgP/kqZ/Yl3LfVvcCRe6+YA0LlPw/7ZfqUPAQMbmm2dzuMYTIWgAyI8xcX9uAPeYvhHP80AM
BBaryVlibza40smRaesiZmVpOFLeXeNCmD5+tfq29aPHDxV5pWHkMg0846F5vpeBMjHhD/HVHedp
set/rsJegguSp5FuVxL7DW43+PAp87+4J7JtSBMrrY7Hbrvv4j1GfjOqjzA9x0kU+4OaCDSflAVC
jPuIgA5ne+BH7b5tX10rc7wYgwEOYnG3N0ggOZboPja5/F+k2/luPSJGkK7MM9TydocsR6qLwMbh
LTUfD9O/eoVTlxqyAwDZ8NeHGpWE3F3nYbiYgz6HPujeqKOEGKVrfv/2pH5s59o2no5AB33u5agz
IKtEJbUhND8nCsslXU6Y48elpsDuFz9UObbJ+TPPmjs2NrAtSR7LXAOkpA1cYrfO+HW2DHVQSZmf
V4QhWZ1EYA66uI8wLOp8knh9RMNOJ1rGE15r+Q/UadGz5e0SADu9fS+7M/QKJXb+3GMuI819zolg
3qElsJAqAwrJEDRSj2AfeW2T6dXQktMYLvfVsKygqURSArAQWHTuwSZO9zftOpm0ZyRsob9UNVOk
yTYtMS/njoJGDSNuCbS5EjtfWwgJLoFrXf3JyiCDpA1mfjII4YBvGO83DoaIT9wqDfOwfon30mNH
sKS17fW28pxb8AIrx24x/jxsEHqvSVIavOgz4fGepseSNMUZ6zI1ERkm4alvj1pu1Fgf57XDcONf
vAow0TYklRg2H8pPHrNKDhow6WKN77LwjtRtSt2OSRwMd6cXX09bbt8Vxri+m7Ee3PPsTGnY0Zs7
9embC9dbuLu/QAJMJuL3AY9RtMZiMDzlqm2NZuM5wK1IK37jhwAsHvGRamnhc5rZfaTe9rN2J638
fYiYmfk3DYSslUhK2/EPkcosMXRRUUVvmoEq8qicodLUtUzYsSVHg/e3cHk//MkmyA9DMdxuIW7Z
TUHgvSY1W+oyk9JCmP2Cf1sURGQlyu8PGfH493ligx9fi9OQTmp/hP0ib2KoAxSGjWonkOqg0kLL
0ZR0rAzmU8UsCoaSf8Sqj7wTumXLpdS9NYK75BDdN10+7y3mBthA3YmcLBPwbVxxmRCYSIhDiB4R
qtmPbTputCnFZZOzIXfDOnwlLmqhUNukSwDNW3DyUq9CfBydsWFqxi1TuzLEhbDsTlS1HMz3BXZo
8IuUx6lvdrDsDiBxw76CVLxMbxs3aoA6d+BCIIbwAVIIEA2yaQkKbVeaghmj0xQ9AAWdxotK9G6/
OXwnu4pv6qx6roxPtYCbbT+EKT4WjTjvUxMGck5A1GnwPFst79St3+yZS0oovP3PNYhSZ4tS37NN
yY0Mu2Um34O3oubqPWVAT4foaxUt9YBIOFy8IsW3DYBFSdj4DY5AmOJCLzCkta4iqGKD6n6hUWdg
ZZfEMmPuvrs9KFQv2twjucBnk+0GXniZ6f2LG3qBUBHkZHGTxkYObiEeXK71pz0N60cO+y8Tyi4n
+Bz1Ijp33gt2aPMZzbd9FLwqyCE8AJD1+9L43xdZ32qUFRv0pOUmRk14TW52v1W/QMgbIekruEE6
HrMUKnVKrOPGRFLjiiEEr8kgIZ3EQRF1hoVXZTLMCpZ3Y5PVYiwyfagxVlRPM7YadGHfOQpUYX38
nuLiKeFix+dLuVBTed2y3mQzNCLeBXxwqQoVB35lPwHO0G3t+e0MmN9QIfdOVrjPjTliCkK/ZmsQ
8vNyAp3oIYvR2/ezdWMRewEDWcAjDGivlLV4DUfLXeZILHZO26wrne0LmuxcPtjuC4h25aOffsS1
xtbD4Kji2iZxj/3xmnvRFStOCWK79k4LpStINgeJOU/z+Be32/2pH+aICcZlNbvdSlTIDvMb9n0i
ZguuCRI7sQbdlgBbyzsYUBqX0d2RnpJP+E18uEuU7JtPrUAOIH/PCdQUR911BJ9qrQlDJNbviwOb
vszaS20VZjs3lzpFIJm0osDgOfGMaGqAijTotTFgvyMugY/nMQazfNtv0+5NnVo+Mz5so3pIHpHw
dTCdzO/+gOh8pixYqK2yDB2CcuzM9B1DLqmscphFv00+/TU03es7rI1LNDVg6ShHWAdH7yF6b1eR
i+wsDngLtNpsHchzIXGoY/9pOT9BB5yysvwMFl8hrRuiHDGw4wdzvLPXIEEOmZHBW3DypdSh8gx7
55Z/fwR4E+MWmi4OI1Nraja8MobtJSa0vwQdQN4KI6DI4wysZ5H4BqmiMpxHn1KBh0SnMpkx/GiV
GWEZQ3KH8UeQz5Ic3LsFos0dxsI85bbvfViEt5vdMHpWly/KeEcS+GeYkT/Kj9Q5hvwqU0Cp0UOq
PboB7mvCAszis7Q82pOwO54VaGuSiYQ+GJpYInCvWjtduzk+fWDEmdF6UbTYaKfNeBaN2lSnlxq6
/01G8APClXgptAih8fp3f+1yOW1E3fZov8WLGCQ7XlaQFYCM0Y6JJv8yiAfxWRyEMtry038pkHDu
lyCQTL6DGIWhrQkVXWa2O2b+Pw+F3ttG9rAs8d0hsvgxhl4nyKME6PqySWpVGzn+Ag0RWyLNRj4t
F2gCgAWq4dE23qEbi8DTzKkax5orosub+OyubKwkrs9AtzYOOQ4+NVVx1nz7Cwsh2XOnerSrDgTj
exB7p9HRNW7gOVuexM5KWyZLaFGnLf+q7xpzyp0Fa6Bue0gk8HvpkJHEgsc78pras0VEJOZr68WT
XbMbtvFbZtLQRo3+pAJN5cUp37l8d1e0A2oNZAt8gyz5taOmzGdmCi/08wmECj2IGRZx5fjtP3L+
BrElATe6Mu6MeoHLQ4eDSyrORIK9pAwkVjKN4MUS2aIgSCKpY+xipaIGJz65pzzlbOYHglOMl6v9
V1t1PIpZEWduP0m7lsgEhE+lxIPvMbhPruzvsAQ++m5CzCQM0zIbcwRXXe9/X/FyPSkj7nLBKiqw
f7s4hnG8c4/P31gXA7O+kwo2GHLBLMJ1PkE7NRHgwOpuXLCry85zjIP2ltiWWbc42fiTfmDxDhGl
6PyzgSpN+7bwXRIXYYcVHvOh05fmJnUvUhlgdbmuDISbhDaoBiUMgrM5mlcYay7UCT+XMcRoOXsL
1Vb1En7Hd3sw6epkmjOj9COU63vPdfyulMp3Hv0f+pC0ruv9OpWI4DhK1DNLrPH9qz9vvwf6Ro+9
2Y+84S4o8GBppZ9AoXaTTJCCZTjmm1anwyTijCRx921DqY6cn4Lr9fNJdepm+iHlWQWN4NlefgW8
CkHCFP7LNHG5An6E6yMsoF+t1Bj3TdqiuX6OwlzFFikiSJSvj3zzt9aX/hfODTmOOTQ+j8EULxXO
S1l6tdZht52uzbJUMXqLGOy95J7C1f0KcFqqkZdY3AM6/XlN6zWkDkzAAW5jC6V+Xx2aLHSjh+u5
k9iSWdaK8tkvDPErt/LJTELqGKS0S2pFPe4PjZfML2/lN9HgOpa8DLkCs/JpLPcwaAHK6dogh3+M
+mW3+brpJsIbjmLdkAcy/qYC9y3AJPk67d+dTfb6AYfw4l83UDqjEo8HPseqqiCjhUz/gp1OIdov
fG0zXhemrmFkMKZFh1CfCN6wyGl0BBVgJ/dSZy+3c/k7oY9uWZdtQCD+NVK1uXFwSfF8ir2MEK6M
k6kduUy8x7N9o/YygSYyu0WcT2yixU8pqd+zoldiQyd6JcYtmmYHISY0+AP/SAKiPPBZNwqpsw/d
8h1d+qVWyg7ghdrBkV/M5x8eZ+s+SaQgpnSYrc7axCbK7HFTWb3e/TPf3N6+aEP0POqntCUO8PsR
K5wgbTR6c2kO4t5RCkNKR1HWXw7xajwim9+Hg3G5pxcgeb/2KjHboRbmkEci6/rsDoOg41cY0n6O
PSG1NhJBn0bPcW0qoMW+mUk/Ib7t3cxm+hwopQHLwI4Q3Nuzwy8Xc+/lZh1Bv0CO8UCAtzVg8Y5N
u1uj9y5tVWJbeTefrZGy+Jrh01knRJrCku44nHOo6y333ip8FrdLCcBJkcqFLX+S9rjqtO6DxmGb
wrNcDAUohdTfIwGsTEzwM0wYizruybiV+oCAF4uLtriKXeeiudYNS7Tj4yD/zJad4X36lqtOfz5I
ZUM6+xTS55nR8CETYimkViJsvNheyinmwcs+04CIs4lbIE9I0OaOrV6uUPh0jkruxC7TwNliWbO7
XmH9AHqSc9q4YJ72aA+tLXMFRuVYP1qlxpIMCO7bSItw+8f+pqa5mlsyNuDGfngULUx9CwH32d79
A3Uay3FIOnOj/Q+l/G6dHSdYGRvKcsiEzS2l544HxgZuUpSVF1yK4F+vDCUh1swAJUdJtC+O1Cot
wZPJ1lLC9yi6jrQBzgZXQWm7cxfW98Nm5x4xYesBzmb9o1XejslPj7VQ1gWtmDJSVCzRQPGMu5t/
vOXFicQLAdh3tAbswYk3uk1/df/+nHw3DZ1rCKkKsHoxIsWytRg6donCDi9PFX9jQfXG12Kui+Q0
L4pxiNqOJJPB9YD4UgKo2irNEBHVRLIROv+/phLniLW1ei3esNUWrNrwO1xuKk6O9baa0Uzduv/u
eVkF6QNrFo48XAYiWUheuHLWCOD6MOHtfRLWxM7uHMlqpD1FkISTKp7eLLNkhYmKD4ZRARZnkFHu
pdyfk0uHt0vmMKZEVbu55BRvKvw2lOlLW+jUXPFCTf4mAl6HABYl3NM9otmhZ+Qbs7PMniaJI20I
M4iIu4b7e7CigwesCLLHVU+Hd6TI1Wxxrdmzo6+f3V8ZktoMzHkRXn6/1FjuM4H1H7MjQODc5QRl
PsGyc7QcPWPwADdW+O5uky0u2HdMYJmDerhhEXdl6JVlOr71yv9FF77M2lCzuCtey4LAURk3mFbF
RKqyKcyVtWCzzEQ4pVnrpBIJM/R/JEX7XceXsjLQTYxv6wt17NI2V/D7omaO4Afxksj8s3LKNn//
0QkYao6cIAkZfTcYBrj5Ur4oEyytU5ioZsQGkrLxBiTloimrQ2Lx2vE4atwHq3xFiocOE8hhqO0e
PH/Gr0eEG84i3bOra41K6iFiK6gx+VAP+qqpr7PkrDJMeA8Md9Vv1i7YhglhRc/tTVYSk4NzrPtg
kzQ7uzRLTKG2+0O837BmPMEu+8YItN2kI6ZDr1LgY2XF2ncLw1X7qR7mC805gJSqILwW9tKrDlpb
l45kCMOFLjkDJVad73XOZOiAqdHo/RvR3fZeht08zXeUxrW7dl+GkP3yp+6wX9h/J7HMTloJ7RmD
w403SETlqY5eRJrZ0QIT6i8AezqUVd4m61UOamj/0F7wrSqAIzzhalOhqHdetGLA7acjjAqr58cX
baZdO4S8diIr4Fx9f45paa81tYFT2rUfDuhCKQ+8cSMpLBxaHiGaKSxZzxG0dIxMz/6rtGbhGJt3
rhBBCvMXBAUrtH9kA0pqwQhpfq2keBHx05j3RBhl+0r1uPnOs19zUnfBIW6ylkrUEQr8RXlaAx0w
0hjus2kNXYyvDnqXNieIeWuGV388qiTZkz6Agnn/WGW91Gc3zb4mxtCR+SWAfHdlYNIxkue+7Y04
/sRYnzdLD8RWsHcXvldKD7irHbRU8B85WHE155AdP3IzFL1CzEL6MTOyM65tvtZc/ENveh6ub+Ni
awqvOWHcen5UIMXFIb34wQXbbrcI1W1tYmOtO7ETtGrp+m12szFjl/LJHEBL7B+NLlR0OlyoKeUS
IYfsza0YxMw+Rd3Rs20wmg0hG6F4IsGNkOwVw2wN4CF7vPAYhOgBOTJ8nvng9b3++zdZ9AZpVF06
+dYQhIbzyDkdpHNe6N+N8n3Vr8sf5C2Bae/VBRHl7+mFEWHv1Kml/Zlv2d5+mdLaPKEo6gibyuJG
UMN4N7hfXLQDtQpY12PsnyzzPLLyHGuH0YSMMd3eNp1sf8HU66bLUcpjHGg+6tXbl3BYmjTccvFj
T/iFQN6yxlKIAfx+aM9AG/zoat3/2to5i9F6Nog0PeU1KYzRlk/Wh8BueQGpesdFZ+k2bK2cCg89
Bb6Qcic+6vN5iIXLIYkinseys3AChr6XPcwxWzN4cm29nyPodxE9Wyh5D0ij4RxOkw/vUW77QLOs
XXu7atW5s2yIZr2WPD0bK0z9wHPEhpls8FOzhUY4IwFzy75s0kuMLmU2YLZUfH3wd+mWZDYx4kkE
6YpGCnJlNAqvnRB5yLYMzX4svHRlgzTzuMpaeBTxxmDgpKNlAbnHYrO8z9Q9dfelhoR+HgJz4YKY
NOtgVM+Sc7SZQ3Wf4WmRFPc/gA9hsGuhlfQOxPx1ZNvcnbs8eEMJJe7H9zz9TK4k6kimx9MswKcT
Hjh1TuSAytYNvZVJMLEL/UkfjlaaajVSzndh3N5HJLaGK1XP/EZy3q2zNqnl2BXu1no9vBSt3WLA
ojK2He7+dSsUCvlts86ciqfB3nxz6S49ybbm4UR2DcvjvZeU5YG4r63jzOg4AWmU12mvhHpFY87Q
obDIBr+2xbTdPa0aQ2WHUkZseS9xtW2z5nXwoedXhQkDzYn3yzf8K/KpFaWJH8QOmHinlIRGRGTw
ssWKecd2TRFiHywo30GSybDZGRwBvTmzoxLiVnUbLm8BVb2jxgQ7ZKPU9YBceb+8wT+JpZBidxZF
x/aOS32sRwZOGYataGxVzFGgmhtIRTIb53Fqdoiq2jyqfyd9frUZ8U19xcB1C5VjWOeIws+Otveb
dLLgt3RQpGUqtGstrBF69gjLFt/nAIq5Yx1iEYLcW+W00zUshcXX+G++Lye+v7DyZ0/INn5m6nzE
XkVoZufEsO4EA9RjLC/OdQZEgj+Uy5EbBjSJYSF2A+RRJ9y4eeYHzZXPNo2kjI76F9W9zRkgJGKX
l8BinFzmUm0SOwPuaCBdx7EjyxVaYkQ3JSSyWTBTM5CGAapgfY/S86Y6bmatlLTm7nnbcPIMo32d
ZxHX+zfMPh8x/N9yvqFJbeOvm/TvWXSfq94eK9nMyCh8LfiWPaDUyO6MdGtM79ygjFjeoQlUwyuu
PRKJR0Vg3ekUyKX5shHQw4wjuS3/Djq6XejQJm8FeMzuF5doNcAxdS2SniftoAZHrz7rmlKJZjBZ
C4S6HwkdNSpnVEO4cnzRwjRbk/DIMLguhCld/ztacidLUtp0YrazwS0U5ofxHseCHDdOJF8vr/1b
lwwRIztNLs9CNkbAnnaB0hUSc3/zTA7Z9RwP0QSvc1a9F3bDSw44XKWVOVhTyICslXqssWSuYj+l
OB9rW9WmKWXCF/YD9u8wcxwpitps7lb33G/J/vDi2gbgFt5a247ISX64BCl7UFD9EpNuHX60c+zM
DG1Yd4DdHzdt2IsMUd+G+UzZmiB/9t0S6ERy7nBHg5qMYB9+K2EHF1rKDtM4htqE6IAD4O8fi74h
s68lIbzJI3Jg+dZw7ll+NbAK0MZouZASsAU4lEZU2q9rAOc+iuBckhnJoj6S6WK9pkVMFFUFddy4
ZG1CQYlyTEStGJm705S2aMJLj5C/KY8HrjQxw/H3r0u1+QXAjH/aS0B0dUVQ5YCayiSo+wwEB8Tx
qFIb82d3ZcsdcfhJGtC7jxSDnXZWDqaLZLErgL1GkANE89wEM1yHLXMYO/1g1/c2ILFgkI8+9cAX
YfOImXbcnRkOLwYUEtFucb8rLFV5fqUtNItwfdkeCop8DcyF7JjdFeRq4rpGzm3Zkx9uUQj45DF7
pfJP/5KawtgIyiH3OYotGOAjI4225uiMbZq/3v0MGQNUSQ2RCtCq3fTYbWrqDGz0D/qXT5Akkuzc
5b0HEShCueO0i6SVjah4yEEe8NQV+46RxuB5dZWpqUdA6gFFCJr3v/EUrfSzhG7aRkpg8P/0OMWP
ausJFZWl9TUEIEYNwTrCrtDWinulr/INE0G2Py6Q1lsxNqtClYfV2WFTrKApGaqnm8vMPjQYtsbQ
hpxvJIa4wOqlOSzIANaceELTcQGD/L15o3Zo25weP+wm9nGeclAvtGyt7JCsE+/tOE52AxyYDZZo
utCeEgTb2eZeRt/wNKk6v7zAPCGmBYgH/hP6dzOG5U/Ulub/Mnlu+iHficxv6iCU67uBzmXrZIrV
kDPPkgb77LNW2cGN85LAhyoYNtm2ZIoSzu1+mhtq1wCElbFAr81GYp6MZ+pr6TCx5mmiU3As0krS
Od8iVv3F/XZTJu6OoyuFQBzYlI+6S2JVvAlHykAdWUuL4PP/9Ggeytd5fz7NfCrYO4XEFeGSHkMb
ceYH6p/bUpgZ6Hv4y6Cmb6r3c3rrzZX2rR0h4Rt6699jGW1Kddz2LLsBaeZ2ZDeXLrtZh67x7HbC
+k8YFCkwDF1PdRK/+4hBeDjr4bxtVO4E7wsrU4B8NnNlypmdur2SsHZRMFUmD3/FPDE/PgfHii1Y
3t4lKKjzEd3YtzORvIDsiKAHcmJThJ/7wnVv7IgFSJ+lv1DjtuDHdH/uk9o0sy9zS4wfYugPrje1
i3SxBK9smuWgosw+XbiKsPy0+jzWRm+jF+xEUDsvckfoOFyWsOOPAN2cXkyh+qUtuTehTHLnG661
OjRhAwArDIX233oz5BG8iQsS9WnUsLSDSlb51IeWg1btZTwXmB1PqisZZg0Vp/OF8sL0Q1duuu9g
JRAeGk/Qgdtzz2mHUM09iKGKTxWd0+UBHF9c1LvM64DAI8iEMPFoJogNAxtf4DmPGnRg8oix44q5
qm51fZ7yeCB7fZUrSreNYlBYBxzBiETN7uA77jhV6DVHXpUZs+QO0c1YjRPsXH209ZKJ3dQ7+AWD
l2raRYBnk/WmbJnN5bOigz6nmCwGyqc8aQbp6OtQ7q9YZVopTo0EOZSKYuJeOVZ+FYiKqgfj2ePe
9GqFpnRFsLzHnO80BkxDU/L97dUQHqKCNa8MqqxyspCA474IQghWyLhZ0jhUIJV9tAcypdna3U3P
8C+nB0itFQcBLcoZxhvh1lEz2SwoYAbZssSlqrJSMbNjFjPyoK7DXutEDoPWBLcZbeMyYH+yYV5A
OQOmGnsb/E0Se7wXb0hpR5Gb/+j09oi77F6uEDoohV7tiF0jbiuFmb59W8nGhl38yaACy65VGL76
FCOazPMGuXCg/s8cqRJCszy6/YfCo04ZT1Hc3XqTXCF63ATn/p3HSMKQVOy9y27VFPC3b4OTjcoK
8wpKDKlZ/+gGd2x++vtKD07oAhiLnpw0snhQrNChAfXwer3DGaYJPUkqteyty3v3jOHK7qmrhE/k
XN+/lMHihzp0zIrs0856INkCViZUIPkiObYTHxtRIq8cPbMFcoIUHwc8Lgwtpi04WUIhM57NhJwV
3rKR2zeJlmY9UAHTQj8SqCzC9CAIgO7EGAZrOmQjA/hQZN3oHijBaD3Y8zsr7lK3jgOK304947AM
87uc0N8CtpimbB++RYuqs6X4Z2Qfp2oWQt5gJYnDRMMsx7Oueclj/ANw1bnDA4M9rHTnWQ1ZZhe3
w3v+dAA8IutDyMHbSrJ5IVq316TP0c4kJu57OnuHNNvkXsWHT2aFTV5VWKUQRI1IKkcQ5ULq8HI4
egCsiuehFBFDsEqKWb+ZbiFw0s7cd+d/9pAw2ZjgJo6rFi5yV80BJF4GHJVeI29LA1ZSby5aC6Uj
00iarItI3/3wKLWi/3YYO8Tawh+OIrz+yZpXBx8oTMDe10RwLQoO1iEJFU44jHs4FfLRUXooqeWM
/awL/+hYV3YQ06JtKLnnWl0H6wsx4/PruR50DFWueOOeNy04+l78mYKZu3t9OQw5Ct8H1t/hg5pW
qAL4s+eRGxj6CCvcE7aTwbiPIkcI5EDDVOYfczl3Wwu+1lv/YaD04mpqCUf16XvAT8DoECqd8cmy
OAIPdq+QnPQIosBWHaZ9nbqatLxhfhO6nvk59WHGuZj7m24l9HFKs+KSYRfVzjFCpjc3iFFhtojC
+UXMnxc6hlYU2eVb8Q/tyrZ8Ts0AZQ5MsniJRRiJTPlEeps3VvHnWqjD9GqEesp8JrnzpNNzYbM9
B88rYdvFd9UP4goTiOQqJhKgFTyGNKmEiSPsp+1EeFPSLcXykm8tAo0fRQBRZI/z/fA5BW+GQv+b
OHIfUGj8V2jpVViCGX7F0OwCfQBkx2l+UTQT3GwlfVaY9R2JVMU3xofTJcmzIFLTPiR3mtARbx1l
ptoxmS2Xbo4Q6jhCstjfPiTmBte7RJlcu/WXTfuKYqE7a/4vXfTb08xIbI/xRzIB+hmow5RImThS
m1UxQIreSEMXtXniOALQd3k8a3UFQyzh/KOEm2MokNLpFo/BFd8hLe5RFF6myPsbKKNputKGSpgw
7R5XDwyHnB9C8UOe/iJEnuMKNy9ZUwzoGWYKKkmyTEk4MUKTEZpsWqKiDxgwPJM3ruVQM4s0Zjem
IMhGnrZlLq0qOvBSwvSVkVF6J+to+0OiZDdKTpu/37bCNsGTXa4njH0zusuCtnQ68OEzhvBmiYh0
CrNWYzYu3XwJp/pIfPiSzqeL06I4bjqlH2CbVp0P/ZsyfcRyayD+2/Jo82PnW+wE42QkOJ2NNJ7c
TNZIdBOySBAIbzTWY+OsBMNI5jYfYmYdEe3AOJ9ashh0pSck2jWaG07y4eCXLcUlqjSoa1NJZNSB
kbLAie2t9+kMNYsA0210BBQJMFqmMnFYY7uuOmEmIVl4AMcRRB2YWaRpY1EbdvklQfvdc68jhMww
BR8xL8jBk3Tv3AFxye2UKZ0dtw3ZmtNcWvZVkmkNgLiVxdKDjcN5fbOdlZbTjbQdYxzWw1tqWUwa
O/XTmgIJlaowcQk0GZP+CmyvkLpLVav+omK4oQWa+Yazj1IXWE9UXi2wuPIECMepB1FZya6Tz6Gx
lor4RwtAhGjimlwtIoxdvqkKk2aEaWDOP4rDP94limAc6Fdjdspem4yUlKBalsd/lPc1mdCJGObN
XHEIVB9vcQGMjmWNb4UQtonxEJDCkkkZVot4GVDtd5LLBXoFM90mupx6tX+lyf/Wc8HiCwLg1NbB
sstOZ2+4XuMUAdI9H7tC/VYJB8q3s16P2O2F1y6H/UORSp77j4p8njOdUU2U8XPtQDsewb9bA0Hj
7spYOTcBHdhIvoVvZQ3bcEZBMXb8cxog3EfBQ307x40Jp+fhb4k1qVi3M41lszc+c+eFp62bu6ra
jo6Ji2ySKtx4JIDf9BMiDbDXzZNuVlO87GRi+yYEL399VD3aIuWJUcVrJzw0duUa50UXCwdMJ69z
V4tHlzTYv8IwLkHrJWsDczNTXxgg/AdP0r9Ijeu3LuQBNV4QoqtDawRc+lsNe2NSaS8F5vrPVLdS
ZFDl5B7K8cN4086MIss1UZig6d4vbHnSW32lAP2urIJLTn8T+RbG9xCAB4qW6pLh/4T8ywmQ+2U0
o1AZvEGcLVbCgJED7TiO3Qcft5FbwSRLhtYhDjfGmF9/6Ntwqg5wB0dBMaOtN5pH4+Moxih+jEF+
nAHfschlgeiwhDBEZyVzYHNz4D05AMtRJJ95JfXu8uowNXx2WmLr6qd3FWk8QEfuBdgLNAPOqWcY
avRxIT4SCkj1lZqnVqwYx+/IR1q3rWjSe/EUHwuG/GbRRZeOA2epNzYtr6/ydzzLTcQGtgzJd7Py
tA6z00JXDu1qFpOfcaVQCFBHgyQumCJG7WrCnKHTy0eEET6eqdTn6MVHe1W8nG6b9menBw/lBQcZ
jk4lHdkdAL9PN9jhFsqxEb6JJrzd3kzQnkeS90F/bhDIgJcZcuRiOzXP6WvbhOm5qngZSZ0hwVCm
C+GJ8SiKTgVFMiALu87YU2e1wteh8WKRVd80SGWNO4Yvba3d1J6DwBuJInFY2IcTJ9fJjXhNshEj
EPKS+9nP3U5y2+iwJb6FW0Gnwz0v9pxk9C5rPOilBYeN3O8sTbJ7Z8W4uqMB3EnbY4CLooQbag7v
9RhsGJ+MRijN041tJ6FFDtl6geRkL40YQBQBnjV1htkiQlu4pDyl6zlWzzLaYitV7Chm5Mv9ghlL
qO+EhLawKBZc+jrbjzMsehLpNR3BFxZgOdYYitpDfE/s1vkKbbSNvo/D4PLDLClgHxQb96NFif3b
B63jBF4QK+Iv4hdgGgShZNgOzRGIslicgibFtaUPcH0s5DW2wjxG/YfKfZjXcChg6Cnj7sL4yzjm
z4bsQF//nhFbkdDRQZ1Ty7VqKZvj8RN9vqVvCJQEbSJJOb2W2K3ePkzjKbDFNqsSFsYgKG9DWcg4
NJkeh6Pud13c30W6d9iAxXDm+GKDgEjh+cy2Mhbk5OjXNAOmAX5QhATu8K8Ue8v5tSG+F2R63hL8
BZgJnsKhfhVmC/4cJr/zUI1rEZQBu3WDbwMOfWnuu6oFdwlC5sDFk4F7UT68d5DsxiPLUes8h8MH
jXaXr+14qKuIU1fO7INd7YxplnxDcEaF24E6lasYax/XjlsMM+xKdFI+rg782prH4DXnSYsbgU1o
DycgKHXfZODIpcthNuXfjoryaat46BuMiX/lCYalPGX6djA+0BXoDp7k964rtc9uRRYPC7k7+U0M
Opcbco+/AkysHtCC9u6qb9FU5fYRYOzoHu2pAj0NPIxDXXJn62/ZlBC0q+VEZIQF9qamYbVXvwZ3
PoykGVks/T0hxTCchT9wMJ5VJsm+mbOecmxsGxr1glzs3hD54lMcX8V4cOw8oZbjKlf73z0Y5Gz2
bf0YoZmtR+VHE/e0F96LJwtTl5nKQZBuyuchg+09KsHK/t+cVRSMBq+1vQ8RpMCN8xRNXzXpyPkU
JPN0QUM8a0jejq4eQxInk9SQ1TFtBUJaAmRcNJ7dJiDT9u9KDyVwmLsubRr/SX64c9uByN0VaE3+
3At9pOPeU8N96ahXII82LYI18SE0cwwEE2HlYbWaaSKPsHGr9rkvlTJOPuTPsyzyzj3KZO18gwTj
uaJu2y3pwVctWHh5z9GSoc28EZm1EY+M0L2NZwpNKQePAslrXkreTD6/Bict4V5Qc+okIrTAH/1P
D5i/mRn4z5Tvmal1sU2B82T+X9L3JP5M3H9TYHQhbQFKaabxO1VZqzBvXQ8ldHec0Q8Rj/VzMCAG
t0eBIQfFg5xpRXORcnnQMEp9DU18DcOYLgCiB+Vu+aLAWU6RUxKM7uwl1GfBVj01Gw0HGjJg6aiT
iAYsJkpFZyMN81bhysylF2mtRqBTZP+XNehjF3o4UGijpMY8s+uuV3g49cacIG85VIgbDWyZfNiQ
hoXm4EfNx/KaHgy4ot2BedXJQb19LsoEX+9FrI54IPZeNUV+WanM1xGOSeBvIp3uJw7hjbMSlu6E
RbGClbdLlv8aiOAG9KLOnJ6jSb/bAQeFAX/elc4mjNiOPj+uM3KebqprRHTBzXEi90Feesv4u5Wl
ZorNKt5CE1LZXn7n1HXUoamc9xDnl8727eIg8giZBLwv6rQ+CY9eguKKOOvrpl0IGZezPSpTE/ZK
p23zqRRtfBF8/IaYSHNsXYdgik7ufDVE3bHPb+N0eHdF1v46yxk6G4Uqnq0gCPWNsRXxxyYt9HXj
YYbMe/OV4FPcVUgRIgrKkh8UPmC2rFFyAsY1hM5czsjTrCvv2D2GuvKny3dYxKo3HPvYBoG3VGPV
kEPw0nhLfJR4ftuhZsDqGQSrBPLbEkRuThxSxt6zFpZKcvgWqtTWQtq8+swnVFpjlGs0tHQ/fV8o
rz9ghCs247QQTszvdpq8gdhnKsjoB3VLnLkxHW//hb1juqyJGAdcHMbSc6hA7qYNHlGAkKkNpW4l
7u5jPsYTWStCnfFMBL6Awz3YgTCQ6CH1zUmp4g290KywhreLQZCj7NKUKTIYtBshjkBIqi1CTSZf
Ik6cM3VqNI1pDzktbNaMDex696ec8YxM0g+2tXf1KrbNVIDHu+ytA+PfKfVH7nO9sj75kEHKll7A
6oDDIXg8A2NTzg1+WFOt2WkCk7lBnfdWhve9u2WNbajM7MbfKa2Sk+agGEX7mOT1UISJXVA+osWg
gCkKMaA6ZK/VdFbXCpS3jZsNJ5J0s2I+qsrSmBWcLx146UcFhl2q+AnnWlRORMONhgzl2tVoTEVo
Dq1/zC87mPLbVwTHgyXqX3Oj6LmgFHkT99+kB1z3HqvqIw/AkV/hN2nOl2dFf8+a9WqRxUK7GQ+W
Z6HZnQDXl2TFm9mBco7TlHQpE1+YGbGfu+dW5HTNOnrDbwot5y2CxwETNGACRC4cAMrFy9baj+d3
9Y24A8pL0gi7CKviMrJ9lnnhZS7VW48RFsPX+rkvsfdRTdJhbGwzKTpaxx4im5XN8EYqB+X+Ti7Z
nYvQNaPFakkJsR7lGAjfP2O8hMVlU78PbzeKbK2kRpvlFy3+bqSF4SZ88PW2T1bWow5uGtyd05ua
BHEGIYR6DqS8nMEWUgRBD9rQKoByM5zvcGfe/My4YECy6MBR0kIZaN8v1VuYwaFyaZehkxclnmP2
WN8YmZJJzkOR4NqZ5aDEQk0YCaP8BOcvGlPMLzq5XFty/fHVPvxjSkK3hxcefX3taT4v5J8R6DTy
jFq8UrCi9GVGVsLUcl/HfwG43VjceuVPgwCubKJUk2YopoorK8VfcnA+0hK615w5K28BD5t+dv5C
pVgApKLqhUh2fY5ll5yP8Ajw+Dx62zGB/EXKK70SZYTbZMz71W4nyttT1i6iUVEKWdYEb3hlMWmY
fpwPUkbn2wrL5Ig+FFKir8RUoHvxJDsd75xyIbJnILRdsXRYZUbSaii7byGCeX4/s0XEQG7weCSS
h8/lTXgiLBksw/U7i0cGmYgNc0kRpp/3YpF/kge8XsrC1ItoeM+YCSE5n0vD75gi/XSFpKVnSHq6
YS7Ao37PtEppI6IOCaA1CxS7EptyJxCTZ5PBA62hN4tMHU8oDswt3LU2q5fhcH3o7KUeytQhMmJO
9kjKA9Jhn1swNCj60gU6fAHZFnwsFnHzRPUMRkfewujgXcAnpy/sAFCpSutEUjnffRROfqamqGVL
F1wi6EQwTmeLxExWlENihr1y1Zwmsd2R31Q4JoGwItSY7QtVJw+vUIWFqqkfu50ok1/qFjaDIwqZ
HlC/1LvqwliS+99wxtkN4tGqc9e7UOuCLNfSUD9rPjaM7by5g8csd+a7R6o5kRnbuYz3HmC796pv
ScWsV9GsnDFO3lzGoFjli8Q3ixH/zpHwOPNDUwtpiP64hzB8KKm3mcG2ISN/OLkVyS1Vx9eWr6Ci
XaQGML7HcS1G395JBib83A9FZhWSEhwoTmZOPsaJ3vFptBoCwzhyJMIebFpT1ilum8nQpLsFOJIk
+5K8qQQ1dNmgdhKPIeXjB68afRhED6KSIlWNKcgIoa5eiFcaeH/DdeM4qwNGlMlwymSvsixSU1FJ
4JUs3Uisuszv06irdTH0+6ZQTvEQrG5Wpgo4BZJW/VCGoFML8K1RwuUZoOQnTFhxQsF8euAiG3Nv
HR2mQb/D0oqsicBrmDDynnr2kysSiLyintuT3lqgGsqWbyHSTKevCMnij8OrG2995NuSSp6vdiEU
aX/pAIpA6TecOLuV1IM4dykVxnsWsSxgpaDVq0vDwdNKo7BWnvgLEkbf+p2d14NZ140Up+ePiaMx
8gPcXIOEFIQ1lXfiLH9atvZE1wuF/5zVpUUmevbHMTjaF49FeH+Kx4JYDO3xIl6paVxt1JkhVuaO
x9UCIfibcWNtsnMRwYV6Y4QTAwFNyhOHn7oQQXxkbjYy4DS/nRkTmealrTrkr6lk5aGJwsH8RIk8
8alqiLnfIZuTBcIsdilQIc4rhRP1sHd3Ku9QnAmMPpBG30T0SRSqZFcR+NFQ2SIvejBJtXjhwnGO
+ZtOBYYkyYVaWXPFeK1o0asTDND2ug7MmSiomqVWxZX5YAiqqF2LwElfwxN5Bui479ZqorBiXkAl
NvjPEJZOWez9MOgZv/pake2YlKV1/4FYPpnSI148SyngC9BYZxPBJot1EotNp418wVGePwljPe+Y
mfH8L0qSwY4c2j0gx0gbCBfe+AvTvpQgokhwbw0o2fc5OvRUJr6P+3VbyOVURsDswcM5GGsKx4bo
2LMAiiWMLuc+W+qu+VAc184b1t4zWJpZaa3Gf6PFNeGaIHfvuV5GAYf8vuGw4zeKQqWolbFFEyWy
LVF5r7EwrUvIIfncNw2zyqpOK/1n1U2Vw0AYQ3aE09jqcd9BqI9Rg3u+1foKdb/E9SWjXJvKVqb2
/s9HL1aBWt9kyV5ptzYtC5bhQHo0vpuidgTo764lHRFtN+g5WJx4RnsmdNYlAK8hcmcOpzev8Cib
2l+4PZcqz5PCVGtHw4xQjgGdV2hD4FEC1eAy1U9QUrJq2hcFm0dxjPZk2I2RyWUq6H7emHKOA/DL
QAl89IxHsZFcvVJ1rc1IdEuNyOoO/vDwb/czXq4XQK1s+2dKBsJGpsH+/CuWkkPi3owtBlxvseKH
JfFAMPlRtnQrfTbUJiFUjQSU4r9BXj9q0nxiLn5yXgdoiPtnxABDzS5OZ5/auywenXM0LzoEcp2m
92ut7MhdvjcQ4bLiwuxfgpxY4vy9Z702S4Iw6yTK69Q7U045GLvsHY6ye314AVXJt0bUs1g0MIPv
kJeHg0mnC+KkAJ1VOLTp9MunygfsZzpjV/hqjS7LKUbl/enDWbGloIgA1PvKgT/vaV78t9lvd1tv
WBM19z0e1LPw+Tjm8w3X9FxciYbOeHIx1VBUKR+fWfueDBo7OTBoXXgkt1CvwJHBknR53Ogeawai
FT+d1S1vqnrDblQ8p32bubZXHh7xKImiT6SKEG/iRn3rkyCSokvJ2xltdnz+jK66TzmmoxbAvcgX
KSRjcS3NDFhrMYgD1PngsEY7Tx7QYQDhxzZskX4tDgR3hwD/4N+jSY8it/072oe3roDg6wpvdQb7
DdN9+4pirKlt692yq7BhRElMr6LmBtJWaBIUabaZcwyChEoDDBAn2am20fAN1Lffq+j4svoGx/dz
U5kjXPLeMJpj8BGl/BelCkyTBuxlwktANoWz07wq0tABnweu2fphfD7ZJKrYV9fC+fQM+gnf/v1R
1dHAwci/cIZEEe/DruLYxOxaW5jffAHexEq81alwZP6rOE+/E9HY329HOukHzTXoNiHzVLVDPkJz
vP+i9E7L1kGKy0p95nXYyMe+5ruFDVaRaqYS1p8p5Ju9ShOurQQp/HpUbVbkAvguqe5p7yCDcKWZ
hI5TdeVXhZZ4CKPusrpSV3ERluklPalb00srYWVnbei3x7x0GLduSKYJmV73DE/ou5VRauAYNi3+
umJxS5lHMic347MXCnLosBF7oiRoffAE+RggPjOwuuaWz4d1oxJ2E/QziYs0dvN+eCIbWvJVMvYa
VkvVqhXFTUoFLQ/mjzMvrR4/JRFbbeYazy7hxhJpFkTYr8gG8qksnihlsMm+PvpbgFjCQjpVf+4D
Fuf7qXKHRnRiXPBFJYOFexYK8N73inp01SB+QRDCNkdJ1qIYr4zj/EGCEmOa9dTPODK32zsayjq5
viQXjTJxh7NMNLAYF7s4noKs1pHOId1LjmTnkRgvCzBgIvGTlpxKNxSau/8qqSdnNMA/HYnhjcN2
uhXR7mi8Td+JWlfFPXkjhasyjlasQvaRjPPRoiG4x32lb26jGCqYtMUMKI8cod9QUF1/LtIcbDEL
yOB/l3hlAEJ/j90wL41Udma4aq5sk5ifjtCncu1SATsWAuyANGZZkFFP52R6Nuqd1hhYEcl86bND
aARh/Pc7xCLHDrEhTHrSF9x4sO6lSXG+Cyl22rUFcRDfxk/fKALRGnCHAJZiPJhSETV6dm1HWLaD
jPahY4Ep5GY3QicWmk70iFuHSg/7mXPFlNpZxBmIexlL5u+UdDDxHw2cO64Lxx4mwpUowp6UumXX
jifZdmkkBSaA1hY/Q857CXMDajAH6lU2NpOc+S2QcnLtallhqRcsn9UwWaKgvhzuuDMbxR2G7TLP
s8BvHNIiH7JRyynuOYaguHYdC9zeL1mONAmKnbcy6e/ZDQfT6Re42FyCuxIjo5cLjfFexrj8EKAv
I42/zzGebx0jMscSxNzFVqS4xpADE0JjpjT+uUyeiNk3982EYdC5h8gI85QBglmSHBBLD2xefYBZ
xrtDZFqEth/wiZIZcy5F/Pr/fgNnGkRcHIunE2dEmDAYLwIa1sPqe+uL1U1N4PEaYEoTabbysJ1x
Pz0noHk9wZGsz3Tj3/cgjalfytdSo3TQnusxz5b0IHlcOPYwVrLSJ2z/32vf3bXVic3XobVG6AMq
bDzmcqd8s2i778AdMbDLNax1+g0QzhcOnG23Qio6SiuaghxRomtnfO6qr5k2km+HzSSS8ndOwX14
foI4DD3ChHVrDuAlZMiI+jApXZT+CBDoCnSoGY4cplj8sm1fyAAuB2uzF3yXo3mv3q31PzPPhNhf
cilFldJWbtfaIiAwdriF02vtQdRQfGceWIhka3nfbZQYV5Unlg996JOyGZTx2cvUkceuE9NYSUq3
xW8iX7vpQvmU2bKDUbNZhcmFppiIZ7DURUpbZ8cNGIBT3INTptygZvRYq3C941+yjaU6QKXEQ8Gp
WFIyG0qwGTcg74Il8nfWKyp8/6a6OQu/Mpy7cvkoW9ndqOLOu/Asu9pA9yXi0kSAk9cxB29El8FH
+4kcv+R8N4l8nHaC9qg8QjhZPPJ6wdCmg3aiOvEI3cWSnf2ioROSub5UoNl/QASF05EnWyibMJTe
UxNXOaYHEMYAuWaEfiuGtYclJOGlpsP7HlFiX+PdM4l48INO5Cgmp8wpMOWhp2Xj6aRC3+10QmM+
+a+jZBCeLh2CCYKZQ/WWFmIxeUAaWhtxNo4LJtA7hetDPnjHqXXt6ZfFz0LUFtPNIOmnHVnz4vxY
eWeqeaTzeu1qcDNjKdwEiZDoPsJHhMf5esKDhAZDXJaRcXINV1Fc3OxSIto9QuVlzevQX2M2lM8X
DVPeiun94taStftpxW+psPUZqMdsq7lNqXfgfSIDRVboDKJbxB69wiRVZuMdbJflO5LMKtEl1Qoi
MaMrk+FoOPpoK/X/MTpPTENMKjYxqgRsjNcDOY3Tl/+gKNvUoE514RPhRtMwjqE9Zq2p8lBSrYxm
g/VuLzK6cRlGGB54j0wvyo3iBy++1Td4JemXMdOQkUUlbRNrb43dt7O2FSF/g05pXL/8dChyI7ph
BKkbQGEA0X/XiwUBhKcsPDRdTu2oUJcQYxRDYyHHDY2AUqTA0QU9cYo6MYd+IXfQDzdW9CtdF71a
D/er7Io3H3iAofFJMu9AfyuVZAT+1vqR51UkddQsPRxeqxfoAHCSj7PiPH6M+NYxcG6KBASyfghH
AAaygmLKho7xrsiXZNk4D6sT6a1oYM7U4xs4/7BOZynKUwfxldF6LUunYK1cHAoRBiBsuBuiLzPr
AuQiWs28e5izsNyoSRFFxU1hwwFXIrHsdDKagKG6yaengVq9CO1jmO0f6zRyvq8YWKHK/2T94zMR
Boij5NZ45Uqow2pKXqQWevHk4qcv3lCwA26KTo+O5iYg0ZTE17V4/xbBDPeZeWPgKRbK7Ok6FL/q
P6YeQss3iVSAutbAVLHdjv4grK/s/PbBT2J48tLH6xXg6/ZsnjBhNZv9HWsIdobGThSo+sncsfEu
Shn92C37NRGYFuoQF55+oVrjoT7gFQg/NAEhFGegWaAIKjcCzlsbJu7Sm61fxogKGaiSZIga2bDF
ruMM42V1Wr9yR3Zu+UAg93oDUJoe6jAugHCkYxpUSdCu9a0cJWkveYY1VhQYz7V55eH+8pK9w5la
ddaXHJBarHbz7C6j+mRgkzHqH3H+KEJtgoxk57EOuU6iH5Cnz+OI4B/WlDMPgSykKrgF1+Ien7Hc
cDp4qaTrkd5FGDLOzYL9sVB7fDqOK/VnHB9EPZOYFrU/ofO5k+fvnrSfbHA/l8ubg9BbPIedmMx4
oahyR0SWbB8gHjRkLy0C5Q9MI+ms7dpLbKeV9jYllLIONZg3Cggo69fn5JAIgtuYj7/BxZZEq+7L
7uZ4bd6ySDftba603709/bYL4LMdaCR2zAaWOI0l6CprkuwpnujeffWU2aedoeTxJmAqPzTDyVXa
AJjc56SNJ88JOlcLzTsqRaT3Vw6I7lS0vHjRb5JLHPKHeHCf670EQhF0LfXtXh97tZQm8bKug1Ta
R+gjTBrvEeeKNmdfyzLjHyTWjhCv6ZbgkwnZ88+h89Np1rF0jpj89YHRBC8h12MNlwAybOojBHVM
FhODIoyz+7qTfJXqOkhHSF7xs8TtrP+6Ef3xFPGUI413L1C03AOG3p6TUlTy/CaQ73PI6cnfHTC7
9oOKa9wYQaJP8wJ5iatziFQCHjI5m0XBi/riY0CMRCMVwFGdDRyXMo/cxM/mYbLY0Ria18lgksyt
2s5i5kF51Gh9AAYadhLB4wO3jt1GawPcPV0S1LRsdWJ3LjF/uUEEi3S2lCRBzjiwAWQ3VvR5guM/
O+blW4mtvvdwa32ENFbCQg6jBJuv/38DCvvidk/4P8ruXkJJMWIAbHlpPz2ho2/O/CkjPWlqQfOa
/BwXgMn2RzlQg1Uf3je2IQEoUQV3pxMhJ5t2xrxuVad35L+f0ceTTeF9x2nd8MBw/P0KJf603FBJ
RHpzr1i4GE7FDA2EYmxE6Xx1jE3mZzE32k279sdZhWeQJdhPD6nNcH7HmVlJHX/3U0dh3DDJAC8b
tz7Zz2p9oZIW71r/AYlmyTWbq+B5MwWUVeRyV48DnriOXIMm/Qsbg1g8CFiG1IxIfk+EO+GdvqfP
DeO6AO6vmX2/qrjkCmQWo2lKHSK3FXDkijNBYaBf17NkQfq6X8fO6T2guSmFDQdF8W3he920IGRm
GDukcVw41vy9H0bqgm7PkdNOAP//5Mb53cHY+jS5R77HpfCkhesKkQYWbPG4wE2viaLqvGp2pqUG
6uLAdB4GRTddgpXypLqn/qRtX9af7xpPUPF88Lm/m01ieVoojkisMAKKTN4piFlDEe5TFBoGKodt
PiR4YLx9JWeziEbgCaUsck0eQfu69f8uVruI0AkKywTUPe1dhCQBEGD/Iwb1EJR7xBydEw9cjlSb
nQfMm0gwtiDSXXBwXHIiaRv5xWZNfu1EyqVYqJQRSxr3i7mbiC5nUdvxgryW3xWnenld7fDVgdSy
KbBipeEVDSDqfT0Nj499UGaoZs8nMzmyTvdRUE3rG7rpPzaWKlM39s3BJhRXmfJcvmXyvArYvouM
erc97zHZz/+pCITUxgdiDno8ZIRHTLsIciJQmUyhAeDjsbpD3K6qnTZIZrj8U+0oHYLJR/oDCpWJ
20Ko66dCmjVA3y69T8SKEh9JMcAPlfk8Sxlcv4LMvccUDNA+aiBi5B2QvLMh96BJwXeLM4VzaKg/
eFOt6NhhDG3DOFKlGiwjeN62htTbENhEBGjG34Qk7vZW943+8CfiBPvTMsyOQfRNp7SXSKRzjImI
+CLuYlrWPzLCweHK3ulSpFLfdh1jLul/kMUDdmjfeLGSr+ZrmqLDpyHo2JLkGWV+3vkakBFteL2K
qr3exc8Q3cwN4VcyokVXbGXqvsOpO/aNZNYM4EVakhQ6ag26sxKBYi2kb+KE+C4zsd2am3YEz9fT
ONe19CPDEMJNGTa8FDFP963F+CWWOwVH699fEIKPGD0zDXR1r4Bdd3uwirKv+GXqXSYgm2kOKTzz
6vbBVkhBlYgaqSXd69elKb1f/hUSDamnKqPeg74XiybBQJb5durx90FWNaCUFzCVrhgrNcy8GOXe
PxwkfJjknq2ANWSIdzN/hDjZxkpznIhdbhl82gqA5O1x3IcMAyemrI7LcaHoUkcGgnadJyy555DA
pofcdU0v76rmT3n8TNLtYYHG9OjPYWRotufhF7BYp4/NgjZ99Vh4+GWXfENhGLVgsm7cO4htEF2q
ISBByzKiItbxEEm6us5K1vXUZq+BhzGpFHZGjT3UOy4/LRIsbm/rJUV6b2DINDe5OFOKmFs7yXtm
qyzoLgN3+9asYhR2QE+DR226Ze0I+Z+lOvkkvH0lmTdOtUc74xY0EiaXKC587dWvrYPqzeZcFueF
dBTi32MFoz5zEjwvnSU1E5B0bcsoMk0Jb7/GB5TJiJmnNmx+gYXivOtnxv/+XNovgx1lDPDj8OCU
JetJUNvE5NCfTwQR86qXFTB4jfSfsuJ67hUK7PMQ3bTEL1xetu9pmOWKDSaTqsyr0wsJV6SQCTtQ
lb2uQgAoAYZetem8kd6fKVCyZP8/bRc0W9XnmuD62mrjMCTx4mEY0jcDleyiQCnfPLIsdMklXYVn
577GNjWlP6VuMDN4WEEx5eWjdQ502pFsvBleQ18zO++Yd8n2wnATqk/7K0rs1psaj5cy4PwjLfKk
MAWLUyR/a8c5g6mhJcIUaftm+1sDfugs6SFzGiT2/jmb4eDtyVJUI62JJIJkfNG58BUpQPTaiVol
jTpDTgGwiuNTZv220Qjp5QXHm2/DK70IKulCH4Sa9ILUHQSunpPb2FKrfkDoksmraA7Imf7RoWV6
Oh6UtB5x0Z4cKIYjAjkFzyt5ifws+bsTpIS0PGO/EBIp563k9H2osUcigsxKqSheUKxfFTqoL31m
amwEx3wcOrWfbWcSX8RSJIA3uu+P0CyQ+MNP189Q9mq3Z+io/4YXaPMLORtcAmbp/LC3ad3OPDUN
n8P/dBanuyo9OSQLEb9iQpAiU9pAb0Ld4WZ1cVlDe2/NoGdH1upEa3jatrlrwI2SXwB9gmbhJqUS
q9md4TWl/BKEfHdXsACG7Hlp4XFbtkmiydajHQJPzCFQ9Lv1pmL2kR9bHVtmXG+Wo0Z6kETEkhTP
wdEi6ufadPLpqD5DNJOAL0qc4Pq4xramJQZYObBQQeuQi48nvPJeDwhDR0GemU8G9k4krkcqC3xT
gfV5IrT0SXfB/vAtHzdO0u9Hjlg+tssMF76ibfIuKqeveQhle7O0MZdDsmX4Hu68hTpxUD3JgS83
XgqSLV3RzgbrWMXN6MLLPkO2kCZYOzZ82CiXfzcLrK15MCA7Dz3UR/Bgxv64PaYsu7Uxc5xExDBh
l8GnoRJzAAz15Bt4CBtZC/GjFdPuQ6/YfiIa0ZXZYI/qEUd8JdpoFJzt0+KIla/l80y0Ua1eaAJb
2YkfdD3fqjnFPc1KS0l5i3gLkeQKijrUNYNqzGyUotEagm5piEIiWuG2yNGfiunqWg3JepN2cG8H
Ix1UwGa+uKzdUDNcpUVeUc5DFH/rVXLGh+iU3YZx6evC5XGHayYaUK5JsT4eNelkaG/O/QbZwsh1
dHFEkkM8+XtmI/jnOsP8ne1FhLY3HkgkqDlr5bGCluljIHzFHTPaCrR7FTThNlpEjGpgdrwhDO2Y
1jhri+Rk6eMB1ruxy+5fGTGSzLGaeDjRoGLJRgr/7KK4pisCwKRkAyaYSZ4iDsZQlSqX1L3O3yRI
MdJDu9NG2JDb1O9mJb2inruqnd0zVicTvcCZv+0fquUswPNqq/9RFeie+QSKWf5lKbZr/b0akl1d
grY7+9vzAloBxrTynteuvRPe6yh6G+BbW5xvTR7Y+JRI1dyoDXpfXHWoTb7EBLjQTv01+PO1JSdU
MPcfmVtYjTzyW15Vr25t+WqH1qdGecUGuVegaohhx4mRZLPpI1pDM4MLT4SucntJMPCGq14/pQpz
HMIveK/1J/jS6QJnaz8YlKfr2xyuZyA6wDohxEc551cFjuXHrlSyf+lMVq1wOL5mVUEJoc/RqVb3
gKzZGrKPcPZ/qcNoc3L22u4UuJktCDfeX2vhfF0awIRKXHinxz90tUASy8w9adAWZyse5sDGGbBY
IkLl3kyEIi0AkiPqWpqJhe0LFqkdp5sFLbDMhhqpai1ve4ahAdN77qrsndjaUn++EjwpJ7hKApop
jHA2Ez21m+S7Y2PBt2k0fNHFp1gMorM60hZKH4K8awaOAC7wKxlkTKktqlOCGjCo57HXQIorfOI5
VFOTX/PC/Ts2Zebs6z3u4g9+6FtRIj7eoS8q/64R2C0k8SRahbNuwXyIgjj8XBPtijlUkdjU3K3u
KJH0P9NKekHDZH9UdifL8ZuTGzqbdlhiHYRS0PTV0+KMVdisGAAXqKYAXu6jSaYY5+lZxNEgdMFp
kQrK1z4qnUZJA6a8XhxDj8Z5cwAhr3cyHX8lx/31FAc+AzoSdjzg0GzgYt5j1OKOXYNFEgnDjTOd
AVUL2HC19/hCdZCgJDkULyJPUCxsb7fM6qFJUjHZZVhiBY47wb5aBAl1NpxP2rrxANKTPTOnDwLv
nTsyO2mEHZ+hN6NNt1LOJd2/p2lMhpoMZO3Rqs3MHg0vCOoTsDma+Yv3gIPBY/Rd+nv25yQi+cBP
LdzsXUIqI+xiKyN8B50hGSaYYRiEjUD5IauwabfZQJrFatDx7WmVexsBhsilelXkcMDElQtPN75V
+HRO0LSb/XNg7kLJU8iMGy4T/qlYpNaMbS9ilSz0E2Uhq11Bp/78ISmbfXHPqoCrQwpXRAztASvl
HDkZdf0lVtRhFo73o/bmN5Ce64v/IbcnZdLp+8FOEVv6e9fxmWvQWAyLrrrDLGmc0p/4xI1yu+Eu
V63zD+G8yIRgIBjSeZRNwCIEZzeThcv1Wajc13jBVYpAgyTkWu5ehdFQSgD65P4sfCpWYfWFGs7y
xx5S2DYqPluQm3+V+K2KZ5fR+FOjhCbTRa2vXgs2QynIIrrR4HQAbsGOmJhYEnayOhApjnYG9Zx7
nB3gViFf6d7oo+RAjHf9lS0fo+88P6W9FcDPyeodiOWM7w8SkbmiT13mZ0kZsNoUDpPWXsrJVDNO
K1X8iQ0vxeWynxXzbSokfaqKYbVaPAlPyjWPHeEU3DRma/eRz2a8fwk1ZEsh+AsVtN8vnfA8Zn6Q
ISJ8wN/QyN/InfZ9zT0JFEnK//A1EaejX8vuJLdsSyqyg9adg50G8Ho7pyihN3nEA2zRDjH+FdbH
REwvItK6wCLbo+lzzSzqhIc+UeG/TLovb51l3xlWae5lxxaV5+ajiLfh79yMj8kyeQSj+rc9Msa5
Pb8euVi8bYo9QShXJHjcN+Fnnm4Po7yJz4B48cRPaHzNv4BE196EjqCZLZTAQCZiLv3ABhUg6qwW
xWdpshQIVJFl+Xvcwt8KlWZDAhvz0wm4kfAAJo+GuYQZrFF3yyhPQt1KrQiyW/7BA9GZeqbsNiKa
CgWwQw+koh4jheBciISZFDvdeEk7iCci9M6e0zjFL2m1bYd2Cqpp4AqehO34LS0V0IFL7Lf6m5Gz
ah4uJwQy2wnpYOcR7BOUu+ye6xdPM3s11eNQ+aqQ/bnHq7gEx2Urv1Rl3ottRD5Fo/uqV8sZNu9j
lw6h7EE7TJJTj7oPHFmL4RqIwYvEx15wSpvYf3rrLe6lbqYq8UQKoIHMTS9yuILpHmc1HArLAKxB
c4MQGS4z+kvruKVvRI6J0Zz+EBa1vvCUWpb3yqVJJXIAwbHYRYXaXwI0y2Z0NJLLgYiaMbDjkpsA
tLdmiajCOPmxOWOglpyR9fjT6Rl0Eh0O5AJEJua/M/6SiUN7x87tSUYcTFiVWBidkwNplWhm9hr0
NzeYwdXKtX56cJyzJqOjQZqVID/V9I/xXGZwBQ994eZeEFL5kvXjagomnlfWW0QBFX1HfLvXi7C3
w9ysgRcPhU5WF/LZOQEupsYqdRNRrnk/XxHK+5T045x0iAwqSXV/Clph8OZNLb6hXqL2LRthSfiL
Uw6uG4VDXHkQpDYu3sMeoB9Ka6MJMHj97Ih0ul6svyp0TaxND6Pp+RQKVUqD3Ejw3yZwu+HyvVpT
paGzlBiWpIvXERpBcZLbOR9i2WsMabDSJzI3s0rj+uprv+Bgzhv9rZ1B0ewqe+159qcmlbvuGcnH
TPfQ2scEDc1Ci8NL8rIKeBUAaSaywy+ic/JbaQjlD8r9XccRGCkiep6PAXbdMOedirv9uUa/EuSj
nWgx7C0NK+tP51b/pF0gdTORPf84372YW+thTWcOt7Naj4fahWm5V0tPEH+ETFT3sWVWx7T5/IRA
FaN7V6qqEuGi2plZ84bkJwybnRmoZ+O6g+ReeEVuz0SnraBd0YGzcM8Z8Ld9eqTl38UzLA1eR1CE
8BzCBJ54c1obZao21Aa4Pyp0W8YHVhvhYUkxQHGRG5aHbcZlgpUGRhSIZaxAHGkmboCZqft3eXRx
kXTZ6QQUyBD78njIcEN2nAgcT2vLVb3w9J31UqzldoeDDKIpeWBm/0CqYR3FaVC9QjloqNTYHowB
8zlVaGyKJx+foE/gebpQp6c+zaXdefcfBeVqEzhgn0WeOe9Sj3gMsuyH7nBZ+UObBa8UfKIDMrOl
Q0gq8YTskxtQA9fx+KMW36x5CqBLW8tG4Wpr3EmR52buo9mHDIOVInWaGQR6Em3weMJE6d9Co4kk
yvbF2QIeZroYZthXogsogEpUlrcTLzDOMK5tKQUTGWXrqdRm142ASZFwTWZTZTUeaMiV3iX0TwBY
P7LjcrhSXurad1jdbTuXXwdbBv5CrwloqvpRCcMD0qOBUcyd6TBDuE3gQ3uO96Vk/1FHQpNanCpK
XAWKKtFnqsEQ5zrJgTpdM1aIntSBE5t14kMIFDnQd1gzOod3tskszm8yzm89XXbGFyPLUxg7L3ii
oPk8x9EnoTK32bExMXmdXbUytZqbV1WcXcE5+Z81Ydz4hGsxFAyh1vBlvPhxx3lV8fKI6cTiiV0G
oKR93YvK/Zs+hZdFrltXe2VixnpAIEiOw207jG0Xb82M0HIIKGIQGX0atBBM7gxT/hvLLOkDP0Gr
f6czdChsEFG+Gr9ReUYWb/wHA0WnHwUUL01+YkHBDOhcn1HrJnNs3dKT1E7kLki2M37BQ/ffJ5ep
1FIAy7kvJbWH5Dx2eBuD2pcIgvYI91WXfZOyGX2cTNOtyqUFB9RvvFMpY+v8+b5T/e6I/hYdU4K8
FK1SeOtubLrEYGrcy4pD39k8wbpCbf9lOyha1MA+oCrFBUSgHGG9k9ZuZqY0QXMNsCor5YWpoOol
tlJBUI7PtZd8JwnN5ElhSPuqdg0dhlsCljYi/nk4MSl6p9saBYtgH9IJqWWnEXA1UJS+Nos1DNTk
LkfSzpSYTFdMFkdU3qispAS6S1e3GTUm/I+SrL4vHpqJXR4i+1oz3hsSCE1BaY9Ob1Ou9q2C4l5W
AZE1FlKB7qJgyXH8EMXsTJbjqqPyzIET1pJnP4uHqaKfHhNcPOVF+FKF2nqh3lw83Jhem3zANJ2M
WGTGwkwa4tgeFiV2kFtXmYBih3urAKw0StPRR5LW0C8oPwEpF49AGT1n6wYRHx6+Bqld+2HJufbQ
q/E7/DuFNlFkN8yY3zsDPGIqi6yov0h+Lk82TAm7vcRZEd/tUpZSddvYW2yiuxFlMUiVAWx7Dqj3
4qpkbHefOhNSmlREhgNannlJzawLkv/15cFx7V1BzkpWYdfaMiPOoY9Vw+OhbE8my301kaqDuOJW
8mgP2YZrHksdNDs4o3hNss6aZ2zWxsPzW37Qjs/gObIE4mDm9Lp3MTf0bLdabgFU0f/4Dx/6Q0+3
5tFPmkQC8lFzRJnwmhXFy1oBtxdpnLq1UH6+lsEpZmrtGqxG3Ya/D2AeWxUFLShzqSSmXPOEjrTd
tWmvSQ6M1/lI7BP+1VcKoxhjGaHZce+xU7PRj+DTPw32B+mKVgwpd0DyQ1rZ7cdRI9Qhj8eIzr96
SJxoMRbsdEJkHYcuHsJNdK/mJf6hXCtCkG7i0br2ZxJl7/bUSlPb1oTlDa9WZw0a9yGd0o2wyYG/
Wcts5DBptepQQZJgJpGm/UyPmFv+t23+cXaQhVBMwAh/aIJ7rVP5tEGJeBgFw5aNhNdIqonJCgiE
15QWhWHxyylWtg79Psr1aeNHJzqz6h/Imj17hQE6Dk/GUDgGY2Y7hLh4iIl1G6lZn9lGzLJEfmiH
mKhlkU8xcUUd/APhOm2lWq8D27m+XeR5AcMZhI1kBnVyDbLHNKckF/0gL1kwhjS0XiXYKbWNQHev
dAogM0fooaAzQG4KSgD6Pn5BjXfZkKQv7rNKGf3pXzLO9Fml9lpWuvqa/YsRYYE7kXzPiDjbAGey
A7vxLDmZxt6Icqv3EYn/6OFBuwptMUMAM90nJnEkErrlbAdjNOwr9l/WRGDbjT21Xj6kzN1/b1ZO
OWkXKBA+e99aaqSLbQ0CPJKBESeYtN0SdpKpTCW8Vep1wUZ2FkZvuX66CDdF8PJi3xr2P2+t8SAy
lhN/roWZEzM6xSECPL5+tv29urb/8WJX63LXGXCjF+2kk6r0q4iHLRBAUVSIybEw9YtvTb+GYarM
x0VwiLgOAnyqHcpSo1Ywn46D4KaWBcf0lbWLXeIm3jkGfIN65iqXJJXdkezk3zq0l3GD6yj3U6jS
Fz9aKa5jTz0N4QxTsrpCNNAd0qert8MgNcuFQDQe7DQ94gn4T9K09wPVzP1CG1H7b+2oTa5F7lWw
w7R4Vm2MAebKhtQ4iQAZCqX6udyIEC3TUmNUTzMkVC6CBbeY/V6QhhMIOKl88IZ9VDP5Z37zEJmE
WAvdf3G31yFP0UsM6550NA2CAvambLqhwnoSZssPt08IgxGUSKeDKXQ3jj9v5nX7WMzRjSBUytsM
t3Yf3qNFhWWbLI9K5wK9hBHcVUm1OjVau5YcDLWIa8wS0Ik+exv47+1kWJ/D2NlH+aCpJssIHyyJ
gY4QSiT3pj2pIsZsKs89fVCpZyzSdHZ5Qo8oV5kfG1vGc+bCaLGjzXIQTmEPdJHmthIBIXzwyB5g
AllKv13sejf7BFmmJ0GC+O7jXKesqEoCPMb+4qGFnTYnJs08Xti5HV80Nbwf++3YTyjR1OFWg5x5
5neVYS5xMP28OF3tZsiplhxRe2KR74R9ThCzXNkAs8TYyFeunLVslK3X3maaAaiJYKlW8BxYpzmd
K7tCWVP1np1TCAOQxF92G3E+WTEx9fYFne7/o/GH56ZqLjX89BaqoVG5Fe9kxIBc8ASF/WtCZBZb
9lPwx1ErZKJJqjGBYo3NHPJR98yw9qRhJg2O97lDdw7RFjbPOnS9kqq2OsMiizgFIZX532Qgwan/
1U4WJgYc1/c9US+cB9YVTBE6mLxCRUXwCIy+yiBJ0DkeqsU2orhXga2biDNyL7+R0G3boQh7uaI1
2lMmAfo/NNrXCox0WfyI9yOZelkke4P0L+0Jhh3O18B9e+bx6ccHyfF9KZghYoSHS5U8/gHOleXn
+wgwtSxRpVETU+7PTFHkknGxr34fBvXi/cYHJWkJAudmBiAlP+F1pSGzMBcod7X1tVsuWNedqfoY
EFkeuWKSqAaz/YURmFIlSKd80GmIO/Wcf6CShxjmBqhc2nnNjVvQzbgSAumdLqgl4iXbUtEB3xzN
SSuDT5uHgM02m0oFGjxvSp3GyzXnyJ8RSZQgsOEnLryG1VEmhy7Ex3PowWpmgq3rwg7nqfo8qkPY
MfX9tM6WETgPhD1rcQ6tTkd5cQq5iEEDBPdDWnk0c4lWpvll+7kpyP5Tig18tzfbPfKBA5mhwNs5
Lz0ciyXtTkYjA87dGpTwydsCJzpRv5K23eualBpxr1/il7uTt2wHE0JSVT+y+JRBU6Ya1ejMn6u5
1Xw6JlJwuUdXWWvCn6LpegFhHipjqmjWbMtB/fTmhXu5QqzhMh+OHZL/sm4/9lsntSrKMJRZHUv6
godfpxrIMSKdulN2QjJtnveGUnTXmKNLGJk1GtqpPACqgcw9A7/IsqJrQcltkDx3bU7r3tl8D2MV
S6wyc5RSnH87C6hENb2BZz5OZ2ImGiQGxK3TlpFw7q93w6y6ZHp+X8tx7ZszvIrsDRoCQSQywSBx
ANVQH59+iRx3M06D+nC1uuasHb8QCbvTqimYjXzFx1YBDbDXOSO41VBCMj7SHaTQjG83u2ljQ3/a
aq2W0EdN3d4NCHmM019YINltQUlNFwZVHCw90LXS60TvDa5PxxzeCAnlQrcvOyf8RAJXIis+nSZc
G7rT2jn0R4hV3z/vFZBOGIuDhkQ/Y3nm4G8JxU+W0owHhR8BjxvI+s+hGiRJXI7bKtp0+Bdef9aC
CoB8UdqIia4EPPyYffbszhV1oVSL6/wIi+GHi9DyNr/bh6IlU6KJCh+zRpmxbhFx2KtRs24iNZkX
GU98+H3fkw7Gas/JsgH6xqxoEgOdfBrhxX7TR5IB5VnPy7NAf7qKXGd/arhdENlbo+zzAMrpgPUz
c7aQYMlIRQS/Qy1hCUyuq5mdg9/GQT7xshhlrR2cNyDkuinBySl4Q4dJW9fpj/s/c2IPq+HyXHvO
el/aOPlXRZcjuZTePAB3Uuz1qSKJ732X/w8OsKGKdORgSzvUUKKkmnWpZSASki5Qiibcz1avKcCv
65/nwT+3W4wM/KRaWZlqDEDk+xDoo7UZDlekj+hqO0YqDSLCaad28yAmBMZ2YE4aqnIRvh5hgd7B
0I5UBAV8NJPvvTZRszj1ox6zNBb/bL6eimoWROld4sdBqRpoKAl3DIeoNrzJVjDKVNg9sTxVHHxc
i3ieZyb2KmQl9osxdFDx9EDAkg/ZRcAv5Fg6OqcSF5wR9k5uTLTVbMch+Yw2knhXRdNEti5/rhMz
f1KFjTUSNXY7BhpicRyk1+T1lCu8e8Vi5f4PnsqxRRGOZJ1N2lQd4JwzoCvmwU1eQHqkapHD6fvY
dnaCyNyC11OG6JYP7hJFAkjiY1otqyFi0VA5YKae1KGIAsCRLd9oSDSeDANvp0cwGLLE5rcxOPa1
dlEYKQ/XbgVbV/GMnMyiEf7Vsbn6d/4j3qU20uUTEiaPq1eZbCeKGW4YqdcbqWihmo0WeL/l04q3
kwJjqyHBsEr8ULzX0eTcqp+UX3agFS407WAC/glPs8Az70vDqgfhfJhkmgqBLdtwsOO5gUS94Hoc
LVMyE8HSUBIfGNc59TKrtBTXx55+z+skMmMVMpccWUx5DTVGRKhlmrTXDHg3SUs/m1Sowh2CyL3E
1TiSeu4b2tdSQmiPVqD+gBDUks/ERblrFKYp2N3+PaVrRqVyolGM523S2bePQMc4VpPaaEctfKPs
zsHDKZxr4Vv2lPYg9MMPRlm+Ul3VL0W8Bogdo3v+WIfQwyZdPhtNGLOUPzL8439uof7BXujqZC0k
bxXX+2NzT0+E/OtDIcPPR64daALcdtbrcKTFmnJIW2w/bF0EUQBJGVJw99kBcZ1zj+oITXGk5KhA
pdsRRQmgSk1hqiqX7I4rEEPHdFi3PirzXSqtemdQDWvvBH0DVstIWUc47xqE6lcpKA3RKSpvevYN
bmeDHCL0Uh+M8DzBAyZcWl1HH6xF343tIn98Vo8fk612Z32PKGmkFkG+VIClSVVtq8XItqVdCejC
s64ZFFT9/eIclW3aj05xiYPdKZb5MSvuaeAA7gXQMptWr0k19Ny/AweJFibqf/4LQHGvB6JCE92a
EcJ4bfKWzQm0xazhIuxjMLV6aURh3OKaWFomHUYofwKJ7Zyiq1Q6eFtrPtov+VFEI2QAKY0nT6FZ
GgsGYnDnlE57v/KsPI+4/bIOhOm91wlGgBePe6xSzHUTUUA9mVIdL5SA7877GVfloTiSPdIVWZUz
tvBu0g8zLSbF1PMyavL0m4one1oKG8FP2EtzDWZL7IqLb4C2fp9E9unLVJ/aqSsCw7iDXTs7SjAt
luT20WxSoNt1L3Fz1neh7eD95cwqLzoF9sJZYOgS4xFgJ8qs5mQLgSk8agm9vCZgQQDcHgHuiOV6
tn6UPJ55QjwLPkvOvTdwMZkgUb77tmXXOVFSYPo+Xu0y/+eK5vgNvBUuA5dDsZa6YGOlA6p+5iMV
GQNFu79Ut1RfuH6rs0gFEdMf/UdJVE5s8hBYlbwXr8dWHBBn62SHgeeKAluyzrHxzU0PhoDMdWYa
GQdzWK1CbSpA4WfIW3uWIGI1WEeLtaxOYeNvFax1SMXWvvR3cJ1lgveankuGHYsUzlYd+TOmM3bU
JS31ykNhIcEo+rtYMHiwnU5fIjp77D5Ww1eBln6NCsGnTFLU4akUYXvD2Ysg+Vc/9Z2riQ7Ei86J
6ZKa3xNHMFuPRPcDv8FqZIylG6i1gLHlIZCwrwqTxUNFE8/6TXZ28/6rw2QCqrdB8c5/rmdHCfV7
9GYAEFaBIKwWXZvO6gQn+d30BBHIO6f2ZJXoSMQmM+8Pd9HZhuPceHoIQDZLaIIXzFtAMnCfjK03
8ZVSX6VhHi4CWlwWU5z8XGj4exeFjXh0N4RWrkRChhI81sIHiQJy6zIma0rj8x4RZZ1VF7Gp58el
Szs6I7OThkCwid5+v5siQgZf7XWiDHwAo7GjFaafUtFkeAidhgJyHPsdEFtalOp2PkMT0HeDcYe8
ZnyU92Ogiyg7e+c6eeiiXgECHs1mHvkV2lVI4YvOfEztl90per1BQ22Oy13AhQtQ4Q10MyC43jzG
yGWu5legCCdo22jcvHpOM9A01aLZ0aVeGWSo6BVnfGwY9roiwQXuUXLthKCcdmX7WhE4bzq8YT+R
VXkvIOfh0nDIiJse1nmGIc9RUiguUCe+7Ihc77oSguz/AI2739m+BQfRyD3olS/2kX4hwd2QaJ0a
XwxwcTRxcqq7/um6MTbO67aPQYz1ZNuIzqw6Zo5V8lssWM+4LoC1vDo9ssLTWBZi7busPkOQomuw
YuBFIlhv8IGet2AzmCRSAExcLvh2izA6IiXKd50ThZyBeo2nnX/uA4QcMlumTjbprd/A4Gue77EW
GGHIR3d+oFsQMX0NLXJa6A096NBfkyNqc2x6PSg46sXoE4IamPh0rU1bvmCGagsm0VNwhBEHcS6p
hf2aGp+ceTYExp4G/37Mw6RBngA3T6rR41d1eJsSZftoVZEN6R+aTXKyHd2TlloDIRj55Rk22nn7
S00WmK3JDSQL8pQxMn4j5lP0j8bdeVfrhutG2kYTLsj6fUiCoTOwL8WdANuqW6bWm3TqW2y86ScI
LLN/FjiSj8j8Fi/Qkg7k5KDUSWpJanw/f1uDG3U6GjHQ6Wyn//5bI2CACZHplF/dC1EKgcxD10mG
VkQKFRFlO7pr7CHRJ6itzjAbUVY/1yUgFpmKiqvrf4OfJo/yF3NMr6pYlyNZoBMhExxe3CN+Sv5Z
TFQQf9pEYcavzZHIAAjsTjWX/EvUJaCHBRigDP17mKxGODf267sAlHF0AvL4fjIRgWlFWpRHCJGa
ntQPoabmnrhJ/c0Nm8n38KuzogHSH1hyVANAm+RtNFj23K+ymVWFl+vFunoMUsJGrwCbniOyuY4R
GfuT0/9Ub6CNX7JvhyZ9jDMboTN2hTXlBBiVsECgQo3ZITU466P6xokEwOnddPzMhbcPDoPze0sY
KPr0dUwF+87ku7/0puTxVFJxyuyXSpl1/UGUjT0I1DxQQuTe4yvuS3qDQmlryiYbD3T/oVZAhmQL
a4Uvzn5fzju91j8ZYfyRPdnOuTJ+KffjV5wRQrVJ50J64M+PHy/4fJeImJS82Sa2+vEPi46LgtK4
D3BCUXRscGVEFPnymPf2iMk9FYLCQOOUdI0Sx2HdTiH844NAdHzykQz13RYda49+dhULb6vRBr97
EbMcrKbZ7g9Rfxx9rcnK/++acdzsHFk8hwyfrCpk3zSu9qd2mSOXNG5MCPNM6dr9YoWPJvYMDD5M
B7XAMS7JqUjqACsKKn6JImyWu5PHTGO7Lvx0j3A22txEwX93zmHzqCW2+69x9No93SJcTuAptvHG
F9J4NFVAAlRtusC3EiT3a5VdCAEG3wjQwclZv7RDn5TfzUpgzNV8bHsgJUQBq5cGLMZ1RNKDPXRN
XuB8KL6B3Gn2LJm9SM2My8AUSj6tIcOGkMoNFlmXA8qxPTGuXW8GymFej2FBN702goCMx93jKXer
PhIv0Irq9i8v91T0GfH8Ua4Sqc54cCKg1gBLChEw/iqrLzZtOxYIl4n2Xi4EqydgF1kNf1Akt6KJ
T+1/hcMu/gNroZSedAwxlIsQcZGLqtDT4bsU4EKxspJj6VBs6V3foRjPH+f/njzZdHkRrb4c7dCA
VMqb6KyvQqgUDHx7D1YFnXtLUdKvPeB3kqRghs7W5pUJnLEdggS3W7RDZDE6eQV3Ur6KxCWubZf2
PyTumAv1+0jaBGeZiB0iljpbznI36s5HtG03yk8gdYNYOi4foXO9IZJPqyDElOwO5GzbNfic6VY8
KwSBBdt9pLTR9XmBuh5ZpFXOIaG8pZCTs1cLa5dER5hvL5C3MAZGpRJDc9u2GpDp0+issxTPzzlD
PuA+lyWYyS9KQvRKjB8VBrgrOZ2I3RtMy19e+zRiY5upUwvFeYjj//lH5ahlF+yCNhUjS1XuqPhO
NXYGICtJZ3ktK5IDNZzjHC4PTRUPoQeG1yMhfE1wvjwtaD87BDj/SBvyW2PsHc0Wd9shv2pRThlH
ehB6g6o4BrjQYc/tMjIs4xuaBR+0IjiN5naYgLUbFOJDyQpeoeF8OyAITAsfJsz+3pWpVlQjyA2u
C5U1Yp7vxS1DydAxr5bUMGG2JzgIFlNIemjirnWRXELxg1v2XOJksWgZBEOCMW6werEG/LrtlUqu
8oPjxSBFGDTe4j9kgeKBtizC2ojkgAXldRV9z/LIa3PmyATCJSWPZp2smEE4DRP163kbmYVv1HAG
/WkD3C8NK4zupA3B0X5SNQDuDBUX2EJRNixsy3EA0peZmV+udNUux3bFMjqGmbmoN1zbwGqCdbqZ
ILGTYpju3+x/eXk3T1f85OV+qYR1rjPkaSlABkyPd++FxQERJ8DG4xdGsHvgWrI1NGKFgTQqtUoS
r9T90tPV458y3cePSeF4Mx1tc4WhEaIX6toTp3Iid44cdgIkU9d8eED/to45VK5tXa3egxsQ8vtc
28nYLXYc0OWN6/Htsb9NUDWH51/nBnlA0LANv7md3kGHKUIkRgRHZsz2VeApP7kRpei/tFd6VLqn
pGc+gyb++iRHoe0siCbhXdHU5LZUHfFvEzz/isbMmowSqX6Sd/AHrB23dioWRpFjxDAE/r6llcd8
FDgnJFHAMcd79brWMhR1rZ/s2xt8KMMUK/ftYECWEa08GjwSIWWxtJiQ98O/nLaIOFT+JYxr1Sxn
IF8uTMdbbzCBmrOYIU/dm33JJGSEnSixEWIJgtDBp+VZVQ6Rdy57Zz9NCbZPLyB31rfp1s7V0VdG
aTGAXhaj9yqvCeEQeoai7ROQTt17JbVjCKbZB8woIdMQ+D3sUKI9V1FUSVbRBysYeGrtqSL8M/EA
SidmY/edtigpfFKT6tzDiQHKrgxxZ20aVXEKzwma90AvftqptfoltYtKGCVcNZFADpUj9zkPdOqW
grocZIgaW8dCMy0vci80PD5dqk08AHX17S+VZPbHK8VZMEgNODJAVjR0IAP08JjIbc8mr6KWgsym
7kIYXdkt6rCxA8+QSayZ7P1kqOhqc39iKlV1Klvto4mPqMXcAEfpr1SoC8wX900mZhHyZ126Z3fC
VeAGHBrcPthO79YXUu0c/FtMDlo1Ao6+4s9+QBr8vF1T5MZvrFLDC8BdKyNll9P2SaKBECrhlkGo
ycSkJi7f+ylL9U5i5wyq5BnzsxLy6KH4UwsD1qLzCfIGnpDskiUQnj3gczMMy932CII7VnenB4zn
L/HGSxc0EJsOSoX1WalQ52y3lP8HHN/n9pTL4pvnjb7iheq6Q5YcH5cHaPItcsIguF4ECAS7sEGU
ZNGmM+6Zd2R68SWm8IYNUM94WElVXS2z0+/pw8Li5024aguSi74fYoNd4Agf1UCpZvpGElJYTbB+
YbLa4ySmxREMJ3BpRowmgDqpMhTFs1zuz/7xu9NizhySOx8qx/oPoNmy77WAT++cImZXnvBHymLS
h+MlntaMmaLuo2OK/4a7WyprOCgVOCwvysd+OgwYMDzKKi225691NIQqkxhXjipnXhStgJ6aIH3J
vRDclzpA9OQK/si6bPGyX/A4jJJqFzcShKZnxXRlgdakIATDnrnzYgQQJuMVkzLSoDbcXO9lOBIC
NjIecN8IxDrY3ZOYt5C5i1Q7VoV30CvLC5s0CBRUSpqBmThnKet+8YzHVpxeqrsKw+LojESVBhel
mwwKg7UV5LxZSqFCzRJNokCKzVI07iAJkm+JmofpdCVyg9VHW7s+FZv/qgrBSi1qkCfri7KxtTmQ
2V6Qohs4r50y9xW+NHpOo5qb3G7uTxw8zWdWixf0O+75jLoG9cNd1S6rlk0QihXzVIkjcr1CSXT5
gmXv5UyCIbgmxYaEVGJfZLTuQphpyz5E0dH0qi/tD+ZGTxSOTynG7L+QXyBvUxIJFuaRZnCkh4sS
P5xX1j2IQXaKRCfxw6IVIQ3CsidTqlWaOvQkFctT+7E6Ygj+HDL4BkGo+tWDULnHnYdoprabA3qv
asf2sW66YCRFVMjpL6YHqUGA7Q71jQRqZyW8uPi32V7CZuwISzTz+K0FVlTWAJLCOFfYrfl20tUr
U0A+2DvM0faeNqNRJtilZWYosvl1UmdZHiTJ3FONZmfuEV0BlW9/KCF6tlgFtOFqFQvdCf8m/z9B
3ohQEGd561b8xAlHDo1hF2VHrIm/5IV15QaM7lyPW84xGX1NJKZ4krpEiXGoaCrQ8YegwzIXTbrz
Sdo0cblJk5z4SrIEqrduJH/Xj00fvoLRAc6bt58RRAq6cJjIvGIXsY3AnJRS4kCC55MH2dx/b9YV
p1y2fA1le1pg5P+jIxs9xY88XSU/xEMrsVxLX+ozScGNYL4UIOS7iDxtKRiUWaPagWiWQHh0Vmvv
H9U2+htdm9yK3p1T+YB69Ks3+0ayr1phY4SB5rzVCkvxzlRRBVcBWBCDVLX/D1Z5xO2H2MMsdTBQ
sUjUtW0O/RlSl6j38KokMIqE0mGw3WxC2pYlvQdX0t2wkWJNjhIOpO1yHY4AtJUGC8BSL+63+P4D
+2Aq5c4Jed6uO/gnandlgcpDB72ZMEg1qPnAD4gTXmNVhORecw3XYG7ekT81ir8LdzEpCu+rHPus
9PXbSr3uLU/X3fKIF/VBTaTN/vhrrwFXuAUlQ2sXK8FVbbiuj6DsdFYsIZwBfaENsf7D734oVelk
bihcML6/iYVaUMq3FmTE17V+wo045wEC4XSslWuE6NbYevRa/C3SUtyjUeKm/1ER4Yf3uUSzEFQP
9A7z39WDYwAEE934j2LUYy5GOAsn+oeuA0SrYdc+GJ/IQpoM72xv3H6rOa91pAEbr6JznhfwM/+q
VKLWiJ8QZe9OYKU2yLubdTq/aOYVnV3EQM0kYyHWYogpMQNsE0Q/UUpCZvfVnOU29SaBrB0YcFcd
ygKDCmyt9P8DHDd/kOLwe7pYY0UFFdZ0ZRF8jbp4YhsApK12oYNNjx1aTU9W/BPIPPewadmE2v21
O/T/XfL7Lqy1J3NZ6Vt6iUY6D8EgqOC+B8s4Ry7Sj9jmGH2mtUDm810eawIKlewIErbzNF25W147
OeFPbpJr/EP6QpBohtDxF5d88cOzM/LZmFkdFlYtl2GVJ8CwJ50LuQ8xI27+vtpXuU5AZe2x+9/+
wpezpNhxZvo/ulExar4m1Cx+Puu4meSoibu3FYUOg8Vs6vZ4AftlFovAxQlVdSsSd188QWh1SDkt
K1zm0DKGZ+S572MByhJtcRa4goLsAbaTBWfXTCY2MW897vMP9PCvBtICDZnZiivETNnCOr/O3MjS
a/UalxRvCmgOZDFXt0vZA5UxXpFuADqfAd7Id8DX6cHWSvVKhDgAi01iCSa7kRrWqZfelP6u3L2s
xDUxUMva8/DYgzSNRFHwx9YNmHapI/618fYQ7Eci2l46tn7hFBxDtDuCZNRMH5clKXbo1ZwjBK2g
6m+F23Lytry5DoegsLclq6jk4JQ/fveIySaSBW/C143P0dnDaxu757Nht+JoiCa/rzB+dscpxwIK
5iXIyU/EM3JOkRT+/PwTw7/f1dGnVTsfX6TgDbzeUL5HdgjQvgo00zaYjC651+10pIRhFHZhAVW4
6bfHgVa2mn9KYpO9fteskAru277kNzlXMpZAgvLpq6rJSHplYt+m3gTi+M5PpEo4ncWZOYyiWRdF
ByH5PepNl8uiaRtMkzBtxrpeE/T28+2iJndroT3hIIYsqT/ym8Dmp1xKQLmSQf7K3YoFQ7o6hSNX
tvpqSpaiJyQsx0vz3JOHycnIGPk/KqJ+Nt3Uo8zEwNzzgTdU+fQ5lwmDd1fclZ2gACKXjKyprFXq
LCtreAx2whF9/XNS0+HzsbR+3J31Yr1ukkFVrzn9roF2gucbjPoWjaV+Qsa0dHDtQPzFVQh278Q1
1FVUHNTmE/6e8TbRBQIOwaonCI0+nrN68zMmRJXuK3i7NYF1Vvii1QGOVERwAIEuqN5xmKUJ0d0i
zg3MisB7VJwwdWt2faujL4Za6rizPdTF0WSPY2uBJtol87BSuAY91OXFPl2Y0Mdg1TQ0bNKxuPsN
vSe9ZYSHO0RkC25WFEhM7yr0eUwOZCwKteWMhGBjn0KE3fqsERb6Ye+8FbDktZ7ik3MDjsto7S8P
gDbDVJnhPsU+pooZDOE9Uo0g3kaRYyIcgkynk1L6XY7uxR6s9lPrAsrt8SpKNLJ4VI5FVbxn+9F/
8O+Sbgm+brP1THl/TIL5i7JJyd5LAO7xg03tFQjUc/2RUWM1z5cQbpquUkkGXdV4Rvb0APdiICUC
4Cj5zJ5pevIfbdVs0vc1iCBWsj7lyw/TVgGwhdvM1SPp3oK1VlJ0zXEHNZwkqtxsNalP14ygM1oA
2jT33slH93GXqEeYSqITS9EnNfVFwGJfGFq/973ABACRgpNkkHoRXlPi8uTSwybjlFjudmczyr1z
MKOn4N92KffOC5tJhn6HvokxHunyEIoxEgNpQh3q3N4864o00VA9W+tJPp27qrAjSCFTaK4Gg9az
NEY/Dw6ITG1i/9sGUG2AIXUW2Z0QMXkoPIPL3KSt5dnWcCERkq7wKm5KYdFVz1LqWKOh4DDLENcD
DNotRDrIaSmZGN2NjEAmgycsVvA+2QoK5s9Omen4qDDAXVwlHNzKVP/apg/GnX1ODr4t6rgjtP9D
gztFLMbcPPk3PXK3r6QmUgJpB06u4kA8LElLIhuV6qK4t4ZH71BK//gfc8dPwfvDJ6tBe7b5VsaD
yK33lMEgcSmMJhwJnO8Zv+guSqYZzPQ58hbSEOqGbklQ6eZqgybMcsUxceecXsWUgZfagczXnoO6
BCMLovOpZ6EL9/xJI/anlobOlFU/l/cPPqVNlFpOh6K8KSyjJTjTgHEhByt6ZaHXIPsPnjlU+Ax8
VHx7vb/46BA0sj15HlPe45eNvjDpGBz16M9AGL6KJD9db/3q14fn5ZkF9akOhGp9kIx6tWHig0l1
TQTzISxerpbSZ9Hy1Cm6IUxMC97B3T/24zngzBq3Vy71AeiOISqFcUQABbiQ8kBhXCPD6kr+ZXse
8YjRpE/OoJsFc6OX+YGM81666SEm2HWiHcvl7l4amJ9JlUMXrCHdOU454P4N3/iwvrOABF+vfAMW
DKZIoXWlCEJ5l5nXrgMOonHBJNOjL4+0t09pjBn0ql+Xzbk18JpEjJF2JS6KkSWsQCrgMIL+llrA
yOWq8Sa5hxuzjx4gGJ+/bQ+ka2Oe6X/OPpTC7S0i9kJq7GxzIlsAfOjBClXqvEgt8bfJJRGZoAbb
uf2WyoYqHTr5IfV3HQ8vLmdoRv6vtiHBkdlAYUZIZK7VC7RLLwLLD/dc8jU9EzYsGwX6g6A6QaM9
nH39onsOQTaPltQnWrAgNJadxAE4w0obFIEwO5ZR1R13JSznrzgLjaM4AZihmyPE4NpnAt1Rclcz
IFtBqjKduUFcveoJZb4BLwZuTuEP0JC0UWxVtQaLLi/cf35LmxG1pv20hgOWEGvHLUFY+PRDW1jq
EAR8C6l+y1fjYnxqddJtcpJV/s0SF6Mz44rSvjjufiqNsifHfHWXduLNHCS261lLzDgM7wmrHhVy
Jy4k7hnxjpFHr7N5uclCBKU9o7nQtmfm8IHjkGsGHPEk5qc301FhdhybFjwCbzbNLpmfyWOrhU/a
XgmWztTYu/Ut/C6pQ3GWgBAd5CdAzNCfLmfYUOFZHB3L4YIXZUsdVv7V3oeITgW4+HGuuDrHtplb
r/ZraeUNgfQRxXwj+NgrJOrP0LioBjQD8q6W3WzEtI6Yf5QIGCgalkGKlm0gx7RCdkrVHS6ro+LP
vJ98UN8lPHHWuse3sx0SgGXIfJ1PNfLwZeOMgSFqLEVUkajAFwKFQCujUpZxU/zXG1Ao8QWO4Ns6
pZK4vPN+6gZIiPyiue6arJnSWK2qQUUIBEwgspP2b4KAU4WVvFklp/LSAUiq0U9j7TJpLVqTsKr6
ZQKtd3M9pmFH3s4fzycfxvEkZctlq/xDLsdU+bSVZZX8TddTdwQB8yhsAutvHum+3ppH0fYPuyZH
ahEpWFD8o4jCDveOlcA2zAc6tSWd9KOaWSO7WHlZmB/fe2O1q1Gnpxy2NHvT2/R7VKPdSTeANRLY
VF5aCf5LaIjqCjytRsb2XbWL/YEu/QQucdufq9FmS0nCXTJ9pSI5pbugldhWhwn9GfW2rRBwEQL6
rS5c1GTkCUmKpLjGJvgYrFB1Yd1lpYpPklxuZ75jpNxp+g4zC2Wms0cfWIMY9ab47WE14ZjFsZfy
aq9t+PHR8B0mxwYvzl94nnqH1l9xNY7NW9S5AtAZ+SiwCjfiTEzIfL42bVjv7didIlHph5/EoneO
8ZM7uhY0NBAVgGJKXez64XSN/lTy5ZzCEBjnNfx1sK3/pu+f+KQaGTAiTFXayQgFAzljB0LuZeIl
npK8QLn6b5GBDASQvmvCopEkB9Z5VvQq9jEysjmrGbn427WY+PVdffSR0zzZCtwIcAj+AWKee29s
ww7VBVztZFEtoMOL13L1BcD1c12UubLuFvooM/lKeeUuoYvAmg45uWpcZ2k8tYpSodePmG/VIaId
gNGJLE71aldfy/KnV42NtXqYD5epKqgqlRefx719Axsf/2QUAIjbeEBdAgR9UaEa3Py0EXSlIyHW
0zZ5h04ovmT0KshehciA6mjomMIrSGeNXSIPkrMs6XghVDq/Z1DqVYnBeiBtpvYCjnVkJ57QY7GK
/Ibf0cxfb4xldEVt1g2Pl6953u6RAxu3Xtt14CTNE20cOS7QiURM8MxEI2zG6ffkxE9rS97XIiFZ
tHsgOEUR1Al7rfCDlkhNAWsv27ArlUJjbqx20pfrtOto57JbMaslvTZrUwaUQkXpvZzn1CZON7Af
OceVJPd0GxSn8w4FyweCaAwrYTCGBI17gT44C7eLmXxzb7Njmi1E06jIFw4VwZ10hu9hXWTvizRX
EKYu7v/8EFhpRXme6N3Dlv/WxR58R8yeECIv9kByqmmV091Y7PTDkF2l8VSAvltoMeyIYQihI82H
DdgrfvyQLLWK2nwJtBs+qkji9N2n0fvsW6TpU5ab+qcFtUr82svVxfIh5Jm8yL6c8YRu8VuQPI/E
NqJmK3tCgPf1gc/bEmiGPYyCpSUFrzwWReVlFi01oQSDJG7XfckVgOAJjSKBtGoUJ79JpsciR7pQ
MJarzg4VtXwMFmga1Boe1lWcEhycBCwbkEIiKQ6Ij6pSpTuRC9B1cK/DZ9BqZ7PKyO4pfvT5eapy
qHGO2xfP5xv8AEc5b3pzOKhh02NkijD2j6xY5cDZDMkzdilx6eHSsC7Ah+lHRxcIVwrOiqppjRU+
/OAMEAXLJJ6qoTXGQNYXRx024GwwP4o+Jd3djmQnqH7iQizZwfomH55rUKqCFgsgLO10gIwPBU8S
94fv4epwGwZS5UKrqNVbUifVYqRbwZcwBiXvuzsySwaeU26J5yJ3cCjeR5xRoyCDpfF/Bx/ilaO+
F6PgzDywIwdZPq+pJifHMbWml/Rox7i1C3YEvuoeLPwLCJEe5OTmvfW7rVJBSxxLxZwuvGsSclwF
H1xFuOeZYC2+oa1ovd8kqyjuTiGaKx6MIbvz0u5pqEWkAMWOesfgzFOV+xCbNNBZX8pYMs3DazjF
tNJyEbS3x0BRfeZKa9f6ZNLpwvT6E5sSa/RkNKx5HN8nZCRibtqFPi/39bImjx4thJEpv3cWoYgH
YbJaQlzDqLKQiyjmW5AkncH3RgkJmGhX5Eo/2PYqFtOInrtm5uexbHo2gTLVgb5euQw7RhzTO+oo
selpKET39DsOsSRGetGMz85Lc1gnSPv2CTwdNToc12IBuOOmePk+yeZJzyCO61l+XOa/RLKco2ve
7lPI4mR/z4iiz2kbPBgeZOQ7KptJG54vlnok8FJDEU/hWTXuAdvolb/k9u0ziRMXRH+PSofqznbi
l9urkTyq64821km0K6zmhXjhZvEa6OuZYF1gYzimfcXRZIkgfJZpeGvs9F//kwfJ24n/Z72efW6u
pabx8Re2OczqT2G6NX6jUhzX8MuZ1Y7qNsRNNPRpiE7hi/sFohcP7ZwlyVGWnviVUJYcEZB8/8Cg
6n1g/4ZMONIg1ysiCOW0lgtPT3PSNjsgVpZ15sc2P7ZNlsVy7Tc3cuncbMWDPYjSpK53jEeO39fS
vl36CiSHmQQOnDQ117bzO/6bbQBJwarhDTZXNE5bATNZtloB+EvX9LLOwdohGBhBJIpCYOfR447r
GVgsJrXXqEiFrp++3eNwTEjIBAKcdjLLVgrfEmZFDNnbYCX4Y55Dc0uwN/OTbgqOYHOVpML8KDN8
PN3U4/4AU1mM6ZyXDIZlDX/cIILRs2CcjfjA1tE7s9n7tCHWvjrJYtiIouGgdkfbDHdOnYo0QeRi
+U88H+eTQW2lA9Cgp1QZv0ZrXl0Mx+J0HcH8HOkVtkDua0eQq/8itITOmtupuWbmNDljWDoptT1a
ycnUZ4OVjovosFSEUD7OTV1bik+xchDEq+PVdSSvF9ZKM8FyvC/5OZEKvTjtD7U+kcUe+lgH46Nu
bvGnXXUZquXsxSomHgTsNnyPWIVMDQMFshSLAJEwRpcuoknksyatAsyOHfwk/lSgHHEV9UH5UP5L
UzaipC+YOpEo3vyzGJ5n7hnG6XF11f28j0KZNJPqlJDhnR1eHGGP7Nv3bDzjW7Yeo51uc4Hoe5W5
oQ9hkSAmoGUHvpcdrVNQKD/eAuRJc9IBdf4EaJGPBj8Vbinus4QEcWqB1oScdFxYxrRgafrtgA10
W43CEtZiYlU82KSqqjQKApFRCxanAXWnfG8j4RTTexJlljdMeMPFkAehdex4HW+oaKEHoTSbBcFP
/IJatdgKaViIEWBg2UJiKMy0UL+3HHRcCZSoUt/5exy4EBa1JU39gN4PdOJMkGoCA1RXun46KCYH
kY2rOBaIDx/9O/PBc18rHAljY61UsJnfsNdEbcbsBKYGQXxhotthpJyJ8Ev7QXlrQnVausVSblzE
rk5liLdkQ8K1G6bVex9Iy3No9stAuTs8QLVvJdNQexC1CuawxJZdWsxam3x/E1ak3jXPq+zWqIjh
sG+JxtOLAW7p+NIrbErBDpJIdIbhMa7yT6I+yhMY8iTRPSMEd+Xil4PBu+XcjSYfrMYLsS7vnmjj
oMDGZXXhS2fm0bpnQTZzZVLNzzNo3jqzzF+TBJPneJafNMn+ahfb5exeVHA5NHRiv+YpeLPS929f
QgOgmnwuFqB1aFG36Cp/Lx6ZG3baQU+9n7cdDpf5WaNrU+O7K7iGYC6tZmShx9GI4+RqPoe6B+Bb
/uBDGTg4gN0IEaVcL0RBZQ9rU8cWONXVeoTLCuUMJuxdIsqCXdWeMUmAiquDG8awLSfJT91KXsBS
QGyJr3Gfbar7tHMsc99vOthNkKRM0rPA58Nl9QxTD1HzpkKGa3rTw3HWl9TQxUDWNF0BXtPJLv+V
5JCdCPyZGK2Sp2c6Jbzj31aZdwjFZbpYVcYXMH1fDKJb4EIYHNUG7gJ45JTwWX+s63ByNnoveLPz
xzd1BuatTWNc9STDLD9fWztiW8Ocb/AyN/UiFlOxprr9WjH0uPmNd0BveQcOf1RLeNjWArYRRs/v
wJK7aGRKmZQgxLTBhZwHktGZCbDoKZnEa/RFSTf9Qcjjxb8sYPUycis8saqaygVydbiiv13tb9Wy
7iN4/9WSjEyXHWPpLYvcok6LcK8FkO9v6LsRugOZaGyW+AxptwSKGXTekWhIyLFFVSYFkdQOkYFv
Z4vEFrIhfGCjj0n4NWxDghaaeE/i58RJmdTjFfxaVli+sEAWh/LG9tVlnxlhtGxho8YTSjaWdSDK
XMzlkOvxcor6m9lWgJHTbGQIxCSkdFDVo1J9viVxMVdj5oaaYTdwEXAFf2qFd1j2Cri66YmCXbmb
GisYFSApIBg5GFRLbyYgIcRC6AyRyFf1ISXvGtdsbgW7oQsy5rMHcTP51tdmD6jy0Nz66WSIeSeX
NgS8QXtDnVUIUxgSPh1Y/ogGxN1Njp7ip4t/xSAztCi++DvILH5sTYwikh37BQerYmMU9F4Gphqz
owEYcTHa5Srr/MF9+BNSN+ujqIQp/gBOdGylqKyRpNZiU0xktfMkHNxhyEmHK5qcnVHJfU7xsTbu
yLREScI1AoEE3kAeXPjvbw/9oTyWObmmQskDnmiluZrT67w6JAUJEnFpudgSYXDoQi9pl+VtZYPL
7kD6vg+Pre2EXvGDuv3YaeWK5qrJjuK76OUivnhQ+Mve9hA4Q3Bt7a6JviNQQuXo3VsKCFqHAYnX
g8CSW6Fv2kebvdzdr2MskbYqzPY7Nrk2PPCSt0aq+6z2fxwkUAOY+1BlwMcwVm/71hjw1nsc3a+b
G4ADlqOkfS0wYuSj/gmVEpxxxR4JRk9j/dRQLn0cVSGh3WANShmNvaZtk0bI+ddkeILgzVycY2CD
iiCZNWrOL/rBuOsChBwcab2zsv113N2v4mNbc2aVYL1WgLlPNtYmD2ubGsL0ciQv+SZICTzS7l4A
sIABbUqYOBM8q9G5/PubMkDWwDYeQCv72wlNOHDH0yJd8zJiRl1FpJXOVwjHdZ4F06eSgq5Sc8HF
ZMJRpf5zS+ZimhydvVPGfPA7XvdzcT4y3frspOlwWUBRdvRniCZYvifGIYp/Ahr3trsx/7/WM23e
8uLqBs7he9GpDSlChTt2xghQieut+Q1C7f2wEhNjcz7NETVbfJWoZXCiWggzQ0v5Rmk9djEcc/J8
ZLInNPa2568DgsAFyfz9Klj4HigarSLPYEWyHZHfbvh+zZiXq1FaoV/NnjI5L0efL+VEjGDP+d/Y
Q7Vo1T8ziQ54aweTMFq2jgn63LWifLvrsn68LQIEbXsjBEa4JIndUb3twhr6OBaNK6uCQK4g66TP
OeDHctgSi+hVIQUeqUybjR7HPIySr9JVmvQZ969Go3yUBuNEXN2eQ7EJNhpOzOcSrWc7aGKRxZiz
oppMsyjIiBJoe7TBykPX/yuu8Ot6N/FmaRIICwH2aqH58IykuC+bvp6aN32Fm1bfToraqpVj5DiZ
eZHd1D6vrSueXRpyUIr6TwHljanhVAzSj5J/Yw13Ni3OH/RCNWd4HJ3LK8f8tNibQHUI/cfb3WJ4
E+2PfOQtKjp27vTB6TwK2zvGRV0E/AgGQVR0Txja5fOTkOBYQfvAQfTH/jsnmL7m/t6Iq0PV+wBM
mthkpgdFtxrQ6BqvnRrWOA7EifLcmmDE5/ynobUbKtdpHJOgaMc6KFhAr1IRu1um3eqsOQFMaJHu
Qm4EsX+S/qxtOAUcZ18+hUgmHIPhHORmXRyCTPZBB/7sZTyphWqu4r8lBSreb430H5N5kyEQn3tA
FjRBbPgrXoyqt0peuw0Vu4VFONxXsfH83zx8RVpSvmxTLhpkExbyfrgV0XMhH9DbWWwrqjsvyC95
8gjsBgOB9kC98n8xXEIE1lXC1+WXro6OgNLY44eqqz1UAln0BZIBncoIc4IID4iix4H/PnjQ95Ja
Nh1MypsF6lpVOVd8kDxEW5hoG4bGfyZH0q+Rgh0ZDgrKzznG8htiYuZnwnFlugMUWZoycq88nSnx
SdDUZE7kih5BzHUVqRqKD4G7HscOqhc4HnLjc3i0LREGEDiLPg3Zxk4/iPsxdYxxCwJH9mm7ksAP
FMYbMkdYwMFu8rbUaQPdRaqHhoA7XH69NZTGv3LUxXGX1V2ZgJ5kkaF1KisvAGdemXEt4rr2gJrZ
H1TozmWDXe+uOgjLGm/AUpN1T69JHeHatqkj0siogXRIraFIfX06n+mSqgI4k08vUGHTsk/IcOZl
zsmR3lmovLo4OL1giu3m6kVuUtlStxMtVRuVj6gZBUdiddP9oiwjYc3cmSR+QO7DTuI8dcd6f8CH
pNvklBGpVGI49y5eCyIQwAHKkNxpwLoILYrwiEy2+Rh2aA9vECrbI3RMBnh2laDxYKEI18tSL8A+
7Ms5N3GiR7+gJLk8J5B1xr+hlMiHsomcFGWSDStuYJ/VFj1U8DJoHP7Wlq/mvpM0A18o4cch9sS1
N0TGjh6Qeg4YY9bUtf+IMJ2ZX2H29rs3mleeuo2vp+jtOl1Akj7eEEe7eOa2jUW+4MLYDWiJBbuF
UsnhHQ03ULQcRnV9Xi8CusI/6bp8Inonosay1htPb8+eUXwHsdi95CpADXHPmtiIPWXZYqylPUED
0EPfSfptIhrtFizZ1ZbTHVvDUVUpQNj/axKTN910eYK/Q5dPRY7VZtKGnY33SGYLYjnU+/9Vcsp5
PS3PxVRmuUuu3TEVNkifDXU5k0O2jG5RVGP6WHbo2n5tRCPHAbu90BvAQd2r/APU7GYAr9OvGD/4
f32ZAQ55GQ4/GVehMnyrk9kDmwJ+jQQsTKwTmEZjl7plS3G0b9WA+YivXUgWSM4Un85kb+Pf4yvF
FWRk2b5M1phO2QUzz3U3QfmMz/YrE+IZdk5j21eTxDKoUsY7Opi22sEz0FqQDx1xYWut8V4C7f45
q6JL0NHSPCIeLnuWO3wnzxVIqs7qjlv6iEUcKBElCyGgKXo2sp2gUy16SufsDNbjr1yM8el6JvSI
m2+9DgUT2+JS8naep85vKco939RY9Mdz99g2MfKzezuHUgsHpVkKbjtbNT0yRZH/tqoIr088muIP
GiIZ5xubPj0RZiyDJUs4bYm1I1KYhWpwTvLiT7YxEha8ZU3J4Wc+j0QtwB9CwNwNRqJ7o8cExyo2
ryMg9YdW594ZP2mrAm2Qa1kXy4TuQAD6V8EaZKNFaqKdwcrLcHwev6wZUcoobX+460Ol3mMhMT3H
E+nsqFxnG/sw3IkETqUdDTF3r/IRO/koEdAZWrHemJdj+yOu/EoTQVmrcyxktQSgne3qlcWluePZ
nPE/dOHR1XdCoa1KJQVJpH5xR6h+R/21exUlPSso08sva6hThKFIkv9+iQ2K4GWeOis2cbx6dnyY
ck6LzWZkKr/UHK4gh4mAd0dP4VmT1x9E0KtGHYFsNDWosYP5Rv7y17Vivp1sNIYZA4QP2ic9PIUU
A/CXU0Rx/+vshnmLJiGRaB6iBDulb0DjIUkuBYKiOsinepbEbhZ4KIQLiC864nhV8ZCf9niBwbKW
rGm78MggO40XrrBDH+9h9qyxd+R256BMZn0QSh4FOqBoTpung+g4QNvdxQdPwaKVFcPcC40ZjqiC
tyRHa+FTacL2oFLhPyn6AFkxiHIKcO4ijbBJh0dg5+ynyRt6OdcovUlT+bq6rJ0ACCM96pbm50Ht
P8F2qUcNUqTQU5i7bdsPdbEamQ/c5kYy5Gm2hy7/CK4ppzr1fHt2E12Lgnh1Glk6bXVMnMAq3GJd
5Y/lAgaNzFZaZ8JFe4uErlXu8XOMsCRlCZCjX4rJmW5iROhDTafSl8eIp3PJ1mMW/BJ360Vkd5LW
WD0lXv3GLXO90t4KgXUPuitBcz/squ6VGT113idrOEedz6kOeAfLZ2Wr+ZUc1LJ+5qO1oA8gxeSR
j/jh8KExG+qAqAnOUi/GTCeU3vlthlqWQPAM6EGTm4tK58Sb885KcJHiX3wr2q9IDo08yB9bpxX6
TvjmyooP8/7pHNPjxOODfopL+HPZ17L3GVrju82cFj3URcGQZyzkYhGgmZiwf5MIC/ndcpu+nhQQ
iwtMXGxMs3xvg0f+PMH13VJZBETxF2hji0lEnhZMqXN9SZfUQNVk9KGNDuX9W6RU8R53mligZ84Z
JDipncZC0C+KGI8AI8QtSCP2Ra9hhz+awlCB/9Gwqvqao2XLRCkkeIH25T/OnD4Og64ZINvUMkLV
tj9Xp0MzqvJ62axTnMIn6SGMXLHSUAWyP9H064GIK8W+WcuHFCq4JKWJuSwagZ2p13/9YU747+Es
ZI9tGf2R1ydULLEKZ40GR4meMxwBnoiaLHIRAe0+m1fVc01QrY8mR0YTrbO7vFb/wfd3hg/R0zLp
/IfXQ2YUqmNbpqS3uuuz4ph6Cvt4KBvWvkhtt66Ka7KD6U8rdDV1VW1r4BhoyIpFjfvQhrDwWTSK
9h/mbNq5cutgwhAifLKaNDhuYQ4L1qJDVXqpHuoKDKE+OiKrnddY2vwh1KbL15umHbVFcfw+WVf6
RWYcPin7inHhDDJaM5WKh0Voy83wfHQnz0yGFEtQqIcM6OMao377bJLUf5HUCu/fts0jBpbrf+57
iFNmIuxydKmnt8//zJ/xNjVAATVTAnj8r09jjjKFVvQhUxL7oxPE9dJhwKQDJMlOhufAAV7UVtKp
ThILM/AVfyY7BQq6kFnrivwOk1Qu9BFnokaiADmMi2+ud6+F7i1JE9LlrEMD7IQmFWI3lz09TqWh
Aahi6AAJxEYEqguR54U8W25NroG6rX5zEp0IhsK1v3DbDvuEObc+ls3cBp53WzogZGqxDdNfA54a
K1cmPCizF1z8VhxhnKbvu8T+GUgQ9fetoSsmj/AecelQ+vmIo+JvTR0G8s1R6xuTHJmgvUKPvK7l
I8XmQ4As5nAFR7MXCQVcE9quhxH7iC1arVo8s+B3YKgmrGGB+8sBFSv3ViBhH2dV0EDTsiy9fI5s
fzfMB04WLzBpICAMXUIQiK5dh8wYtnsbmZd0yB0fr0eGDp8iFeclD5kpJznGF8yqHD52r26NyJNu
t0F0qyqnV09TZM/KIGQczjvUICBPuLASTwgZItT1VezkYikZ1FkYQIaF47yTeZiQqhS98GIUMgQW
PEkuC9bmD2AgyWC818I5btyYhf/5GPFwbwT/DlfeqCvZturwpr48zRG9gXpCXs+0U6AWwRu7EAvl
BXC352raK/4jG0cT+VtX2prlmgVloIXyarfAD4VT+Fdo/oxGBJ+M/kxSOWRQHe35Ji/YkPFVAT9w
JKoUj6JVoyVyjS0IUSbfmVCRFX2CGpxE0N2M8k+E7LJsqGoGevTy7HDhWoORQtgd2WCuDiZze+PI
m3Q2CyZUBzWsZbbYVePffmFvlUNP0gDHZSsZbrSv+/kiItN0wDhwUA3q/ope2gcTmUl4mkAR90uo
1MaxClQCvmT3INvGQQ1d6jelYtI1++2ILai1ZvVke5Sr3ZDqxi7aBWm7DhUn9/3wNRBeMv4yGn4T
ulA8sYnLh2C9xy40agt9/4CHzYkHiccUTg2m+vKzoZ9BnSTZFJt5hCduDZ+NS+vwPLs3Lvq9QAvi
iUcQ9so0CugrqPUoQAKJ2mOleeJa50uzchqStwM6duaf4YwY4ZNrD5gttnZfQxuUPrFBYv/pjtAP
hIaxViGgXucQ3EWuzyoDLunMbMZI8WHEjV603uJIst4G5KN+TUAl7suWnmqxaolVulXdDJMS4wZz
XevijC7FW/ERbv6c7ffPiy8wuWAm7YFTnJOCAZZu6GeBpEE/m6pfKFMqKpGd0aCzkijsqPcY8OHl
HFC+gX8hwq2xH/uMBFqu7Ww+O46MWcm+a7FYeup2z4fhdSWBupYg376Ol53m3eNlx10JdpqpwB5I
4ITJZGzzV0qINVgcbTdHT/wNqbpJJDf42pK/snpyQDc00QShxXCL8wgHyLeCeqftAKh1N6Dtybje
Vm+CCrziSvxtW90KPrSLHyx7QK03iIh9hfg2r/MLzApXWv2Bubh18F2+iCwPtaI0Hj5UKwMzle7i
lVMOWwJDrJZh+bR1WKH2UlH/mggUmNTBxkJ3zDHDvqGfR+zkQizBidJcXSbAQb9B0K7ML+wynPFL
DRbzUAY+L6kzQZwhRj8xHsVnNK6PP6od3Bvy+RH28GUs6KtciZuhWG/gI3MMP0x7xfcmGExfSJTO
mUU8mf+ItD6q1lNptz3D3nXvjuSFumLylnd0vHCVc9Txuua9aHZTg5YiCdSOl/rfrfwU2QLU10+g
0pWaiqPY0MataWvMswfmTKq1EIMxPS7UO5pRxyn6COA2lPAIv9xrmYoD2X6g/lKhW9MGkNIlB1rb
pkr3nUA/xA9rFDMezwax0C3dczu2ApataOTzv8iPphluQL6JYIdvT/s/mbnCM3C0HmCGOOShmrF8
U55OO9rj+R4Awb9IEs3J+hXfV4txAkdb9CBd/mMRllmMhk1HJWeDQFWKbaEbyaHVk9BUt4GG2tsG
yRDcYxM9hrpEH1vvZshTtUE8R+rUvkgRIwnbbFh+I5qYH9Mf2nEDE1gjq5w4Q9lpOCKIwIZkxhsp
4+px/LUJNTOZtzw/2GYaz3W9W9GHKtUoaoNOPvckpbXnglEDI13ysvL/4bNMb5rMwMuZPw7720uF
hD/C/NzJ/ANZrDPUfGkrIIcK+bxBctjAJ3k6g9KF08LxcSUYSfd5AZxwqf0o9SjacssbPHYyc5V0
MJkXZCmDQArEkDEVSbfeVeY/raQOasWQwiEoaVXHkp/auq1aBKBIEkUKy3CAVIT69O6zJjjqx+wG
4bWXRkOoFEEPN3aBNezPqxdPYp7V5vVcwU7PSCAg4o0ypRlGjdUM9nCjtTAYAK9qx2mOcUXKwywS
UVepbifK8R9rIFp9Jrijy2f3NRw2LspAvq51uI98jSWWojEsNwHmM56VxvRQPnI5RkozfZ5wIa6o
eJsSSxMaw6pNBWEfC/7/2r3t05fdf4I1AO6BMwgg6QYgT/OEhCvMf+46+ETtPuAqLuPQlaxVpEhm
mmtGwJUtYnPdQdxmdsP2nEfpGoxcfnnrFNbocfTYfKzWZ1IDuJFetPDyTAgMyUSt56aI0Z5kFhl5
b2FKw56E1iMZ5TEhn1I8o9UG69xPi6mjeOntBH+ayx6/ByAuGJGjugVbRuA+ORDOx1gWJrYCMPdT
DAauZyEAt+kKOTwhl0EQGJ6/ARB6SnLBc9/A0+oqgooFiuo3p+pSJ7u3uLNgn3Y6IhLK4c0LOK+a
2m7l33RwzN+TYB1vErw2Jzkjn3ilSmH4zYb5V/RtPIDbZ705CR2SOZttKSCfjmJGWjKc41ep0BPn
2qkeNuTxiFWTx0C/yDHnCYZEAkYwxgPNTS+c1Bcl64OdPK0LT7R+65hur34IjZXbxPBuJ4zQr/nb
zjla/SnAq8WgHYEPJni6enc3KzXwMWEz8J9f0DMoUHu0B1sfTQTKISVDv0YSy4nIaan3Ac94yep1
YSEwX8b4LK6fhN/Ss7FFBSF0L4VzfGMgBaWOEff/pxdoXmbc7RkaMh4V9Lbf6HNSVKuYK/4fFtlf
fss6EQPdYGxsKEbuFKlAvz3n2+LK2iSg3iDYvbuMZgKkwCB8gZzZH3ZMY3LItzMZubWuwB4AaZDJ
8bMruOZAK8W20nYRgKChUzmGAtXuKEZ6hjWp1+baSckdWgOGo0eXc0uybWIIlfeUXNLXEVAjlQ6o
N0mKwLBrFsW120g/h6TnGYS2tlGTJ8bj0QhbpaN0xw1ZEti4m8CgCXIzDxdA4HO5ppOzcgzx/H8F
NPM3ZHn6b6isyK+z8uLIaLjpYWSEWAyvdERFQ5ppOuE717TYHm5SKPpWm2Yg5aOnKyeNLhivBEpf
g6LIXmOJuSCJPZgrbCbeZpEnApTccn+rn9ntAYJWxEL34eI71fziHXI4s0pOt8oNf9sAiqmxDNIC
Ph/99SrnZHiDdekDHRcvKIEg1JJA2mnFmwHWhCKg2Ei5LoEnMzAODSGsccIh0UO/hjG3vjpWpuO5
+/ZGsKd8hec5UOQFJ1BvmdSs0bSVz3/+EPhJTP0ryunAylbpTlKMbsZgsTSs1PUERwdczsdRxJ2s
Q3S9Z6FkbAxdJLknSc2HVjsyCYsifQw/gOK0wX96fqet0zCNV9ziJmIO7XGkpujbt8glQNNM2LCq
knRn3uMmbl3ivt+nSuKohuQbRU9TshJzwaOCyI4qKdZk257IOZ+bV5YLGXMAYLnxB6NnmBWcvlcH
WUtNJ9tY6wMyBXlalRpAxjoYYgh2ay99PdWuOWFqFW0FlO7gfFrx7i/ILuNZgEl7bkWHVSiT3N/Z
8BPd7OA4Xa1W1wrfvryjHYXAVUrC3FxOUOe1AxprUe8U0FvpkdgNgZVXO9tLgWmggefTtGBt6YaR
aPBqyySUK+cafQMepIje559t8oPLj9TxCQ0G9ZzILXQasNCjJ9Bq1sZjzh//hHWiq7CpVIoqRc1k
TlmZsj8sXmcG8d1/3cqQ6wNspQHyE6JJTHLMPbH++sRT0MsemfLIlzxipgADslYcYTUE2OoP5JAQ
EmKgwWI4+GB6Vwi7KpocssMNG81nWLEAGWVMyr7y8VtFri8DzU8ccASuB1mOsuggMFa67Ug9UCpZ
NucETW7f/VSggBg1+GNT8rpOl7ezET9eZLmsUBsb4iJivcJzgt72Cuw40851FXf03ELsUNXTthe8
KHvCX4aQWLXSWtkJAtlXhwegXrbf1az1n4jsJxwzMvjV6Dv7Mpm/Kwg+jo5c5osnyN0s0AHpSztJ
aWrCPo+bvb1a/Ml8MNen7tgeNscrPvQ7E84XZ/0oLOWlQ5ZjZ9Rr0s7KSE49vyErvd+ud5ZPmJyB
egFoKKebKPjMOsJcXysHnLP5edKI453RO0rO+J6sQeKsfYPDcrnFMg3MeVPkzNXaCZTtc/drm1l1
QomWGfwjUyGWbwzVD6UGFEP+uB5MkF3Ou3MCTzi51Fe7csiUoHK2oPV2wM/nxSXJz57vJ08dXQZE
MU1trkwuUnrrCxinAWcHLlMw4AJTkNYvB777p1ugIbQuu9bGzqV45n3n3rJnZ1CvIaXq8d4qdFos
/i03rqMUdb6bBAH3ZSTzN/bqvvNA5yhsuQvOJawFOmVkfESzUvfxkX1gBgYJL261Q0uIUlhxLfyM
0SHKGoaWVIq2VN692IVC0vIIPqHBUw4WBARxtgNK02XbchTfRKijFie7PLwbjFCQHryNfRsN/6Pd
Jsiqq/WDk0ZwcLe3mB/ohOtNVchQcsNXnh4QW1PlkYOODgigcC15MjZzY1CWaAPGZvD2wJEQquge
woyuG6G4i5KMyoKA5xKxznGos2rby0Cgag0y3iPkY+X8oemKEio36IceFzxos2D6XC9RMJSZ5YYM
Y/HLjsW87liXOI/XXarh/Ld5de6y7IYGl9Nv9PxLS7gyEPtEhDZfNd5p2myQbvoQsSZGj/lpOJ++
5chlKw1AV1Ep/oBZ1rgUZ+MeNOe30CzdR+cB6SbpCYva7F0sfDNPZWG6ZQyP2bysawlgffB/yN25
koduwYIKLDqF8O3m2OtbxtOGC6BiWMto3dohdJr3tJzdc8kvu1rPgvtSApldO7m7uGw6J8DnuAxC
hO8FgU/wzzXSUCrgEBElvUHmXmdloSL5kFYiuL/3GjBv+6DL52rygnSyl+PsUEI7xiOSpdWQmEl/
47abLXWz5vMTyxdRH/w/uggwVJEmJCJ+xtqjIA51PPV2sdp1Fb9GuAVHYg9AO1rrhqp0XYf/qkDD
4R+/g86GsIrSXlurY02nz99wPZspfARpYLbbPJpPMtvdNPmam0ya94G75w6XwobnT5YkMWy3fkh5
YpiNdHzVYmkmAQ3a2zhq+S63BytqAzGRyuTS8KFDyaWqZh/FdE3LSs0647rK8Ql401sA70ZJz+dS
FqhwmS/0FtfJv6npYnILBmYSpLyf4k3cKUkwD2TWCP05UaPOuWJoZ6zI/IQRJSIVmqjDDJ4bh3Co
Gbw7TYOcez7Ug/E72/1A1LfpKV4ouKwDoKf4kQlcKXh1Qzd+Jjmrdbm1ial+W7mdv+MjDRVbqc21
M2VRE7/qT+LJKTIei3JxUWx5xkp/aubqSBNKyiBkM2JZ4w5bxxR7iZyUf/8mJEL2IrNt0oaXXbZ8
DCMDGYnaZ3Z9GyMqLMgopwn0iVL04GgJ0LbuSzGgKTkZyc6v66UE027hkjdwZbTj3pvHDUEQkNLe
5T7z7z7Rk9Movny69PXvJciZovETVwSCGIs4pAnkG/okYzVkJaV6YXnnMoHAWv/m8F2h/T/xvmSF
B1mgzECSPJueBRpxuJRjl5rv7GNvSfbeOHJW0+LraOZuBakaiZfimfP6KhCS1yqIbWftn5hMdsQG
ILjRWEtbGXP+HFmTcdlUCG9HDF06c+IXT0YGRjehdlaVdGpLAICXKZsN22wWeDkoOvo9q9hxfyoW
9t6wdF4mcCM0cfPPulgQ+nG8ItiBjOLclck6Lv6f/N+1N0vn5/xb42KQslATYpcD5EziAmDRXbQl
x/D5j7mYM3UjlP2x7VsFBvG1vsShDi3zkGligXX7aWvamx0ivsKzOpQ9kb1Tv4OZIiYvo4OhyzLW
1AtI0+ZAv/EakclXKEX70fHbs/EjPI6hj/hDIFb4vcXvH34tRJa3BC3k74fK2BAO66epseJYJ/d9
HKHo4yDwOXWdItoh7df1g/EU4uiw9B5tKZ8Kc7Cq+C+oaBFTapRyzcmsQ2CSGIOt6xobM5H/lpN2
TtyF/7q80jk0nsfixeKndYhXP0v1AFplYACWNMyEwXieOF6ryPvgTxJRlMu0VGwCHPQ8IENAOpdx
PXlFfLe9FYFFo045mvxS0uPa0KD9bAXj8J1AyDqMuO5NjcpykdE5BAq/2FIN2eDy4thyRiLA2k2a
A5PJNcPcan4nhKp41oksahMB/nk8vXbUxdbTOaEMCs+lnCTUPr+4HLF+fuQ/FePujtpbjyEi11jd
BzeyJidZrxEmQ7mM4Ed5v331NxqPAERtbzcdgPJOiLWIcW97/BsVxm34z9ahkT4M8RXkj6L4p2gr
9RZnELjaM3eZr6MbNNHb2RC2XHthsdHZSSxunYoeQKMeHVkza6d3hXyt6v1G0r9+dbGpfdoPsO3l
kRnpG2xXULUjSDgsZGtPfYkfvLchA2vLGmzKBPSttIMlJG2USiQRZ8mT7UPsvJYkgHB6AQU/f4Gx
9KtXEn2PqUaw8n5Rg0qefHvqYQN4508kaM2yFz28NJZc2Buh5aCMt18HGpjvZ+iFKwzq+UawQ6VH
a+XRMzto8u25JU8LF8M8vAOrLsKu1A7MPMfET56yWXjwhZLLXpDOM13Hs1W36XsI/eNWjXE7wNsz
H7FVBKVDdLk5cC1wo+WHqWbDe0fmPtuX6C0lPv4G38T0PZTsPWASF/+4GnQqiC/Gf2RacJiXFGE0
/XYX+nw3ZkoEY8vnSf6Zqs+XoTugoKE9wKT6KVFDRHwvYsv2rTj7d+UYODDicmnSo4tCgvCXPHxn
ATy8L2NTeU1p93WrcMZzCgkUTs2I7rQpF0t4RT1nVvU+YaOG0ECdrD3C/lacsWu2eIu6YKYZUeuK
T3uGVHo/6d4sH5q4zebHhJCrD0hzvWDPKuCT8BujTus5Ei0OQCOkbPi8ou2jr7NiW9Y0IseA+R39
cn0hV2KvU8JezCdy4Md7/krLMIvCSsY73tzcCoXL3m43lydpOsv/+CZbiOrsFNtx7SCf+NLBlo4M
XJ+F0vc8JWAKzGYW9wz/+6laMp/WB5AYQGT3Smz1H1YVlvJJ6WOOmhPjrd49rQ9Q6JByv4ZaI1Uk
x7a/1n4KFxH69gZB3dhKPQHEF0tCBePR8fGL+TsOJlD3lKwAOz3lG03g0LaCt/m/mc4MVwi7R3vc
l48WyyyD+zQh1SL63uwIGmqm3KTtGNV5RtAAK+z5dZKkSxqgvV6R2KtH1qExmpH48yEapP4M5cqc
+tZs+cmbe2qbp/j4VJtxaUTj6TbH/7eBpnnl4YdBT2kpyELdPbb7lC6Y0uGSiIk7G3KGqemWNPdz
I97GT7pQgb3QQMkjjC+1Rl3UfGp58Ks9N9lpVvMBYzGQ/mfszu8Cw/WGfOwFzQYZ3FI6aNkZR4ce
KT1OT5M7m4W1r8L5VZS88OZuGHKEKP0DSKaAdgHSUQYOD5gY23fsoIg+ux5XCpCLRPe3hhziNqSy
UMx9AVnQvoWiyPFz9HEgUYDoAqgWA/WS/0K+/JDFzrmL/VdmomTM6Oj2dE95kqUrG5jJ1CAjjZCx
kISPyiB13hti0O7rTXfdSBGnybtniDE7/EQyh04IMqMwce5CAhyEDnb5QeQRWe1ADM4U/nPOgAy9
IZFI75gNh8jr9oYp8lcB306icCdaefp/JVKaBMk2S4H9QY3jgNo3FnBspnYKtIFLRfR/oaB79XuN
d/exXcLt7bkcWOVfC3+lIFuTaWkkkx/KdbEuG0vQ4xXLjL6vo+2qJpwWmiAoZZjkDn0Fbf8Dhwgk
H5DHsEeQ8thKpJ4ItrcRGWMWyyvmkVzqXkOZMt2DsiAoeEnsvIBU+LSnbGMH3hKfCGwlBho/+FR8
OZbg0RpcEQUX9NWF45HyFqogtxj9GkjQniuVO8DZJU4+dG+8n7gFa8isGQy9GhlMoPgQHTn8QNgx
VUsbdHhHpPKirh0zsDsOgvhZYuNAiaT4ijmYvW0nRl9z/3Lvrc5M1MuYC/SUXP9D+WRh/fhnErWA
3p3+JZoSxjeOLHIdzRLNwTPXGITP1oMfv35mkxp93riZX5qbpqFsdYN6ceUxfTZTvwj+Cw9xSiQt
xlYMi9tt+ucdOYpPxsKhcSRxdRLUxlqghv2roE3dkFxekOzjBqfCFmvg5kdt6X1a++3jCgpJzacd
fOcoYZSPiBn/xjBHHupiELCM/6vHDWIFqQqZS2bxYwoqtDi+wcyBOeVdVhRzsp0d/2Ruqa0tGPuj
zPwTr1nHH9j9a5rsLPOyQsnhGVqGooooVRmYMtpHBndmkExVccoAeE8WvVA4gz0jrojE7O0fhy4B
sS1CK7XMLqtZCHA2YnUzXHQ8HOT6wHBTblW+ka5uYSTAPCKnU4wtgrIXfqFE7cqEqFCUBgPUIVxO
4iYLLQRMuVdOQo99BLkjpNH25gswPuIim5SuV7b6kCdzJDsp/1us6wYkWAPO18OubOOye6FHNQKI
1AcxqawRw+Du20jRm+nKY6zprzryQuN2JyaNML+3eNrIrWgb43/KizgdbpBDyqhC5AHNpWz1DvBm
2SHXSLo4FWFf+vj8/M1VZ1JWI6Mukg5A/AiGc72CavS3OmJ2wIU6M0JoLUelkDfexZt3a2zJC5ug
OOd1kceX3BU5Ga4pPOB8H6peRi+DXlXGBmxrfk6RV/GCQIFNEt7hzu2CX8nRgp4ohYE6P5oSVsJe
6qfJrRDKiNXrWGF1k6NDBYoUC2KravwI2FNnkhfBxndsxNzqWgUxdZOgVl9RIIggiCyiMqMqHz40
ZEHHWw5OW7WS0/uHQWqMmoe3LCNKiao6992y9mTVxoUmkkRr6JgP4MU+6zBTRVUgGfHggZ/3UOIO
Jil7905dNHHhaTzYNvpcxzoJw32dSXai9BmpcID/rV0dhzZlUwGNS473pjTRHGlK8Fg1/E4JtL9r
Rgh5e7Hw8MQQtzONMfpaEpxkFEbKgH8eC0RHPCtSF9HNa76r8rB0N+XPFS3yhiqVB5l435e6pzl1
98tiWczSq6qhgRpKK6BvtOgkjvzzWySkWV+LqEVAXeqsqWI/bvtmFAPdtoH3rUDNi09U2NydBfWl
0XCKSq8WELVRr3Lp96GwXI5WEOpIDJuJScbFhyD9ShD5NFt2MPutaRETSllQCHCkLZm43/2LziTy
l297XpWYvrrDc6Vo+kpg+5jwMUtSvDnKo8fFRqJEhzPq1O5m6jdGlDgJDc/xlYtd5BWPdQ533mFN
meYiw5glCtBsfcaTfjY6sR0Qmfwf32noJO7TaasGkHnwffnRD6owJ4g4y+67PF99Nc50OCBH15dM
e2AOdjRlsBBleQtz1uXBTJCOkVdGpbSAWT6wv1YSSJyyIbX4IyUbhTLhljYoeo8JpPGMPCC/zvln
XYOszwcFdckXcYQto4d25212KhcJkPamswfgarNt/dTuaD/nhzBdZOkp8lTsjTDKPFyEW8P/kTfm
ISyWrnDg4OfDyicRAl7lkafGMJ2+xI+0HfGjhRhxR7LJ1+1gJidEjMYXpEA9ikFO0HQrPF9JHcyJ
W8GBGnyq4AyBTmr41zyPnDpqTW4i9+j457k65ugZQA7vZHaTvd9hgo/4ntIQNnhko0zugnREIWmJ
mwrg3mM8ppgkfFw+ig/4UIp5nuzBkMPlxqCr4Ls4xk7GP6KxU9JIGJSZoJ0zTgTxbccHMOsu5Uh/
Y+JtHNgDMkMpqbGkMeSi4w6lRxgg+zEQbm3g2p247FLjStDTwYqAY8m0n1AKmYOirAS0bvhOq289
MihOsV/pvmeW+DgbvcaQw6PmKkG70L3oz5flSpQvUTA4P7jnxskWCkkkdd6SXNdQSOe2Siexu0SD
UDoeFYtpKYKzlTlYSjT+puEhoBi+VvYytxd+BOfwFjpf3GlVT/f7r9GZOifyYrpvfC0YYnCmV6yQ
SGoG0DS3we+CNo1s2yikxNI3F2kd5IwNsv6bnQLWWWSEO1aXMRYREkIhoQbeUln9EaN7o3IPoU/R
sLY3kyRpqbVTQW56yoMaFjCRgfcy7oNZi39DOvjgEOSTRhu0DwKx/5cuaHPYbP+SNMSxpMh4Nx9s
7Tal0s8LeXl8AN/lJx5prkW6h0UpOic0pM2KuhiTRou4rN1uMWjTllGxFhb+dMRhWJ+dKSSQT4fs
Gt1Jz4rpa5cx60eL7yfcUZY6BfvdWcnfSTmxfLZIIztNkBE+su/BITuGfwU/ajNAxtf1wYxlnV+H
wJWthh0YwEoiGaYUdAPBTWoG1YCUdFq2h/T3oUmLc7QIRgGducocArIggTXbqAwHB12rsOOd3Og9
ZOB//jmQK7U3e2J+npeJ/+ICvzsPUNV4wy53LwfKhYfdyrCXLSoSOa8p/9h757ExpNoB4yeoGrWH
29T7zPn6vVn573ofBvu82dNOYa8zYF8ezCsSjM14ft2PIAAh5z2r977ZTDNYUvywYZUYFWBqy2B4
OQN2hv1VBLFQqQavUHnvakp3DMO3QaMxhi1V1ZJpDHrhVkqDbrrnVl/JD3zogtJ7IcScJyb4hfTk
0XrXI2Rdi0vcqclw7Q/46BLqlNd15nttTxT93mgPjJ7vcf2d9KW6jEeslXzp6mBh6Q/BqWjm1DMx
KDfilfTV1/Jby2XR6z3eSlUattk/vdtmlvetnawwMZlhL5m5K0HI90oORZAcRXAnKw9DZRqddVq1
ziowThufv+saTTzYZOuBB4+FXpoStsiNk+lN4jgEUVpI/tkZtFHnYht7sddOxwMidWB7VcbiGsYd
BJAhCWX3JDX7e1R/Jrn9WXI4YcUHwrHmDGR08yVtIshaB8VtV3lljYtl2qjifgnNTEBJinQdD64D
bvmpo9xJ8ehpHSysMfXI+ZIr4wL+u3CuQCVBU9PNEdPXu7t5874C10bzLdWwxMNfVHENDQuxKAEo
mlkQDZiwkJXrMbEXO+r2M5WMbBcK7vr8n2tEZI26NWQEyhdtXz3qJ8DLjQWBzVjUaGVMiD/mDGEm
KpNRAd0L6OF0KWc/+8/HcON6o9vSOuW1YjiOlqWVttNYf05rcnONiwDvMSccE/2J0ThQU/jAWcKz
7I+zDNbT89fAnKc1iYR9jO6MAV1bZ0WN0wdRC15xGZkjTTyDvv2DddzYCk2SvLutlz+V/eAYBQPy
ZYvkFlorQMFI861v+OHZElYT7/PZUgftQtGsQSWLHNtRR0laDZhmqVwUdEJ5EN/KXnqNHq/H95fq
BeDua01C+9fy7FmU8LNaHegQ6tJ3hpYYMT+zYD7LGOkfU+U4J5p3phGzQz/qo+e3MmT88w7JkdXX
5rxYTrPZupyBFuglh7CndmMDO9i3NrB2sdl/TqVOaMtrYRqPYJbB9jvn1uzVRPb7W2cvqvokwYc4
EEC/tHYCUB9vA6AzVJXa6Taussq0wVyijrzazj2wOjwFX+XckdSPbtWlVZqF7U9iuhihqnd07Sj7
67W+++X2MJ7ZZncjsx5iTNs2kgu6EyZwzLd+zIP2EYI3A0eeet18QZw7gbDAfZzUmLsY0dZtNbwU
JMjwe6AsWQ10Hfzb9NpC2s0n210jo/RybkCM+zvPNq0fTw364+/Tp6vmcEVdBC/Kwp+lUw2Uh0pQ
6jdszPsk9rlnJ9RXYUXMnDwvcYHJXjqi/8YHirGm2m3SVn3TUen9xNj0IVbv3PVjsmjEu4Q5+Hj+
86617DxK/JDC03ZWS3qv5rup8ngOxvnwkeVnMV996Na62w2JMUN501T8yfxJcIOyHXRY/miBKN8J
uH+bbhwuctYFrxEGJmNRJhTwBLcJkV7bJRwyG25pQjfzTHnzXG6aI/zNlTiwJ5WbS6VoyC1mKB6i
cz+MD3HZET/1MkCEZ2jXPvcsQcV3tbN4Uud9RLF2JPWgufnawnr4Kl2xLsOVIlQoqUSEPzcHT+8c
vTJQpRiIPGfQQRcLrRh2xirkr1szMxyYFciU+SRQR36EkRtFDAcznBP8aPzPE9RoiMTFs2o7z3Qf
mN6/ae2ttZdt2ziV3aegd6ZldteqnIUHoQGmDRXIP5m6EzP9tAofeCsu/5eAf42w0NDT3mWrOL67
uhUmU4XpSd9Gtx9Oeg+ZpKWQHPMlCQ9PPzqK/Nj+pPzGc2C0tH4Z9JVWQvNTX2oGEpivPxv+wjGa
Nj5TDPodHuNakxKzA6I9n1j7Ws0LPelKxgomgHcOfz2XqPlwJL545OY+ZMdqNNWBa0gQrbQ6xaCT
Lon7mmfLHxSIPNiwMpUl7lsqyLqKK42eQvFJ4MmGse7Nd4kxdIEv9XHVz64qvbty0OiUjpkh4xqp
I46vnUJHmpPUezL49DboEl/QbrA6sQIyyNCUeUaJdVYDWkeEpwsYou/8pYdpTzl4YgEG65adaVAF
53FlRdioNGhHt1X6YcugwVJn6b9azW4oOaET7xPal18miyudoIF0lqnBfPnlLYbrUnTfiyodHk01
rp3pizoUVE8LACgb+HFQXiQ4d5ZKF9OM2pAQ9jMuIbo9tlkkd0qzLlJb9gAA36QPkOXWZwotawMB
lsSG13L5CvWrYimSHQIl6Ck4pWI3VKqziKUx50fQZGcpFQhD31VDSd6vRmmLb9Dv4GOyO7OdTIHt
paQsap9J9/+jucScScKI2sdWMNI/g3CDvr3hUBn7zmTUhHbGTwuPmRCPJdrPQrHxrwZUVVr9If0X
Lrb4d3UBrGRBjySeM5+9ww71Gcfw0gsAFtBmzcZqJQuOAce8+k8jZw6EjjE5XBiTJOPQFjT9EUg+
6ql5xWwF2wvuNhkWEuh4jJwxtnlalMFKVE7aBjQlIIrgKvWyj3hTM1KCwG5OyBI3ai76zcgZvDhp
pypUZAKA3gcs+Ts5+xG6gUjFpvW1EWlumgX+VgKMVXZ3cVZbdQIBh2vt8c9EDZ9C4R7K6MVy5RnY
9hu6C7+hrIjcb28QU0yAX73q8lBfzbF6fks3Vxl4bRjEYneIjMZwtYfBRr/sEGQg7hsWtBLkvDil
cYj0z8eU38m4a5jWyDsy7++sBdmC6GB9tq6N99I+i7WH3hho90dNsyngLrWxHIND1VBNdLRo7pwD
Hb3kWjkeuh0REXf7Q03lH3TEkAM7z8O1Jwbd+um2fizQqrgyE8IbK4VD7baXCqkm1U7Jeji2XutE
Zj1Q5EI8NTvNQzDrhJQr0U/x1vBPejyUpTAxvRFAt57J0aVRhuiykbTip4CsQRADSkjoF1VS99zu
OUS58Ve9wI6DXpok1VqkTZxjcvuykQ8GG2Aa/Kr0Mw5bYDG3GD1bKvgBDZy6+40yDZmkZTN38BcJ
xZVWXLOi9bzDygUmEHlW+8uOjJrnK/ryt33X1/yc2s5HCwXqyUYPUjxf28iquO+bzybqW+gOpzGS
5nTa4HZAVfqCwgfa2Fw5E5VmrU0x9UWtEpn6r9fubkCKbQUQMMEr1EF9hDuVUx5XBtRNeUoTDjzf
wCzIkybMKZkxhqA/ZicjRldoJT2ieqllpYE/ZigNHN3KR956Ocgu2U7Z11v0WsHUmnS7PxbvLnKa
8R7VsXMADb2APByMlY8dq/77TID416ERHwmInYJi4ZGAvnz9iTPVg6A3TpXtyqpvy9wGPX6NY6U3
OXSXg93ykOTKzacFEegMotTbRv2dgI/koJzfBwNLm8aSdkSxNfhLNiasjUV1noreIP34H/hAyclQ
4HDJ0a81gA4f4Wlsi/qeNDU0hEE/I3/bz0ffC1E4Jgpk9oiDNEisCcmce0FUEnbU4c6oYomGJF3v
OyCuEtOPRrVdfreYXq7qW+3iwGoBYkYC/J3PZdBwDaLlzgVYrcnHsMzTndD9axkw8O351RE7eyxG
RNHQm0hg5YHXFyDcxGAg11t4x2z22HUDOVZV1ONMDaey5v4TxITgTlzx0VJ/EwLjfm4VTzWhPWEL
pTUt15QkGU5IReyLMcCaHlyFRHm2WZ3tcW5fDwxeHcbAD9myblt9RVudsOBh3uAf1BHW1VPOvSOr
uhE28pfmzBiBHX0dt5AZPIO3P/uEvXkOU+7RuBvhfRB5SNePHik4p5Ujp4W9vUv2LGjGU8Pu8YVF
QwxC5Y5EY0vAGKRQQfw1oybA/DQVcoOAVKs76ZlWIqtB03c70kJaZABZJXQmdV3Cx/vdVW+FaxRj
E62WNUJXLncxLsBWJ1rZ6e/TciKIL08zjYDBn03z/nFzJsdKMyuopIwEaf5rOmFZGneDzTvNX7ot
p/HfCG9lac7v1wpnzPYsLNBYg5oJNkeEc5x72t+3nWBI6pEP1EOu0CQ0K8F5YignByKsesWIBi9H
cNA8WFtVY8ZzrBE8A74+jklzD9xpcWwiJsKlOhj2WiBkfYxpUcrvw5p7roQYQj+ZHrkTa99wJ5ec
ZxDFfvVQOocxQnoWe7469eG53my5j8CRL+EX91/z5vIKSyQUA0axjfAbWroo2vOydx7qZvEbaDjU
5DguwpDd8c4h56+yTypO2U6+JQTl046ArWhl/LR5aPeGQQoWMCeYjiIzawuQeWCq88R2AC9c+Ci2
hZ0mMc/r7qQIh2lr4euhlRIYdMw9UjTg3IbrNmX3mg9rWK/o1NqQQLWioEDJa/m7P6wja4eaHLSq
xqQY1uS/Fhm8AIRj5c+FZ5FAyWiBhRDhYPbiqPl6V3ZUzCFMwK4JtcDHEy+pqb7w0eZg4J1TfXWf
v1c93OIVJ/d2kgH1ooHOhnP0R8tAwL3Wf1YMAYDCjKe6iEKPkQ1gBQpS0SZLCsd4cQVY+1CowWiL
9F6/mLe/+d1DICYfGmz2mLf4tGkBhTPEb6Z6C9D0Evz9cjhOoD8AfY9QT3rIo97SCEePrgZFmq9E
3nk0QsBvN8gwJmndbRdYZ2wctZMU3mtmpFKbapwuApYYNphRtIJYlN/zxiXztUoKFQ6P2jjFlAlt
/noi3RBTrI/HdqzaSRLD4rq6mK7mYr8gevLV3+3fkZizBVHyYOg+q+y38LXyzfTe11irrFb7KBBL
twvOiEZQvFwNhoLC1EjbrNmzmuEMIRN7eZNerfzwvCcD1H1LnE3k9zb1vpcIaaz1+uYQV2ISSEBQ
XrD+m4rolyMEF0nz3x0JZzexNUgwhwNKnqDGkavCgoEuwhnGZMNyPUmgI0OW3/WHP5wZwa70olPI
OBcBl06Cw5SUGDvW0rx5GOQJTStpSD1wv6o6pVWEkVkkIlzA5XD1fHifDxbOIa8AA3akFNZUPgxh
7QkmmenMFQETCS71O/dMijL8hXgLCdwsSvxyYCmRAEqPI0ItR60DOcrYP07HFVwkZN/+LQ/s5/MI
E3mcO35We4LjNEO8XHSE3y6RbI9WYISUUSluMJqEq3fbhL+DDEsC8M+M9PF/i0sDUzpSovvQevAg
UgbK5HIeCC66K8CCJss7KY+ZhyvABTLwjn5dRb19xhpraVZP++kJkDrpvMuksWPlQla2DqETd2sd
62QTOkxOqf+xkoTeykrcNcvzGJT1xSmsQIPzeyecZS4VOOgfHpxWoP8WVdTreDC/drJIMxBU9vld
R0ASPPoO1osVLPREoMiFPUHEsjWXzbYdDGDcMvT98wvX/8/CABAgQuz6cNj4ShLcybTobRf+Uywu
HuoNKeUB33MgmvbwNIMR21XHZ8stSzvoK25V8D6gV68l0dVcN6Tf/FqNv3Qp05z+Pgx746bEjgHF
PxnFbNaw9rkSmkcYr9+N4Pj9CPIHC/tKpWA/Z7SueoVauF3UtMK9XOUQhTpUnBPmpIg7IC/pjzvL
LJIq4oLrk9c0/AVRB0pV+6ARK27NtxTR0d87mxX2wNW4h3HIvp5fBK4npuFVo6yD/2gaqvUqmbvw
3+tqM2+tWNlLKd7yR3jjql1MhDdwHVfZxRA5rIhxTizcgRBor50PocCFH7KZkCu7uOlQ2YEEHEIi
E+k1mCBdE5rfwuzI1HBB0O4Mho1672NF0VW5ndfw6t4FWd+zfqR86tx+gP6FNsGwPnA8yS3d6oZv
yo37300KxGU4+BHNLtlT4hnl7I6DhNxGeoiBPkUIL3U3CSp6m76vSoscBeHJ9VidgZjOeocQfM9T
KnaoyJS6KcJq6aw3xtj6982WAQPxwCa+nqDo+olEPBttg1jyfACHXCKOpifcAK0NpXU05LQ0dHoe
KH2IHt5/PyH752wtrZivrmN9vUfjBbV4cLVVFzvvgP5NgM7Uypuq/pa+hy4uKYuYW6j7r5it6Drd
d+tiIoC1x+9MU+6abkTZQ8pUOSWXYNIDwamU+VgbX3ErYdM+gT3ToUSKpiGgnPSGzfC0fm6MTpkA
m5wuBI28sTvtOxxjCMsWjfoGrLM9mJmao67x0Mwihryms2YHju+oeH5KrG11Ca4SbWkDsi0EKUy5
kU850vMlCjBPDSgE1T7/P0Qmi+g8Dd5ZmR//i8SGZoKbPvnW16hib8toyrerqk7rdvgTLyt3d1bB
XAM45tTpINLDpr9RY5JVEWYPbK7VtJgTAxP1b7rSq3GQ76SwlaeH7FCjN3N85jrzaCOuKOBopLT2
PQpBuXk1aqbRtag4lTxyEgiW8C6ro8wSoFqYGlbKP+8CjT5k4zIYQBeTHOUxASLAIi/BoRylrZr0
3xNjVHp8guWA+dCJIFZqWMSddgvGFC/f0tMVv/skIMvIlb4R1o7QT7yoJI9s8e/3/6gHP1NI3K7c
q51CgXAzzf3pzoO6/hs44L3E8gintoLbZGJ4QEktwnWbSura5yhq+Ii9mcgPRKnFC2HpW6yoV9bT
RvrI64d2NnPOz+PN2I+uzStQ4auBkIc08imUNexdTU9Mj9y4HtZV40TV+/EVnhxZvHog7dsXWBE7
hAgciTUpwf0RPHh78vsZg0tdSRzMmJaEAZP0yfZjMg4+VVOPumS/6qULOuGKG1/7y9VoRjx9Vq33
wJy9guxMWJvdCzevHGShH2m79Emv12W9kQr9BPPmlgcg73C84GV0+hZGiLvWp2AU8IlFOpU5FsAC
ZQBh8AG0NlsRqfYLH9YlRPt2aXRZ4GFzi+8l5Zh+ZYs7ejXRgt4AbV02ADwsAhW5/vs7W2mIn42f
aFr2Hplic2Ay+OqD5oO0EGdBaNvrfilgm9Qi7/J+GAq87SVk0hpor32s1C2Vh6iqcwL5a/Uqjmh7
DqO/XesOhdoiYNAN7jOU80f88GkAzycCkJ9dZihNCobgaxVk/jwuIlsK1D6ZMr0iEqLuoCWw7Hu/
lKHZatWekbm4Bw5+Ddmn5Jt0bqOEbBThqY+d5ja1aNYYRI/Kt8q7Qg27YPmJn8eIN3JAm6LBZGSn
58QXS6vlemruIgyrIf3isDV2Y7RM3wChhOaxVF2zzMgNqSvrntpXBZZ9uMBN5MJqAvuP2qYmuLnV
pJIm3cQfT9l4eOKHcRK7z5yP+0UwpyVirFUGjbKAGBuzSxhjH4kx/IAcXZjvE323QBhnuyUey21n
LZ2pFfVkzON+NuWrHFsCKy0wDHvQuAklaUOhf2pkjv41cf54kHD5ad7LlyJY15NAbcmZIM6gR63H
FzWO6sykrotyqcNTnpE9NLbMdVtf5v8U6xfryrBt3hNbDEtTkk3x6Ze4qzW+ofQQNZL3uVmPYXcl
ij+0WAxmwdkyoxOjTXiqzeYfzpzJuGky94qZhQclat1x795Y/F2F8Jiwlve0MsFloOG97U8WlNFy
i0zv5wq+z+iUcD8GVsfNL9WcdNDRAezPlCOL9uLV04OEwkaObzY6CgzIxH0YPkCzqb13UygUSaOh
RYgdm79vD3OIkwni7SYC8QM8zunCyRrEPjbCWOO+Lnq9/JYw/XPYllHwgYsutMNxkx//wSgtl7l9
jpyRdHzRMIPjUfbVVA5yXPKvw2MFxvcFh1y6+WUgsp1lDGR3as+npcpOYUEZwHgzTwIS/QSB10Kg
sXARBX0ic8YFc7SIwZSH7RhX+HKWzd7k5dN9m87Jj/vWWffHPovphQHj+v3sgdN/cufKjvNk7eIw
86YKOMdU73RYUeiA/12oPPIJoaMv1XbwUB9yp+K7YZWyN0Mv/WVV7Mp/wwQLatpqm5Czn5sRfyCV
SPqkOJvtlrL0keW0fxq13H7B1WpyTu+4vXUpJf2bPD0ZbRTPB3qF2zbK4HyZEEJ6GcyP3YsCTMIm
G+cAq4TQIxmc+YJaNFwpzJJrkZGGR+s3WORk5W7vdSjYHjUQ/XKCRdjixXOI6430v8DOjgQwvH1i
HFRS6GPiKUyOE3DxInHhq3KpZSh73zVdkQEMelD7fEgmVUbNvPX5WiHOg1+mlUvrJxh6QE8/rvYJ
etehN9vZXUldjg/lGP9Mej5+fSRRQLIAPEtzSvEeKFTTCICFXTx1es+0wtDhmz07cqylJr3fz6fV
RbCu5zdIhN6cJLOEzgDrZxTMg0KX+9HdMrkLDBs7zkV7qNF2061GkmP4tXa6aJRQ/3afdczS7DIX
iepsG/X20o2nkHdFwHlznttsvNRK00P7/Y2Wkbj2RKh5+MMVKZnHktRUgP8GomQkVp2Ho4SBo40M
o3mrSihMSYSXBaRGDkCMGIlF7gPWbM2/3LvO/fA2R3u1J5vBBRBn11tRZ58uTWjZU2IAnHlbQTp1
/zAwsjXyiEzCky/sh4mw7XpH/nYdqsXOWqeSguOblVJaBKELXFeJ4qaNA5hu9AUQ0b4PD+YXX08V
s9m7UAIHaOgQxOIiOQ2rEqBG+EhyvlQ2tR3FOvVpfZ3GpVTSxtWFmuibHqa+PeJOnZyonzAWo3cp
b/7o3KC2eVBT7jm79MfgTmgjC4iIDXPcsWw/Cx+VU5kRPGUXecjWgWho/tomD1+HYRsAeyf8LpYQ
j+ow+3E9A5XdH8opZEzfnhfVScI+KYWlEuStJ2u1eDZBKOlzDOB64cdvXg1qv4Nc+CL7Srppq8aH
Zw9C43rCzIaumhsMJNaRfbE5E/gPOSoAc/wn83AE7/Rkoh3jTMNche+FBvyLLQqHH2WrovEXyYo/
n2nZF+8ktLQ6DAOwvdpdAZdjqaYTTqhLvkuQmbu1AuwwKTUenorIP3HaF3kud2m/TkwaFGcNZ99K
wtnbKaBNLBczSBS0CfMfuKfO6EZmDzqoNF7gB3Q0XisgglE2YG4jLJH4gzv9ZwpGUSIGW3ZO/MTH
lvmXUREMIMzP8xqcEjvcoW/WXzW8JZ9e/hxxKrgURBFrppc92xaLhS8warMOi81O5JZDcS0nKWrW
bQf+NLyHLENb+ZR5CMwkv8lLx8befqHZdX9tQOEOWqEDhFXwe1q920oSgpYh03K9qWfiY7jkexew
gEu4tp3PCtVRliD22ZUsIqfRBge93N0czN9rCtejPix/nB0BONLLWs2Oq0QjwoMZxjp9LecNsSkP
KpHHpFnJt0tPpauedmqJYgLDPKLqC0PvsaBSfHMxG6VOXwJwSMerY7NIpJz5O/5j8NcZPuBBDum3
UrIRtyI98N8Wp64O05GLkav7j6a96NMzrry5WUsGMcQL6RSdGBIPRI3L2Dj9DSrwiWNmWDgDop+l
nWjRsvHQIzHeDwNx/WCS5/gH7MqZbOwYVMTqvn73qyWLyQW7kZs1xxnKReJuWsg/A71tVG71CMCW
taF5E8E7nAYLpyyRGWwB8I6LAkHdMzCm1syJ1I975Z2xPIkGRUlsQI1gx5fK2muK+suX38CKc294
WVzDI2c53qZ3nqXve5iHIs9uAF8ioCHUXMQQIbC2wHMjEijTOC/HVBF4yLVQlL7uZPaNrTjFVjJ1
EaeNjdCISfS9a18Qu7NIkbAoqVofs+sInUxatI+RpA4Arzp8VrMqG/6e4yzZl/Ku0iArlZXtqAT4
LJcGYyP7uh73jYIE2XUVwwbm/XAQbM4qz3aPDUalEOxCV1XU1ms/tA/ZOx5TaZK/MjViSCLU8jlt
KARgt+KwXxPyh4NvwMV3ejG2cn1WbLo8FK+JJXKAxnLPF21Nz/uSDkwh/tnMFf3jRrwhRCGjgav/
bmo1jOqJuC8VMunMjLGs5l1BRAfMPQDGAOFume+h8PFZ1H59/XKRU4nuSrLCo8G/wv+y+WozSNum
geAy5YZHQ/sjTRKryGauMBJT/7yt5f6rWKa0PLEMXhM4AZP7r5IO0vIx7LP97Uj8paEF7CMcQOuo
SNu/dG0Lrl/Lh5/6GtX0DVRCzPJsKAin8puIKOy1MbuUnPSkxcYbEJWWwY31+Jp4+M+Jo+/47jDb
zYInzfzHHeZn/UZbW3KUE4RgVTXYBHD99cFkX88HAbCrldtVHDsaiYSCLzdvQfavjwT0P19wReX0
0nsZsOmR1IE652OmQKwG4B0eEOZm2OJ42o5R9SRsW2ssNC+x8/H4UdwOEHHshtBkT3aVgHv3PQFH
s6XywRvwuT7Qk1YUdo9JTxuQ31xJgwxkSaNDyO3Yg8/Jz5EBYk+gZhm7cEFVf4sC6N2TjYsuyboZ
FVZlu7bMCZjp2oY3EyjUYztTI0vuGDwmSdSc6Hs7qfn0StpATpodi/i21etNF8efm5bggsrpYkNp
EFpOTH2H6/1UyDauFO3lhJXcMI6vDQAC+/iot5JOUs/CLqIVzMHbsq+BfVnOo1bzzSwgFIYCJBYW
xUQ+vhr86I1cw1+Ci5Hh0e3dzM6k+fzlpoGpJ1sgfZUUFW7wKnORDdI3aBxJytvxO+4UiucJNh+z
Hz+H+8mFvUC0dNHurtdmWX5zkkcKguZQSMG9fzOF6Rc4PQp7pp0neTmI+gORWnNd+0/J/RPzaEz8
zMTiAci3encTrROWRkdUpfLnzobK1K62WqrsOB5pxSLIvnrza21G17fx0bm6PfkXzBZecUTXuhws
k6KJ0J7LUhdKJY8/00V1C073cImxOPNoSl9uUOaLIRvwWpPi7aLm6c2N0DdyWYcX0wYfytu+ItB8
eZjYSWjPjq0rdWlwKCcOTOYMS0a55NmEFhOl7XmSddwXulu5pjsbhvz6yghB8vDl6ELJdlhE5Wy6
msZh7Rvbzc2QhgbSdBros+NWKlqfdeg7iMdXjpnGIypSzn5NGEU/jEK3QBixcQmZi072JabRVSOb
jdnjb5IgmdcSIOpvXYU7xE9J4TKdcvGu9hIz4H+iTogmreMUsrMM/IpSHkAJKn/SQ8N7NHUiyNNc
PGerg0Cot6kKJc7ogPRir28CSESYRrk8piZYe5cDmxAB02oeka1V28UZJTxkhGzm8yEISQHFqJQL
ppU3qM3fd6RGVXc2LVTRXulzTdTC5oq9M5Hk7H94m6LwIYNNRIBV2uyXrr+/keBYEzP5yrYrbvyA
I2VQ8fxH0oT/oTkJfSZUq+au29k7V54dILwSPHTyVge9FxGf66WEgvkTw1+vSUETZ9gKnUUQ9Hy6
NWZZFIeSPl8GQCQet6g2guIby9Dvr4i+69C5ZpsV54RSLx1FxdEAP3LCubfGF0NAAdi+xt25zoo+
mlD33s60GkNDm4qCZysKDMrTYvUv5sHgvxDWzMh6egmhvlhlGp2XQBMffykerAHeiE4SNgADcx6L
QnbDojdHc34gqiMZzZhEq2pOZw/uyOz0TPLrGjyXHbecFE3qXA/5VHjYqNr+T3/1kXmP52NlcC5U
gosP+IPSMW8RDwmFMUFAuF/a8SbvJwbioebQ5Ci/8EC66EaYxgvA8iQxnZz4C+YfaeKx+73zgjJc
IcblsGbSlMe+VPzpX5GlpUw8e4Vzn0vatgfxW+/EBWBsjNci8YZSWxA5O3kjGkeQJNmKdUerTIMN
XPP6AuKgF0Yko4U41ZRzCuvQsfBep4OeciMFaXa7wozZ+UmL4yX6FePhW0KbRGzLxJzkCLq4ADpH
y3FpIdzSklWOe88OnQj8xyZevNiT/onkCZX8oeUMz8hn4Hrw2rti95qeSrUEdkpO48hmTeMVmygY
dD/ZSjMFu4S8shQJi96DPoeGDuBBDAkcK8zV+/JyVyYySzMEOnYtQdU/2eokVUTL5N3abuP5zdWV
vdFYwIqp8ic4Lld/VK5Zo07s2g9wimdqyconVKfS7jOxYMLhEp7mXicFvxLuvVx6ppKQd2R+VB6n
9M3DMkTUo+ZJhlTc2yJ67LjrwzwNxMpeCg9dhMin+RoLKwShEkIbBHqOBeh0DrbMZjzha1kULl7G
UDvxJj2m1cnVf1BA2wXBqDibqHXaZdA3eFiLOR2CHfaKcFfnGGvcHo53/JKesLi6Fuot3/fe6THL
b0Fv4fyJe2rj8LHH/7vxJlWrNcHEezM8sUpFWH9P+9xg1Cb0PnZoVKv48pkFPIvVBe1U031Jf5xf
47ual+cKb3jZfgjX3+jMdESoR9tafMM3WKSi7Eavk+Gv3rcw5PQ1YVFtiVqXjkEY9RO1E6bXr9h/
hhwgY874Ioz5V5zgvuVgQ3Hd6OfEtoZ0c1AQm4vS+zB1toqaYKLOxNdLQ+WrSHC0XAvJhq5vv4QC
eJmOc2XgaI7tbFLvf2yrNzJRGiBy5zcmPKKxSVOMPWovczi+fDPZhr+Ax/da6mu+OyOHtLAWBRCi
qJvtPtYYNCU8Hm+mm9j0HB/JSh1XOWwxE9rxgXf4jx11++1wOskbuebBJFNl3qNg7V58zQV4OoDy
zC5eiHEiCpZdTStI/4ec7K3hntHoHC9C/r/YJdtU5C7Q832wSEvupBfVGjY7myiabpIWLXI257Sl
oGbFPj1WZCJn7VELr9O/KT0v09oSIdibiyAnbUjnjfbIcvboT7iO0brOaNKiJ4AmI5mDjLsEsEzA
rocWUTdPukVgn3ZfZ+Iy/oy72cI1a+2WHcFR48vetlnTgZZAnU9/vJLqEeBNc4ab5Q9Gh9Lq9nWl
721v1WfJoKZl10Ih+zIlajJWS1K2gM6+3ElYou34qXvE+Nlp2VYp16OLZ48yq8mGRA178ScnxCDq
9fYOpJLgi5I1uxnp7q0ZSOjEkX2e6LucGgdXnx+h/gNkr1VusPZGh+64X6//mGO5AOfUVMyP073C
S0hxku/Nr3tZurMbwSYqAR9PAeuRD+GQywwJiXDiHbEJEzN84u7c6G17T+XAM/1T+7NidPvukWX/
uIZx+j8hSyzhjFtbP3COj0HbzgR8qxb6O7gaUfrZyp2eiIwJVAaGmTm3Bmv/UoQBEvYT8lHRYsek
YDHI+7FQhWG76WkIt5axYAGBwRaYYFwbUeQPaBGcEvjnjWbzZwm1Z/AF7TCS8On5hCkeK1egoTHJ
wrrCvv5XWvkzitMQ4JM8PwIbIDaC2grQwYxrpbtdZp5d4fy03weVnjrSKveO4NNirC4xu5htNdaE
O9mToY4lgmGtn7wa0PqLIptSCnEt8CgXnr3OUUaC0nN7N4Z5BA+uCL0TSlcjFlfK8qge9qMu1EKb
M/BRt6FrDHdFxnaP7UDnneXlsBiAjCWMm1nk4tSBeuyOXVtCzwyFVHwtoMC37PCippCSuBNYeAi/
oKGyNDEK+t2dRKTqDy9joFhW/EViR1I4havcUJ6lCir5tij+HTaSbQTYxNttuVbWZxDnWoMLt+qW
NN3ezq2tho2KywVMSbcKmjaJbY39TbkiGMUiROK2JW0wwO4Q0u9G18S7egWe/axNlT3pRmH7DQp4
19+8bOyFyA/99TsrsKkAPVBFAYc3ctinL9W9pjMUxZZKKo+vhHg1ibCKh9nDdDD0qAr4ESM9ZbG0
jpDZMs4mNY1wMmq5WMSI0Tra7u9D7/C6WjGNdmePeXPQ8cHfPLvPVgCfYzq82q/YJwli4kPEOzWa
RsQ1o1ZDd+KSLCBY7haNihXsG0pKY2AwyUsWBAmSCxSKra+WYMpBszuaVbOl0YDIG48gMnE03oIH
6kvUx2tnwh5hBt18XS3dEr7fKKiorJGVgIcyH6jWkhagr+/19UEoHDWdphOdwtzbhkye8CRt12da
JjAJ1bHxkunwthV38hd+jApebkn14OxggvDRyFywJkPyRPe/GOXu0j+U8RXlKbTTE22RcH8n1YaT
nYl1dzUea9W5qg6bP35JrduSWfkDGHZk1s78e61pez+bBGwwo00XPRNKXQQ79mbai7gO6dZU43Cs
UdtqjWkWpGyhSWcvHXVAVs8I0oa4SEbH/Voeq25D0h6fI1AmHrAnfjnwhgvNfwjdpzKI1BYW419f
BqpFzIvCahByJmYja3QQCjfq3KwPdvp+x880wzNzF+PnHOUPR7Y25nwkWy6qJFty5YGKBJXuk4Gq
Hp+te6RbbKZbjTtqjogl22B/HqzLgNORGc30yKjAwdyc+xhZh7MncSTTQbaIgfSU4d7br1HS+Gpa
YjAOeJKu+HTlOpG6z3ONhXX/t6xMG3z2mi9vAlFKOUpk2/DptPNYu9gJSNq1DAdxWphUXmh5dKyP
CPIBiCJmWDZfcZFieLqyl5eF1wdC+KmmsMeZrfblFHiFFyOixAXxzmYLAXZP6C+s1PssHkNLrzix
g9SYHLAw6A0QYE8Kctad+AFof1eZnyTGRuQFZG02gKumH4k/oiHooQEBYwrn1zxM1UUcT2qEd/++
oVpCKnqhPtmi1ZOFwGJTAKaSdAUc/HEmoPtoZ9VobRLBqtvjnT+fsVulpIt9D2BaoWZufkX8OBU9
hxXV1E0JMrJYAxJisMoPhB4ieUAkFcEA7dPytCUiauvn5VYBgih7r3ZJ6eOp3SV0RyRPNlpR1mih
9QTQWk/6cjtKGS0VbOpd7R4ume19stO34xXvjoHEkSFVmM6nhEv8r8FjtM1S+MMKQ7rvNoN6+2aU
bGInDiu5lAiAcv1YZ7pWPGj6HImSllYuE/QRp2vQyeq+8CGn7CnGDMhc8H8vz/QxcZVgNDdLPmOq
UYwPxWXTfIFDmG5hDwBpgRfO357Dqp+EkJKYI12IUUHRfNTwFK/eRAfWCVrYA4GQUHLLUIrAD0Y0
aIW5G2sfwL+vNFVoioLJmrtphdaFrJJXzzjCA8l9KA4BFKuXZI1FMJfeslkQVWjvXsQjr5NFfC2B
aC3hzcjA3izkjrDq5oP4mcUJiEGjMDNFBZ9xkexhDKSbIgzviNv+tybnsnIoRacrZn83UsOKcmED
txbKkOjmnMfglyF1sKW1B16DvEjF7hUGT40B9nrDsSP5jwJqJEJX1ceSmukkZmRZivercaK7CsS+
UN844+IUcwK2ELk2GverakPWjT6SDI3PD7yJVfIC0CyuMCN817Oy/3WHN5786ZpXSK6/NoV2B12T
69AxSpiONfBiz9LAYcXGItykLHxi7vjT9+c/i6szV3VIkTsB3BsZKirSlZ3TJ2InVAKAJbHYFjsr
b4h8jfJqisy6prQrC5PcYeDOYwyB1l/6MFkIp/6qkF5Tzekwt9SRRCC/oaNsR9TbnNOakV2dHxMV
SvPqQKGk3HbM3D9OqeKAIabvPiiVM4M8R9ahf1YLTVD51ASknMjha4FnKfE+6kNfPPPwyo40xO51
a1OmqRa5MjBX4+sccQHohvb4hKl327aUhpXjg8O5M0Go9bvpGfvYWvq22tYegjm/05vcc3/hgJFw
5+sBaD+19uZhWi+y3B0Hg033i8OhqxJ4u8X0UMb33qcDyvXX6K9L440MIaybCBuxlB3CcCRqevhS
s+/bo0ZlKFnt3biRQy5U+yr9276na5GKkf5uNukNx5320GqVakb8zV4OJQ3d723dQHrVEIuPT50d
CA+680NF0tclIGsdhx8Gcm1/k2Yur1+DYKeBVBXMCeirxXPWk47MMd4PRjIJD+Qo07xAyunQRrvj
MKzNEzWHPeW7gC6EQyyRNQClSjAQN8aVQsmMKKNme7kC7U04PSnun4agEihYpTCOcm7I8UOBx7Wi
CNktVoC+WKWh+aWih2K65ieMjKaWsUptXsY1b5xzwT4wH2fW8oeo+CiaDzdALDbxYP598PWqFWSK
TvWoVmFlvQuwIJzZfXHzrInpJQymO+4LapWXHs8Qsh6JomnRa8E4HejC5/uTNXmb6h7fAJ9LARi4
LzMRod8P3KwyXsKwpDm50wNkhFGc/wSSECVEg7px9cG1E/fApV4WlQW9ICsbZOL9WG49lN0WeSvD
ELPWZOgDHl+Ex7r/G7okmAi9xXRtkQicOkNjg55K2RPviAEk0gctR//CNNsETOG0FnCMQdlKce9G
mfbCSPloXapw53iyTFYk5lq/oQ6+c0KbAqO8H5eDp3JDIzylsbU6EfaZvO3zr6uBUXM10QfPENtG
+sQAh9enokdqk7BW0HeMwbBH7S28R2X5kNae4MTqvlFX1qIPXr7teRXuN7MJ1Tj4F2JV92WzF+O8
m0J/1nKf6q/GxVfbQyCdRtviSUVTrg2RWcfNN8sNykUlgSF+UAUyRV5xQz4sKwpES9Behp2OzBBP
rheCAQHutvp70/NnUQ/bGN50qgtR9HAjyxe8qujT82rvr4o1zjBDxKDsGANQcOa/hovXcRJAUmLj
9FI2k+m82LPbFNZdN5YEeCe7bAwaS9asRLeDK0Pnw4Qp7oFnUg1BE+WXB4goY0NXVFp6E2O/n//L
G5nniNWMVstBcdFXyTukIIKCN/t1zfinjZ6YNO4BP4kJqrB1ji3hYgduYnO4UCKhcUhvbPmtMeer
HcYwwkJ3DzkrV21TrGFJCHZYQHjy5kxktzrP6p30n+e6yfM4oJYoZVJsWvECYthjvAK6h9BWHR2u
Oeug391Gy9i8iEhYfPpifKQkRiOZXoicGIyTQep4UvDgJSoH2WinRH42iqZ/GS8MjpBiSrGhpVY7
gho/qrdLBn86dZakmH9m2H1g+un2nX9Q+Z5Cb2q9wBD83cgJO3E8mOMZuk0r9n1rIM7ZIWmJClmF
N1L0YYbiFp8mZVNuyh6baVV/XMKdprnvE/ntCLs5xvjuy2R3B5u724OLdFrCuYpqioe92S5djSp4
TjoQU/KLTYCF3iMLJ8WmMXASm3et1/c/23/pdCx9af9QrJPt+tmGqO/yWPXen0dMo6ADfXtvNBFd
Q63NPWIUAf41aMW83bvTqrDMMzjI8i2/NIdpcEqW+lOm8Cv/gebcWGxgO/r9WOMbsEKrY/Q9eWlZ
1N/2+UUY8l9K3sTtUSMLCJPoXwkn5Hx9LCs/loWz6dJZobl4W0vClCdvzldwj9iZACOs4/uK4Ve3
ogeRa7XGgYtPdzy7nf7RfpxPYuk4OJlZnuR6PFRBcJaADwWteh+z+iEREy3Q3Pp8eF4s/d8coPIm
WtdZQUbim7hmgMr2H7Le/jNYINMVAjVSl+7d0Y3rDeh/O2d/NE9SPBELhWBh2lCo5hWfVyOQ5apd
cVjG6uwFD2LlNRs8yUThNaCanksr58jcpL/ZtogsAQxEIeZILmR3m063ZBQip8OWhMz9X80hRJ2t
6ZgwP5ie/dnVjk9IPHU0iuOMj/zSelf3vEPAygJVEww9V7nnWF4f1kKh5K1czadzgsEYFIeS7BFM
TIMBaLyU5QaWvLjNgioJckhL7bllK12sd170M8myyBa2Yc9FR62lSkYgglHd1Wc0Sz/nM09aqaqR
2iwGx1Yh0UL5x89sOwGCd2/8IqVlj9BNNjXq38O/eSGG5XO7xyOhzYV26CSaeqqj98U6g5OTJirX
8wgxx8WJlDRlMfigtV5xwEAbcjQwyBAg4NlAJTxgEGQ6swmYuIeU216D6ZlTD0+KCLfdwCiLQuJY
6VxLZjk4YnkjHsadX9wncv/KjL7eCvh+8edEfDeiuUgBz4IQcxVFXfUu30bgLNkeVXMZLoAsaqgM
i6t0fGd1xbfSC3l5EaidvoCB8BXsHmfMCEkLfFCAoUS66iwYCjAQYeZuX/RRHUTEAFnTAJvYWEOJ
1QwAtiFs6vk9IZ0u3Yli7ofRtQ39kzqNSEpxxqt4hK4XlibSzpecD3BQsAPfW58pYzZla5cCyM+M
wM/C+VlAjX4Nkhqnh0alzQAx9Wvws5dh7MWcwEZ1kAM5RI/9mlgxjTzbAygf0Cy3dYjXam1PJvpm
FC2AqWVTRIdk9TGQMvfsL/CyRB1p4Cds+sewCiX2k4EoXRKVJRBM8COHjNnZF62BT9d4gXoa7RVI
MkYUhtqHCV5NQIvE2bI5gc7AqJb/RriWrBjTZTal/1GOvzTXbGGgtvOxECFISHeS2PXzrgvVZL25
q4C4Yuka2x/FcKa4/ilsfCaNQcEenwluqGfSMxffUHmO8VFD4hMkUIdXKleets3MVO3476OijdAf
CTQXqE+FjgQDb5RpZRM60MSoSOqTV+3cudlntycYZxLTiaciHCCMl5IkZdsrWAp62917U10gmHVC
0fqIVsWfSW7qfS73ks9pyF6O6Uh9yK1G5FnRYdHIwzDlA0SzZ+JQADO8NKkEVHdEkYqTtKNlpJt6
KK+kidL+sUGlCy9QkDYHByxeNEXO4wFY/rlCiQUUNy8Lx+MZrSwUIKiapW/865LzCqnlxLFDlBQT
xSF1c4PY+OyfzJtojN4KXoWqwp1qWk7aO1P6S4BaqDJPySyhx1HWg6769xagfGr703LZh1qDXKcj
FIsFqGpwdl/tDZvXTklvVruDpOwCMWVH57quMmK9Fw4ExadDg85XRRk9X10smSsbRazQow1zluTA
DBgt4Qjx1Diji9L5xD0OBWoZMZBwRcHghX124gQElF/7lXeWcsXhYOdTm6ejMA/hFhdWh5NhT5lB
ppiq9i0sDLy9D5HKWY3tauPOOVzuzbKSY3NJNABJIDe18WCkRCjn4d3p9EjtS4RmmtRa3V6UL1pf
jCMAZSka6JIY3euUFr4TNB3Vcso5DNhf+UUReJEVSymA8pZLTW62vCPFP4GC2o2LA38p9xeEo4kL
heDOJegjwMEM3dyX6FhZ+5ltynfaBbKBnSPFIMYq6g2cUYxcGlBinl5QbjDIpQsxv8ys6D1+Qiix
qTXQImDNIOzCgNiC2UmNdtQ5/n5JOvvaYyDG5THIIgoqt3CSmhAWrUeQM3Pv4EsQgU+7wMjashd0
ZRHXC8rSLpAvnkhttwqw3oSqXtjD6ePZ94yUoC8nmQwKTYep3bKJ6sfEf6OgeTvI2NvgA5vtt0DI
lWhrYJQjwjNH8nZa18LRqkqKxoJPoXqEHlO/Ex4zyFtH8vWHjp/F5Ol/dwcgRGdlg7nXfh8hrJdU
r4rQje3cmW1ppz8xuOf82VWmIzO/JRe0wykVyNUW7nQy4ZqFWDtO/k/C4//gbOjTZr/VbeGP3DrL
hMte0fWZIA6AyZFpeeZ+EuttkQz46wXnoeaSDwHr1Q8CjxYsbz6w2nOA9nAZL9FohllZ8K6s2pc/
RlsUFqrSq8tvKhmrLtau48g8fLGKzMJQ0edrF8QOIgy+Clb9+C4x3bV70oZ5LQN8XPebkHabeqvf
eLfKCJcny1Q3B5goDac5NAvH1p/57sWUjBr4LEVJtn98nhdOAw+KcSwaIEXRnNGzeZMjnI8HWmyf
//isreB8NaF6lovMiWJYWrgffy82q37HIND1FfUDVIe5lAXWx9kNvp/ZyKMbJOZlsRd2/DU4e/Fj
+Nry6p2ZLh01WCSx5TGtOq1xmtWmytAddA6fmMdjN2OXNC8J74HRph3DsquBSZIc3KyXqWCmU9oV
A0RF922S7CLLaOzgcMnAg2thIfRywLVMywaYRTlSDnj9P7ZSr543j0OprD4e6vTm4Cgj6bvAiFiz
RL3L0W/evXdw/p/rqrlSyg6dHrkuEORwUBgbQCltvcsiT7o3e8/IvAtbdrNprTQokCU9Z6RebF+P
ErUxTTztvW+hGFliuKmbRW8wCbFsnQCVl1kY3w7UAOPkiW0klwcpVyx4qXgDjNzGSIvgyaC68WQ8
nChbQQ+C+FyZAB6g6GGnAbP4lrq0kdO9an5SiQOdsogHGhwuwyqFLCkQt08Eb5TOoPxHviz3Q5FL
1880txXWmBVkApodefcD1SY47mk19WVtlLFDoZ+92g0e13BXzpcrpP5IGQDTHBMWFETzusYJzsmb
kYjHjnb4wBd77wk5YHuCb5KxtQpJvjSwepbqwx/bz5/Xlkt9AQ6EkiW8DfMfyDBg2yGazw2DxrAM
z1lXf6YFbqRpQSzOxt6DadZoxjXJ1jtK68VXbiEZDNJCNKU0LmFKu1aXcfEbgXinGkeMB+L6Jps7
BX8iAhwwr2vv45sN5whCCh3h4eAd9slJWFCPnMAcKKXoEqkI0S3BryR52xJkUB5b6XAVxpiPQZ0K
8jQ+uVfopQ3OosisUd4O7L376W3OWips2/mZzpnShH2q8hNuR3KIw++gCPpfBxUlwdPiJcDCOqcS
zQ6fSQ/T9LlkTd8uFT+0rfmtMzQZbhnj35G5Sk7XHBf15EKAO6lOyCIfdsmNw9RJ8Klo14+bLtut
43zHyu3oaHse7rV3o2V/aQi0AAf44SR962XGWkKmm2VzXlzBvHoU5LJrV7vWrVL+6CmX6AXFOmr7
RA+185Hc3/KA9NUUeYqhB+a/pgA26fQH6RobY7z1BN1aZvGibZuSO9HbWTSuI9pOTojpmq67QuM3
NKVKuyBKdAQkAYLCtmiItkQrWPuZe396LQQL7I3ZbOm9dGSoMu+wxPom/53SeslAC/917RCgZ3t3
na9EdybealWEucs2Ao33SMb5M6DfwXDyLNg3ncKplJZx/3XREExQ9iX4aFU7elEcCmZv9yFDo33K
iOYxDkYQuqZ1ZZbxUDllBbxZTNSlGcFkdnOaQ4w0PKLJq6dAC1cx0Gyz+iZtWJBgUo/jS9NLczG2
busme9DLmeB8NChlEnXZSj8d+4eXOtrmVHFkt++Gdxw0+2gF4/lk2xSa2inx6a1rMybwcqbfGN6g
8QI2bM59sc7toc94kN+TdcA5tCUlsoQPcKZyHAwVppGk7RD2XHqiysteygQPBuTGzFOgrG6fq0Ag
uRRumJ0d8o5/hhWkQIfOdS5+A+Q0H8G/vIk6QDSdsuik5ZLzLKM1jADryJeOqARMtBAR68+Z+0vz
hjrWHoFscwjA0+2BOTsHNa7ZDaSV9I4K57TLkq1SEl88xXK3kvEAbUUlmuuuHbojlV8XCanfxN4u
DCEWXS7Iyl1Mbj8TFReOmwlsOGmkLIQa5vZBTQC0iGjeh6u0ebdVXiDb8Lnr647oYrDjLPzASXxy
iVtE3UozexqI1JqMDPVlBrlsQ9Ugt0vH9Ah5Q1r7TWiYPHNU1tjiz1I3D0ZIOppegKz0w5OiQMe8
D0mtxYBGnGdTKoYIBljUW3CB/hoMYXOiOrMPRdA7mgGh5hNM9Ilu/qc3OVFcuPTcOdkJcM9EYGd/
Sm1fEYGjh0zeXpQbkX/lE0Ea1tGPOAx7SugOW+BUdXk3l73RgJ3sbt6+d9IL4JTYmUbrQ/vy4t2g
uasLXAFsrzPWvQzHLSnq/6vA15DlhY2T5Dy1mjOa2BMSrYzv+cZY1YZZTm8y6aS1d7ln1DL4CtdF
oD8QWAV5ujekbSq/w9LS1Uk2X0z+fQbfEutlZBWxqVCf1qJKZ3T3nSASqOqxNT2GgpKW11d17Cba
EWzGkjDB0J5FR+xPmQ6SyckC/EtAkdtKW/UbLOg45O9R0WFqTDqCoPrm+30EGuWETbGDXp+WR0b8
4sx7yawIqi8ESoUErdqak/oP8PANRcRE6M1SuV1mhaPHAHz6M0diVpnxrEs3iAJYf8973iHjKuS4
NLZKZ4vQRH+vE3IfWyw4gMuEV2wPj0ttoZvtY2ceuUgayWYuuNkUtX6Joiw9dqvfcatL5MTzYD9h
LFy+5ZMlkt4Dl0lKyATpQFCc+ey3OLM3kKppDWDiakJ3fXzi5vmai2Et7LBnms3uxGq7zhx0mPGn
T/PFuymXZ/q1RaBik8WvJ3zftQ8BMYcmTt9lAJjWO1vMESyADuijCzHIA+Ap807y6PAXDeko1uIv
7dcD7QaXyNJF7cDY8YE/VgKVc+PFZPawaBN9S6InnC1ZCKKTNf0Ohbe+H0pnKC+r0sBfpRReR2pM
JHeJZeTEtdTdNkJtdFIHVAi//9JZpdTnDhdHuvMI824vc7NONDO0q27LcdrOLkoN4T1THrDJiQoA
z9OfOTY0YIz3RKxagm0k3wmHjbu0nXCzXClY6Bf1+7jstiAevsbu0brfQpULfDAX+JN0+MwwlvJi
RFth8RZbmWFCm70I8XZSJBnsm2Zp/eSsdwVRPtajR/+H62RTFRxTgHw6gFAwn9fiFxajiuYfcMIX
/GALCUw8yx0+FaItSZCwMSgjKBwb/+JsNDsqxK78Chr9C6Rqapi06hQbPBOJufVjs9zhofDhHhaA
KoMqXPiwxdOLGknbHjFStuuV2CJguH1hzIOQH6esxmh8VfxKMbPkgcxPa+ac++4ZMvjz/Bss2QnZ
EfYC8m56JlvSwVtYyh+8mRtl9GoPwrOeQlMaPSuTu+PQJB3NrrTOjdV2RNR/9tZpWogJcrCyio6u
qSrnJOZrBsvQ1XD5FPdZoXKIthaJFaqgAT5QCxUv6shyFEqoFG5tLoknYRQUo0j0JEKnd2uX0/iU
njFjzR3aAgWAe191rU3V83q5Mnby5YA8HKvUdYI0gvcn4ZZvGPTqMq5J5oda3fIBIpTpVBcbzfqD
T2tzsMw/Gl5h9ey6mkra395Drw14v9ldhHvIdiNKsogBv9GTM9POmrHyVAAQW8ttf5ibmcP3GeAe
Uhjq6rHFMXu0AI+zDOwjqprasy0yXENuM6aWFKmlhwau2eZKgEyXoRL168R80V2ziFwCGsVw+2ZM
C6ry38we/hzsvXjnkOaXwirkVu2GwQ+oSDIhgIaYvXFikorFnYrYMTQrN9Oueqbfo1kfrXQpNLOm
P5VT236+JyrtN7s7nMxYJAD3bh1h/p6r9bWTankAmTLyvDLrl6FkkbbsVXwoPMkZnGGptuzg21ND
MxROYNc+iaW0B/8qzIdlmHB/9vE0+6wq7EEk3oAvsWhQAKki10hyzwBfHZVQ1RhajE1UU4QfN1Xf
GCEJzZGALlKXuhUU7Fh6Yr5vZ2qAbHgiDkr8AC1MRtU3kDQRMdIHMWV8u6f+xr/II1J+B8QJU4Gn
Hrp5yaHiZsbzRrnz4V3LDBifJf75+ExaFsLTs/E3o2CICz9TOV5cHiNsWnrW3ygx/oMZUafImm3/
JTW/ON4OY9ZsxXvKnpA3u0OhaNdc/khJnHz1zHsV9mVUY3zbr7rEgzuNC8FNXLKhgqOtH/Tik5lF
6AWZs6FomXCgin2CsTT/P7VA5B4KEP70S4h0eHXJ6gE2Ux2X8UwmmITFzsste4j7jH0TbeiVTuPk
DubXyGDqWMv70/PKScnEURp2+8CObeZmsuvxK6VM09nefZ719jp2iU2QG39rWm6UtSvtwAV1cJFg
QayL3v/bc6XMy6zQ5suge1LVwxZUqp6b4P2kY62HRyB2TxuCwysNiFNhPpsh0kYuvv+o0iZcfrC2
tDkeDH2cyjld/AeYEsP8So1q1+6oVWtX5JMEkRMFsqRULvtatEmG1lhyj1CTONq6OweWTz9OBtxF
/jaW37T4AKNwIfyvch7Iyh2QljhtJxsegXolzjo5OpO9N8a6Ybk8MST2fPgvgiZJcP/JC3pVgnPH
FA7U4s9R7l6lYEVuw+t60ZnmuvAPer2BlMvtxEMbvgKqgtwyt8+nMJw582YmDD+n2z+DmRofdm07
hHFmnwTLw5dDeTmeaST4NQDuodzlc5iX+awAuOImId26c2hcJ30I6dFcHrXWIJTSFn1uYCqwNPsv
a6+YlANaW75CT01PfGWnIKtEaFTChTE6k6OXGLpzUX75Ybp9xxksr+0SBP2rADSyurU2BWR/UGGc
MKZwHDgwc2AWcZxIFN2HH6v4FhFQdxQskhkTX0bAfjtH9sY2F6B2f/7BlNeIcdsywnZz+y2f4bwi
ykgbFedW61gX5cYveQ0fe5sZifYYqOjwdPWdOSFmYa3VIHxJNQYfxmPiGnYyFU5801i119QzFJtH
PlRV8MSa1ClrxzE6KT3zxdXiSUjBDI9y/IM9TasZFTu8yAZOd+1YmMDroHSZV0EMD2LRlZWd77Qv
sfYYg59miYHk+O7spuGWZLfbzOKgJ38OcH61l/iPFu2dlZmlC/84+frWGySNwec0/mGesB8DWURd
4oTw7PFktnEi3Fp43Kyf7TZutmZSkTO3IWZmgVYZU4VPDmPRTvawhuINUCo6tev3elczfwT+2ShX
BblQyhEJlurOR/hPVEUtR+2ZIBEUObmrHyJZXm1uzFoIUrQ2vwuxIjCerdjLd7IBlxS7Wono3Jv8
Kd2pFrt3PVQ2cUlOJozp+3ReSy4rstit1I8yBWm26KXHuBXtWuGVZff55RrrW5+y6mAHrXnhLwbo
qLy8CxOYEg+WoLGR0V9zT7O2Lnx7PEwSY4dTkDMlBNzwUhlvJDSYf313j88pxKDjyXIV3tmozDFI
miuzkY36fmKKeKvphtbeIUmNzqOoDNWhVCyd1V3ga+Brz0P2fT9heydyS6imY7y8wtcEVpiA3/JZ
qYOt7Ww0/FdIQAsIjCWMBEROd+qdB/hANpzz1+JHZunZ934UziRhp+jYg9OUMIir6gcQM823fovT
gx5PhUa1Ma4cr7XsbCa9VzRrEEE5cmVm1wzLwrHYFSh+eoQfwPdP+bSaqdZbdh+Fr4ZYOeOFNEQb
Qx625poLu8HnwzVbL+7jwK8WiV0VowiICjirl6eV+0LCaYEhj1VHp9AxOKO0tJfGpZGkO4N8RhN7
RsKtW2wo14tpsNg1zbpDqeBR2KG8pS6ze2nU4aXcKmOE5ucu2e9Szi1Zt5sMhYjGCAgh4GM07OsR
vtzvLTHo+84kRRtuN3inWnBvy9DzuqTc5k/kL5saiUUk/N2nY95Oudll69viXDBW4Ew7OAsnmk9S
G8SKvuAlChY524pssluhYGHR0NnDbkbsTyOLddasgPpuaSsfHzES21YxfDPjANW8R3zc3cI8FYAL
BhQ2kYp28vFX1oEQKAvI7Y1THo8ckQIudZbyzz8sV8olKCLsu0k6V3gjshTu0QgdfnqwDVVviPA2
YHNR8Ss6oNpKbTkQB4hiV57RUurWybCpT/eKGcrpWbvPhTIxaE8lE0ZWJNdtdKvCUuvEZ5+/3e1o
IJIQ3wFBJKMmxsEOfH9+NbgAFYtocgJhd49xn/C/8kCSNpekOz92urNOZGOHuuZiFW8WeNeJjUzf
9Mm+Z9InGKtgQ78jEggGAeaDMeqNSPFiS6iuoKDxfPv1AKkhJ3W8KXeoT821UZNQXWc1gbzyLMvx
UthKb6ye0R3wlg0ioGnCa8fMZ2VyjAYbZN01EUI5yyO8/R7NV9HAMoKkwh3yHaDbEYvjcV4Loqc7
NN96m+Q6Qhq4wVOaPWiT16RRFLwlhaqAg32jORtj2WWHfl9jt0PCpWwY4lNZwOa7Nou0j0jEUmc2
2XGJXJCajS3IkWeLMAhKsaWMa2rHiJnSrGo44KRbrPfPfFcPsvK1fbcsaqedHNQnDkCDq//86Cli
SJog4GQBnNQ5ORLm1vjpom8m8RbmTLXXm+Zrd7JsMdEnTue7Z52YlPCKp2wYSV8ZvaF/cY0jHEs0
ajOBwxmh5vc8/WuA/O/p7SQ8C1uQKJ20UQeDEbgJH5ggOFv6LEP7BvRH1hHfRSm7oE5ACQU0uXFJ
1s1R/vRKuXQ2tBOt3JFltonidPMRubHbtR1SwRapEuEN4An/AhjC/zlfR0LQdBjvoV76afxdJgaS
rf/DYd0T7RUn0ZABd7zDPVY66+tg6pK4mFAW3fzisUIcLVjU76sPXF0ZhCWlda+jjw8CRFDYxADP
9aRNmFALK5TdhR062PaYnNlvN7rqZnOOgW+mA0XlOzYkrmUaiZlIo5a/nRkPbFgmIMQ7XkNUcwf3
L3B8na/8ZmBujZ/PMkn5Oq/UeCZnXNPbGtEWjIqaTFx9G35jaWPmOW00mg2b1kxdWfnS2o4YLuX4
03A9lNd0fjDOkrdFW/zxIDHvtQDGeyZcJkyOQCsf13HB4eEq2ekn2U9pr1f8d2q2CDcMSkLs9HPd
brD//LakhS08rVdpwrJAWXyv3NDaIW23LWa8A8EaGqdCTAsyCmKIUvSIRpnmr3z+VCS971g5lYp7
1IAHRDozorECrNUDSjKp2LG/oGLSPd8CW33Xijovbj/ZuHY1hMeSzIm485istuS27yzG8BJd4jFl
3ITmh7jAk7e0NptAT0neTEE+3GPsU+ehR05yPf8tNLx3PXVx/8vmsRWm+eeiF1p56JgEX34NeMAk
40VU/wOc0Fq3kYDHJzclG6k0zaXhwiovvQNZ1H7bHexziJU4WGrRtIfUWj09mKginZ7ZT5EUYjy5
xs7ZcHEoKvAGxlJnBFU7iLMxLnIfFTnD6RL7YrMLu/dzvyI7FQKykaM5/5QNM/BBLW6qBGDW9rQ6
cKnjqbJObZMjxFgsIJKhIMGekOZKFlIMaXUSvIvd4I2kPMCAFNq1b686+48m+TP4ABmSjecfjKqs
2iORt/3b+acSHTB4nS50VePdmMG9z9AUdxFEfNIyRL9rLa6ErOAtqvit74mqe3OJ3MenSHRzBlAt
xPc2kXaCALE5GPsJ3jmUO09o9qcLMsMiMeg6418F3PP93gX51zvrbXvsP3UYuZdkJ4wPGGdeIkrz
0SQoZwvMVKivhcZSq+QLSRQsKkqW6hc61FhxAlE11+20QUqt/iKhKjrXhFQWDP8doFUtJMj6WWEA
X8M/Xaziy032VIl8689COB6PfMocVCBpNPiUbGwQsBSFTx21FZJ8QR4yebXCRIo3ZvJHjZM8HAHM
8IGstZasi0jYYG1/I3TwDMT7cZ5Owmg0Rl/+9A5h3W8B+41Cx8Ab/MRV5qStO2VmBCMjNaEKKX1a
fxIhI+Q2tLgumQrXyeJpvbcx2Ku9Z7Uj8zv/tN8FkNxKbxONeiMHB1fNqMRctNzd7Ilb/LFVTzZF
JretmkR1iUlUHT7njnlaFlGhKia4AfE45BshbJTpzPOyElyj2vTqDl60rOb/MRtsrQR+NAR0Oard
cXeFWSq/KfNvl/XKH9k5a4VKmqHPkITUe8bLFKk8maSsRDqDixSoppZ5FEd9Jm6efL1JWJV0dceJ
R4xT6cJf023YdXpvTVzFwCTKEyRQuOfuhQrxrnT5ERi/wOl6FmzG0mJs0+lyDC/+AG3WmeKp/y8Q
GiBMSKHseJ8kicJggoGSzR+e9c4jikMY1jtquRoXr4ziSpG28Iieok0BcWTjDXKxm3DZh3ieGQ7U
RS1JoL3kyuT4zD1E4crGpmN5hw4I1VCCsYYnjkpzIRaGb87HCpaPP1sfBdellRrlnu/V7xBj0bzV
XVuLWQrV2STZ/+Dpqdv3ymp27iLY09pJxz25n6gTO4G01O0TDLQ0yQsqsDo7CJc2TCQXFbdD8Nbh
2+otHcKiLdVj+6//N47ipMxtqYu4jyiSJfFoiBzxw9VUhuD6BfpnCgQl1havKUsXZU11NFpTclob
+KqT4Th3AXAkogKDl6vgFHbPi4AeLUFK1o0o13YLC9ddIacaQ7FLLyDvW0TpoU/i4zRwWA/po65p
elzoRmwfbeI3n7N75Ta/JXfegoylpuh4XXUqnL6HheW2PL6Jhko+PmCA1P9vFeUJqUGFNBO/c18R
5we1cCIUKY1uMRzEGQdGs3P5/x/e5gmPypySO2xHPCIiun5f6qLZoRWr+CNYQ7yYEK6tm9fqpObq
vR3dya4A6pbHhFCQ49mP8v0lg1C0XiO3bYFMtyqe+qdPGAtvaeoj/ENFAhmnvsJhaBDs9f0yGNwl
JGuGso5ngTgbEqgZA96jzHMajTrtBgjt8Zzo5cRfW6cSgo0lzajIs2yREOb50ysZDWEx1TpiULGf
475IjN/DRNyk3Vy82CceJeAGdtjNQgUD2c3saJn1IE+UwwGucPxNe3pDVko/ehi9cVvLrj+gxsS7
n3sMhqtq3W4JndWw1JOaoFDnlGetsdz4NUWBCezUgijLOX6SMj8zoeENIvmCMiGY+aEzc3yF1G+7
d+f7vBFAkOuBKQWQ0sfLVNqAsF3Aixy7O+yD2uZaIkxQ05stIcy1WIWY3RsreZH2MFsx/TBxcbbH
/EFw4GjCiPnLa14jQUWwTUU0XVyArizbb8iUKgQvKPpq4tbSV7e4Y1dK+1eo7sFuSbrjghhg5dNg
VV0l5E2uoi2sD2gLD+XIADB+dYoPYyBKGBQchW122q3bZGbON6IJi5D/5sc7TG3nkEyn7szAmkYi
P/WOaGD0Bmvgk+I3RqQ+5F3OwZk7BMud/w1SE7Mm0LYLhXizc4QrVgse3+Jyfiebgi9MZV775uIH
7TSNknnqhkpjpGv6g93DU5aAQqxurCEf/VzP+vkA3DG/1OemvD8ZvtCA07DKg7yeNEfGcRQeP+4z
Eh/MXct7+DT5ncvci4Ii5dj4ywNnsBrUDiqF00b9HQfiUV6LZrtYnDNCcHVTKPXwBO2wLnyyMVPj
zR17CTOASwvRmEVIHrLZ5k9kp8r9mL4vZN0JAofmpMG+wvdqi6N5Cj5Ovm2F5IkvVyOrkJr5jDe3
dAQcKWDENFI6PYczqTiCfxeE1d9A1WKNWpvN8CcGgEa1etpDDe6+CeUWlggkJL5m8wOUR0kDs3eM
1c2+5WvWLAXz3aVh0ZDCg3RR4zkpyz4bkt2zZVXVk+7CvlpyWpvROjS1xWPcqKxxQ5+pYHEuKKO+
RuDh6zDoI5/MZuHFa5qc/J52kCkaRjIDFik2jdEvd0q06QWKQOV293Po+RrXjKtKzWGnst/bqZ6p
mcZeprncEePXE9cCAQe5t2hxG6uIpyK2DCnnSaxZGi6yF/S3CcZ6d9WmxRWGjLujZsXEjdWvWNkR
dLfvGKtqtdA5ZkU0aEQr3HaCZ0q2ddjkwFju4ZkqT8JLmX3vzjbd5ZlaOKMVdDzxWYPxvI4rSeAi
A90JwdcP/oNyfN2wy2GmWJTyE8HqseZ7gyKNhISFQQKa2Zhi28bouvNB+iihVa8XlrbtKiG1mk1B
51GX7sxIiYbt1TeSLZCzAEjyJspvqZKlYr/802Ad6X2TZelgzkPCJLqMUntsN3rtOuTvldK+jt+0
mPnOJSUuqj4wNNeV9QanLPiSty0CtD8T6C0Bt1QfVR8TThtUa/My0FawwWtu8xJgu6P8Adf5yO2N
DXAUNY8Q9dEOfhyttNl3tu33iF20xQpneSAsufGg1jgAMbuigRhxmzGAb9YD6cyTHFnItig2bivT
j60n8+/R7wQjr36nAF6jtwNcXqeG2lBwCYbxV39YfXGBxUdoaA4olI07LJUGiW5ttzaTRpbuz7Is
X6tBU9FnTf8RO3wCnc4zINjOdoxwa2Wm1vyzhCahysQXYZ1nORci9Lckz5OeH5jvyyENElrKr5bL
yEi43K4eBdXECCdpHCWb96LiGw4rWZZQhczw7YHxkI/w9DGMoOfbb1Z4lh6nb+sM5nzDP9Rss/Sn
EBXDYjrIy0y6gG2FJ0LPywIkD3Q/6RPlINDj3UVakue+CRpnt9wvCI6lTGIVYb5k68FSka/wyYhf
iK7/5Gks7APpRLusExNH4Z1CtH0fZsfmHeM08kP3nQrLPDTiTbMTX624iCzhg+YBPDcQRlT41ZoH
GclxyuR/b4id20+Oi6AVSMT4oDPgcrY/Xybw+0uq1BA1EGPBSqYwKLaEKeLgAfXAI48Mq53bHNXN
ZmR/F2oQohYSj2yb/SO2WG4Zh8ZhpdTJ53SP22jhypR22ohh9qIzXN+sml9KTZTjkULhf0ZYHdPj
OloFRNrPPOXmtqOnqwxkX/2R+HwmK/8zKrqv4biklHG8IUk7KXRnu5d4OD+SDTbkxk+ZZ8/512JO
UBsDNHdU4JgJNmYQy0pYEDzR7Wbsnb1pU5iMxxV1HOoZ1/SF30IPlZGxGT3Ek+D8m+jREoFLtvCo
mIPNh5jSp1ZG0x7teQfoKEbgXfiYFVEytLaq9xIsxhF2TuiJgeig4U/aMUIYlhtvrdL+VGwKdtmO
cP9UTFhh5j46lj4zsHNgyTeohe9DuPDfHk5HUnl0F9ZU7umpQj9GqKZYQYuVoCdN02NxjTVtpjvg
SjTKWZKiWcGsoPK6ZywX54tUafHzgIH/AAhMZdWAJaFNQnKLbwtAFalaIW0PGPPrpj8cKBRC+CAc
4TmGs9J4l3+xgoGEgzYxiG+uLnQE0LQrBSLQ5XwcTQ4lYEUTd5sR8Kb4X+wL8KXIqlk2sKV7f3lD
oscw5Eckef2FhMvI8FjhirwRay7Nu67V1GmdH/K3PkGNDIbBQ0sTjlGbtD+gmt2001MEOS/SiZWi
4MR92mkvxEIZ0tRJrMqWE9qE+T/SDnb6TmjlpW/MWgEGaoQfJvQfqa9fYKBUtzR6NnnXG7olnEyX
bE0zDoOZeEHFmC5TMRXLtFPWzqNFrexY1SCs0eSLHUROFkuC9hKQFWLwmINKWxVrtQL6TlVoNGXr
B0ncFBfBD4E/1h+4N4SAKAq/a2JFxjLxB8NHI5KK5Kuj3ZmDvPfB4iTw4cgBfeGOdOctYVmjdICk
w40zX7pmToumGA5QEvnjkOK2vEheKpiPfQMiRBP6x4RknnkkqwARqsCIgg6Izwb4eW8s7F/7ZuoL
TDz5s+pHCTQSBHEUhiHVWkJx//XwszgzMxXZxv/O/m3PsZVH+coMUGXRlxM0cMHgIWicVKMRrPAr
ULmVxJHuZL9O/PmTeaHr7ipYZ/55c3Jdd8CBU01ClaOwQJf1UquCKYtJmbBxbr8m9kHi0ADKVo7C
Supaj273yhoLaTD4UISsbHirDd++9Mxb8OTW41Dp3yppRuhTbO0Q9/0bVMqM+QgdIddSQQly2WEh
4WW6ZIV1o1456Ni0u+xfzQsBTDWiOcrkekwmIj+giaIMns1yrDH2No0d0XoLjC/IvtCNPBE3rKRI
5DiK3ykZLu9JP/g+iWEhRp2qFvGzC/Jkv67PHhsnLAQ+TJd60H8l4gHIgZe4wyu6KZWZt6HvrI+0
4gewhYODR/YtaM4rLx82ykixzikY2FI7Yow0xnKH05dNfeo2e4+Yy/MOdqcitxkFgt2jlo9c0Cwn
r7ZD/LmCXKrRycMrrOe5iv1uGwXo3j9hIEd0lVpP2A7tIgBP9Cy9TJELowhk44bks6YcXbqUicEW
u2iTqOCxuIvm+PFcsKjo+Klq+J/lXI9FZkElfFCY61ppgly7zvw213calwJJfkr80rFPHBoD/+yS
kd0wGh9nMlSaGed+NbxvwRfOtvjXr+/yeYmvVRhrX1MDLLWcIHWtyP7T5qhH6VwsBSgwc3sJPa+K
63+VtgUfYx4Tzh1B93DIZedx6gnlO9jAHDsK22f2vmzYx/FDHIMvZb1m6VUEt2PPWa6CkRBHl6at
mNgWYSP5w4jQK4dSNTJxAipjw1fQCDTPmF04KMYxz11Egm6CloKVNxfN09fqXMrqXqF6sDvpfxux
7BnMW33iQH7oTUYXuJIKkcI0pMTHcIyPHxRthpPaMJMM/epu44JCM95HVe49h431XScRP/8bEiXO
IjrqeuOWEpWqW1GvaMai6yxHk3X9FhSeVR/nbtVnQXhBR7245n/l3+5YucVToFbx50MImxV0QP34
wqLEwes1MMWfqO7EZR5NfBX8RrvEMHxYPP2BCzOTYJGGFJOIXfY5zVYEcpbBlccq+mdUAxqVO8b3
7P8oDS+smYkxfpoiKgI9QrkSa8YXvcQ22ON+vbc7KWKa4jLe8HEwnLf8UYRuO2pGncZkYmXPlOPm
Mgk67gPtCitZNY6weUxPyA/NduSI43ApbE+O8i+4NGyKURy9soOCpcxM9BIYGfcACDUHRhEZ6xGw
d7pg9kniBM0UKS8E++FD5NzryaDiERq/9T8RI5wXVcOhuwerubLI+94dGdeOI5lqfOyEmkWav5PM
M0VOPbH+tF+lMEM4j96wVZxakppAksOwKXmIR2dnwGoB16lQ6+IfX5NE1RdZ3HZXtT+8qT7Lf16v
jrqYd8t921f4koz4rUdjPULxPLEnEG5TRG/BfdxdAu5Tvfo7/RIlVyLt+c+BueiZksjTW5ahZBD0
S/mMv/qXDCXXWlyNtTQ/uidjLEKMNEbOXj79MpAfcZ99iBc+5PWuFm+eb+e+Nupv8G1ZEA8ftWx8
rhgFaqgqikJr+ReQcGZWUCR3VJCmuKsfsMfHsP1A5J3u/XgUVOcPODOx66N4qIxeZJkWu/8kUqKG
Iu0ZJFhqV9hF0KISM8oMK2J4R2gg3xxChFlmpjwW2OJloydv3DavuCvgf0SMq13kKQau168GMWW1
oiNi4mzZfjs0lgW2Iq9l65qSOi7M/mv8k9dFmfio21Fbtdllq/DXmrwYvPZV0j7joT8odj/3ao56
I+yp8b91GyJQZ/nUrd83En8jeGDr5iAQoF8emtUUkLrUYCUMeO/HWci2sOE730gVq5xIXtO6a7KR
P4fYjGIzm/4naY9bBw/zU8wrBD1mcINIi+yoWQuVFfDIGKoWshCvcQEC++fp24RRUZFxAj64CcAZ
kHfUv39F8F/lMGB/y1c4s1Huq8/pPVniRq8/NRAzLRELRXBW1+2H8pdHpELJiwK3CaSQChlw+RYL
dykdYvTQJXiCMoxFycxbl/TRTC+BZFpIxt46gztSnBD4nDCMGHmRSwQOlBrKkb/HOHxZo8B8kv6J
KV24bsOy/0kgS+Prtzm8HAF1gzY+caRCqGFtZ/zo3ViZIqb6KL8J6sAuY/zW4KgK2ecJMZ7U/Qca
vAF91iWAfW+L26kEkLXUpnJgc0oYvR6HVuluE8cj0eak4D4ShUFoWP4gWb1GxfzymvaQiGHvPKWx
Ywp5RM44uLoAP8hMEWXXFkKByGnjTEbRdf64UmhKvYG4FtKhmcJwMopwbfR7ZgrA8SQS1kFalt0H
cqMRzgim3LPxjARSSRVQQAc1v5mpmiCQ4tcYZhSDX9cWMzUKxtuI1MmyafNJYpdzmbLTbzVJmwZl
c8FUIrW9Gg8I9KtSPWgJftVWERqwAXMQaSETzNwi4xUGUAWIYkco/feXVDBITDHbAKBmhRevUQE8
GFAUL80PrkBbmlwdPytX/LpARsc1FcoDFPYFemAtX/CqFDyBMkUt5HyLHxHmfNrQMYrvB3YUq4dX
wSYpGwwpy4w7h4RMU1Kpv1NJD2onK+QrtAr6LD4im/m4vFtLZ1rw0Opcb1hqiVss1mdMu5oSkiBv
IAI5+0JFU9I5cras+8GldZKa1c7yX2S3xYfETSXZD6iL92ohMmbTs/rUruIRlE+slFky8irf8PtR
yjyS9BoezUJyIhx6zs/bYqyBQbQCw7iMEir+pyeiIb/1EaKP4aoZV9ZL0dO0QbRch66YOkj8xiaq
xfIo76QtMEbHaJvcp1wMTijh8LFTJe8/GtX0w0gHrjbxDXadKGbVKrknIvCajj+4mKZPzAvMXBpV
YOU100HLynk4DErBcjr+hV6kXDA4STVaYS/m3/sDKxVGX8MYnx75s3bx5C9ZrSXPIquI+jbSSvwi
BTV8wv3COm6BPXL2oi5D3MQOJhGh7sgvt8meueyhY3XU17VQDefy6bSNLz+1RHn8JmM3MYPorC86
IQtEi0AU8MKzX00sGu76Pn7wP/x0oaeY0t4q94biGYPg28TqwlfX+oahUJIwzQd7CBhvzweiojJ6
R2R2r85X/A8VcQmroHRWH1mGN8FUPt3MyyQIsFYIO4jyrVLT84+Y9O9tZJEq7hfplCtOV9DNIKFf
iUgK5Y9VeOblUrYAd+hoqKl5DaouiLZvYW1XzX0MUJw+Z0EskiwRy9nIpt+zF1frR3Vt9Ugkx46l
5y4NNpF+8golmrCS+9D1Hjoo+4e/oc0xq3IFrKuNb/j8c3P1qv137u4jpXIbcHYKrtNv7uo6xjgm
0o2ZHB0h6+5ShoisLiUr+eDjsndFV9xUadMC/6+k9lfHag1KtV8aQufrD8PubXU1EN2pu4cszRec
IDkdd7bB2V0CsXhQ6NSTlpgehSMhYixl4LRhHtODpmIT1yqf6Tf9Oo0Vk5D45mldO1boe3kYEFdc
eR4ZH6Na1Qg4ya5rSxZIlgnGBMuwym6dNE6RL3RoBUewsqZOyUWRTTkfKj7ctHdpZIAU4l4KHKUF
3+Slv5qic3fGSm9kv9lhEIu57YM46fDLTyvKKwyHl1Z5ZTTRYJtjUy8IbL622MV5+8eaJ5sUO2rQ
ET+8eIs4Bg1mJFozGY6Bv3jL1s6u2D8R0b0VxSRRoCW7DQTKagaBibIcBBwkkkt6e2AjUsRM225y
/CNNZ8go0GIPO1dhwDv1Znw+48Z88n44P/71SwRMydh5FwIGWQ+dQU3hDKI5lyjlCN9WKAVnBe12
HbTFLKrclUjAVb/tIkvSwGhPnp64hQT8J7qbuarfQ4ZdnWIu8W8xHd/TIibMcy+RuUaNWQPS4uD4
1GyZhoBdJzO0tVzv0WgTX3IgJqebdziP/m/i6neCy3+iyBLiPc1DMxvkHfgxKBMvJCzBN/bdPk6U
85lZuaIBDigsEvVe4qZMIQrZpEnT/QQiDlGyT3Mv739dNLh92WgVS681qOCVWT+aeoMsLPORlC9H
3QCtdgaDZxI3XBOjT/wN9f36XZhl7SYZLj5svW2VpHAtwHhSE1H/QhFjCVX56kfVS41T8iufcIKf
y5/VZeeQwP1jveOw/XuPYAqSrvdXyHDqezZ+xy9HGQHzit2M/HAUT1chjzLI1rv01rzXcD+mmM8i
aFW5teAX6r5imRAFx0IBBNyrg9mCT5Bpn6LwCjEwTHpNOYXFs+A+oFa6Ki5Eu74nL6odRzu9rLcX
zYzJApMC7p26snVdEFHD9B12df55Alpm6NOZvt1/lUQxNRnI3QkU1lj8cr6FISCBEbIcss+hU9zM
jwG2KqHb0LC7rl4G1YkRkSTnoLW1szQ4R+0VvDGtI1DMTnIDNe0+1V7pvySNiXF71bXGdGB1sg7J
Ij9kumb+Rug9SabKPsLlxqS6vieILMyL1mQ+M9ueIRl2lXejRHsIDpmqI0JPyIV4hFda1icOiPOC
a8zLT1IFNMGBi1SWFkZnGDkYhG+mu0AEh+L8uCUa+Sddfr8PsbqZCsvIOVfs/uwMLKZySCSDHJND
XPCERG4U43nhXkm/kANBc0VqBS+6bCA5bKN4AN391NXGCfGaUZs1iVYrMEnssR5WJJP9wJBSkGoN
E9CHPuUxQ0/leP6OiNam7SGeq0bI8899zYeZTiddOIs0YA3K5nQA/JzqMo9w6mIZYQlhjoZlt16U
o+ymWv85lLpRcsrlZsmDp7KANBq2JnWhxnxcePa2vBnQK1N/pUtoQSFHP0iXn35fmeLwsSnjDkC+
PMTbZTTSEZqBvWEOqpsEIhhW7RLh5WOeFxDkQBJMMPdo8VHuPFN/i8jB50aJI5NclCKOaJr+KyT8
lPUxSk1KXKXr3ZFuWb+gd6f0JDwDmYXGrdxoeVbQFC5d/qoLwbC2YUv+V4HomccHmubd0xt6J5Hg
aUmpdPeGdcseDaZ3igs4/d9ECCWZs0PDqc4mCYjL7Jn4AUtL2LmISY3Chq8bWhgyMse3DEXpUryZ
RvtSXE3vah55a2zo3ZiYzRUP6HrysZYS7cX5R6EuIfxYST3e3OYR1yXPZ0aJZcIKciOdWb8hvGfn
hlKQxdCoZP0iOMHMcMlxb29QqrvuLkR0hjN07KxxI5VaMYzk/bmdpE9D2gsAWGyPhBtq/iySbF2K
lftUZGwo9C0UmZSmsZqTdcZPEP7hvE7RvPdZm5kERjkMnUo6dltgPbs6VbR1APk+xw+pE7UVccw2
7Z1W27a/dFz0WpdB94bRdTCT+pi2+OUW1Pd7MOslHNfu3I5Y4+hzh/dU9u4koNFtlhso45t0nRw/
sqJgD1BgLO6v79kOJ6TesdYeMD6mfIc6WR3EZjkL0laYi9LuICczQJmJ+sVYTmA/Rhm36zMfS7f9
/dAbawSPkD27XPNDoFoR76ZTIuybkBhPTq6SsH5kYbZz9r7+74j4WAp7kj6r0eawUJwqn9YEV+t2
468Q1hYlVO5E/QkcXKNSIiN+86k+YArI8/gkFiPWALf97CUx54GcSHYsdwqNPsOhjanCyW0/xulZ
yC9ubk/q+mIvhJZi7lEqPM/u7PNY6B+EAwyz5HK/ldoa9GgXgFhe6dXEe+d5pJkqZK0ssv7i4cB7
nnQe3E2An7ImmdxiX+b0Miz+3UF6lwVD+gFXH+nrITgVFFzNpOiuqKjpEU4ylMbb1KSdxpJoHXU3
idrAlgzBBuotIUb5y3cn1uwUNDdrcls5PKeZ7BAvcLUTml7JkBy28HIGKyTS5zLLVjcWd1iFtLhU
+dz73kR/3UAXNAxRN1VD6WTmUeRQS5pJFKkiQEkmHOccBW6zAANKamXHF67qOJd+riN1wl8O6Oln
FS6Iv8Q24nGtanKiMmzLSwtowkNbDLi3LaN5xfYKLZr4CCZbzgi0qGXak/F5unCPbZPqUlYcP/Jr
sCAB8wbWv1xy4AKfpMSpl3mplLIvzfGjBcxaRAbnSpPJRurUbdhoHQtP0voin7dr5MMd1ZRhNjFu
V8GcvyNCklEUn6kEZMXGRRGmBir7//+Dlf+YDtNrnbcxHG9tyIRkQcNFRau8ilvfGuGV3Yxur14J
EQ7JEVq5Uvr6MN1Ncc3Wi4fuGzS494YbW8wyK2Spe4ydp1oO4Nruol/dJ+N7DZs7SpmdoiYCaI8g
fOp6Yaet7OBl+A3/odGLOv2Cl2enU79Swzyv3hNcagUg/8Wzol/jFBu9RzAUnlG8qD+02s9Pa0kM
4KogUCE6I2fJoA0GYR00766LNvHE2De5xhi/22K0TkN+e3SBmgmU6yvKuuRUVR5UnIQKBBQE/qku
54QIJPUU1D0oKzRqWz9t7TOzy7N/j73vJSQAgRgkJ8ruPR9Zb/6fksojBxn9BKiZHfzzqdr2lPaD
bbbBBxIhqRhkTfF0rmX9Ufh2Q+omQNMuE+tx2JGDVlWFcHrGomCVDG+ZfK+NGg4X/VZot6i+0X0p
zq07amv1jIRqg/4+R0mGj8zUerUgyzhyZtlhLG3JDJuBh95Ew+fVNK4t2/2elWiwmD8Ffn038UfN
v5UzviLhrhp+sQR89+D44fewXJ1rGKIeTeVoBzeoQYqXk2v9pbFPMk4SltB7WZ+gYjvPOIMStrqI
9AKJ+mjlIYKSqTKmMeftDAyz0CeLrsfFjSzYT4lQUlTM1vdHSDhnHhYZ4yu4CzAgwxVEkZMm7PTF
/Qt/zFTKJNofTsCpmFGMeHX4peYiqnXzKGoyZayx+w1b26K7CckMsn8NH9L+Y/XlNBmrzLJirmAR
R1xeZwX0H8wjj8ecLGPHe/l0cc1f9XtqBv3YZlY08r6C9yXo784tUChNfHki5RbDQJs3zjkD7pV6
7/hxCH96Vs8/Ctges4Qa3bBCZyUKDZD9IVAL59bBQTEFSMRZQbiXkM3cH6yDTBmrpXlY4Uy9qhIQ
GSSjokgRzQe/qU6Q4fAqC143jtgUwR5SozLNOWn27pVYTSRDS7JBb6r/Cfv770e5iD/hLnJNYeTt
lcMcqlX+moi2JK/OZZd4Qh+pA3zqGBAuF1B3/8ZwDieNqYnrNdKoO20rs4gokdXEVyNDgP+Rs+Ea
sOmQQnZxyG/ouwXrUMT5mSIyOVIqTaRrRX9PRNgTgG1AxGp+lqwpQAQeFdvC2IjT+opsNqa8NDbj
VE8pa7QWorrA0/0eYFB//xzyzQzTAYLV+bWJOW5yeRPnmOixiHMqy016zY50nKdK9vap6kMe1dlg
XyfB8c3fvxA/+fP9fIVZXtBn/Y9mq7wc/JKZcKJLzzKEy+c29Gkg1NNC/p/LDGCc39KBBHEZL/pQ
h8/MwvRMS8uwuTiB5gUeeVUne17RGDHlLlRAxPyM5uqV9SgpiCxWWBhOhnNfuBOdatoo/0ttJi0S
ZxralT5yZO16IBUDRC7fqxEfqe9ekJz31Tg6SVG9V5VYIk8pm9WzvDTIqVujHN3FC5NQF6nMOVTn
v89rBhmafDN4ca2lFI/AdZMiZA/cvwQmoWx4Bv1EzG1AYZuFgJnLU2MLc3GSa8OqZ2u7ilXnSb2d
z+oixY4brh3aXhnGin689sRFmCepLqJRT2sFMSMdqNVcDQ43gl12HXewA8WPTyU7e8vWBV8eHyF7
1qBE+2AhEAobZJ6NzzrmAqPApGO9Dng9J991TuyodsDZvykdXR5iC61o7OvbflyLZ3WIExfRNRwc
GwmSj5O87ViNzgN5lSPAQz7+bsCHV5/SdSYHT56JOrDc4cmZDQ2eF5LgaXNZ1VV9Kna+tvoHkY51
lfa9uM7RmKeMVf31ttMAKH52DN6BAOmwZZmYsTOdDZQpKq5Mnd4w8/cSSVd6Wy8l8a4OGZPnzEYH
S3TUKt96cINaLj8ewy3MAXR9G+aHeUXPWMSAczwpWAvXqu17zOSMCOx9mXpzZYteold5qi1dSfsM
peF8JrT/bZwv4k4ts/H12egMovb72DoJRBYQytIIW8eBVqOwfUJT8LoOmGFDZlPcFNMgwnmCKkC6
n1hpCyw9gYtehCK9x59UwKE0A+T8MWbCdhJZQ4FMpo1j6usloAr34lMfIHfX5LSr3/MiTHWnVYyu
b5qGlP4yCZDiaF9QHdT0VW+4ezRC1lTcFvbHo0SuYd1z9B55nslAm3GF/VwGvW9cMtpXv2M7lXfP
Ob61UVkafNdGncRaWEJXQ5Njn0kI7TrHCMBxVWUTSNdf230b4vYUYOg/4RBoRg9Prhs6Q8iJJr5Y
P6Bz33/BmCV19Wt9MSfpodZZgLZyydtzNGrmyXngcQPch88UOUBrIzDPI+r7BnWyxItejQCcNAX6
s8Edfibd/tT213YTzys58Gqx+m0SaB4nXEEhgjzyRFLQDa4G4frHU13+hDa2Ud/5petlagh4g+Mz
Wt6ouV6MVUrPfujqnt1Ng97udCBYZ9o4h/DhlCyKM0WyEkppM/Ki+YVqKzQ7qN4FGAe8qb84SfjF
YWzE20+iTPwbPIV0zBLwcp7RDCkJEhR7yVj+fumELZow9OApDOJzCNcs/0kd1Zz8g8NDuseGODLw
e3wCN41JwZJE5SyJM5LuK8WwrXkV8HEnFtl7t99vq5MLsM9k0wcOWm82vTlVBBjTakjiXGbZKXx9
NGup7FVXq0ufmLHVS9hSfamxbpdeRC6EgAtF2XgWVTZ8v50vrtC7lIbCwi7tyEO4kWruTgvvHudY
1Qw1EblfnuXw6qAjfYX20nH5PjykrBFS145dgdApBakQckp257wCK9Vbz1vZb3pMdkscOBDdpyWI
yF0yVE1vrhwiENTfR84BDm9aGlJE/9rVn+SaN0/c8hMmnbL4X1JKWTEb5IlMcSqAZ2hmw0TmZQZ8
RngjsweduG9jbxzzXXZ/aDbMUcddcUkrlY2QW2N+xZjlDcH1bzpBfNA4VuHTGILDNBAKuLs2wVeo
ljGoH7oxJX9kZ3xgtbRzqVrbUFGT5ABoOpgg2Ffx0UpjmBx0lVYRoOt9U/z5hJrlXYT8HGUX/9l4
O1FWr9/nk/f+So1HeVX9KuZKGqAr1ao9s3dPKVtBSfwz1YCOEDE/6+TRpJZykjwnCI9BPLiHuyKq
nRnSJlzaI004YwKK3IkbgE0EE5jiqzWodJwdizWz7KpCmURXAaOoEytC/FUOjQ6THTlb0PCs+YnY
NgBTLNnolOg8Nz1NNRXtj2QCjUPq8Fa3fNK4v0Z2AFtHnDOQUdbqLetMfYnfnZqOhIbIYvgkhFww
I7XpJGOS+qqv/qmU0GzEEDgWsNEw9H3l7NbqfyCHou4eFrFW/F+kvWIm9eq6xyH690/O7TozKMOd
hJjvc8y5aNwx+kRp5HDD0WfPkRhbs7VNo2csZlVpLywbhhRETrpm3Vq+x9Q1jlbZ40rmknKApfZO
GJi2OwADbTabr7vDGIwpZ8gDmbmuPVgJfzUn9NKk7z10JZOTj61WP0MLmt7VxU56HbqQnaFtTvFc
/mozJkWuv+aMMIdWhNdag1caHcBb7mIJdsPtcJ/6u+VwETl3Yb1MPv+rnsHeDtQiYzYBqy7Xw4tl
E/xo+1/mZbSWWm3BpAPARkzgLdcRcXsZBA7hdVhDSeP3kxuvjpaBUapGIS/UojbuvCs2VVeLKmna
K4ZwoL9mg7qqy8BsprP0TJfj5n/EF5sfek8MQXX7TfliZkVgETo3vBmi+RBDUD9pTdTHu35yfTnx
Z/E9xd5NNJ5zPY3FlB09FclepYOc9qTWuWJsl6sCQZyGcwLoeU4UZMOgKZxF/kEVTPfaaq7UxX3w
hMZwT9CaRXVL3epAhwHVejnCNYkL5OhLB88nC4EV5MD2iR0ChbfhGGxHM2K7AzXVvOBe3JdyRQ6M
i7hbERyLTGnjE+fyojIejsaAr6kek0z9A46zyFCpEnQepITwQ8e9Dq4Yp5FnUfaXLoYx22r71oyt
t0so2iKEZyNOvIyl8MJadsG3/8JktGBqIwqqLvoUuVbasUQ1uGwfeg8v4PhYv4ouwcYJh21UTxLT
F/G88CKxX5nKQ+2QXqrbZJBLms/fOzF0Z/dxxZk5XobGMTeKIoJxId2r9ByNy5pfTag3YjNPmhPT
+v8hplhWWMSO7BArcPsd1SEVSHKaZ2xhiHo6QfIGH4JItjoQTqUgk1hnpNkGT72mc5jXnJ3np93j
oWZH1qu29CBPailaUlJYK/naF5osgRzevaUuZuzxGqZ0gPfTluT2/f6L5BjMzSy/0OSjE0XwC2Ne
cudCegZjTY0DkBJRtD9xylkZI0KqYnWjmHSsXyDd6QHqbkDq8OqdMbBlPGVVUzbRnOrUJyNa6smE
y4iysribBWJrD/kzadYR5MfAEKeqt+s9FDlEkalzeJkRfwo6u01sQw0hBXCq/67CPmxPXtc1mwBI
yHIKj3Tf1bIxykeYiFN0dyX6obVuF4cDBfJJlKjludhc+8ol8MFiFdPe0jke5lUt66OW9/g8D0/F
8Znp3Df7zLCMsUUbUUtvKBYX9K5mY6GfpDRTOTR8s35KwSQ0/W0/HtjGHrIGexaMJDUIaVcNwBAg
X7cVfg8Y/j+utuDxaSWCHfmjWSdZa+LxMdjAzYbBqH1WMHInFC3Soezk8CioP+nZk+ykj0ZIMkYb
jZEULQzD3KFjmpDFCZzcgrcw7rM98dgMq2a+BDtNITryK8xC6rAuB5g4LBXhACrlz8Q7mJFSpURF
x7dbK/ePoLj0xdZQTNV9lirAQaSLD2At1EL/6Ol98ydqPP6NZNe6LbqDQaaGZQBE6Spj6PUJmN87
ifYkdgLq4g7JBW7qjlkxHp2DNFv227mO7J2cpPJGxNQfpkicUGaTPRj9PQjkHOgdcaItgG9bHSi7
tPEkQLwdyxPLYAzX3mNoDAW++8eRFkry7WZbiqe6qozDej8/W9Fe7TvNoAEFtqzRpEs2w3VGKgQT
+GFu0HbiRyW5ki1jHVADJv06qqcEk1H8Hqqr9A+Vizt4qQvwvo/SJvGqAvAFgFQ3fKCIiQy+B3T9
unwzrotRHjA4h9so2506bEn5AbEkPZ11NQ57bwuKG1Is5g97zoxCshRDftReBpIk90WB9U5F+lN5
AgkGgq1k2iHjFNzVwRic2PZQNA8Ts64390YNN0n+dUFfsBtu5LDN2yu6xe0JWU26mWwhOC6eBbgJ
FHNRc5OIkAOCQ8MSizC6BfU9GrvueGUOzi7lkkNTAYPstTky8Mv+HnU2NNrZcbxNdkjx1Jug/a5U
MOUgPCmRe08Fakg1EuzqEy6qxXF6xxfZLIWn/1kqKptXJICPDxVLSf+a9aksCFiiDd0BiyYQ/M9N
Ap7rbm7tF6lvI6Axtf0PNj0lsv9bQydhx90Sw1a2UayZx0aFRPsU0Ejh2qO2hSvMJ4C0t7ywWjmU
k5jkWM7tgA5FARKnVigNIW/v25HeZi+50ZVcvTmWVvTRGPgCgS1EEUgYVpXcM5sb3WKkCQv8SJwX
+yV2FUSkwiwIwCmq9NVXlgU16tmBn+z2dGxG4xy46iWreYSYKiAn9GuvjY0sj5MlRJmhmXu3FaIQ
+gx9++so7rOj1Vi5W9DUkOiz+hDq0QtTcKkk72oeik7dJ2ViESscwDLjaGTXQQy2LNtqJCwporb7
WzCkztAswDOu910q+FGXXeYKbg7Im8ZF8WuIdwBF+2NYya06oj3u1g1X2yFw6mstfulQVyzDPg5M
fIhHNNUKID2WYT2B9UsKnnM+9XTeMD8/MMc3rrLPjCQiqpozxine+7+OAgz28rFIT5Zp67oUXVtt
Xn+aNZmJZqF+aeOKgKg8o300t9P33ZVq91xl1awISKAku1y4OwM42vagUyk7NHfWBKOCju2uJTXO
/ghMhpSIZtyG22Z07tp+t0O8Nyfzi9B2C4dmxoWKHT/mtuQ85VduoXp5a3J47C6CpHfMZeXb/ZIk
dtFfuyjtrE019qPDzk2lo6Sfo229zlct59h+LGuVvyJw6mLLh6vc5Mpp0g65mGv27j41K/0AAdfW
wNRy9Yn5+nNdw7qs3pZPUOTsyZPJmHQwzZQ2xhJiq4yRc8CY2P2ZV7wrFg4yQplJ4nJ0sggTQObJ
ac3dpGo3LM6ZuM8lPbVE1xkdgEKyrYGwWGc81LcCyDPdOECBCbniUR/b4yha7/8UK63igtFC2tmL
jNYCdpVnbFwGiWYRD/jJNH8EZpDtr5qZ9xlzB7Ik4ybbQ+giRG15DrApGk147zKFq2d4gu6rio5K
Pf/i6E7T0Wu8tkOSENwj8C82Abas3CY3mklKD7+VDhZx3SIYVwC/1o0jW+xXrTiSHxQItChT90sj
U3XDq3uLmzjKnz+nZpjuEmFBFT+htLkHWxsxxHlDYTe0rHh4YNvMG8HJqo5N8H9ISqEQTMBa9RNc
z1g15tJxi3VW7VXCor+3UIhbbGRjRkV2lrA9h6hzpIN684WrZ4/LI1mXg2bZoG4rgTsyoFCouf6x
z94rjtjDt2BLHcCm6z1Fq034AwsVrgh6Sv8SPuHgYg880I5Ss3a3aezeGnq7+C1cGB2MUaGmjeJ1
NmgAKINn8lR2Ft077Xm+xWxhZlkxXXSehpgoSLOdlsgYxxDxJfvl71MTMUzXFWU1yKxU3Ml9uCWw
7qXmvwRumhasGbYCxwzPx6psgzqGbxtRPPB10/OeRlQtAq+OUDiitZPUn3JCio7iCAh3E2vdeIO9
CkGpjVzf6jAGlwYFm7LXhtPXKHB6/DBSvZP3NmsMOLaNLVUuY5rpDpAiNVDzqDFmbXLPEOauqL5E
ZFNDEML6a+lwmkjeKUj5VwP3uhxIgN+s9euOQxUb2bAPnc1zk0DO+KtCb1Tg+PA/TZz3ZO69zkm3
zMwwzoo+o+ZszEhSNFHwzStzUf5dCGzN6Az6vf/clg2ELJGQNadXXo5NFduiQVNcUEgokdQlk5Cg
Gexndzh+mwMzy94LJQMug+ak4BPiCc6qK9chsdNRpfwYyf6U4GFVcPElUQKGj8LGJT6HvbOIW3XQ
QHl0skPff8NznqMlunVVawnfravYBOKUca+RLgBm5d4PvsX/edgzzT8X/2GXBAWbbP7q7CGXvQG/
WWd6jzexKTWjNd7eooB58NEeJYnoYB8zyrOeX9jCwxb7j8ZaERRXIvOTO5BF++JurU+f5Aclzd9T
e+ko+KtsI5JL3FbTsaOWkLrPXIJNDr/xPXD+O94EbrOjA8/RNJHerj68xvLtWSuW/ka61anS57sZ
g+YLHZ29b2KJVV/v9PDNti2f1z+cR07SMH/cFYx/5C8gA7bnfS5yr/dqMROI034sWOVHS6Za5bEx
TzZrGjOqf1muFMYbCzdzJs6uGGkLEWczzZ4LyJC711fy2ODcdMuMTpv3afS8C4xLIbNxmLdKoZQv
t0ZeLL6vBtEZaItb7JyvbskbW49GDUXzbQgud5nto6O5VvSgQdzoE8/JUqbYPGRmyZ2JdQwzbrg0
1Gd/plom+Kwy3LSc6ulNPU+YnH8565xlg7LaED8Vi7pCxuPSW//E8oir1YpqywZ89zWZXuvJQsW/
sj1IgN0N8mwQahgMHT8naPopH+X40OirxgESDyMiYh0GLagtlxM1yqpxXfpY1cSgR3MFYh633xE4
4l4WL3VffN6dthosxGJ5GrU2ida/ireEpymxgofeYDsGrYBVvesYYQ9ClpxJm80mCgLlM3IhfwIB
CGjz88vYW1ZrOmNcoEwPI9AN6LPX6jSh8HBniIOHvcVlMAJbrb1Pw40RAMEFOeldESI8XJ4iGRRd
D9MiMABYhlke+tW3o/cuaELXoxpCUvz7grZ7ulTTgJ1/p4X3Akl7f9jfvUjzEr6TK3XrPZ653Iow
ii9/erJqqJ2KnOliWcg5ZZO+Z6apxW8aESlj5Yw9BLR/heim0Pm1dQBSA54mOJ/LMkqW1F09u3EG
60FZfqcp1dqQigzIN8YJPG/VYXs6SdyU9j8KXaPmgawr/qi+6VRt7xtbLNS72jN8FnavTL46M8xq
YieWlfgkSoQp2kkrnruBFGXSV1slkNEFfWu3Ghl1MLKJBlw4f00+KR9Y3vfZ2f7/a41rahMEed79
TSqSYgcr9vpGGvoqgOdBCGRq8p8htg+JPv8Hvz75IkD56YNC11Z7OiWb8QmvPIwGc1CS4S2KrL/q
6sdXpN5JGFL9LdC/mDApQzxqicgXgYELuMH1y+MtXT5or7pWUspUcyh2ZDI4ILcz2/+ec80Mn3dl
OuQAZGGybsrI8F8rWWgyz0NycpHP/QyG4gt8avO8MvqEWNql2F8uSHqBBAQsocZgsTcCyG6V3LJ+
h+YM3dA8LL+VgrRHhoSRVppGGkpuXap9VgXDiFLfCAdM+3aLBJrKmjVmelX3IQELH+aXHRF3l42B
e1K1DgyiEWmRmdggkyMhB/7At9F0C+vOZfhCbcuSlJLfJNCuKJW5UYFKDf8ufG3TtzbVxIDdn+UD
bWRqmMXbQgGsDJQFqYCXnMtEAIm2zF9mMJgpr901sKj1k1worCU3jIAlJZd0ZcqpagZFftCct7U5
MstjPXv2KmZZwqOZLGae3Mgxw0X6eBt75lGVMrDabN/JAKDeSl6YX4lxNr439MG4s+EdwPhn09s3
JlmxiZGNx+D3bZADV1uf4hBMtI/ex/UQHIv6ePZCcWMyZLE4i5meabrOhyjEyJSFhvGmotD1Jkoi
wGPj0O42MwtOFg948v6q9ZpbwSpkuY+9tlUwftu+dKPWyc/7Skp/+PrB5A8hDQm/GZkOV52a8fJp
FR5UEJJ8iyYGwgMrMOIpIcwR5SxpgNSE/snxxdyyInFALVfC0siJfd2Xm6oQJkecnDouI6EWF9TV
FN2Li6rLUJm7RTJ0wk8YOHFeYdda33+XnPPvNZbLH5vBjSxCNqzU9Ml9i+hy1JGEw/cUVCHt1xKx
+iNxQDAkO3PWbrzw8xPoJJAdosra8MvuQNFOG+E8wsDyf5MfhntcwLkBI/tr4KL5G/N4KMA3GNxG
2mFp93wh5uhEgK8+5lnl1/9kLu6xBAb1Z6lCRKs1W5AmUZGVB/lHQg07pzLNIgV78kEmOF+0RpmY
/bKzh9VRL3ZkYKFH8IeN3X6fPC1eWYO20NXi0N0UmR27ffx4ICSf0FlBQ+1+J8x1Wl97jh4WfZb1
n2IKGt3gTRbxAkLET4JItZMJUZQ31epklCVa7j4+c/SAVOPsJHbuMrzA6kjFvUmkeD9lgTfxLnKj
ri6STvbJMPRSIDwbPk6Q01KzeJ0tMkKv8RBlAlJ3yRvfzscqK0usfaT6tUmgFQBqmJwwBfi6cocV
kVlrsbRz61WNgaRYoO17B0/NnrbNdPJP3PxI54dAYP7oqHQ52LG6roDdlshFHsf9NhB4OTuAQEFg
UyZ0h9frexcoz0DnNCHdoek9MpDeRsDdZ9C4UrVFttC3rFdsS3kgWXQOwtNhTmBpDy4W1gPlmJPz
XLxO9hX7bdODvi8TGgtGwakmpaMktCTEnrmSaFGwjWufD7LNwv4PPViC9WgDLu7mezmQ5xJyOhNm
c2G1B1PdefmDRqMqxK+7uR4x16YDoSjTJkpRF+VjrfNVJRhQqvu2dnV3OZ6Q26QMioKXH5crhzrJ
JKXgAsontXR6zGcxJqK/O9DNIRxHWBjzyJLala8xmIN5gojGkEifJgC1b7R07SxfPhCcIQdKybi4
CdtgmaXtF48zCog6FUX/uhpLGcPrhCToU6tTWTlToqg1PefPXSiRxIDpct49Rcgws2Mnc/f6r/7P
dhH4ntZkuhU2TvMUOx3udrn56IziPEp+mxiLnj+5YJcIGHT/M38zReUb5io82Ek75u29oWqIJIJx
LSK+CEeHFxc+kntMNktRfZB/VHNwsZFKSVVbTQQZ5MZTX33+ODqhMsnXl/NJd04FkYJIiYhigjnk
snJ2BWetp2S/4I5NoPr63lnKv/UfHoDLJ48D7fY2SotVYjJXOq7YvKdGBviX10OoKZknmuC+3/KZ
+cgNg0NfRdftofFZRDE2cnKZfdo8dXK62+Lt9eunCwOh69f7+E1L7uMJc3MvrdKlLpCnagNFUhFt
U7OzOFyAROfPHS5ZURPSH+JxHSPNZgCLNhOQ59ui1wPrwhKVxqWmcqkIBPQ4hJIEugDZRbSlHDSz
3qNzKBVW0sNpjHuDYGxPCiZr5ZklOP5I2YrE350EbcoDt5sr5mXo/bm+chw66xV+o3xP6B0aCQn/
AiWHc+B2Bg38/5LdCJDk8ejEPt01JSQ2s6iG2lPcx/GgvxxC3TMn1SI6c48RYS1GhQg6zDHq8m6r
RtEWaa7qPx203Mc+lbtuPxVP86xYhSB4qVyU/5OmBFLT6IR/HjIMnux32wuKrLf/KHEGwIpBKb3L
dQr2mDJSOLIz2hJ3Bboxl0WFJrg8nf9OrppJpPvrDk5BAUuhbUPw4s+HPIfhTs8CMBhiFx1x8Is2
tOZNLUZfAEcEkrsMnFoSIcX6MOsCozRYCpJLsCebapArD4ETyRHpYWlJaEXkJGvg+rGWyQblblBX
fIVCrQaoEsa7iXEG2FkZouekGtzTer6cu9oqjiiM74OF1DlJkHuMi6lCvgGnieaLlGpuM8qrruA9
WjYYyHo2PWCf4NFHrP+E7RM2LFX1aXmy5dXkktsVTdG8qjbWKczfcLRttpiaS9/Qi4/3hI28kRQ3
VqbikgwE5p8QdQ9mAWZ4ERYDq7hMIw8Qwtit3ucpnEFZGEiXk0x1pryj2QwdgnuQfQBNuH/M1CNm
n3iR/g3j1HsBz+EqecuoagmptHJT8uWNeK54kIpof8iEUX1NLOAJ9F2fjw9rpQvGE3AAGTcDvQUb
fYPj/9PpzjKKamU1DF0ShXAa8z9NtqZ44HQvYw8WmaugvpyJ2lem/K+PB4t7YT2249GtAvlWcCzj
ea6nN+403napf+FsGc3JQMMf18VJlIA1lc33Z3gOmhmnBFxxc7IzBN9ZrFvHHfPX9Hl/qpZVMIeN
4zjx+NRaohGDwFpBkxYSV1SV0tjGDMWQkxK2W6s3eNwF0Di9Vm73SkvbuGkb/WU72cuFxd0LOzFV
IVn5lPH+w5vitVYr2adYhakfxq8OO/dPh/tIDMyeRA65uD+iNCkY0WbAvyoxQ7F2oMLaxZTRsbZn
4ZZ4YpacyHGNelyEMzEbSzeBUddXjH3VYaAMikHUycijv1QY/56RobhhWnDqZxh+DPz7uDjyqc/G
N+RbtihfFbSePf2ReLtNMyzA6dOnHxQWJqEqv63cz7qKhgUocEOzw+LTnV/lXM9UbCSwAi1FXJ7w
vMlZdYVwYytBHRi1AvdgYafoLd0CpYDt53j/ZMX356a1bZ0mFZhZIRgUFQmruUWDsTSzFD7tl6X6
gjfr66mr1wiVXhi+K8D7546ZyaAp422h3U4981snQJ0WOHX8Lmz1/3fKMUYgezSqifyNyz9uzPQy
tdrZlCA4sK9WgSsOtoxQBqpfw9DQ/bDZLWycB3dcf6PANo609XoLkYfikt2gDaQXdkBYqGwKJu4i
KPRALWlGNAWs/tCTLnilDfKgCYLDnTVM9ib213yfIQRf1k7T/zHdczY7LuJdwltzEhyTTWa6CZgj
71flePiaudAdk3QmflyvEBQAX271TCsCRMiExW8hOZ8zrFKOLbLnQMPMQNVcKMEhthLg40C0GTAt
gHxl5K6ILl+Harg+Y1HH2vtM5RdqoJ/fghSQt6vPXFyFlx5XTTHcQLCWKzdUt3TsoElF/JOtK/D3
KxdIDyD4HDmALtwk2Isw3NyoMQ4GYI0QPrmqtj9rNoaSqXdqbGJm/d0fL9orFPai+HnZM4H6zwkN
EDz8SCXYmN42DywxCUpINeAkK/JTht801Fv6vVWzLRgq4rPoS8grl/B7V9O/l1yZJE27SrADZYfv
NNGHkqtFneR4C3yDyyqhfO9VyB6dnJEDkZWYgGIKxLQQ+P5zrj8OFBunfTZs2g7aILQtM+NeapMh
me4QBN+YnGEWuYEXbiFvTPdqPJWtvFcoKKDUByOEv4CKzQy7U8ERDLSZmtIN2Wri9V3YQE1WKwaC
CxjZiHF1yZsTDBmOUL+wB4xVOoDYQoXhgyXy7Rs8+qLUPx+acK3dhuD5tRv/4G4Ic4nthE6HBWJy
hQhHibxGbE8JDhjhfwvTQAKip9m4+n3+EsMmb0gPF8W52h2K3lDtgYKPIaBgzyaiWEpzoQdb79Vt
4NiJUmTSlKBwdgEu07p2Vc+LyCTRGErAYBDGiAvJseVjeEwiuaVhDz+9OZKF+EyIcPA4EfFZ8VXD
D18s7F7GECiJIjZY3ynYhho+poWOSMg/1SjvBFb0waiDwp549aYGDKkxVIL+DwlIBR3/JGUaAI+P
8WhyWNyA867YoYWjMv3sYhsva0uyzhiXwjm1MhvaF9BRLx+JDQPsIRC/UxTcN2n86WXcAgRt2Bi8
GEYyX4/FaNrW3oGJtj6vFaQnYxIP2AbX1FW156EXWvjodA+hDlzaJETsHOzsdZY4BsXy7+Ln7In2
fTusZFQov9RYIvKcXvzJinHmKG7TbYXXKSfjlVPuWGuiR+MELAWd81LSUqc6FSE9n0aFmknkp1Er
1qiujg9EQSAs+9EKcS+AqFJ0rz38e9mldovggsth1BuP+A2dB7twdc3U8XfrvQfIQLhQ00QCItVT
uiGj6x1dPecK+qoUPPiGmnzLGOK+PE0x34wxM/aa0a35h7wAgLIGFSutyoWLA0e4q6DJ64tondPa
3QkDbrpybmvS252VWf4hdpPokebTpjMr+golgc6wUejXO9hgBJ3ao35J5Jqp2smHN0gF1t5+aY50
EZKAcoce+uE12750edrY6biIUii7HQpiEaD3jsdgPvLNo/NDNCJNoY7lgNYc4522LpQCAEdOgxwZ
43x8LIxAX5iHIptWuVQn1+ats5L7PEmosPzrV7FTI62XBq5YmeVmedzsyI9VW6jlUmJPMtmK+dJo
B4MC82fmGWq0NfHk/0D5oTaSSy67pPzVA93PG3b5jkajJ88Wy3mXFe2a6bUnz1mYW/LNekPJFWw9
7o4GDsPfJMcCO6OEc/+mgNFj/UYTYgn6N+YuQJlQNyHYT1tfKs4O4Kb6zzHBMz5LfUbXkRkp3aVm
7afDr82ni33jdCXxec0kKJHiY/k1kcLItyUteRsnqNceYQGMHEnhry8YIHQjqk+niNYlg7209JIi
/0hujct8e9i3iNj8p74XqbrKSasVKjt4bbE/mNrpyptEdDFLLoXiOVj/S0gNCMf25jRsL7zLJReI
uCoBUdHnUIrL1er9bz86mbclRKfgSRd/0htc1FS7VpqHf5lBjC/YSjqOY6Gxk8TeJumPr0ebsZad
ebozIh1U/WlT/EeWG8MgeI6A0xgIyoORnbg9Bk5U1iWLAciwhtdU0peEpFYApCx4kHmdppC8onnQ
uDD5I8Kpo+T32Qyo2+y+psWd9OFqA9M8+R7GiwNlpR9CjgjOMLor4oLmFeZpp+cGEBrGEOIQJUT4
DJKRmAzWBiOPA/RHZfcBDtxKdSP6OcFOY8OUbNu56XNYhmvsg28CQWCFgYJoMlQlSFnj09PNKymw
/GEd8obEZfheIv0F9QEB/PpXpNmMBDSU1GtO9HsxJu6VCD3KU87N21DN0fIIwlEVuY1OEDMR7LFL
GGAJKc29EWeKSo70yAcWBVfU6pFpM7baqYS8nMe4+rWn5IOafrOpYh22MLywrlV6/7O6KolZfKHc
MBCKcE0hr0l84IYISFIUGRgDKju3v0OQKscX/eaj+c0naHc83A1SZvNkc2yUEQjJkUtCKRvR+CRO
u6eKJeFvipRyxtNhpz75jK6doTgjqLQQYwAHP+q55T/w3tPLQZL69eDh2OnJqx2NKOFAFUOGV6kG
byMbJtcxTShJFjDZNliiotKFaqYYl22VMOl1/LUK16MB8CIcav/owYoen0SBSJuoSJufWtEPK+nZ
v7cYi4z1QtynK+sebztHpubyVcGE+jYuyukpNdQ5HK6039qjwr9fzULkWmAAoC3FgezGEuUQftTx
dRkwstCHIl3HV4haJIo6jBFbgrOOCtj4pj1HV7S/wYZ6b949KW/3bMVaUHAo+EZSrYxffVRAip5b
S80ex2RVtq6giNL4HJrk24Imgqj2bxGCP+w++t5hFFz6gADRkZ7e2lGolSGdI/+a7yRR+5aO+TpU
h5ZUgSDzQvz3sxkcBpUKqwywHMmJmaPINXiyabVw42+qnLd9QrB/5Sya7Un+LF/rj8i2ZUulHR6p
Cc3EzwY6W0lkUZuxIB1BUKXjDIz25lkJibSE+80ieHsh3YLNeUlDYiG6gEABPIgU2HZCj8kVM9X/
s4CySqd9MZYSefmNt/hwElx+DS5HBG3vzOljb3tqY8v3Fpz+/z3ClpRZBusJqbIFW4RW/RLhWgpR
CgZ679xP9HM+WJpGmADE2JbvEyemp/7Bbs6lmfOQHngnptmydB3/ykuxz7wHR1iEdyIG+o4IW8tz
yrBuEPX+ory+nfUuqYwC1L4SBEDzlsMJuHdJybwp+Zxk72XrjUYDYUi6gV4jffll3ZWWmPfUDae1
7bJPy4IL/3BLarvKJp/wOLDVIncNFJcoMfwZaHS26zza5rprcGAQKzvyNTASDvv/5TUGF88zFMlg
T5V1383U1vCXlHPQw9IP/HU9ln3kh19M+AT+vsTDsB/IRliVty4NB1SvxGmD+yPxmYyv9DohcN0F
qFMivvWciMz0+agPlYE/r+EyYignf2uDLnANuMH1hoAPEj+KoMymWKKGeI5Oq/2DN0hkBkTx00C9
R9D5i58koXSITP5MiqIW50Kj8v013s//nVJpjSCoOHAX4W86l4AV3d/5pRE/gXLrYmsCr9PiX5cq
2oBTO4tcMS+A6rHRUIoAgVd5LBwdnFp58VB0HNvC+LVVeVSgzIm3lWymIZeTvSyuX/0VHFczA7vV
ex0Ua2m51ZK3jsKmkLHlTbnm4Zh6fuv3XX5xMfDVsGolMMTIyEYJZNWc4EICZGUydJL5ahOerSF3
9yQ5HpNMjDxxlcL3fQujuRkqI+DMaoJKlF519hyoHv9mQI0ARu4B/CI9n3OFCJwDC7hWxcD5POXA
MXScXmTohjuXxJTaSztDs5BgkE97dzOQyFJbT8wv0dDtBhCdpM2BR/a0hchxHU8byzSvOg0/Es3R
FUQkiwLwdYtBlXzhEl+U3dpcooPOk9Smt9tHkPtM+evFRU2pyjKD9VzjZNd+jnUNLUiPo4OfA0oP
Uos6un6cJr0+bwacTttj4m5muRnjdhfyycs+S1aRgDpqsssx20gFHfD2By7hR6OlPuGvU5CjL6P+
A09JUcvQoh29WpaTNeXBab9xPZ6Wa2XOPCAmfoDz8mcdzeKDvRCd/ce8+PpUhO/ffAkc2/T1cKwX
vkklivp60TWxZ+zx/nXV9bau3mtrxmDQDzc3doruVdcs5BoWf6PgcsDNMAmpIH+J5wcrjsAg/eHN
1wXlGDfOwB4RFIHsCRf9RZfP2jNQtZvv8P/zB11pota46fp6OCCFPzedsL4pFHzMBJX1RDEfSIaQ
Q3c8pl6Pg2TP8icOVwCqCqAZRjIkj4e+ZX1FA7Ul/rxLoAvivF+hBVKkLv0+So5LydXJoQxALSHT
l3kcaj7X2SdB1dPI0kvihTfmTY9QE/uyUfRYAKV07GBplQbpTDXmluqbUeK8xl0GBpmS8bKEiD3Q
mat4WeeYqUw/Y6MyzjpAolp801gncL+yr+wUz8kLjC8wAOjArm/ZLi9qQyJR4J5bed3PVAgKhHPg
GD1hnle/lA9/CRgTumapzgOzw4FWmT961Ejb5myiAuLSsQoKY8lUYhQk9MNJz/G3yptjNIYIyJPu
a3kdTh17ybhqFvrTBjcf3lJdxPL+4JdVn0Hd46oqoiuvinAjBXBXE4TB+mAxU7H+LiTE1CFZiPAa
pRx4as4GNcgScFfRbw1NJ38dDHQvfiufemDGHa0ckMQSBarZ9Uh1Fq4vBbs5PCHZm1ELOJXB2Jj/
IpmuvmXJDJo85f97anEmQyu8EbZQwZcAkbwGzkTc8ctwLXUj+Bw/wNRddEM/5WocF2P97mm8OXx5
8oV66B/8ttswSDu3GUyJY0DvvAJaruqX/RlFZAofD/LVFdYyxxgoqvYgv/01HzPkrxS4goHHAJnk
XW+2Ma+jUDnMd3j6nBDgPA5y8cgbCLhV8P8v3QqYFOCNkk+BkSGjyKua/LyJsfh7iGv6KRJAoZs7
rZWcyzplmrBVCS6YUgdREIhOmQaascP/f3IJioe5jcJYKiYOo1ktw7vBBFd+D/vzQJujvGmWpO/u
nZBf4PBW6kpH3Wl+/dy+A+s1QBjld49D6CBCcM2Hly9CZKfW/iOI6J4GPi9/2Q4o6Ky3fhgRZFbV
jhrtuCdWT8SH22LulfgaPSlqKJ+M7H/MYFZqeOJKI5iSeqxK4MTQ9pzK4liTK9piZmBeH6+kH5aU
a2I0icvd6PskVU/H2ZPfbkvvrXzbXAr40F0L3MbtdL4WjaIcejcyWJFCrlNrMiFIW0CMkam5j2qe
Fs+q7plH6aRlDZbyVS346FO9L9A+jt7g8+jPNp0sNGh2oItYi+fAvLRR+A5EIyR0K8HCb6Ct9uNc
jeC9wEH7cA0D39yup6debn8M9L9mcNiyecMm96zonROfT4MK+w7niZDs07TrjB3+5mclYrFpA0sA
gbcTWXxlG1RYeE5azD2Z+FsKwk7OI+rYkl+XCF96l+6k7xHiF0TsrhI+yiU/i3vhcq8Ang8wi1AT
jvEOVlsJN44omSpNIrWUBN+cLUDUZ9Xk5ZItUht8J3QfB30rB/EMELqy0ym1nyd14NQ6ug5isD9s
hyZIiGN6bW+pum9Z32wHrOWgOL4o8dtG6GRQuIJ2O1d9ocZLCiHUWZFD/MIijKkPK3IgsSnf74sW
uppG6HJIRog0aQHnIp/CMmJivOMZIhOHPvHgxBPvqm+r5MKWEWlclKJzXYTaRM91s9rR1+yOn+UM
77JEdM1zeGtvy/FbIHhbJXU04/tZV4F+rVxmqI3oO9dXG4U6l66q5Beu2q+TunU8Que5PNpZ6LuD
BI6Gwzi6szQscJs/c751wMKtbQK2v7wSUGvWsIpeghC7e9U7RN+GYkWMZjpO0qDyAqxCKyRGiHiy
tbTLdb6/DEx1/AW5DZ4KsO6YWLO8wYzGOrHg2lN3htu/1gDwEC7eHmkRTUZr77gFBz7yuGXnukHf
fK/gYp3WBZDST+2x2WKv49dSaWrZs2qYZbkZ1r0dVmgMvcZhFFKOJ+uaVszbZCqA5NbxbDLiSVHs
WW30FPSuK0R7ku1uGJgWsu972XrZ9Cs3QZ9ev4laK90PbBAPbdGkgeWLRZViCvUk1C0Qa7g0Q3fh
xIeE+BC/5toE/gm26cgIs12FI2qZFfvLjVo8XlWON0kWy+OT3gxp0Wo0KkgGTJldHh98rHgOfWQF
Cirgl4mF9W/kK5fxasBPakLdH8YBYxQOBQT/siLWchvN1SpzNB0tzJOwi/rKirtiMKKKfGbJZhMf
4OH3yy+D6UrKtSy/jPAJiHtIG7TExDIP+scKWEGpEg5DIAzRvf2Oij7Wg8ko0Cp2Z3EDn3ZR1FxM
2XrgsBo2kKimNRZZ4Qn+SwJCDG3Qfx9juGL+x00iKrmmIGNGm2IU+ZHpGVJv0yR3wLiS/35frDJ4
NTlkCSpLEzQ/mAI00gyBEeVmb8QzBTA3rrunFJo8BGJsAl2gPxsB8zfJ3oGUEoFY7GNtgNyoWSxe
iC1iJkRSNpki26TldHX0OZBa8/iuab8C9h56vRzcJdaBqK18t4wWcR/reMu01wHsvq0YnUMClaxX
ymjJ9VP43uyZT6guaetRSchLaN2AvdCFnaBGNf2tH/vf6so5go9d0C71o0uIy8WBHhnEKb+pfk+G
WlparYv8WO84z5eK+U3lDBO3rMiQGEDWhoqXzL5x7q+WBnw+Scc8RZqVUGyzBXEtgbuf76ZwAhKC
UrSni1yWDYl9lbTwR4Y59Mfi1EOaWhL1fQwaOjz56yLnS+AFtYFuGVwRw4YaZAEeKsSiSKbg7h0T
RpcrRJgRe2XMtZSndj4bPhtkrR80xTy9Dv6zJtYgqsN3bOYVkt/0DA9MT1k4CP+p1NAzDbxE2OXu
6B9BbgW+I+jWIMK0GzFS8gpdzAQ8YXlcJhCu2dilUPb/yezMhaLPXNnRVyyaPUuI3e0MYOqsfhZn
V4o/1d+eeqFFiuWZdgbgYRGR9ThytPtHf2v549XKtX8pKn/OBt4xil8L14aHi2o/58QAdreVqp3P
i6JX88eYwO8A9VHhwJ8FEa7fH81nNknyq3Wt7WvxL+QIEsilMZT8MgbsXJQrtiD8uR0OtJpRk4xO
6SbfQJV7c3nCx+iNWKFAR4zCgEez3hX3Ia4Sc7FjPLG6kYWiAXxnyx7PWqNlYJkGGYb8xJqJbxOg
NocHNWxN9ux5P4hP9qMHPYJjW/YeC8tt9aqJHM5AgjoruSjMGY84B9P/+o2y3TIAn4hbx5AcGQhp
5tPhL/JglZxh/8Re8tpUyla+JZKafQ0nL3YUCXdslkRod7XVl2YF7ZdrpGyd/FToV7k9D5T/cNBj
1FVnLJRMEXMuYYPkkkn4qc6iJnenvvW+deDNwU9PK0vQStP4Ykjx4eIebJsE7ejJecYe3AXNcwMs
4moK6+pVdcGYbTiuU2PXwrX7TDC1QKQExhMXClcaUBQ87q7tb1xr5eL07QPKvO9ZO2ew1qtAAPsa
Xn4icRg37qxeSW2HE6vHLxykWvwj+f8wMalEWU7knb4HmM3FMZNCvRwhCAf+uXHG1kJ4E6tBTp3P
6hzh+cz/bOZJ6y69xYIKdxpHVrA/eVONwJbRn6BwDQQpBawF2FbhVIwRPr5tW3QcS5sVA/x5yiLl
tNls9hLwNq84jYpZxTKLh/GqvQYC7OdHilkK3MrLgwelZ+zFenB1Jk1oCu/TA+DAWd5329AX8Z3V
lrqc9n9xY8uG3XjxORPABk21F3CJz9mf7AFw+7CS6OAaXdUSt1EshaX4C8hJSwwvhwhOneyBhDoT
lzBcD6JHr8SDquR5274gJRQSnaKbTlCFLBEiNJrdCW0S1xXBuevgq0+edniRYF1DZvzuyFgCjcuT
1kNhgG4CC5IG0Om7N/kcKDXRtxVn7MtmSM3GFu/8/atSZ67rp9qTmCrrS5YHCy9VrWZwhb3m6fCV
d3ZaiQ946faMLaxJs5vlHn4XpXVZjNBaIM42DSztCphNTkj2GCnvqD753/aukQ8RX3pTTtSY4v1L
KG2atvdj8ur1oHA+XgtogNro9/ilBGTM8WYCGI3RjZR/FbDHQtjaZQ9ZBUE2Tuv4cEv3q0jGLYaw
y4OLSTudaKIi9cUSy6UsZx+RAySORkilxC/0ksp4+4DrjgTwGyDk17iuWsxmBApmbbRQS2AfAv89
kJ6IU1MNK1W4Z4TSgTM1qnrUFiyEhhxCi62Fo+B/dBZnpPdwqwBsuY5vXpLLpe7xpC1TgkqLTo/Q
ZORLBftpwGQfD5jYWQ+NIoo1uWDs+WU+WaW41AeegJLu7OOBGijOAAEzFS0eOxbBXbG3xlOQG/Ef
ZeqD/tg6LLwHNt5aSmI30urCyYFhQ/fy/I8oaP6g4Sev3+AcXWhUQfJXrdffhZQmDm9rNsya38vQ
hhyLmy64QZk32GOGmyds97kVVvd9vthGtT1jwD0EMbpXhf6z8oATmT/QScqZYLEuxilmsBSdGB4g
r2jcq704RSEvsKrGykNrhoCZKQkWL2Jk8YahpgYvkZxuHqYVgoZE/1NBZWKwozCo/kMDfATYlons
QCP4xb8mSXxLmojV6sGVJNUcnwtuE0TSc01so9yrqyc7yKbNTG2BYQQfsktIH6lorG+/s2I0ZPfz
nVMWF7wAkLCYgre4Fnn2GaKjwiyBSLhqfr1pkudO3DGf2+xDTASDCxNFFJutf5zmVcOFdVHFnO49
JdScUMeNTB42f4KwiBgBouqhVRXC2CvhYEpeMuPZ+E8pAGtWJvazGnwoMGjsYw22Lo6hU/lRnfSw
XDVU23+NfUL016jqpfmkarHx4Pb8trIJ/DmlFurB5IsIhdzsgObKkqSAtDzrf64nWxM/aYx5eZoy
v1UHa0oRyWa8QMxreOGyxamlUobiyZgLzy6XPxVYDa9EaopViGv1GX0RWBu0qiyRUJd38zqIUglM
2eouQMaYpxfdcdQr82rZmJfFLVpKiEInN6Eged9R+6OXPxFRqBRfdx6RmLHlx84QtatqdvrYE9/G
1k7JycT3V5dyChm1cTBRBfNfjWKVCWUp68Tvewk3RGrR9FnEbEBvzccYLlNcob/e7rP3gKlvYgxG
cF6AnJUi+rQFq0rFPAOlUGzWEdp/ChKX8wGLDuT3VMTZ1Zvqtdrc5XM6E5YaHSvcVRkS8rwiVLXu
PAcJzYjSwywzNT8FmPi3wMmOXpXOuoH13CJF/j2LUyYiqifpH0gRCTIfjUwNlTMrUzmT0cQoOqeb
3tZun19WyKsm72Lj+Aa7mFIAEOgpATzozkQML9LVvAC+DPCVi9TLCzCRSRX2bP8JbMqEo/fY995L
lRhga30Q+Q7D6zwuESSxM0xPtWNgQl6i6PnjxgFoHyFpTXWbduMG9VbBRhe8cbPDu0/KfFUzsgBB
t/4hDn0ZrVnnjKV9ra793wIz2O7eqMK1SvBo4gDZ7JW1W8V2UgypYqQmEWnsDfLo/uWvNAWt9P0t
4+lXIrUd05NSHQrZxdwxPOjfoeeUQHzj1AQGbWz1aWVovVphZe41SuzHCMKRWEFuCF3Oq56EGU+l
OrE14w68qR+mxPqpg7wou8+HNLjPbuRbGxl9re42dmi8Jw2AhfG6KwrRbUMpV5M+NvvmkbpMJAXo
MsYgZELOJfqV8qDkbprlSV4/nwEmDlkBRuFeiX9CLepYCUWa2WuRcOW68DMIgj3LOLuLhIs8UjVw
6VNxhCHqoJN5dB9v80Z/HTymuFcCeRHXu3MZGjCS+MxyxmY5HPcuQXcxgbKQlEwvXXBK1kTRPowL
i8Y1k82u/BbRTxDZw9y9dlzpkYadeFeK/n/7cFAB4sO5A1GQ/sCoIVacNKOO06Yf1J//4GTTThpF
7h6aA1pEuoYj/jOZXDLFReArI36k+x+5llSR5b1Uzk+WM4LvVzRUewpXbOGoZzTD1hlGV1hh2WIp
KHtIz/g0dglT3qC5h6jDOyGinb424kot3mQFVPoi9sErUqsBQ7tyJFBoPUTWY1pvkNBjuAyfiwbm
4k/kYXXd7MQg3zS4tqPzuDvwcpLdoeAFvPFkZ/HEJFEhmrAL9vDa2Z1VbMH0oaiUtKRwyQIkB8mA
sB9MQl9yUncoaMtDsLe07KEn16o3ayEYvGelUfFlGV0e8X83R18DlFSHFIAnSL9kG1BwMdeR5Zk9
qcnpVtPylg3aPcZl3fmGRjzk5J5jj8kPzAiEe9KCFI/pg2lrF4Js6Z43QqifOvbitjD/t2aV8u6M
wjTZcYLXEVQXBwDNFmcNfyZbnONyGNqzTB0T0ZefLeINfDrTJjXNa5eh3RKTVsOSEaTB+6k5EA20
GKaHAGx30b2v3XspsWQV8iO0wz0zLueQCmDRp1/YIcH1v/VH8UpUm/wVAmWn7jK1TXIVVgiB4orV
PXauGonWa9P0mkige8QeIuMl6r8/KYGJBAKoMDXDqgxga8fO/AhIZZ5EY/+d6le3uq5FlchcCZdD
B/rxQQ9i3pGzjh8lzsNgZiG4SqPMe5CSdcxv5CLFTMfKKDta3P0IAQIByVfoGRLj+m2/i6Hkp8SZ
qcAmSQ7aj89K03GEAa2cqdA6pTT62ck1e0YvKH1XCarFAkRzbHScFIryEgxJO3iblebGuQDVEWB3
GCY2ZhLZzqgwpW6EOwoYE2IYBePJjwOLuu6tfId0n+whnxrgZQissmHbp+89C/EMtW6m5uD8lAQj
KlvJH3Y4/RaGaRbtdK0UvWO6WoMCBsSEWtfw35b+0okt5G7bFOFz26IfFIM1ZeepGxwUaimdSadb
R1tv6Th9BXRppFpn0EGQyxpo3tkB3zWGZgAFJRSWrzWmBIWbEfkyqmiBBTid6E8yZOnpIttFYxdU
41ggfSi/TBrYD+iT9XFAXlTLntns93KUE+kr+Q4mr/rXdnNvNzC6YESLnkMkqV+t90Q9sUWo2jDe
/Uh2H3b6102XPtqbSExKVNHQsuTv7UHU4qlFwZPXjaRqZVsKgEJDjSdmAGQiH7ZitC61B/x3783A
lJPPcqLWFpUGyPyDSkxA1awm3HhU/225Z5fWwqIXbhSyW0TYeamY0PozqJBxt5ib4Gm2LSImU7It
aDJMPYD9COFxB9VzxA8Z1R+aIFPlAVKKIwS0iWXVkyXTUzyGLO9yR/0OfbAVY5x2+ANlWAiSNDiT
tLPghhBh0ZiN1DkEqw1V0uTx8ZIKIIMOKJ0lszXRAlPVZSHN+ybYaVb8qMYgWK3oXl1cq+VNsWWa
t1u05GcS8FQyd+TAIcYmg2xgOMnMH+9E2nuPk91coFEWjLllye4bbhuPcrRn6DMzjI1nBvLGmkk0
cFJ1zky2IpyJnwjYSd/Cs6Vo2TPfcm2OMO8IKaeaENfgv1tLtVDHt3Em9nR6kypywZHE2d3mpHqs
1bxmb85HA3jP9jxIH1jJ7WMILh4bkIpmUfQOceP0sB9HYdFDBpuXj5ehQhJV27tFwhquplKJ9nQT
Wi4RCt3Ytmf9tRSA1F0Kt3kwX+SCw/CrPEzHBoiLNhMsmyg+0AkqELQFkMpunI03kGSYZEMlOTqG
QW92kEJlGNroLPziu06KVuAB+hnDzyK5SJgzxlMFKcoYXLK9IxHxEbUMY5hYZEXnplnb2Z3bZ5Hz
jYEMGFDHnQPvBdIn6BqEa9tX1Mw6mnDjxyhHOroICmhpyFvFoh2GxY+nQ/tPjGWi5+bECCqazmi7
TJFuQZ8Wx8ecEfhYpaSF1EWjOf5Cy2tvh1dw/a0tATgMOaUl8gYbv7CEC+Mi9XAc/PNn8SrBrIEf
cAyGLmL3uMnpO4eHIFtDkO9AcD23rYC8ZKyjAJmlARsy1H/8nnD7JrpDxqEkQx5nFj6T7AT20kfe
3f3AZ9utd5fV4qXT27UHlJXYzKhflxz9xT9NV829bShDjDgCXbjVT0gmocP32NhMxAyXoMPJpCnh
MtKPxN9FKkJxAnZSH7mKe7v7rwdLGdfFkGCeZiRHNvEqvu4QI4Ie+bQzNpnjYIoSoKYzBwya3TeG
/FiSxf7rt/RKOpCyDoh+rw3nUUBBnmIs0Dl2xIPBQ/WQ6wKxlAm5tISmzqEWDd+gccxkMnOu2bjP
DvdQbhnOY3WmOQc4jvyUCey3yBL2IryKc5dNxuO3CUh28ynz5WqlZTBekTctfCy3PqZ5ZBX+KrlI
aWZcL3dIVQ7Sm2sWJlVop7gNB9Bju+9Um0Y3kqo+749nia4GSW+Usmyaqj4TCzL1yxIAp6xf7cRr
jc8lZ7S4+JwsoQpqKzGF1NiH8M0+d3v+UYHoRd35xPcvcej1fYntCmeLrkpW2c6F7Iwp1hTG3mOu
XSTAkrK4GmxWgECzIDDC+x/2whFtjGq4kxGHZPYB2arhIfpMjjJb7zAo+zzhYGAgs59kG2Z2XHso
cdFIx4lkXkZGXrzrSEMjEEgiHLHa06jNnF/EoOwmEd5SD0cEmCmINEDhOK3U3dI4fuQacZx/mg1N
FGrsX7paLIv2nppBVcVn/gN943bfUaHwJJzedlnLEkZkSzR2QfGSHTJH47sutVKLJBRKH+DOoV/L
e00P+53RW2MsiynOP+mRp9yzjndKi3iGVNbJTcxOTXRrB6z8E+b5XYSdYVrti7Um8PH1IUXSCCAD
WiG+4EPZhwIcFbo5zVM26Wyn1aUwWvkYG3mk7g9uGgZ3DC5Z0hwWrN7XIipFZ7wbZJG8o2olVmJu
Jhi8GhVNopON1yxeNuJRLu1glTC2+p2pln+JRSrftYVke8cl/hDPiflyI2ejh4+mcq7UiccjpYu4
1Phmro0pghdsHZrb/jt/6MSQQYZRoqV1YB+zzRcLvxF3Yz7yiEHHZGvzjNcCwG5wLyn84SvnC8Wc
6An9fa9TA8ijCYJ4iOllZ6isooKnxMM5rdxlsZYScN34hC/djMO0r1WKYdiFoVd21OTliQmuaJ0o
sG/q4WAHpo3ycw08xpGapPFW8PUE7drMmwabhVcbLorCClUJ/pBn0UprkdgrC64qgUohcw/CEYiK
rrG1jBpmEAzMo6rTGMvbJQqfb1sUjhTiAyig0D91I20jH9tCaz+boC/O+dYdNyLX/TLh28AIzdup
NLtRd+u127rgarERfRQrKTV8Eh6tUd4aCcYVjOXAchTwjG+ng6YjMi7BKNcpt4QaZ2ovyKac7NW5
n+Yo2oAj4e9TMYwun3Rj10WYji68Aluf5ifVrG+2t8lyBaGlWOe68JeMVofdToXozr4p4urx7/b7
6CS2PdK4h4EHSwXAl2WqaK7W7CuCpggpuPzn0+QmyQ/SNZI5k/IEgfsko2Ip9UJk6Y5EQGa1nW0n
P2cA4KW/DqlgBS4OeeZfY9RPf0czuU3lnQ02CvsICIlXmDyUOMMJKHN0EshtHdysp1HmjemgBXv9
/i0fGftIiHV/JkZPfmqt6AUY/p9XwbCTfUbMHIsCqqvbdBSQr6+jJ25uK0IV+Dbb9obnsEzhIZsN
c2S4K5l78yiYcYkJvF9/02jdVsPY4L1HmFGtJYD2fkoVWphDdMmQrEn4OQOKK5iOV+SLoFQhY+Xv
vpGXARmcYIWAz+MqzCmryVyBv55gkslO3MHQLXgI9+jw5a5oNIrJlYvPuCsQ9BL37A35t/Uspi4U
eYdEfKwRdYZX7SYY+kJ6re2kB9nXZiOGM+ONQOiveawXYs72wxxg7vyOtBnQhgZM03lFVe4ki1eE
9Moj2CWqejyLYTEH+QVTGQ6QD5ZrjXLWZVCXvFGRu1NK459QEUiPEM4oHv4O3KveEjLfCrS5O/HD
QXW9lvcqXvCdmXa6nHrBc2/32nAeZV+ZmrdAmgYpMb2GBPFVy7944b9PIONTf40sd9tGUqTiyPcp
y2IZGMQEmL6xD7mlTnWFaEaYl0Ql0cJFBEmglYs8fiGNbVt9fpWmvKcxCFZCIuuJvNiAbUdSwuMU
ZHAzrz/Nkqbmum1aLxJ14cO26/s9x1w9uAKz76n3s7gTC49Ll7Gn6/MC7ZDhdTKPZyyci2/MPcCf
YSK7eywMM1BDtq1CaZ6NNwjF6cuGbj0YIlBhniD0xBSgykGgk9P6l1DiC/bDcROU1dZ8pr0ulAqz
raKs7oYmm7skRDB70kXMILcihRGSC3ZzmSQpfqTFn2sToVjStI4jh7eUT9mwadC2iMTFxrgMuCOP
E0A4s3/zHMHo9p8mtVbHw00sOuyGWTE+hXk8MaFmxfknrjnkODMdcC+7tlFUwGts4xFUbaOou7kF
gEsnt24f0N2wbTF9A8iubuml9Rs9UHJ6b/4yIyl/cehrMz4pbwyDEsTZnnTRJLINwJYNl/2kbXll
Vwe7bGTnlPEvCVoZ5Yrs83GTcRtVkVwZkfmD6jRxdacV9E59MIh7G0/OW7+KCmJVcMTAmWYZe7FV
GX0yTHh+OKgWvMFOOTYeYH2nDeFEtiGEV9onhChxyuoDXEhCZ9wATLe09D2zMhpzFiedOqAg4V72
v3pXz83LJtfpF4FYfpyPLQyybGBa0ZoJmy+kCgbW6tLugpjU5y+O9HW4YZLtTKH7prAcVbw3oL4a
khHW4Bb2r76YYVnfEf/zfQdAH7DfYKJyzylKnOwlGpP6nHXG/nRVsA4+g3Z3Zo+y/iC/PRA54DL5
sdVCZAXLs2Cq8Smj5BK7inYz8nmfqTl8/Wg49mYfLFkW6i0eVul0rTO8Dsglh7UU0aCuy5bSeY6b
A75n5OhuNaK/XPfTBIlmJDmPHQ5QipcpP9rq4u5JtVCeDTWHrbqCCeBhBMh+AFJqHkUfTyRz7kq8
jViuFWXun/cyaOZ/zFiUSUqBbXA8ZHr5FAR86X9csdUqzflsekIqTlWngpkCZ2W5uAB+qRjslZcP
8ey59V4n2YC3zeMa0exFg3jlxn5zLxj2HQsHp70FTthDe4WCr79xw5/6v5LYVurqSSn9ZlPOdCTQ
R2jCLgcDMoqL2rQego0+Tdb3Dmm98RBb7ZU5/cfEC+ASkVfqwwWrgyp7Ydocd8p1KEmVeHoODqqm
png61nbxVpN+xKSl1gOS/Hjh4fSpvUtxs7jQr+myQVxqf7bAhypqtrKfMX+v3+s7wAHCxF44LWo+
/NBsznZT96VucpdCG0WUrhHqpzj/HOAsPLgasetgldsONCi3jRd32JbvYhCdrQzIOX+ZB/tn1UKn
52Bb192ejFPlU6O4LvrGMqtL9theqy8U7x0wGp6aScRkoc4IRBKKuhvO9cMedCagVz946ujdfmNW
1y7m2iXW10yWEB+LvZJYuIAAZKH49eT0ZvqC1PS1p2wcPcEYQ2Lc7ji+5/eeQLhrM3sa3zOJVj93
LDzb8iSyW2hQaj4oBUA4MBq6xpAcltv70807rgIrL2IOl2ID6edRrrfK0k2bJWAey7v8AbilXTWu
lVoD2j+RZ31cG7e/hOHSzhSuXcCoQJHdbVaYnHYn6fUfV4+qi2o8uBpCwCWgViAFSyWKQu3NIwjM
/1ahci9PvrBTiVazrW9CyGiFxUFL1uZy7m+REx0g3WVBJBiLEVFc0tz7ZtbKh29QqmCVna25kAIx
tB+sauuBbDQvgU3qeqGlK5sGzkyxi+rKv72ykTi+avMnP7VIJGGqMq67IjAk1ZPEbgdstPzhYwhH
VqekLNy8klymLvvSWBNwWeW5UCNSEYaxoU/nQCSJLnwCu9uxmJl21tU+Qeoxhs23AceG8ChNoqkS
XseoNa+b+xOu2MPXAC7XDid9XHZS2FPeNLO+Ys4CYnURUKJWDxg5Ih8VQo4tJqjNcg9r5Cs7unF8
Vhpw1fCi5JogKBQQexeO1JcaALqL0cBsJVm2SKQoA4/MazZyTAlzt2CABnweg9AmmFDyjYL+1HDt
6NcwZa2XjEN0kmStsXayT6Rp0ipkKMK0B1wXHjQY0Klkq7wiblhqly5dyFkgC7jePYi5MlLCJFkx
XhFbv5x1wh2W3A7SOtwKiQD6x+HcpEHTQrVOGBiPsTMFuIYINtngsNdOUtRy3msErZcmTvFF8SPY
KoRFZat49JY3Vr5g161GgQk0BU2ovRbk4E63uYsx49b0QjPgwi9V8sc4eh/WGJFLEh4YR6VExYkk
l8vakiTt7VmWbqDhV6KbU+0R0GSnbaDxXn/IyOk9WH66AmRFYYkYqrJck9sdxY/gsolHoRyojGgq
VCHvkimEv22joVKFPi2oabqYUqT2IpW/hNIccXax8L1MVYGFjanCyqeTws2pLXxYoOK8B0YSvitR
8LatA5wV55HjyqV7DSFRBcwF6oduAHGWM0IDhQdXr1zC8svMgbpLoMuUc+Z33xZ++c/AqxUK/xzN
+bqdBGERjoDwXxo9XFkadnaQvHkk4i7n9bFBIPTZVR4F7c4wKrmfbZbsrIzHpoRW+MWZAxMDG/tL
a4tpZ3demwWmXosuE24Fv6P9l8Yxrgc1dkaAA9xalriv1Cok+X7hkF4+hSc+pU9gKJ8/hTu9EcKm
+kXmwRhzJ9SGFL4p6MRm42+da0/HHA1fUiEdExdSgWVQQdRnGCSiIOVk8ElC0YS74gTe0GMlAypy
Ou7tpXMAwuk7mEtZTnueCY70xhdfBIuy/YSeWGjgtxtNVmVWYzrGkh022lxSLuFZoZmi33EFa35x
8AXO/F6Afexe3G+ozx9gaOAz/x6/JbYmz9NBvaZEb5Gk71xi5jrsR0pUMG4wUk+kS3QTuu1QVJja
NnjstaKiBuXsJ0WTh+n9mALsIGtA3WR+t1duwggm9RSNugaXbaGto5rL4jSJyicCxYLoDSIwveVI
/HXmUk/IqmNLq8qHVnyOR7Qk0P5t0tbwHgbHIopHY8rLnssbcoRnHd4/X4SJRDqMUjgDQ438zIvr
NKMQjfGkGu4QFWcSRm8vFcSG+AIEn8Hq+Snhqd0d9xXRHaXEIFEDgCnhgazCM+6KBYg+aAsJIWLL
B0F6zI5j5vm7shXWD417Dp0uvlH1Vl//tbcnFOl/WuULUazyaF7e0kKJG2HMJE9u/eLoJ055GYnm
qBOHvFR7Oynjh013GDSSLXYz435NZpiytaE/P4u5oxhWvwHkSpsNlhpXguwBRcxG88zaStoweNyl
QZPsWH1AIEt5D04DFcs1wF6p7N4HC/KnAnTD+2iJgZIQcBlzpnf1n2CGjafJ3ttQuqvO9Jcc9Ahj
MVx3UEGvlo4idJW0DBg8Pq0SGGcjDTk+WSivLQjFrqKvuDqvEoGfmz6efebQ8alHzcI5vWR8Yv4J
eLQIfvUTiWNMukHKQMtQQe+4ulicftfdGxgcjZxWD+sh9AUOasz9Vh0WGq+43J2LZybIaEqEwJ23
q58A+AJ5ZTLME4sKLzTt8cFdjZQYXEKFHyf4BHmv8Ph5a7NkrnuJWMxh6C0rISJsHYJ86v1cgCyE
nlfAxK5knjkism2GYGw/mlnv/g97aRYZ85yuT3WGQbUn348epewUbnID4fn9oAsJ5gTlLcbxnMbN
/x5PyhePaAfJsOWTHDIDWuXIpSVJBPNO6AJ2bZ6nygdkoglJR8e9Le5G2ysrSYi5NYr4w5qP5QRf
MPX00sbtLe65rqNEtrk4nHTEWe5E2jTXVPSHahoGmO8DRr2trRxXuhrn4jn/RQOyqAPX5vVLxrYO
J2smFudxVif9QP54kYbxa56UEt+JVYvad1UjivndZZOOzcMxGsk6I5OYJGQTAG3do8JyNPWyKgSL
fptmYXqFFctktPVAIRuSUKBQZQHU7Chr8Vl9XGOe99wmMiuJrj8WVb5e+RbChH6Hn5cp4KQ91oij
P9MHh8Op6CjzsVlO8Q2JGYJk9fk6PnL/jaX4WzVI7V4sx4YLBliaLKYQyW3Yv8niD+phFG7yhhJN
BrpP12p3avE6/fgkQ2u1wKPWls5ENB6WNYQ2n/FfNq6pimMrABh8hr20YflmzS3rDY/Limvw4dGk
QrIukmUwCBvWVHyL0TV4KVxrcMTD9zpW84tW8p6Po6xMO0DbUemixQywfTDAt8wJ4XE0kUYll+CI
JMFD14m6Gp1kMmdyLImwbs3nzIgtzxFu47PsxRY7dNh8iuQMuUowhHVM1dyWprP7S/AmrOoJxa7j
gYew7KeWucvwL56IQGdIujGAOE+DA2h5VhtlanvK/M0ZBs9Raxxn3NhUkLkBz2bNAN7XhEgKjHHK
1wndU62bnBJ12D79tT0RSfF7p5CPUCBg7e3M7CusWtFPWyDWXbFKwRnaYX6PCO6xwaL3wp0sqzWb
/j7+ftu0ILO8omdevFiPgam6j+5BdqxOo0azwcLUMcZ5h0zsZW2vhzA0yasNyx0e59JMSTO65RCF
kzgDhhtxkrpndlZw3e2sLuNsFDO+5utNLDhEQdji77n070IaYF2zcpEn9TfadduX32W/BQWbdzgu
2axyPtHfRX+gNPaoF49qx9QmQVTJnId9npqMVJI2pV9JCTyX7ZhXNG71ZOEuNGqaJqCgR8SxtJTK
Imtc6bwctwKWEvGXhH0oGnQJUef6eK9Y4HvX6pkmU5M9fAvGekO3opLTP5wnwJy2TZ9kl7cQxopG
DgMVhLcTF4JISaLFtK20q27Vb2QItB0Nwet4Rq0siDmEayIT7JHEWPfMel09NrgRUtFksfDQzEM7
Labk8gPcJ4c4/Lv7P8Fag4q0XPAtlSA/iWqkhUjbD+8PL8h0TJThR/LF6c+NZphR0LeJWWautSKt
6gxq5a3Ttg9AAzbbs+Etqkkf8zOiheXEwtt5p5UGL78OrenRLLR/vvLR8uvf+qKRRuF+mvffyuj7
e56otcUmDHrDE0cTlfI0yoZlwUxwF2Ewl4zIShbdxZl11SGVV3Cjr9ZlhOZ+2Eyat9MYuSBVYCX6
hh8wuxIBMUO/QmYfEnyQeN4a4i2AIQjzlLmXdd1yOu3hOqeI0TA+0FgHB5RmwrR5DAQ87w68DyiW
np8EY/LX2Gb3nO/sQeMmN24+IqSvQxyQGNpmGUuG2xnUTOqgTDkkG2YfZ51tRcD46F7by+4uM341
2w/j2hU8yZiwgbYW1TPq6TVk9PS22XtkNK8BPENpmqwu/4uXwIAyZXHDN7qEZ6aYPAd2LOq1RQcO
hM8dagffe01X8h54Md6DNYnbUPONpxqirpPMKSvRLp1TJAtEJ+KVvEkB340N2GfxDtwvVfgJm5y+
OdIzSnalD2mxmfcLecTRzV138GPHGNY6AYxhl6x8V6wuHSyOF30ul0TBpID2m7YJcUIkeqStzCTO
vsBYSUSyEljRXkFsbwXUK1uThCSKOyxxmYx+9J6sTcquaPuPnXp/22NqNDzMp1UOLQgYwgYujMAr
hDYfWDKOwt02pCHBG3NYW3pRZEBTecKlgWf6c1A/4sfZf4Ad1QVpT+0ynj/TKzeW9Hw8NFiMoupF
JCJNaMJw9I5BGt4zVrm2/7/xpSiPG58IsC4nqsGNSAgQF6KFV7dvLJs2MLwYAZF7P9CE1jsokiii
HwhiTApHjS/I+ALFNGsdZ1nln/j1cIQHQiDALuthEzxhjjxVTjrSKGVltLdLv5ki1oDFSvhgENq5
j9shqRU4ni6QMokla4LmQTn0ihvlJJMq4EVTLXiAwlTwR5waTg3pq7p6Ucj6MGAVgX9WGhd0JPBx
quZxDRU4AejoRyQLiKFuQWeLn6En8UZVA4/T9GVbfFGaLYc+WV7PywrsPZoM/23v4diS+PmTQOz5
K2eaZ+Vo/FAHK57ltRQqc2J3PdDbv8XGFSTjJJkOGQgR3jZsiufqN7Q6Sdu/Ew87TrL4ha7g6PXV
72UAozNI4WDnZeWlHcxfZFLdpau/qlF0zmHdx2QAyXryywrw2CcOuzA3EaUrdsKn2dZU9Ar8b3xK
vQJR7gwbPvv43eY+xiwzxDIu8HPOaa2D137nmOCeFIqErlPdpIQ2qnoFmqxw6ladrdrrsi5a3tDP
aEUNFRi+g+38ITu/wzoxCS/1sXwzyZF0v3vxiGhF9MFAmCp5CkY+A7xVLhIOKxEvVY65r2t8swZe
1GyhYYK9JYkbxPZmZrSA4VYLl4HZ/AV9TQRpxL9fKTV4i1IfPqClLMyV6CzweOpZ79QcOgZzwh4D
4tgXscKBLXIyx55HedJW39lbZunb9KK2Ea//ooMxsCmCoeS8oc0lrIH3VRwu8aHqTDa+7VMyrWyB
ExmDOjyyk9ii/1/ruoigHZKMbauE78kfnu6ZGNf0xtw++5G/zOxII3N2vn9ZxNbhKVqGKrMlpl0/
J1EF/MIwwS00DbaFDJ/L96FAdw8GLy4HEeltRggERv1vc+8A4+ZcXuwRHT8P+02NvCmLY0HK5WOf
LdxxlYeLHZmjNITMgbmZ0gzN84QfjpRe/yn2CLlbZ5J0owVJyY0NwY957h1OTh3cRwxfNSjZmV2Q
4tcerfguCZbkvbQjXLFHs3wAchsm6AAmlCMOfLAPDe2Qv92gYsa88cUAfrb2gRibBplvqeYH8FzF
6BCf/xW14bgjErL6S+slewayKo1VuGZ6X6vv9oEMTo6dcFA80GmT3d0KcVOD5u5UVOa1n9ZNpIhz
tusUgjdmlcDmuy2XKwygcLzcvP6JNryxW/N3UmD48+EU+uj2EKfFUqCjtzxttc6frAwi4L2Ikfeg
52NamnHmfilix3dSAq0J3k9h/kaLciX9jeHINSHJ8zxSskfc0s5VYCF7C3+lVUv0WZ10DdGk1NIv
mREeA8U3X6UYXnE23zuEBMVlhxNbwwxMPgR4K2Ohu5vE4gd6hU4r7PgTfS6TSDE1mmSD3QJczv0t
gVLgUafioAHItQZ9WwPAOcnekAXYHkI9pnW9ZGIiSNwiX2T1tpzteLhilv1xBGE6265UTgKqURga
QRsFAyFohJEN8tvJGGEdlniujR3gls7nj0NAzqKCIQLR4oW7NTMIHPkUcgGIVgtiTT+aIFytQ70f
bNn8J9+1L8VGKVimemi6hlZ+hcblXNawkn5BK/YXGXSnNrMAM8fvgpsEsSA7PFwvTe2uqaTayw1+
7TxzqYaj1PaOjXTUaZcdsnH0ocXQ8UZ35TboZywObl9GVBpn9Fw/J1nyhJq+I3vm77Wr+Ezk11nh
y2UtQlr76V/ig2NYe3Vb74ykKNcxlDExPKfuglPWzcHuEtP6MinMuobIvof2MLi2aQuHjgDxUsEj
rxpeFRO1W0OY0jKZo8u6Hk4uT68jUZdz9tXcKfIJphvRCZ5E+WOPHRgqRuEroZhS6qQYkabQPmDs
NlNA7Cz1I8Lh7UzIoY0T2orGzOz/JLyc97DFC/OwjuDCYIVZg9t0wUgPF7OK9RJXW9CzB/v6od1m
TON8OGv2bToBg+LrZrBLd3kCC5khXm46wL1OMwTmv8aNV6PED87aUsKAQhHEOnADRLlf2k4aVwE1
sKRryD3beDc2eF8WvxXFqeLeEVWNzinUUA666kG+uoa/WBXXNeg+mwtg/lbR9X4HmydscUYr4S0E
O/jS3s6dwAhVm1q5TCRb62q2Yho635oaqRHobbiq1rEFBgwYItdWvCZ1qZ2AiNs4D3hD4Cg1i9Pn
VZuRYSV5ncfOnTIRasvqk5uPPex2w09jGiHTA2CufDmD7w0cmwVAAJccp5v3ugxxEb4UbbZ69KPj
gCuXCvEnSG06wPNju/4KXZWqG+ah8ObgGRiUtsc5d7zsnwL+WJhIx3btheSqlM7UeClxB3Gck8j8
iiBwhVbTfh/GbzF6oJjK/8ryfSX0vejAjwct1dUqSC0wLSgL1x8JiL/kOBKsv/hMI6doXLjwLzj9
pDygG9Pp25U94NSr9cbgjOH/qw6ZJdS34rD3ySS+DGTxp/LIOb38Y5NGm/b1DqNxVZk+AcBsVovC
he/bFM2dQnngeb7lLVa+pS6Q4ttZM5Xbu/UjHjEGrT5Zj03D01K9jTPxZWEVJ5RprKcyZWtZLvK7
iAfbRRqualvs/D89/WQLA/avVjHfaI8S3lwspu9aFw3SSSidX+Nd/rpkygzk1+tuFvh7EABNv7VZ
L2SObICVKbcMGLxXpg0bpTpGrseEHhHILRtFLSKTxkNnLzS9nv97u/aYTpoQN6rS3YFOZeOq/UfL
0Nk2CBthD3f4JA3adR+UbvoJvZcV4crf6luCYMrwOr7wZbCYV+TTHXuYhabQRfjVq6TwT3UZo2Ts
u+P9oamKjApGOsfAfWuedEr4lcBHXA4YrPTz6e/2dfTngLfeEF6wSBytmxTtAckhZ6NYu3V+olb/
4TJUtUnHqWBT3nCSSQCv9OCKWzeHZYJSV95E3RT7+jySshhah1w655mD/xv6fsKmfFnL3JYN1MJs
+0E6b9nQHSVtfqGgtsJSQRiEM6FG/+8mqONsw6c20lkiBb1N1cR0Cq05MYP6duN0JO3672dfHoKM
o770T31EUlCb9X4ceTXUYM+QOcGP/7BhBAm6S/tI+IgaJWkxG/2otrDsH7lEOrt5Bpp9qFKuiods
VmXLWflgd2s993oLWoxeBV3WpGf2uXx9jKyA19aOUdnsAzM49K0LFkt5CX4jeazFSQp1NBzlZwdy
BPS91G9JUHSlzihQW6bVf5FasqbVTkvcTWr1dC9Wf+0NqgykLQj0pY6gRK4dT9WbFlu5nB7iL2Hn
IksoeK3fmpWU8boRFNjjd2priLMKMo6LsXMY3aj+6Awc48YExd3ms5TyF0l5q719Q6epF6z5O0zB
4v4/yz6qIg/z9edaczRnbg5AmaAH8pDgOUepfTaTlEAEJ/ho1wKI6luU6wA+D9ESKBHicvXnFrt8
xNnEX42BhDUslxLkkmUpzaJrbAVBaT4ohjt7H9pVJdd5KHxLob/IKP3BCsYFgF6sxucN9ULTxJde
EVWun2RifL/Q2xcOiMVJ6FF2N51WVLllahyQVHuDX1Ow+dRjZaAAEqJHURUOyNQK2Zj5+jKvx1HB
MN1+pe/DA7q6EgCmI8VDJMYxKzEeUpfdCVXkNfWpGTF69W+SVBX58gO89XseufxrT4wlmyAGElxX
v0rfcTPPJWrAbzC1s173r20qEzv085nnaZ7bUj6gspmsworAz3vltKXHpWGwgb4IRkUtTORo5gVT
0Yzjp5hjDiCKa+kP0YrMO7dC5f8fn/6v7j1XrfIHEUHViKuu0BazlP32TSsxr00QrO3wyiovKieY
crHnzD5eKqP0t0krApBTLoWRMv6gNp+081TZTsOURmhwTmUThXqdNqxwfYHSyochZEJZ8J3Qf7vq
fZXBhmop+nzyBKyWlb8vLpsrzDPT+pRTE83L6DzflzUZqLoxS6hPhJgGr7ai+L+TOMtuoqR5yvt8
pjax7jwVDWHsK/zyfk/Z8Odu7uWhpdZcSTQFhwuoSb4G0YdJ4K7cUkOdtc5ux5KXXv848Hp/B2A3
FVqW987HVtp9HG9zQd6dv0xKrfsEj52lwL/xeHgZZk46M0VlTPM4Td1uU+qyBuaEqfyjr6bMZrQj
vg2R9UPrvlIVuQHJO1OzSNxJJknAUvILJga2eKCaQi1WUjhNAote1J31mwzU66iFWhySikFHz4kZ
/1TO+m4SmJ7BLJKzUaj2wWUF5E1p+Ox2aVSigxgxFKbL5MVsohKIadC2p6tSXVzEWvy8/pUnJ658
d8FXSZI4i/rbnx7LzRizli62tyZEYb7vAIns6RXP7sBQQMWENO1c4bltMP6trQKgeSq6VYwC6N7R
MrgxNr2CcBA121Rqqr8y0TBEyh4/R+dmHQUWc2ZBizRoqMmLsW5lRbWSVWLot5Bb72hfcUc6AJCZ
KQAOYLxxxSkj3EEeBF+huGfSFApzRVRmKelH6a5lghCzCxzw8MkBA900IkBlbru7+gTHbGGGJZP7
Taxd6cKPbVp3uY3EMatYcwvV8PN8TFToOXixG8OAI0Mtitr22mufgd2awj64BhkLXjmtm6JrG+8e
/FN7ivIdnfR0nnDeMSMQXkNFWP+D1+8gFWZ5q/SRgiOBCn52TTanazj6Cs3doSGa2qdYQILswsFl
i4jmOid0BJigYdY5nvSzHAADEb+OKa7vaWUIHG7Hjl3yWPJjHr0bpQVVjR6f3n1UJJ/7b9g7V9a1
/axYRxhVUe7H4vlr4Di53PLP6O+8bW++K60HuotP2h6x4Dv0XVFa0dJ5POZS8C4crzjBr5/3gZWw
6bG9oM3FFChCY9DSaejeAoWALPrzefodo7eci1HaSUXLQ703YxFrdocFDVt1mkEMqt8wYL54Ns+L
/RbycgXC1odJZ7bizvdzdcg4Wfa+8g1b7TAS4uznqqW+u9AhboLd1hjB3OQXL+ICRoA2eZUn2dZ0
V7HpywP1glcpfRgOUon8HPDDg6pd04Upn4Ev4oYmNJIyTes4LlK7MKRmfQpqT9YCYX42bJvZLnzw
naSwEuiWzT55y1U9e94wN3wIzcToElU6h2dDAi7Jc4NAcCDl8KmX3u4QwdZAxVEFCd25wEX8XHV2
nY4FoWL3pvCV15nXQpDyyT5anq/17I2U0DfvE6cf7t+45HrmmRtuXqK3P8qhVl5aH/xbzCtm0JMl
QMDBT1z9xu5lCC/nS2b+aFgjdCsYMvgDg19xJ//8N/DZHQqKVn/BW+AjKE2mSXGf7y4MxMkRi7fD
PSO+83C8jp/6NXuk544VEOejyADv2MDZ7tMdeX1bezpdmzjYh+SS+X+f/YXG8KLl0t3l80iC/8Ao
4t1lhGabJ/nvd49H535P8SbVnIxEfrsYLpyUkus54XVzuLkxr2TKKWC5fSvBmvSFjGMMTpFEJEmZ
oP8g1jK2+n4GcsU7Md6/5qJ+3Tk2vqL9Dyu8hsogXCsfZX/tqQzKZgU3YVjAEm7HX9IAHNSNLA9+
lnZxxE0rV0mj4MmsOYKulu2FeG6b26gHqrp2kT0oxrjsR60v1bjgCaDaGY6yfwROCENUzfuIH+oV
CWPvp45z/7VTK1PBv4dn+mQEZVjO3nUrqQzzcL77ulhfIqHRVefsoldL7nQYGLAyJOCf+lfoB2i5
W55EIds+H8l/r9BLCCk7XZm4H08cS1aMHog5lWz5UJ/BZNVgZuGS+7LsQ26HnScBYikyX/YmlpKX
UYNrSipVZCx2ABFov9s9ljWhNlMUcJKj2JWwXt6DmrNURS9VFC8jMA6HwzzPrJiIKLs4edUTz+9E
jDbNbqTINPAOqzVgU9FUnaYInq2nhvxA3jU9hnjOuJhlTyeXf7mpOpA/uS5HChieoatiG3Y0WIq3
IM5Ez5Xjnq+G6wV+c+JbYvk59I5gcroO2P+KqQtP3FNklNQ4LMwwrzFcpzZCrAD42GjG7/LAF5sm
4sRU7Cr2rf0oZJrVtB4kXQsQ2G7BmZXrAoZJEN1r8qeeL7K6h/Fjs2tqt99JFUwQdYf4qibRWaml
VY2PwAF4HTVEdEheuqibB6ickrZY257qljeT2YAdB+clFnJZEg/gCvTD8nWbksJ2BQ3T1xYkv1Sh
nY4X7pTuH/7xjznlscV7EBSLbloxXAP0WcyrGLLfoU7dxpbhSyGKtHIffzQ9utnqYNkB0TTgWfcV
vbaQM2xzNeB2zd4xSXUKRB/mAyb4qbjvAlMFcxUWE8l/Y2V4xFe96j43RyaQ510GB3yraSNS1kpg
exXGfhVnflG6YYa8TmOkgf1aFfd+zX02nLYvIl0AdISsVbKU5aULvLdrenI5iXFpCZZsomMfquqo
Fidd0voRRNDMd1Vf9HdyoIZf5o+BsATKdeQ60CXBfVgGRvm1iLFaNWOYcF3WRRVc7VvwCrh72cwj
AdDZR07HNMMCsnPrTUvDKvKHaAatj073Qo1dRbks6sbCEtbsuB0b05uXQjdk07Anxbv9c7WNYHCA
Ff/q8K/qXGAVtlOT1C6fGZ20X0lJtfyGEyWIC/a7EV/7rTgtwS1txcMOqwO5nspeJmwKtZTcr7S/
5ag18yXehE/t0BMwq9k8NxheGr80w4T04x/J2ax0I9zqrzYu1whdmzyqL5pe5ZFH0UTXC3XXZ9Ml
x92/BOIeLlQDyBGq7SlabpbwHimzceFBoDjhhbGUUbDeAeFAbJQbdXOaDVjkqX9jcVfsQXhW/FgE
tWIhGfgxKeHj9bAXl5AvfD2eUKFmnzyxiK6gnt+dze4+rhIu2dFBZf3Bx/NNTJfhfjfBd3OOBcg0
wlOO4aLR+aQg7tmhxiCA8JWcBlVDqT3PwvjkIcAP4k3iCBfDWd9TI0UY0jv80tkG93Uy0nrWe2D+
0wrRTCsIX0T/1dfSqSlOP+iWdRBLypAJrlngH5laFejjKZ/H/SvP8M2mc6kJzKekoy2gdIEOcAkP
nsUuCBry9hjS96VLs+GVsHrCQVmmaKIBtO+X/n/hJhZpg2HFuuz4rXub+518NKKWRAUTUQq9oJeR
7zLNNuJkGpBPqRIUBlEWpd7SRTgWpEnMNUwH43jQ4XrEy8AFx5Dmi8hxFz18syUx7gBDUze9s87V
sVEnypmOZox4K8a1dT0S4FdyG0G4RIXVmx9es7Mm7A4mr2+ia5FDVXfxZZzwmhE6CccRls7rG5/n
myv7KZUCAMy6+xDuro+Bg5nmuvLcO3r+vbn5+/bo16VfhCV6zCh08VbUXjg2lmHhrpJteHuE73bC
RFSPFrisQ+4XEhWrWhz+0bRmfIkvDWAJ4btFIIsEV0leRyRZV/oarqunz0STuDwUvIh/Fvq7Xe1p
3wyHXy63MsngS4wDICQAJzXM1v65fT0x2xnWwGKN0sU/ayeLYkK+uujrlOpcnZWdZo1O3DLYzRLp
6jQpp9ANPgQ1j0VbwMwLPHsCHpp8nsFmXaJB7XUMuTBiyvz1xC232isC2arSSQ/ekYldAqnWNVJV
hhkJU1CDYLWCu/dFKFUntZePlb7sWZBbsixaoJK6IMm9XEtGv+X8M9XyCK4P8LRvDkR3q6UfjflL
fLUNhEwZDg4Q04Hxgg+mytqf6Q6EpymNCmqkq1uttUKGT4SMUOibo+PKcC5u+51TzTV8iHAltQnS
k/3g6+PxdlPLE2EwzdEo0W7inTTCIVk8q0obZ58L+i+N5p+rL4GwwhG1E7uSv1moembhsGfls6Si
axQKE7TAqrUSGmBWpDBilN8+Ur8RcHyi8a7TZv8M8qrdjv1YpuCnLP9TGvgnPec8phF8UHojDOdr
INxXpQOcUJjrfEoBDV1+vshTq/SdzYjoaC6VTXs2HHufUJhah4vvtCJzmLFATv2zBDKehHmBCIcG
e2rPHbgcLIKgz08mvfUgB57nfyvzxcwIN7CaJ/bzWnnD/XcZjuO7YPvttRAIKjEKcjeVzRXSshnZ
YAh/g6EY7KfAM+yaftIXTnutpsElBad+/xBGsSEPIrfGoSXTQgZQZqup57zwuVkJzgthQ57bENSV
daeVAUIAOUvZK9GDx3H4kZA9G8LwuA/z4kyKLk4OHq2GW+rJglYCaupdPP02b6SabimNmKY/q+qo
vcHLtUfRJPGH2qdCIwX+FGD0yJSAj1w9JR1fUTxQTxLTYxZEB/3SQ5jzlmhWUnDjC5oBn1N6oF/u
HmN+K1YMsFdX0V+z1XB5FA9Boj70MDQ16GrjXvcTaUDTxLjHpXJ65fz11UCFQ50K/rJ45NgZiXCS
OD5fObJKKSRQDluR0K2n2y0v5oSX0baiKJpn82YGpgUW+VLt2c1I23wS/irMd2/5Crn839sxxKRd
0Y+qUa+EC1QBVJBtw9HXxHlF6QkJJ1pd85i7TVLWlaS7fceSpYqwVR1RfglXrC/Pvu0aHwwSkfSU
wvwu4jKtSR5UTOfzjU0++TtHpOrUAq9f3147zdtHr6wDv0RSt4NQckxwVzTrS7F14ELW/ZNLitsU
PJOFa+3Nos5Fcu0+I1vOD5mHqmD9KjIrSA05926/rWIa4Y5i/2kbLTFCrLbQFaf2haw6EuME4+kT
jo78pi/DrAVz8KhFOFcNOpqP6fTOvUzrtGjjZb52JVPzR1I+7j21xpukzPbqduM4HEZRZ0r8460v
HHDJ1pmnc8UleRPD3g6YhavAcQXEf1+7DIbNO1+hFaqbDwMyBLR6lSC+59Achy8/KN8MOv/z2p5Z
fBP+Y9erDcHnWl556aGMfy7c0P71rpdM810V8InQDpaBK1BtOzfmiLl0AGT9b2adsopKdT9Yskov
pVw/h3FrRowi0FGUA53oVI1NCOubYPByf60RprrE6b3nvxOKewEtpWBmODgjoL34r9M5vqh64pCw
8naVEoYcNZqUg4FpXJqDVvYz5ySBD8rgJrqgwr/LfUpREbeqtlNaXoxD4zoiihOcomSWsfXe1ary
X6dvKLFRTtWO2iRuNsPNo7D7T4rkqMiZoePy0O+Az46C1Pp4vkULwmqPu9Ue4NfR4jRnAXvY1kXv
9+x3UgbWQNG4jQFCoZD3VDreuQvY73Jr1K6yu0QHWXvO6AjV88DvL+pmpHo5HKRgI5//Tr5yPAVK
VlbN2CZ9VHE5pXxfdt0ZNGKUwB+AZmaYcQLw5Sua+EGzxu3ThSEgkI5OkNBdY0kiU35/92IaGEHk
yR/hE1t/TRkToJ3cgTWFjQNWOjJsVMv/JaiLKeMYVJQe+nskNEGquw4AjfW+wPzaJB78ChRCA97y
UAozmzaJgBcNPfZS3e1jSfr4/eOLF0SE+WZI+Vhc6zs2ij6xyLXkipnyTnPRsE19Pw2ASaYFqJGc
HllIf9S2j0/sbumLhUM16Y0720R1k+QZ6i48v6IRNdgvCRUSzMGRK9KpRwGx7LqA63bOXzA5M6/Y
UKZSVXQOHOkNpedkvluLPZdwAn64Os35PmZV5xeKWkxXZMzvClf73kH3ykTK8R0mdrJ1RJxTr2tt
jFC1rLkdmVBUr12l5qpX1mnbs2/jg4flKUQNF/R0YMY21guyOCiRhX9frQoX+Pfyh1yibpsQK9FH
Qu8EGCFQ1hJHfRKUfexWIR+oBFey2Zj6wH4q6MPls72ESHblj0Oo6USl/HLn67PvAP9k2BXetVq/
wdCMJAxRGCSIKpJ3AUSCVJdtuYXZaUUCfmqdyQvZRtEdeu3rK2TQ5YKc1XjDA4wqk4WSIH8WWvG+
2dJzrt45GNecwJwvvVZkc/toiNZG2gwfA7P3tJ6Pl6sWeTBvdSllHSa+OV8ZcuFW6oD914YivYvK
7hrabxi9W6S/JNKTpX+5lKrBpisM6eY4bUImr5zeR7XoXDH++qPWaawQvqbHCtP62Pz4Pm5XIIbx
5k5vUUahdajG+1IKc6XhFqYJpoZjofUvYl2IRYVbIu/H5RIUzPbY8lMa4rgWpB1jmhC8XHp4hKPS
uFRnTm7WEEqaTBpw/tsF+Z4JdMwd2qtVWO3nzCOBQzxdAwoUMSXyJS8meeD2FsVQQGL6cNihYRdo
Rth6oKVzknrJXXNrk/vJceV3pRKNS3yUXgp/ZHcIabCNG7bq0iZnld/Ilh2MYf4SETty8LHK5nyb
kmzoYYkPWDt8tIGZj5AiFqEWoEglOjIE574+g4sIjrWxEWTJ/88U3wzX9+tF9JsITsxyG2QcFace
3oBXXXKDd3uVN0ppFvBQDs/6T5ZJBNp0CEOhiyHmawnvYTu5TjzWkSvaELef20uY1kt5Zj8fBEu/
bH8dB0KFeL4Ykb8PUR/rloiEcbXAQIWqVmfxKV/XyAvErDf4a03gikl73ZPWszJJj6jEEISwR3CD
PdASXBbZTPX5uRjrc0yq7niQK7mFpPsNSqFhG4BqCXlkJxJaowE0IOq7zJcwOpSVacsjj8zUtH3O
741mgBrwLaOq9GCSKy6wxlUvVHNLDpenhCDwDwCeRau55OVghOTAFPnOYh0hNFSgZsen6t7UTlka
r2FTfp1pGfDFvQuLZWlHxhb7xLEkadAUTIEjZAxPny7fzcas9yEcoVHqkXo9Kl8ZcJp2HMJYetzx
8nw4B54kWBtNNH7iLDM1z/JzEEstSaRgW3zk12A29W6T9R5pvP6OLP1IW/kh1XRjVpaNcI7tVnyu
LUNE9Q/XbLMT+uitKpwsGsrVqACpTSkwTEdF0OuTCoBg0mEsXaaekBAa3h0IIp/+2QBaOyF0RvpI
2S+LnjlHVs2o0hEFNSw3OADcxlLm7yZmr6q8LgkA6EK9Dss9fu4NGqkZiaNoHfkz80//apfyTL8W
FDZ8DrawiCZNREPZ0cTvzrx2p4VJB3lAlo6uAZ+fyNxW2y5ETZzBwlXofomLf1BsF5OknT/CW3p9
4chEd5m/d39ILnx9HSxzEZzbyMOB2awT1Weq2yLLB42w+Mg5zAuXubhSDG2PHJLTbt9vj/YyXpP/
iCiVH/7S50n+qBzkeOVUaAG1KBlPeXDdvbDyPgZoK4TRU3yHT6UDUV8JlqFdZQ1/WphT9Hn7IyrT
18wDvnjFite0ZTdtau8iXxxVAJWZe0kt7Q+mYquHn9ShC4MDTRJEW0dgHj1bRzEmHe8T/iPu40OM
aPs9/huIK1jsNjkVuokk4gG6Lf73AwM5+L0h/I7V+46W/YVo56G0qQMY0PrbNm6dr/yBVFhbjFNm
M4NapYRTcwKOGeRBeYgT+wnu99sXKnfaE/nurqYplwy7zlI14eZ+gsGpbFzmTeuf0YU7vLJ06Z01
kNcqHYquaG1pZdBUQTcl6YYSjEaL5mfEpeQpYUNvddv30syGQSX8c7/6GcqA/vObQfc7BZNZCJvY
c0ZYtD4FAzjSQTf+oTzUFJtMgtDpydEMAyjLMI81Y40GtdcSrP3Q+Dj+nqee9W5/LCtgo/MypfEQ
2g0c25qqgk0AFKp7eXDuUCdzktSesQ2i32G/VVszE7ztHieKaefr9QjmuSUjiYZE9rsWV96zFfH7
I28MWiG5pVIKbNcXO3ZYDpXkwDT/N9SslT5IMxOk9DwdwEUT3ko+xjvZUBWzQO3ol7ZMMreUNg4X
0xZRImzwQkrmySBAxe1bsYpGBDAi6vqxLzldEgYLe6CiAE9JNji33k9xbFEHddRm55j6HKsw/FXq
JyAT31hXy/kplAAMxxifGxfvOWpHK7/4qHc9mGMjWJ+VxguRSP9Hb5oQHTtjFoUatTb1mnExONCZ
IuCTXLZ3EDYRM+HWjfacS+l8uZTfJguxR8bGDWAqC6RANQocF09ViKM0hwGG/lOaEe+cseUPRJSL
2GV7hIen8kVnr8rlE4qOfBJFYRAK2nty9uxY3U1eQ5RfSIvSxpfzCMIokRtGCAvBjhwHq+AeBw3Z
Xwyj+y+2Sz09RjebHMS9zFm9OegaaJLJl1v822u9XYawpt+ODB7nmOnHjIMrVSxqVAPn7FYDpWih
vmalPb4Fw/sU3z+PkwCdeQdumaNy4cPxwsJUBjK9xmpKi6VdWTu78whnwJG8sfgIxqZA4wWu9HSV
bMb/8VIl65CXcjZ5mVl7G5C2/9xuxwr9jabUVSQy7Le9Mln6kitGOJpZT2Ef0HCydbKYXLEfbLoI
fkJsU2jJcWme5bYWx6hNrzgpUan9WxVFP2m9e8x/3b6Mrk4hZAWXi61+fzBfsNn/ATbsfbJgAoME
fqVihDliJ+icNeGAiUSULZ7Snhso5sBtw1Ugm9x8hQn+Sd1QYFEXJWw8iYSWxPdv2o8+2q/vUx14
wX6rxu5PKAR7fyEL0Os3VtlmREjpoYw8YjGcRCMNIvhAmdsS9lbd9y+45DepETLtolcYvG1TDbae
bPgVOGX21yDq5Rz3FeU2kJyi/eIVCk450ClmK09//tHLZF8x/G8tcxEFs1jVTbqz6pxNY/ztrW11
5ykj5dW8qoxQK1Rpf8CaULHJvroXN04PZ/Z72JnItr7FBHqfnkjFyvP/Jiv78qmfPzmqXhKAGHKY
RefUb+3TX0Z5Iqjjiqov2Pk/1GBGpew/kjW+Clm1N1JbQUvZGax3w12JONImXhfDMKG2aSM9Ngoi
yb3LiFQPaAX4qi+WL1fUCw4CuI+QcFWeDVvokjzQuDJ4UBlCm+HMdn6bsYxxc+RqPYsIx46Y02st
Q375SJumB59sy+/9C2dHlrI0uBC/zKHCiCiCq8AKcwT9gDLWNKQpBHcbdzubqI+4qojmIobQ5zf7
YOHozHew+Lb33b3vMECFt2ToV2XTfCV0tJxwFHz8o9y2k0wLdjWpdmrnDJ7DHbYVnkYmlRE5D8ay
TjPmK9RB4Nepc6BoT2y1Uo5CCdym/f+XAuufHdB1pvOcp+cytPjQaUBqCztOKAnVMdVZEfg+PSNm
ijL6riIrC8qn0+4AjEvkZsb4WDHMJdltWtD8naH4FAnut7aSmiKA/ufMcH4iKefFnNIa06RcyTrv
oNWQJ0ZUyxSAG74JJDozVC6SP9RMdfHgUgM7hArC2PnAWZxBCTqzSrUQjyoGwxD/OqBrQG22CdJE
+0ytCCkJlzHKzGYoTYv5MKmmSV298ERqYR9Yre6GcuyZsjqR/wGh48JTdaHVNB/zfn5oUBnyh9Lu
tkGT4hEXowLPM7v6r2r56CIjW/a+KXoe482FQl3kTkUuCh9UB8nz3PAtBuJ1y/ScD4NCnfo/5u9r
alkqKEb1VjKE6eak/tRTkDhmLrRdFe8JfExhGquqIzaupmlTBNRPa5kuswTsGEkSZevOINgYqpNz
FApCDYVsVEXQh97DIPjhW+oGCiqm6LRjTHvVu6A1BYlzj0czAac034t59zeJLKcZ8CxNzm/ANuz9
9vODREZd2tDxQEtZTlqYaJUP7GsFv5CmNfk8mWbtNo47BWmxjoG+MXWpuhWKXYAUdXiwci8aeuez
GeyjYmXZOHgIf6S1me9mRnPZYZZjTlN93RM8N3YI8kWvM4r6DRYMDIB+Jne51chnTRagdj3z+/c5
I0WNHI3lBAu0nXvTKAhLYgmhrH7/xPy4/yW6BGs55Oh5pt8fsIVjvIYnGV6sPbKPUiTLo/Y/VNBe
cACASylo3KHEk2/36I5mOV2iwjcvoeW5D1VOHFnE924GW3LDM8rEywqBqh5Azj5WPe/xN2gcKE7I
kw9V2UB5GmDw9nJr4rcmiEsPlhiqoO1XjtwZ5OTb2qXOVGBdilTaaaFMYEkzZHc1maHcqAqEh4f6
wJ2x48xv8y+XLC20/KWpqo9osRXWJ3YQj4hctx01j/23hnTq5bTmNsSnvLMRE9Nxh0+ZPRUzIsNy
a9TWWCvAktqeevYdSOdV+9r7682r8TKlx7KDIWzwDm2+tKch/AUKACXwE/iNY1ZORS7lhsEmP+0O
M0EEqFlYomYlMeDn1jeGDSmrKThVAYi6MbVuGAmFlmW5HIL6O4czVKlU3f+ToyfPxBwRZlFMzZ/E
plWe2i8XZSI0nsQH+C+Qamle/UQZ8Hk5A0V5vsV7l9PRf0J6Nm+WVhaMuYi6IwT2M1O1SlY8oGlc
fhmA2rXBKXTTCWX228QuXBwd1/zNLbnMSGGzLBWFIPbT/VYAaFgvQPt1UabhC+pJp3yg0VkDrTY9
tPPge/zI1MElEWmriVUsyYBroYesTk4e2mKbcvCm93IbmbT6bnONzBR6LRcbDOGZiBNKCoFnD8Bd
2gpUUzHJflwUq3iPoSnjFhXcMJoYxHhpt6xVV00NsxI0SY76YBWXTCGJu3+woQMxF/r2ZFBAbh9z
s2LtRubx5NoPVZf00b13+zGke7kviB7z1X31s3xlZoBz7vrz7+aNyOkSV7Hv4QoHvF0OyuER+9kV
jCAmoTtzC1zEM9B3zHv06+ZW2xEqVVLXR4Is3YzbeXeaDQnwjiw1Fy8Fov7+l/vH3ab9HsadGn+v
yDrViZWLowB7PZH1kDFvgI6eLYEoEoPouLClBN4vb81nL2W/iqYLzhXURwn3Hp3bWvaIqmlUTkhx
Mgf4Hrku0Alujh+rXKU5SkrOp/TZ3oow3jRoCjcvP+86Q96C+tOiPcD8qsoZhHrVFm1AEf8x9sBN
OV+n5z0uHG8UyMa+Bd/Ttng/SwrOWK5fQgVGWVp1xtRp8TzUqDljQsvJZrelIaaZ9te/0dwpG0rC
AyhfHtok2iqDGWcZ3THYsPBhadKxW/fAuKezhTvAncLqXNIOUVAtdaXJlPGiDUeyDy4MhYAswBrA
dildy8rWQZNQaTvNfIwSEtytDHNbIkrPBwuOWIJFs+lfx+GTZ+pKrFA8l8B/tdfkZjeZvCpI9oKW
73LuWqp4Nd9LnfEC/D6L1QztcTG6cbLML5bkK2JsjSHb2tKL+KF3m+IT1JtJh3+ZLwle6+gpXEoV
S6vEOfSHz5MdejY9SM/mq4nExUyz73enIZqZU/rzIBxSaAZj0qoDB8anNWgbfwwyhoKPpG0kBXK6
t1/tSPOw1SdYc8RYlSSCAwkJL74SnlOoQhrdc6fBuYsaYk3nhnUY6xI5FYAbZ1QLbVnvuml8p+uQ
f4PWb3m0OTF+TMmSWvmJ/R+qQdksJplWxWsMQP4+R8SwhTu6igKuo+YRvnGSgc6rUoXuA3Y6UwPp
5Kxo7Nn22P0Y0L8W56AQiyaSChU/zwyaDFww66PscqfNxkm0jqz4yTCjHE3ed94rkN9DPo3V4aOJ
zHAcgqXDpuxuwBehEo5Wg9MScjklab1Q48OwytYuKGw3wCE/i1N4qE9eKPrD4g6+ojJmaWj5l1nG
tcprD64EyNmQLbZtS7Bg5m4xcU88RuhAC3YQtTjb8iZyXYcpIjV2kJChLjnuUr+2whQ6MJWWSZYp
u23eTSKud1fnFTTXcc0Miw4B0ePnYn5R/Kc8WLfQAF/kfrKVBhleMVlp7kddPXup7mDcGkQdi4QS
ilMsE4m3kbrP2u+OCrE4E4TFI5EG+BowRGoIorZHI6AyjNOF8lIZrOrCsXca4FnfP/I7wfoPei8+
zn7mAqhFOWkEtR8dFhhXvBLhwGL0cpnWQ1kXDH4JuUcoVZ0ZKQacJ7AHzrVBYa1pJU0Ny7oeFbFg
gQ76oVf+dEpvrmp853Zd6fs8Rfe+6k8l8eFWM3g3xjM+q8Bdn6T+mMwGDhhOMR7e2eWzMFss/Fqm
Yn9pKNUJy5F7vbGjO7WpQm9VfvmAWOYZD563aa2TqFpoTxLrLrrz7QoU0IanR8vZmlmIn9CyMlBe
xQntFIELdPn+rBvCNUnuvi8Ri1fhTHwHPEh7ashdpAlzMd4OAh33/bWt6Kq6oKlLPhsu/FJUohpx
JujSKlGUuAc3o8YF53nRRnGo7spmFNYDU/qyjHpA2lTkmu8fiwi9h3/evvFkkzQVmVJP8T/M0Qht
1pX6y88/8KxyNb7L6oIPDfzxxTL2Pf2YJDygizb/n+NKddS/XrOEuI1R9fGocjX/rLWVntux9GoH
+cpxj+NP0RO3+xTozHNzqjyyC7hOpjy20n/5RRDLLqnCei959cxVx/ma9d5YDZ3eQXgfZU55tnku
ZVm9Wt1IWiQPwR4mSMuOLndD1jIn2x+m4xsIsGbKKpAazXRnI4hQqkZT/gJeLa55gvGo4U0ZXWE/
QrbkupRhm4qG+MQC5jIRlQP+VcujANSJ3SLDWkWk2vdWvRsp/+HfPeRbrXFh7/Mk6yIatYOcgcJB
UP8/Hj+qLKVB9aTWYbgxgkrfgBjGYWB3tNtkw4j0FsrgWn//S92+v4FRkFqqNEHorhA4H1q06HLW
ZNrYIkmko7Fsr8Ba6Zo1tk1KLbkg4+GafObkxVNnazYbRGH+aEW1jh2fYeFiqA/Sj8drHuAcNEC7
ZnUN9y6ANVgBZ5Mr4/f6jru0vPQJsnTOKxYt0EGEXiEU2UOG/0+ReyfFKq7nR2pu9MXz8foCrAJz
5ELUP7yIJQ0X6NNrMSj4pji5vRSnr2GI0dX2mFxqV1WFTQVDUa/7rnDbCUyBHQEWxcm4JgcCYowo
LOpp4c0571hEnwLomwMQIL2QMMTt2omFE4eU/nbhvRu+v703VjKVYktxqLCmALNWY72KZL7oq6BD
czSNJhvIpdpM9xBWLB/OjBbKCe/cIgCdr/oXp9vFLB3Yc6f3Ta8J0Hp/vIiIGPLRX+9SdxYfLm74
J4aeDsOo+B5Ua5v/pQNFF2vxQJFMABK+XZuAFhqdWBREI+73GKD6/hWvnBRvxHT0ks+gOEXEIio3
TPNWePAW3jEVibPAGzfXZ/wfdiBKCopu4BDVGILuVhNiv3vrvHlwCICwWP2n2120ypJgvKReqqeb
PZiXfvnHcgr/vgntFVY8oEnQN71ORv3OvWgvNPvzJ74a9lXHujfGorGRPrXThr0v3Kqv3symjcFs
kQKl+V+M6V6fzANoSyiI8oDFB1XT3wQhkOPhERKORW9S7wXWvkloXWYbsl4bumNgwwPvziDBvu8W
NakyqteXO6/BxmXaTzqsRH5JNYgxe0fXXJQ5lqyZVpq0KbPoWZy2A+YHl+1WcSXVZPI6MKN/HD+2
3Eh0FP4U7PTcur684pDM/hJOMlOmb0OnUwUQdgojT31ww6X7mkqNna4xe0nHrn2ynGrTirPlhdhA
1VSADVrwquHzFKLhfshjHC6Y5oQy0NLxcQ+pXNyyhjF2tKl/zfanpd5EpWEeGQ3KOn+1NHTXCDUw
AG7Ng/e0WSGSPJP+4dpMkpXNRTemcGXZbj1Jq90bnANAph7MltTYz/CjEMqXKbXPlHUsP06izUyv
e2BSCN1zoHAUgMmC1fkQK/hX0s6DW7t3gt0n9uJqMWEFLc3SLJdwT6KX68REoOktqm38ZuzpdljF
beRZz4jVUYBPqmBuZEiJcKzFREmp5iWQe0bFB1Iyhy6V3gtdqBrwYmXUSPePvj4OivU6v5yqlCFQ
N6bJv5Lfiu6a423rGjyPL/+APxBe5wpB1dx85XYF8xEUa/zRrZVzcV0/9N1w7mCIxJuHt/XINfuZ
Tq8mjzyeTX5/tPoUcuA9VOgn/1cvhYYWAXO/BkOcBLnWfOOlinnKAFH6+x1RdsxMWOnKNEz/aS2Q
bUwbFtov8AIxYBGd0UlCyHhujkXvPYF9DX4JofOZHamjPn9GigUsWyQavzp3EFXMPE+Xw4bI9Ve/
eHH2W8awunuzAgL9HIcFkbJsOoVHqkTP6kxEaXJcduXfMuLZTT3qY8sgos4I3SwcnSuEuBXNG4Ql
cyfqKUK+5zhDkbBXTf/gq4Nzb/lXXuKCRQqTJ8uPuuBsLpYw6AhQ41n/o7QIBeJi8HUTD+v6WJ4+
ysgIJHTPS9FScyOFCvH20WCdhPnhT1ZEX/xrC3zvdVbRTgL3dySxSImKAWVLcY/2/S0sAAFlVn9p
iksGCZ2Fp8Ih/zIXYosCYWqSVkcugOR1nG05tBqEafIh4lf9Ypy8han5+XOG6zbtEv3Ns4QJOXu0
SGDM72Tk/luS4Hb8nIyTWAdp2iXSMgw4F+vzpM3PADeFiCdbH+hn+6u0WX7Jny8S+HaP0eg1haZ3
4IIun89aKKQUaV/+byO+P4Kw161frK+S+80HN+xTSwdpQB+M+XQ45zOP3kOYKe/vL1v2PRZ9b8+J
cguh4iT+YcNEGvDXKrPNHGSHB4d2fzRj3eLCjDXd/ljIanrllVUJ2bjwjhw16SL+RSYdZ+HOi+Vz
2vedtGSQXWzjG0j8g8X9L+dF5LZ+hmmUGBLFG6NndqzNr9MIRF1ukV+d1zdyd6L+a7pR735Mfvjh
ijGbvXCTCF6BYsg2Xi76KjS7Uf/ZUq6UhJ4QGHOIZ3Uyf2Gwb02bK4+3UY2tZTKMrLMDs7b2ERDr
YnX3xT19PaY19eW/+UsAEdPG8NrLtQ0M7mCvsqlwo+6G1D7iRh8nHE4IYjm/aH81giG4jmVVM0Km
5j9dsEeRXXWahYWYL1wOCocwW8EkwgDDIMvWHbGE+qhrcA5p/Km2XGHMs01jgO+vKLkbkpsBOLBR
GJp1XiOCJ+YO/t5xTp5SFSEJJ8Emd7/0+gxGJ8vMDU7HPXwuI+LyZit+zxOjPlC/3fCdHse5KbVm
CtIaGAUmyZ/CFcQHxvI8RSb7aKwtDtZJamjiFTTXbSrQmNTx/B+wGcxynmI2efa0h3mxFwgECZRX
yrinYurs2+fhpwqu/r01lFTD90M0fz7kj/BlP6ecR+uXsOCecEQT5MIgtT+QQECNogcBZnF/hrsF
+VfztXZKGnxGWZAVBl4jZlgDUIGuYDf9FVF457MFT0bzaB7atMOQISpJi9PWNRmg8EVAbxEpLAaK
5lI7kYroKJI/4dY6z4o36JpPijCkipCkTAruHXiGMaYLXkX18GtkQYbzLjIeceJjeF+2oubIw0kH
TMk873XV05NRMov9fbqJDfxIgwOKh85UDmZtQ9M93LJs1HNK6SmEfTP2L08taA2517DRZ0C7bqgm
SK6VaSpVhq9yh/SxfWtP7T8W/dej7Nc0BoVMK41ltrKEWbK/J5VgaPWxTbJFncOUCWNdcvvcMotV
llujVCuyJGjYURQHvvWwIBVWMEs9VJ74ytG1hSAwokw8EBuLVUTCJLViHHkHN0yGthVNJTWT+1NY
PKV1xrmlaQMPq/cEosQ7YczTL1ozUDfZ4DzEbi4uI3b7SGuV+MSRYJTAiGXKE1uyJc6m+fEvdbLr
3m5dQCMN+JWCe0fvixG0+ThrwQhywNk0q6jWu9hDfCYZcuoow8os4jPZ60SBYtI365+qW7fVMM57
PXg8CJFsYUPLWgb/FwHh9SC7hppVSfOyckAGwvtII/XZ5uELSXgZwDvYze7mU7PuNUKJOdPZ4dZh
hi3INjEVIaD/VuLEUiFoIBc9cc7s/PhV02nko9RxPE0mErdbmdUBovKdUf/e/w4p8BlA+VJBjlyK
Gx/C4Pg/i49eh1Z8Zl3pxH8L6RHQZKAfbKNxltxwyw1RGZTnmBGJsgHLl7zMfnujQrXWersdRYPC
CYIl9f5FNfw58Hxq0l7HwVXARPSLFK5sSzLVuG/gVIuIgKoJsdHb07X6xjwhfzE4IBGmCRX/0W1x
H5CXyvwI3dyqCj5TWFDf9MvkeleXeZfaI3v/qTor76vTVXXyei6uDY+ssh2oOhUtdM6krxv0Dl4V
I4estNlQa1HqueljtABkTf9paSgs9ofl2kY4dLY6QYu50Xaf18+d3JUYPXKEXhrYMiq1m4UQsIJP
e/TimJGbdJp2EjkDb8MeUHFGVHwAVeg9jE2lPxak3Z6Ha+L7FPji7A0LX9Nnelxq5w/E6eJnS967
4ofcO6EZW74oNhiXkrvXdl6NZ7P6OFJagCVSLGWa0Y6idHU2MxKCd+an6dfBRDTaj3BWZ+c9uzmH
aikvMoVyIvzqX0jp2TR2PW0EJKd5olRnVr13jGPVVk+kNDUB0+6Pg1eDom0u5a5LX/iy/Hf4hP71
N8Ek7MyVDzxUIdx9t67LnkvS2q2DAwBJbDcqJUFIvGLOrHhq56RbvJhO/pEMY7dEer13a2KVVEAb
vVXN1ky/x74u460Txs/LiVlqaBMgLydlbncKy1owJLolyYTiEM9O5Cb9TwBBTa/pUenXI3fJ+cSV
LjnXlg1Gg1KUNzy9DcyDZi934G2jmYhbT1X8UzTYcsbc6MoRohN8Nt0Sh2T3OoMoEfhh6SG2LvDE
ri+2yGyMSWVyizC+60nN9V5uRgT7r0VQFglzMjy4773vvaG/o0BAMoz4b/+vijY46GHiwFT0dJza
Zf3c8bxm5Hej1exQyoRC+l+6r9SCPCQWUH8kk0L80mTLyrEnW0/bruKIkwEtNFCLKhBTKb4m6Glv
OHkPXK/LNR2pB5HzsT0+qsVyAYQQbGM/h0iCD5ITbqqBQsWTkEIYB29xytn28UylTTWXgwfOAy6x
4e9oV813dkWm+OO0l2cfjz2haaVt3KhZQH+t7nztxZ6VjLJjmNYds2m5rBXQmAWtvZ0hjFHhH6kv
iWCmUevMgkKtKsUTYLLcChWCL/qzoC1aeBuJr201mCIIM3ux27gFuAP7Go3PD3WR8DAuaTqI8XIg
xU5VY5tbTVe4Wlhhlm2BDWdWq55YF2mNs1wWe3/5qBDZjrRxPqVhdtO3pSB6pnIHrRfOiPjU0z8r
kDQFK7nG6Rz9xkx6TeiB5pLEW6UcgmfqI+2Ksfe4cjFDjCFUQi50q4l97t0r/TS5qQZEUMnkTLlt
HYt7Ht8YFkEjcQ0MJsmhGL2lnscqU3LqYQG/1JVb5cyi3j6kLWyFBdJ06GwrQ7sWY3fAJz7XT8RI
r2YafkBJZajEu+bMJBbIk81oh438iy/P7m935VLETqsKHg8CAtsDBNz7RkZRhzdQICB06CtFXhO2
UlBSc82twK5fCWf6iihTCO1xcZdEcaQkv0Mz9s6TkprbDoh60rxqm6bwoyNTNw/d7gb1ShPLSZSv
PZuVy7VbeOJfKCsOPr54oNWcc5wF4FOH5eNs5yjzWD8wdS63sINAaNuTnEYAhLOHALAIS18kQSqj
MctYfM0g+r+MGVtLZrJJfD3dDuor+MPbsjjiWCRqCx/hIsz0maiWOi6HAQGDXrbGaV2Ew1/pLF+8
o/Q572w1RLaXabydx2QkXUSXUcZX09pxGaQn3sX7hk7WMGYROkOaRXL1dpI0R+K28ykWPbXFIjxU
YoxeA34c+wiROidXnhRxcN18pn0Bk5pZaZwBzmcp/MxWTEPJzy2bLvM+9QuPHp3iDHeziCw3sg27
tOA10jnyZ3nH8OVbvSME3bGWp/N0r3QRHAdyMgh1QoMWclNkD56ng61LWGZrwpNywtB2AiOm5E93
EHd2nb6jGT3f4LL4VLm5/Au7/8gZGLsJfpUf4FedY33ctGUItN2QmB7QqP7YJ5BVS2JQHg1E9RmN
8Jfrzx+dRgMkornVgKFf+T39NKzqjItQncFQRPBBRw3wH6Iu8SqmokKx6ybvwy7c0H3MgsgDcelP
WlXFBBnXOq0d1eIPRUy6UQrMEMRHNkplaK0yrcbJO9JPVSdyPPE1Boi7HK7i1KGLBCS3scSDLWS7
oRHy2rxXtBXvxZ91xmxrDhYkMjUcITdB556Y6dCFYoSPSmNsZ9gj02MkSMRHAHVam51yhn76OBIj
GpZt0WMntw5fhvLNbuEqhahLhQjBcPU/3/6udhVL6V3RsL1LMXU2Lo1Lama6l8ft4p24NRfy0qxV
9T6cY2jEjuHwOkuWY7VGCjubKw9H+/YBcg0rAc7PoclEZUv7ut4zNJFlqD5mpatfNE3Mo1bIYQsK
WuNoyB8BYcNVq6KT1fyePuDOWI+TYhsqAxE2VQ1MvDY+WUvp7PANz1raWivE87HGBeET213fFkYu
wTOYhyIZT4S+kMlB6SRsNLsV6qSYPVFLjsRp6gdgaYtfYP9AJKrfIIMEddBsXBF2GZ0IJLYDVZFR
+q/tEJzwUMYNz2fdwq402WB4lRoxCdSYs1SHjIifqbDFHD+p9cRq0zuZkrg9o7k0GimdKnYjYnVC
XtZ8Yp3iB1CA0eQAZNQeokI/r5DXz+VlASmkEADRzID7Fy8peIpfk36Hvx8A5MRrAgfTKSP81C6h
XCId6D+q4HD58p3p3NTaGJI7lP5Jt/UDcmsBCJuARnnR4zVDcMe6KbhUuGPx8jyCvm0NONmcC+ak
LUo2oFZvoNOYydOGmJt+yN8zkL9PF9owaoJWP73rcGVZGjLPWQDB6mghyltHuJhRahA9JHEnJwy3
ztsFjhvNOtWp/4udPDNYZu1KIUKTFHGQcPdjX7uU2IeBEhEROOKC/LbGm40UPa3joxfmsbYXSnBj
6hNr9EfOElDazauUMxbUDX54C31lTY2Wkxsv/X/ugYuJyCcPLw25ToCFsJhWuLHAtZDMAAPY7HXH
ZuQre4R6Oj2kUEqrONGsKVPuH7P5dMQVb+IW8f5aRrUaKvHnh/pl8IqWjMT3LlrDOzC+SwR/rtKa
VYGrMcXTIP2nVAyfj1nzjjhiXxPBKBJgbWTdE9yM5l1e8mqMveQnRS5WHt+aQDYTplN0n0dE7Eln
iBGcFiKp1Yn1QhjDqd6NU3KaWL31FDfOpdRP2lt1Z1EApq9t91MRajz6u3d4AQcvairsv/9wi/Ri
4Ycn3XabttyyjqqQ8lHjrSnSzoFXz0vAB7u8PxxaM5XCl8Vm3yQZzPIhsZ/lxorXTatw5RHFG1w7
JLL5aDvrXI3L1mYNw3/MXpQlt+KpNr0KXkc0sL+qqq6KcF8/mC1nNUvN/g2BXOTybiECBXjDYiTC
Ex476BxvzWDjilfBh4WADvO5FZ63UJNS7YdcSs5ZBzxzOfa7eo+Ja0mO6c5TPnVohzKnxspSGyZF
esK4V9M3Mpe8XCWH29GFwfkp72mmXDUen1q+xCpowiwQ+pzQGfq/7YNEYooekJRFYj1a/L3HdxpV
0Zw/B52ZfPRwT31rQZc453SMuEFRJGkUd5ApSDnMMtgC1ma/XvLMQJGQWDWUXq9XxmFv6k2/vCzy
hogdftZe9LOPY59lcsYw+GFIPz5kpj/AohfKjdlLbt+NDK7D0XKAFZdEy0sWQMX2pbEr90UPBwbZ
XO4KRJvifWDaHKmEpQ0JBy0+S31wZZlmpZnw0TmvgRfEfZJmy17d9ontk1bRUO/aznTmyN2s6dn0
CvONwIGvj0Tk5BHWvq3snoQUKtGZheqSdg6C8hTgUKhmE05assjNNPTgYpj+aM1zgGfQQyEMpBOf
03xuyirHCORPT+QKc0AnhFhbLLT7bvf94jGEizoMFfhBHW38gOXQRmCV1tkzM8ZKL5ZW7hVxgs9Q
cnVQYM+tfIMDbPaEcVaA6WzjM87jWv43tQeKKj3LpCOgIufhd0+q/au5VjBPEZuET3S9l5GkdCxk
XNGP9xa0keBPHSLIYk3LTU6KaZtevQZKTm20hg2z7zSgEWWHP2qemVUkMzNbSyaUmEn/4/q1wx21
rzQcI3lQ6ln6xsvahKWur1gnP7qbgy3uXdRy6ONFioClfiM8yopAGnRc41FsQV02nPJ6Z3zC/KMH
R/Voz8GIUpWYW2iYAFrOFMFmeIiBWJRS38Fa2S+us+LCrXIC4dwdOZGi68IQ4oUJBEO90b1H7WCi
3kaUXlvsfWk6hpV3O1Y/m5SDKSfUaXhL2W55OW7eZFfcOlJS4OiMejjAdKJJwMuwfarqIHKjX1Lf
UL2YsvHJ64GaqH+lyDTOabncoktLSiJ/ZGza5L2SBr1ysf4txLgx+lH/Ovq753IP5/m8FEpUbHa5
7z28x4ngBrYiyK2xEJx1mF8JiVxDvU5vIdtWsBD0H9mIaxMgcNnqb5fxYco38eJLtLNkA8M9nFWE
kuEnypeFomeziSoQ1/gMBKQcFAp5o5h7R1Td35O5JnuJjb5VQL4XB9NEUuay/7JVYtYkfOr/rJ0X
3O6ZWd2V0Tv8xd8aeOI39kfTJ5vS8eUzC0qkaaHAIO6dJrMF9zWmpYVO0krYBlo5IZHnlRKhiGZq
tsRWNXxr0okGXcXMbVl0zeLkM8bCzirVcXxYMfXN5QyYifTJTvcni7n4/FY8ZZzRY136lMzHRKod
DOC6YNZZIaz0Qt1h9DgbgtTefW5x4PHrdtyIhYr56eZYc2kjIoCjY+dlDWXr2dliglqXPj2tw8AB
5WUm2pLrDdj5o6IpBld/ERZ9deTWMcUr3jfkzSmyphCYg/elDJ69TDc8nk8Yuze1Bc7FL8hYsBKV
GxYuennV5/lMhCjATznL8tJx+Iq1ykipVr2WEZ8UAcXp5W3aQXRFqhaSKwXlCibs2uNaVUvf9Ndf
1Z/StKSpR82gf9Ez9NRR+aWzrR0SaZEHFmpgrClphwKWUNx9kkdrz0LaQlXlQofqygEY+sHf7nvI
4Iid/TreGEh5fWeS7tN4FHdchyp2K4K6+X2QR6K7TVFULbZONAasyoxmeH+dTOgVk2BEzmTQuuW7
3sx32RJ9I9xBHFeNHxHiVoaZNSi377q/8F/jIMQHRCDGm7Sz/UJMuN+Ej0o8kGlwrIjbvl5+kFYu
U8Q41Qe3EvXsagiJdluiA7weoqrQ09JMRAQlC8OxgI07z09jIZeONLjFi2KSDYbZQeVOF1U6kfsA
eQgA3/l1jL82U7gIHTjFuGr3DmBjvNaPF6mzJKSzfVUImkwKHJi1zMKFv4JwSlvhtPtnuT5v7YcR
6O4UcY1vpnyTpiqTOmU3Y5xycSanJamPOV1AMBx8FDXEJh1KhvSUOl0LlKl1RrOkBjITtSRIEgnJ
O15lJXkizj1h18tb9kk8GEt//ZsnZW2s5/Fl7n4MRpnKZE31U6KDJy3tEf+JNM5ZEmIXTFlhUovB
es/MmwJYSuOVPhFxfjKVI7vhmJCKPVnlzFGr65HVR0U6Z05v4iO35Sr0sWG3rje8ci4J1C+p64sH
PiGi+r9/ddce1UFBH9V/1Qq/ACGChmtG6VNPG7LGrJDTv/PPetQ0G9VgJUpIf5qOGKkqrQFqK48Q
48IidCn3NA6JXgQLlbLJVf7bbl/VeuRo9Cm3Raqu8TxgL35TTiujkSE83pcMR7H8xVCQY513pxAI
8oT6P6MWhrPN4rd/pi7IHR1eqcPyJa6ZrQ2AjI6eZyPZkaQeoEeeFOpFR9OoJzY8d9AY/jfRvbrx
6RdQZ8LBI93l+QZMjYZcGndBsf7z8an76ZMEawusfxYGsw4Dc5EnAPUhnJEZONX2q0f8FHFide9I
VNKoLVlaAs/Jj9ODs1Y1xIVChqoEcYMI0NqrK/00roB2nEHvJYoVIvZ2VhYPc+eWCOueWXZhD7wW
APPLE5oX/gTciIE0TXSXsBux95kXLRPTPLjaSlc3EJ6ojuzyJGQULLsDnz+0OCum+trs/ktMsOL0
FFbUVUsaYcRJj1vSwPYbxuqzUOh3vhnVD0DTH3u0hwTGcBhHyUnHoRnqUnLqOrhHtPasvfSmRHvt
WpPth9RyXQBDxfPUKV8+tnaBbxiHKZZ4UN15eI664ykw6ruJ6cgIrRfBRe9F+YLJsW51kuxM5XbV
CAGJlZwOqSLCKMk0PqoE8R9CxE4OGPSsT7gYFmdb713a1SKvgLxE66t/LwiaACCXw3Dew9QM7fuu
vZnEW68Qxr9vKkGU00gK94PAEbMdvHxK2S7gdn9biOQD5b0sP+YR+s3vFUU+U5ACvDuhWZxVV40s
pqaSSazKU/+gm6Sck7MFGP0xVXhGZq1CNJotIaHl01vEl2hLcgUJo+zHI9dXW9ZsHTxGdWSbLvkC
+0h/RUm+4+kVy4Txy4DiWQxl2mXLmMlpXyGWfwYcEjywfNvO7Wqi6P4I/jevWPFCBR3FKcGcC/5+
4+OIagihYhBql7FPlGlP6aW6y/IDNlhmwGU7SRUBu+11NCuaEmVk4D17uJ+gii53s7mJpZ3y84sD
8fJWEQpo+p2uaVvMrYzRh58DdZnIOrem2wnkDjoloRsmb31+ny28gX7OhGvylqi1IaUR2SUToHC1
s+WX9v2Y+gwZ2lUF6UDjZ/r+aX/9UiBwXqXt88/PmsM2QK59n5aZle0OsHFJIWeT44Fk4JWCy76b
rHGELF+mUFBRHWs6zCW4p6iY77EOaxgVSAtTdmKbHRH33Tke55G8b2xxPI5SFjcL87wRhRwMyORw
YUk+g2KZuWHT7miTJULyIOskS7Qxs8D8ZV6ZRdKEyxnMsAkK48TdHSvKT7XY3SfFBPkVz3O9K7ie
6/jWMQP/6HjmDfgKSJdp5Se96DAPk9T3af6zwvmlK85zgYcLyzxrWVbZa4a8IszwiW+GY3T6MPld
RT23U3jY+6AsAYkTtGUqQ5gTI86sVbzLBLXiO3kLeJ7AZLJ2948r99BvUdazzl5CB61blxo7w3v4
uzxQivGxCvQkUU5h6p/ff2FsqvScRsmZef/eHqefC+k3n0d2E50BSWK5JwpFGNsP5nwfqipycOlw
RMdPIu9PhFwbUXYifzxem6CumdEF1Cu/l2gZDtKhWEg4vtV6fxdMnR/Bksex50JuL/u9O5n/95pU
DEuxyOKjZR2NfhjhjTbB81qq3AOti6oyc9sjlY1IG/LDt4QGfKB2D4MTypaIOq+U+0m7LZRNAD3C
6FhUl8q4dJTMDei5JdCPBMgRsjFgxLd9I0M78oyzYs04cyxTnEk0WqxhSBg/oue3pYtgn8zKiBcp
4CXhrCcGImfo9JT3CFEAn1QyBaG/BLGPMAcG9MX86U6ezteUGIam3bL0p95OQsjR4saZ5LXHiewV
yFw4cGCWum3d67k+0zWb0WMeMspRkhj29kr/rEG4M80YC/Kns0b6qj4O7L22OT2Vvjy5klAJzXS2
pR6OoQR5goIhBZTng39ii6zuyjYOES8aExn9rH6AV+XC1lFuihO9QqUE31J61SnVtBF3JHXXEnjc
xc/+nesbhkRUbgoa28BafWppFTQKyC34DDVcxFKayRdQELagyeydzYvGltSZsOx7KoIwBQjILK/A
gH2pPOc9/90NZBYqAgtRgQvl6pOTqT3JduFSh6v6F+YzgtGvyTlUEYTbigOQ86B61ZRBQNWhrZle
RQU1vEtSKeLqzp5743sYGWyYPQQiYXx77jqDD2zv7plIRmt8ltkW+dtrNydQRgYZS0eIRPPoTzXo
Px+lpWNQN0uWHjemVQEKqJ5tMGzumplU2MyhbKDHLnpcMrU9Edbb58Dk8vgE3EAHBsypSH4uGHN2
89xucMuzovkNiiqiDr7As3CZr7yNd0sRCxqrHLZcz86af07KEmnaWKCLdgxZHzEYqjIcb8SRGuED
qYT6tsKf+AyQoADD9EA6BvMQX6zS9TYPNQh+o4Co5qrq7jNM88NJpsvcUsJpTDXPVwVkmIjL0lSa
fKxeMrxRnInfA0n5gj5xzT8Ut3cZ/Afj40Q/XcXXtGjw/5nmfJfAKH0FAbgisbsJDgypg9tjvVju
sSScuR6EMNWypi1DYOC68Nx+ZDjSHoB8FGexzhWgUYmfuSjXVkrtAI2wTiaSqDGFYKtQd5RwHrDV
KTQ5oW/1Ksw041nn9y8Z4RWurTyjw1K1wgb5UAGiYjIGARw1GA4hhwbVQl8bH165OZYwXj44G97G
sxnzD7bNm9LIp+5rcRbE8Cv19PUbmqQj8aNm5eJAN+HIY5jWdjMSVWS+xslU7ypN2fnuMiXyBeVx
GoaI+XWwA7wZs483qrhEUXCHdNuTmHe/bHOSSYu8b/sOvhtJta7GEjbUYcGo0O0smUlFyCzCM455
+TGC1iytmS4Ec5pOOMlFYMDJQWvkIoXbPhPb1KD7RJxd1nDrz9yd0CXfRhh7Ze2iaU+4j2gHYdhp
rI8tA2ec4tbiqb4fLcGqyLHZp9kIefV3G7xOPEwcF2Cuzvytzgzi5OWlTjCdWGrwDkMFCWSqWzwD
7F9f/2e/HK4hmIhP95uIoTVXGaWHJgnTc3/ya01K5H4Sy9GjHv2Z+AOfozf9oXRAo8GQZqGaPS/l
obvvJgeThnRbWDl+SyXRhpalT/2Arwv4jDNL8vIpj/6QPoUgfDrlzrABI+ycHoa5XnSOZxU8sCtY
mxThrSDpbYa/ekgDrhXF5uAwJ87dkeFMD5aXlh1nBebp398kiUAhcptsWUX1K/zuRqETID9YSq9W
yW5TNwCZ9F0hKaxf6eOU80gNE/kNsq3tN6rVg4k0GoJuGyFpklErmj+CIA/DrM26mNemNqCSuB1q
On2rwn/b1pji3GUGSbwnENoZcEZhgh00sJkqWqwKI0RJ5apWxtgH2VcBr9R4b0ipCzuLqcaJKV2t
ANqpGq9v/o8t/160gg6CQj0saBFibi7K6l6R52m4OI78TF14nx8J5FH9yz/oiKBt3Uyd5haT3jMu
R9mrQH1tPkIyviX/Fs8pRbZh/449BHtHAtplBeD4UxZaiksoHmeHAHUeejOVfCC7XWzuZzTwAc7G
jIob4+x0ti04t9EGUt1tjSsSryL/ssimyAZ9/M26DxQPAVcm8kPUkxQ4YoAW35Yq3R9e4LdIyA5w
3qYnonqA+FUUN+QV1juP9O6raoK8vBPdpEA0ZJF8vPSi/HSPYfuvgOX/fTVvTB025x48qv7fHAmQ
woTNb+PrCraSUkYGmmPKLV+k3KgBh3rst5CjzlF3Nx7NMVLUgaSmCGl9TT5Pzr91pvCCPVMbSGd7
bEqSUjG6/SJAJrjLmVm+SpfFVeW8zQ5xRKKvHK8Rag18g0gW0kIj0Ge+JtgRtTA+l4YNZD7wbGz4
0bWADWrZjFZNSRZS6ZmoCp8STOIphTAwBfUxh7Dn+tQH5zYebtpWBtqZXjZN6vEjNCM1yjX7YAHe
wkJg9vlzLeO0Xv8lP8ZXEvsuU9SQPHZbv1pzJgaOHQe/veeOg3+eFmE8zf7nnWo9TavAtOV3xZ83
vNMaECxDIykt/3ooV+HXN3+17UhGTCVz1zUxfVQy2PIuBGxDbywNG7+ZTaUAt9rwwERU3/FRO9ME
qyZ1v38E+nCz946p6x2ZX8uCQm2eILOkmE2IxF5merDboPla2/ysmHU4Mog1l3ZhkCrol+1P8OiG
sTUCzZJZxEnW90nEFaetkCUHTqUw/aDpLuY5Lc/IBA0RWN1a7kZlf5tW4dw/Rt96kZe2suC5VL23
DizsQE1fFM9H2Z5Me8Xt1BHMt4VVVNnYGNn/K4sY4C77JpCJ30UWG979MMRwn5O6KnMPZafBr+Hf
g3brON1NvvIRqYwwPI4nsJPqBLeZMRXZJK+K8ypogra3jVj/CyXIa5A/+wZ1hADLVXS6M+9+2jac
C3bVoXyM1j754aQ4crk=

`protect end_protected
