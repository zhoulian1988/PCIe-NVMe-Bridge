`protect begin_protected
`protect version=1
`protect encrypt_agent="FMSH Encrypt Tool"
`protect encrypt_agent_info="FMSH Encrypt Version 1.0"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2017_05", key_method="rsa"
`protect key_block
dnGab+xWIctP9apqshQ9h/gBLY2s87YgD4ITJ9z3iozNmZU0gJlVSrOY+Ddp2Q/ZYpkOYvQplTN5
yvLy9a3lpEDbsk5XKQljUa7UzBgoxRjIrb2hDktMBqdMqFn6M9dLRMlxWyPGkDj9+TsiJm1J816a
54uCe0MfWNDd3VZzgnVxHGKLGpo7HfyiR/sYmm9gwbFHvbtr0G9vk2sHavZDMRhHxlKcM4fbXKTB
59sFGRBTJWY27Gp5j7VGP3rIlgdvfJczf412LM1ersffMe9kDG/koSXzdMse4IQW2SVSPk4G8b+q
pi4e3fAytjM5Dsyq8ithsg5fqC3mMlfjovYtGg==

`protect data_method="aes256-cbc"
`protect encoding=(enctype="base64", line_length=76, bytes=132672)
`protect data_block
hqObO+IAsdRGWY10Aql+I5Lwtlp2osIXkEyTwYgbN71wDq5Sz4SBaePSJsHsfUF40Egu0HOCMMy4
Lal35aFXNZYHFiLd+gkCasS2QFsBw5e+04udOKzbsmKN6yDoWU6+PX83PYUphUESAryj+5RCDEKx
KQZO4VxL/75mS56PSpZZA+jKFfIXkEzU8Scal+P7o2seAsqYJVdqg/KG5lhdWqhkAkOCJlo2aQcx
F5PD1rs21roFqbXC8c1CEwzI5BgEtLAvBsvIZn/HcvRHVPs7kFJ66paK9hXGxDZRjhLJbeXFvQMd
g3waI9HV5/K7mT01HWWTan9u6dLzSFjhwdZhMYBeu6E16Q7lpkxHv5H4Z8UwPdToDx2oI4iPnZRf
4xID3LEvcXJlYz1MfSda3g+z+g3oraHPjuLg8aVZhIjgJFhk9OE3IoDkwSPIXuL1RHJNWbI8mh0H
TgBPqxx7MASQgHavV8GLHwkREEWwpo+iNk4jcYyANjHAip2Qh3KlBa9tDfhDK3ItYTGsE/EmjwNo
1ujaridxaF2ZL/ypl9lTeiBZqn+KE8DInDTaa3iq0NtQycUTJifnEtE8AjJ5TolSysB4mmb5uCpf
8Mra1ZMOMCC8td1VbRolYHePMDLk+fQdiihKXREC83U9ARKTCvKkzYGC+3S+PCHXOLJdDBY/NTQi
nSqAycvSBa3vYUy+XlVBUlQQZ62LNkM2P3mOywYE3ZpvsdSqPcmHXUJaOZgMo3ruwuz6zoJsqe6g
bsA0YmoXUgSO3aOBIrI/ZRc4Gx71SYYAZdDx44p570c21dJ0Nxu2R2igd1om7L5DXmsUkfwYT+I4
BjAft8+kOk0ToELZ+N1TN8mQ8h9GZIp9LXwWl3I/mQe4sZxn7vs0eGY9GTsOJYZ+n5MP9woBLh78
UHsQiMXXgnRkj8VC4pHHVqwqkuB4ow3xDFzGeUXhpbNVNoVDRDqx5mRaC703QdRTqAHBU+sZO1Ki
IHRI5ZS32RTwF+nl/Zr0eU7ifvBGIs+aVtOOVMWzdGjhVaaytk8TDTT59pGMwa9Vv4H5BWv7yMwm
+piFpskRZDMEX1Az03Dj0xbcBvzfjKwxyOS2iaNRA/XHEMLni0bOJ4RM1UYFZT5EJ7Vd8YMDk6f2
Q1kmniLreBWHGnjci6sHkPKPI/t6Gl6+6abjMuDH/LaPz3pCs5jzDrFE1IrEC2eGbwHitl30XVI5
/RnSJhhY9sXribyDyHsHQ4AjIb4XbXa4cIEkBwvjpprCx8XQRoaNZ38w2lXW2QXS4To0XmthzRUP
K4N1df5okvCZ5kMg18ebnENUz4qUEshy29VfN45Lydl37zMyPnnVwFrF50RWw2EIvsHI+op6HbLv
7O5qJ1lGBxRNq1nLFIYQE6HP0YebvUw1X3j5vxzXqdyJyCXDMhnbAACA277seWIRbehRlFKKrnLx
6oQ7qu2zbA52WX6UdIKvxwRQkIE66Bii4njrkUtNS85grWwplrfpWkssldQ69NSo0abArFmGv+Fj
ZMzyeV4JKxYCPB1Ew/j7kogSGEAZiPw4FZJKQTICzWHrPC8eUsW2Mw7KzGf/Iq/webiO/OeQaubU
ruynMOtVAQcMLKH0b9gfwEIQEPvMGDOjA9NDm1njFD9qKVw3EOdNGCMKLOBfmaQkhhJSQextYKLJ
vcOVGveu13QaZBTbdPZgjfzLdA/ENoFGYuOvfCxQLCysNIt3IQpfhFndMawS8eqSq4lts+cD9Wbl
kGnQKwG/leqDOAqHJhBgyQBs5x/4svZZq7C06kLJFSvueKWHy/gnIBUZJ7dcx3dTwj1Q224TEjA7
VkWKg6MnxNd6KUAh2eejI4MNZbdVfhm//LFcu1tCyCpklszIc6W/NUIowOOBBcZt0ISM/bDO4gHB
/RORxGXrDDo6qrYlhm4ujk0L0immI/cBdgzUkXrorTMuP7MLAJMrUwNssKdRSpWpBhP9h+juDIVx
Uym3b400IzuzEr63RxKG3zMynUryXES4ML1yLgOTYtrl8pY3ihndhBR8LJwhiK3uw+A5SbayNb4q
8TuPnmjmqpWaZJZMKtAv9bvHrVfooItgDCxiJFvepYtdKlhs/2vWxsphcoev+SDYcuYCCO+xwdYm
oM8CN7Oc1MeAdvQkcE9uIW25ehtdxzK31WVLvXq/B4AXeKlZC9aOeRWRa0sVXc85drprrXfr9VzF
mh0vu04tjtAXdn5/EILXGlfenQfEUWRn7KFNDVdzhtihKzDdvsgdWXe7+tQc2wZV+QYE3C4cWrjG
+mTdo3I4fAC8pFqGfI5BbO9Fp0lwMTVcxfqna3p0doRET87Lj8e+gYxnBF9Hwp5mXHRpCX87rI03
Fm86IGJKctMNsoJSlBsrxHrGiB5CuFUZD+aTIETWBy/MfC4DJH12gTQxysJzg7kHJREVhWYyvDxr
W1neqoVEXrGi472wIWgACTGFxCkvkarGb9ujqRiuoRyHI9tN8CGYDGJPQlpWZuFUit9bRXwcqDJL
oI5wWss/PORfD3c41gF7kFn2JpqNFTaU9rcYR3Tv5lFaUiv56bhJKO72aeqRgKmYetwGJTwwr/Td
n7PirqhaahXJR/xv5Sbo1vzpEE+Cz8N6M2DVA5nYSl12SsmYQstaUEog3z36S2RdOVfPRoG7hmKd
r6rNUqv+wfQ1HurycnPvkqpPZ1mVpcmG8+R1/abPT3xU3MXcmonLVJ+Gf9FYi1BtT0x0mCh+buyW
CMQQ0C1L4Suc+PQgL6p/g7yOvyAKIA01nfyIXiTSMKKNCu26PF6kwd2PlFDgMre2k2c5s5ChXUfY
Hyv6AvBqDtQpe0A/ArAFSOydca4jm6HQ7j33yOMHYgrJNGmhOaM2U0P0QM0BL81+/XYXJdNkPCFh
ctpQZikWE7os3GH9q0FVAHyU88A9LZGSBR0JR6HwGSHAGmyB3Ma0bBLtmqqhYhn4zKeAqqHS//Vd
RPqhWG0cmUDxAKdAzxzh3mfUWRG6iwRMOU6bLVfbvmtYA5JsR2TK02mOBkxtP3vlxZ+Naeg+qQSC
3WiHKoE4OLkXmZ/Q2uYqMJztZlc7r/Os4yJiYWhVIBjiic1NUBEMHp3eFDly/7IXP+ppZ1WM+i4Z
dnLsOcjMpdkBtc+mzpSRWZlFMetFr3nOPXLX8Rd00QBlEMvIzp0ilaTBUQa5XRUhpYp4EZG90y7H
XDDtyn3nVg9ZVExWA0KMZ8e3NIuefZufW1V/x2oWl0X7o7snLiRcB+nHsSGy7+197v3Bq8M4v25L
yAsSHqb9+ldPK1qCCXHqtTrBlaM/QTahsUeoznxYnvXXA5E0nL4/GfdmmmjQjBvdTWd8zv4q8DVc
4q7WYK3S1Ho9/Bl33f6x0xF8i7ILqZrJz1Il/DyUjzzv8FW9q8XGQfD3lQ12DAo1gzVGf7R7pCuT
Bde2P3VXWUWFq2X1b8FP+o5hO3w83LT92W+N7w7ad+2KuaVJFvReXuuDY5Rt2g9aK05/6Xad8tMG
HvpESpxb919tcznlMNGru6+h7J5VmAojEehz3x9Bk6fSngO87Ilg7qjPlFe6DFP1cahwVVbwYlFr
CWv7Qc0/2HsY0ymg2A80F58VsSlVctxh1ytEKKEXs3AC3KUTxNSdAEpJbNbMc4wb9/Ki7XKAXM1W
RTOUdrnRmjyalxOrOBowK0zDTW+vbs0HnnM1b0QfSGiNuFs7KWnhNKQvMVSCsTrEYZWVpjDRuMqW
wMpevm3CoWm9ycebtetWuLFzfrR5o8yGEmCGNVQD7a6g8oqlLhRpFdLIiEDP6Ufj2Xu/Z0EJd32k
QUxBlwjNY3sAH2G8+GyYD2lRehn35irfhRpAAlCUSwk9gCpyrcm0bn5f3veyJDiPAtNBFPRRt2h9
KOjelqbkafHhoaaKKkq2dpTnD4Xoea6+QbxtNNuqhaiq0I8D9l0j9WQkHMLujfXtz5CaPFHlsmK2
IkTbMLYJO6uHg5eH3JyLx1wPTZj4DDP1VOWvtWpise0rLL/+1kWC+0HMVS0sxgaukNtemNpkD7f7
ko3UlqMlYCLKLwDubaGDDdiV0ntEpgmOCB7nySXEmyL+0eY8kmlLxzW3WR3k60YKdY5RGAn1I++d
bpny91Whct+oXbi2u9Ek/mdjDeNd3Id/4qkHauvWQocc4QSaltfPp+rGdZvBcjQ7z5GTS1dNo/Wu
7RPzaC1K/VyT5YIGjLziEdX52KU5xIFzt7d4qhP47ucFQy14KhK9gXHXLjKtCj/Hk9iVU/qhe1Z8
u0jdCXA8NABvVPsFfgDBhoWbDGWI8DsVZJwydF/qsU0FGHHwLZiSLlLkxLPhzlxIVviMIoaZnc+e
cJA0WUl+wRXjPsrRXo3DvLSs2O10FkpZkhyn79zgTItCoKeWMl20KXg6PCH2w1o/zSYxny4yNe93
jsLqK2bL9AznE6DwyCTuPuF9BNzZmqIxFXiDjEyHJKuDOO+T7ey0uihVBr+ng69FrAFP3McOAnZp
MyT5Y9rSqlUUpjwd4xzUbw2mX0Iy6lX1/5QT6+N6j/DPmMKsyZ+kVdTOUdWSBY5x6dXZkl+wHd42
jeDCHTVGo/LkorrqdBU18rG1VfW/LRXudQGN4j5bLRJ/RFUwrJRiJmuGXaKIZpa6DlptUXkpsnM0
FYbTNfPKebqqF8VRPMxGsXmEl7sCRyawm//fdXhtBTCIJtfvh6zXh0DIXCXqM97x+VqAIHeKhCav
cFu/WGO1VYi/2EO/aQaJZUGkiP1ne0no83pybQ7tSU++jAJNYk6HTcqnBllZxhajjGrp7asBWWBz
bdUVx3YajUS+QzHeeyCh1yjarnGtH8HcYTu3SncgdHw8F/F7Z0UC00aMVh8suUfEg7Qs1g9pHdkb
0ONvZEcJIsdq0hQPiZYPIWj0yZxoW8mUb4oEq0ndRPT7naMMe0NygBXuykV0GCakxqjome1wARYt
unVyU1Y4lCKKdCzH8KfRgO9lvDkhzSilmiU2ijGlUJHksZ6OrPajpDoPMPyasWKjxBBlhnVbMVTH
AlM8mFEG5E93pQ7YhemidRQkGvgw3qjC3rGCrqSP1CJN7D0adKClwD5+WqcCWoQPsn6W0InJJaqX
Gj5lwWUkgajI1XSBieuaZ8bFZ+MmYecUU/WVweDsEu1Q5W4K6hpgsGq40nwQxQtansVD6RU6zJ8l
ngTrx054xRCb2rYDY3vEbLevCQQCGtpjiLNFiRGzljkXiG5aMQ4U+RVmoE9TVqAk60yycRv7GrKh
3WPfVN0k9WkCEoaW1DpWCOIHSsKtqReBDXDwrG4VpFxp+zAzuvX73eSHcXClym9+1mZmEdtzFnyu
soZ3aT3uG1hONsyh4bjPKR4Kqdaws6wUEl2hOBB1q2/mm4hz2EUxqyEq7U83x40TTFP2y5dWLLVF
Yw4Fdcd0B34fLhIA/qt3AXBnOEuIeIBPgu+evQMicG2ozWhT4vY/MFO7i8ly82J1VX4SiyX2hqQk
PoXkvGhCTVlp0ox6WqLFvm8aSbKzkaLCnj0tWRktvCV/Lx6GWOI8xRReQA4CumW5QTQnd8wvri51
Q+nbu5M99Kqao/uWM5Osj+m2GtbjzC9+kMY+4I8m6QsNazt343U/WW/ZjiWjWQmluJ8NLVTH4+EG
3+rPPIOVMWbYLEeiswKnk8Z05oAiYEX4vBLWczGd3MnmJy1B1crkJ+THFJqy7SUo1Tvq7ywMudjQ
D77cbbJcY8lLM4fzjrEfqoZat/FLUQm9il3j3FOc0qVc1m7smolCkVB0aHyxM8HBNoHBZP5vjM+G
A5TU4whaVVA9dLJNAJ+6TizIn4g7OHlkSz0BnlAAHaDjoJvZvoMZG4L6hr0QuKSer3tc+MGatUGF
2vKY7OkBDnOaL3JZYA1ExF8tJj0S1Ss7d1c7CpZ87vflxQa2TWstP6NdKC/VCk6xUgHS0ZJ+4XfL
uroUr0FsaaX03AANdVqk28mLxpYxPUR2/Oc6vK5/Ia5aNjBkfUHSdjiEI+7K3GOPgbFZr9/2P/R5
DfU1NW5BXvAVUEljuGPd9cskIrE8fh+FwlN+8Rws2VSf7D3eSmFQrEb2ZgJ3YGxJDIFJ/oETTkVE
HyR18WDlxo7UVML5pzUNHBbf0H1Cy55IS4D8ATkq9kc5LVmluqg4O0YJmb1LFOTzkngN3yXN97g/
K0BE6a8zIBODyxxpvfzOWEO9KtXpgzJ2UluyJKOyYnX+dFHbRPwMffBi+gWx9W+O29j/dn36ltH6
RV55jBoEN6xkg/6i/PjzeGCsd2NjLQwBWc8ZuMCcedjbMJwG58Ve3jBIeKoR91ff1RLeFgGn1lA/
980K3z0zZHac5kWao9nqFPtgmEx/LUhzZ8JZZzpbBYP+4ArBQqWy2VFMyVgpyH9xsBRntfpqeLQR
Aw6ahv9XhiZ0K/lLkFE6T+t12sa2CKv7eC5gHrt/MJMOkL/iFRkJPjFZDkrMFidIIF4jKZ281Esu
vxGsaAhYWVgLj1danx4kAJoXatC1EqpiiQ2fS3fJeBFZfRWJWeUkoO9/mjN2AgztlLrkJevuXYsN
17vg2uDmx3M0HxvlODK8g4k0lwCBsVYysHzJjSP97PBTMDSDFQgQ3IRMmgi/IK4/P0kGf9dLRNkt
9vGOjEOcJNU/synQ4sVpcKZ6nDolNBGCM+BydNV/8qpv8haz6CYjsyVNbT+I0Ikn9jvPEi34fH42
qHLP3XqL3OO05zrA3sS32pJkSizjMdvmDkK0ZdrfqN+4dE6WCsRvPb0f59qsFmRUAXdUhn3AY7SM
F7FpJMUHOnz3/qED45KapxwRF/88xkMfHiUCvaEfIGCnrk/Pc7BX2Ym4uvEBA1ORQqG5Kq8hvuGV
Vn/27hzGo3i2NAMh1iBj9ilVdIj53CNn1Pbdvia/vaB8kzlUC+D42m7LaLcupBTZUPM7x9TY0fse
6VSjzmUGJutqHV2B6XU6xi5Pqulzt3PN6QutoyIH/LTNN9nmEhPHEpARXhY/BU4Lzu1vadDuDF00
46t25mjJOpxgXQLKYMykNYcu1P6WSz9pR36pLptPwf76iBNHaPUFAO1h9F8gGwl1o2IxX1viu/gR
OgOmDB2jccRt1Is+XExR2MYIDXWCLAjJMgmDvUb9YrIATG2Or45nzLShtpEj4wgjN5c4YmDaB4z5
NCU76rQEmfS8IyISG/N+aBTtE2MPSVl3L3EzxXZGTv6LBP0NSlJ8pvheTt0oQr1zeVIkfaCPgCEY
AQlMgQNBGkyYwPa742m2huKcsx4+MNaiQn24UUU145z+krmgBIm54Nl1WQNN265u/MI2Sg10S61v
LDnaQrwy/Os/dIPqQBtZABV7zEGCdVnRQ7D6FNd51sUfmEu7KbGwsnqti2r5fGi2dL98TYMNeS1w
yF20TrIGW38vzQBp82L9sQhQUTrAyFuGPb96SgBp2dF3oAF+dUZ1A/pmwFl26WdMoMM8fhZC1/M8
Hekb1yYGsHlAXtVjR1DMaie576ryGkMiQRAZ6963jih2BCekzjpdPYIwOkL97jkXTpsRMrn4hCxN
bNjOG3gHw82+haAFjwQKoySoaPtmdJslys0R8LtEliWSgM/HPKXaQr6ai9UEqVO8MpGHSlKcIr1z
bmkMq6/hthExYUEMiSIibTE4ItkNzXyRwI1rKgB0rqbRs/jhqcKqF2eEAHeE9lRIqwgyJwsT5CS4
Cw3se5sBCbS6Two3ctxGNbZaeZa/zU60GCjYQ8LN+Sj4w7B2hX3mDub08DQ0q+wubbpaZKDjLffV
ZXjXj1QItRQZuM1KpqErl13ZGMM2aaAVnqXYIPvlJzforjmSQGYr1iIuHlpGel4nTt5bnLgHP9Z+
c1jwo8UOek/+cGxEU/wwEZKONAppuba5ZVyQtkvx8tOPnCuTSa0mW+hCgc+TVxua+//Apk34toDw
9Fp9Q7KgacjyjjHXxqEEisQ9IFLELkUlRfWOnUj3nBr4Kp72v3jy0cgpbq9Qq5g6OL5vOCWNZkHz
7m0ddqn2VHziQSW1Z5L1n/T2ueKup+v10+tXF2b/yfSyVlwuRWcnCOxSrcvY9GU/nDrvm3l9W9CV
ROXoTWTuklsxUurs7aOPjL3EYBd0epnjA4M6sRHk1GzxLXPn+MxW3Y/FGqIcizqdX1rijXwhCHa/
ZmOTWD0YtaU1h6auQC3G7eq4YsNjGIeQyhUcgh6bpvj2l4l3xN6SjGWiz94m0W6e5ViLI5WiISCO
TpbOUYgSZFMG02ezBP50UdNL8KOZaSrVYNdFD60nWUozbNY1KrpB1rpSJ3VZHEpLMBQnF0O4R787
XUO8HrVRaf9cFVfj4lhKIogG5PPgmrg3c6iaUIuAe07mlpeMIkWZz+WC3gggBzmyAknhw8LACNFn
2vB1JYZOvexg7fesHRzuBnvaZBgVytk/Sr5f1wJkdCvIyBjuwD4EteWwIrP8Z2EkatNUp5AFUbNl
vqyQzl+KPJUFXfOYgogfYtTJsJ1b22Rkai1Yw+Zp7ToS15QQu8ZWJd/vYGenusbZmkReY6JcXzAw
wt1oYT4pmY1iPGyJ2UBe8LQ/aHRp5KWFCoVHB9Y4WNowgg8mK5nOZzlfe7b6x7b5zkWDUiF3UQ7P
N3U6n2gr+Uif2UK78qRFLKR2e2KJyBRvN5bf7GybrM/wn1cJ2694Ff7/tLZS7PV3i5qunbvEd+ON
vNW28a6CQqdNcsROsgeObLfxGJDD2qKd7W8q/YkxkVabhyWVGBG8KUe46ePekGSDxTkSTAbqet7L
PBFCocvYfPAW9nu9dXa7c3tvJ8DkHOXI1w5vYdIwoGBEoeGozsoRWfE7VtSvW2j/0G0TOjCf4eEZ
Eh2ilQTylxT8am0qo3n6pPYrTW1tR7WcdnGwy3Mc6zF9CzuUDVs1DwOM1lxYga1YEfSoyT44aHkJ
4HQ9OTUts64Zw5QbIqa86Lw5KHk+ySzhcIIGCxpKkxRL5x028mM0+2izvTYqf6JpvcLBqfk0efR7
5YvrzfYqtB+mTqE9raXuvI9g1hJuR19EkrdgsZunOomMGW6C2rYz8Xsl6glQAOA7FjRB8ZOHrXSz
knLImuuE6qAgjHA/1XC6ipTuN+7TUjSVoh3ZGzaZX6t03jBEmNGWaaalYNSrWFSCXUg5Mm+6x6xJ
wQCVg/Cpx6akdgDJKwmkOba43lnjQV5SOoFS3SLEryHKAmJjyav+ns+iI57xPE/eqkJsk1EiI5Xw
RGSs5HXktj+K0RXVriEjQ4u56FqFK66WvuEht6VmKgpbTq0iC7hJesLOSSoZEgcn7YmM6KfzBzNZ
kxUWs66gyu2pqXzc0HswyJX1YVBYBbMQWTv/e4zfzvw6r7wejjSgMHJT59cssS2PhTFIuPbQ6Rzc
Uj5SkmUQiU+APxUKW5Ek1eCLepaXP8QdELyb/icnwMpRKh4uwaaEHEl7iv9Z4y7+2AnwN3wVuNYh
sKS2Zo3au6HBVwncC22CVU2k/wjW3NztmF7WKuWSq3G1q2NKHOIlfFO6VJZBXcRmc4KMmP8McN9U
uzEc9hf1Bx5HLNbkTzSe8yKYy+qnbJqfIc3gkbomQidwx5pmURfrUbda97JT5UTIOXwbCCx8YDkR
yvGB6Ic3CNn8r7g4DJxQjRZmw8AQ4WDibfwskzAScIu3axk3fX0uypyOcRce5yYfPIhtJFK1pClu
uJqTr99M31Z4PixyRN1+tEVrLgnQEvQm/UpsSt/kw8Rn+slpT59Hm7KljY3E7U042wy6IWDLssUU
TJto5leY0PwNvA/eruEicAD3sZmxvgij6J91U1JyyCpBhxuS7nxKVL521oj1orhbUagykijaQ0ti
qjQ5kHxM0ZeU7ZmnIsXwn7/LrdEdr2+DNn3jGuvKrFoTn2YRxS2l8wZm0zH9pFkGMhs+spcToxqW
yJMXzRpNtg7BwqtV7oQaFZIdqeyfX4MVmjnCSkQBorATQMU2nT6mZbRZHQbaczbk0hiO0dxltusN
UXLd+VDLjGpUyx5dvG4/KbW5+w6B2lvWKk/536kWTjMuvzW6HAXUsQQVmr5+bMKLivU09P6751aR
CJBE+UtujTlLhMJqWCskbSALZLABib7R2C+ljOeoUvdODh8aopHbEB5ghkniwmCKE6K9h/k5pl7o
EJPgG9hyz0QV0PDSLrEHbQYPQ7I4NcdNH9hG989RoFfTKLQ33+/Vc9rs2BQmh/qWxILw6UtRIdAR
AQCaFchVFkprJsv60CAlITIQAvrlrKYNTj8pnpp0kgJpopeS58/2eR8UBJRtOo2H/xFvqVAlNYRi
nh6KG6OshMcMzmUyA37K0yKWNFJqG/wCMrOsS5yjsE/kJJWbsPY4JBdCdnQfKEFtl8OwCsvcFvnw
au6hs6brssMDU7U/E/NFay15OxQbjo4nq2Mz9ccedLlGr4fgE0mK50ue1oF2YZDnc6/pxHAwde+k
d60khtnyG7cuGABl7mxo9uyDXyMJC5j5sCgPcgs28VZS4ErsF9z9trkI03MYnwpNG/uenY4z4QKL
vkJdEWQwrvHoZvY0QuriysycWoGvQVWGo4lUGZM9/sfdBOYV3Tz7n+QEBhK5hjtcmygy5zdnWaBo
P+UxXpN8ikDgor5/LBKtLebGRYxe2THZp5+RtpdPiAZBw9nxHPHOmHChQnXCoAW3e1Ih7Sk8ypuv
hCiN5TRjQPDrVpQq5SvznDdPdJ6KQy9i71GPmL5h6poTTJBSk48uoZ2+iiJBx76DvNbMWnMUNT7w
ndRQTKwN0worLBDHuh3ROj5BC7tRFotz3mhgd7GX6wcX2Eid1Dc1/G0Qzhaxq9YG0TTmQXAzNrmp
fKTj8LT87DI2QFY7j58TwftzyEDZaOfISW+hSnznSpm7bd7jf+qiMYo4jGco/yIrYkFe0S/8OVVv
OV5+7YK1bnsJ2+e6UWCJmTKuxVlnGp/FPxRgw/8XPytj2jIDtLPJfeVQXgEyWvKdBS648SsDGp3p
Fj5f5Ekz1dw1+1w82ncr6mCxagTpJ+lm6hba5vF5qVY85yR33FD0STBCI0u6tlXL0q5IatpV4t6p
GJvNioviRLVZpIhxt2f7lpxn9s7QMjldP2tjkhaGvq8PlFvlt1QNVcbc/OQhvduUwKasPRKc3Eov
AvCrbqP+xahANVzGYIfQk3R4z68wHBiN8s7HzSq+Fn85A+h+1Zwf5PawNuabFc3wjlvx4HMuXwSW
+EjTKKbPQwCFsyq5WDvXXspY4WDSUFWnMQBzrlxn1XkGbVbUDG/tnrhusfJP13u/H2U+1etcj58s
WDHBZM1B0XmGGVGUvoPxzSQu6Ab50WXZ4FF6XrFnu0UvYcJPVC1/7kJ5TMoMCqP2yLkzi7WWI9Q0
LMESCuNWkoEN82qYt0wxFDrqf+MEnVKmc9ntwuurTRgTRsi/+ylZILpZ9+ARszxwsgRHuf5c3B/G
LHFUKCVCo0/OKSPBY7JQnh8tTOy0Rbg7ZfewJF35roYlw6Bh4gzOV6w3u9CtyzL6Oi7d9Gc7XjLR
O6y4+SryPWMpvNc/gKVizYl3kp+1cfwWJ71oqGDJClROuzkDO/aCwhABWjbnaE4Zrf3jvYP7kths
dDwuDAllfsp9YzY4qez37Njak0AqHMRFl06JYGo46fZeowkthZJKvOgHdbtV2rTRYWWXvP/a3vDs
jVcEfmtEXdTcAR2W3waB/6wPFXs+9mtuuEE4rliiJ17/hTlgm1rKM4XrzN8UzAP3P1nqo4Bxelge
Ym1n+4eZlEHN08zV5p6YLxRSeNcfnDizJ4YHQIbkPxrXfNVqJOtuXPBYP8Douizoc7heb6WDqoBY
ExdGgWGyMFVsfmXUtsAN8rQBOQuPwp1tKANKP8qXm20T5b55nutA/g96ZS0OGgX28vZ73lngOgaG
wlZqmGxTE6n57E0GdCFKVSejxmB9LXoBypJvj1aFdU+0utJhkLWhMqFv0Mr70fGGmD/FQ+4HrbIP
xiSHipdwnxYleqtChw+ewXQfUOOb5UvNgjs/F93WTd0QVn1RbQ5KfhSesa3TCmCRE9z+GgQlysWz
uZkvRk723xwGi0djplNSkBvy5TFxtoFGj+X6naHWT12AfApt4BwN7UL+SW9m7g5DLsmi71h/puq/
Ge95QftG85CBGVjCnAJSPsWwu5MR3GzIf9zxMQZMRcdorRqGiJD1DcN7rokNQbcsdQ0YGwcB/o4K
d3PX0oYl7RnNlHwX+d8WMrAHyDOWe0NWfGbOgJWM6HOEeZTwl2+MKuSqsITiDrTdySvBZ/tIuWSt
jTEbv/5pAMDPshwRfV9GeZjKdU0UF0BG8Dz7kQF+O5KmrfkEBIj54f8WKXsFw6fnP1IQ/h2fjFM0
/R4K/cCflwTzmGqDxMnEBHAX8NBGstOFE5414pCODGY+RVkSq+PltOgZ412ilE0X08bUJ9gn1tik
Co/xqrzbQYS8LPWzoGDAlkdxIs4WBf+P98mKYH4FlNTkvZPf5TxydzIx8tsAX67qn0gtG4bAVyQS
XfZ50jpmi8OD+v6PbjZ107uzb7OVcSHY9eE2Hp+IDBgWGQYE11MdYnO2wTInIIMHcjk/cAFegmH1
wvm3rmV72cri//sH3MiDPuI9/C+qZaGpjrj/Kt4mgTCQV6WjgnH5c8me6W9E5V7xp45LOMb+bS9V
q7uIOAQPOPrmJhAW6O46ruSLJivOlzYMi3McZhNIW1ymH9CZnZxxwGVI0Alyq51qD0V79J7Dm8lW
Agc4+uwGU84CVzA681VY+ylWdyPBRjCp02VvWP58UpWlvtNmgfHSliZF+l4cl02ixiK7o5FCOPup
6O99saYLd78XmcdzV1+nFgqg9vJQQmnXcNU9sdDOXC08kg6xelnTN9ga6prLLttisISilqvzey+n
cMnKzuApEgQiiHjoQ/XKft/Y7dkxLBm44gcJJJL71yKPoc/dmw21t+uslQa1kxgWdgxHvyZcLWwK
Ad0NXhmWMVrSvxJyuCatyve1FLXA4E3CZLpfD0mIZqS7k5DuKi0KubAaPoKBLn6qFfCfaXDgr+wt
fTpX0PIP6cm996BqzsCplWw5vrVF28DD4DU3fK3PqzNkdtp7bPFscLkLTX6ZCvK5fb6ymTAASKnc
gNWFcWa5BtYLfaKn/fqYPFZu0YecdHyIseRA45ivGG8e9+IC4tlsQH4bTaTAGLLA72W2dgpU3bQE
7FaQW3Oxy1cK0MVp5O0LfUty8y6aXzuKvfVFQ1/dRKrfdptnOAXhjLSX51CZP1fdaJLuJwHif6Ih
eQeB+99kJlR/6PIK18DhTKnBSOEMPdkzWlVeXjJbziKqpdCxwHSsmIVPzRCoeVlYkvcf4MIS8j1P
LDSmHOVocksexPKlrnUDdAmx6EBIH6f9fxb98/DjDHpEJWxP2PDo9grCddUrFuN2QgyNzi30tESt
lLVcYhFqii0dsjWekK0BynWWukTcLy5nUN4B6OTgyRuT8RRdiwwxOmL8ANbPc1BYJOC2pzqHIVW7
lk0pneW5VcsqWiwETUluEo7A6FspjHo+d/oxkYU3xv5znp5W4JP96G/R2tkH3qijDCLfI1m+4qw1
HjUKubSbuZ28ysTvmqpTnNRNeBkJ4CvgrrU6FnQU/KArQCTT9bkoKSt6t/M0Sxpft/jZXJNHlL7Y
cd84qgasGb6lJ06omD4Q5JLDewFZdYhSf7qrVAZ/Kl/xIOXKby3PFWnP4hZ5zsKFHrc8/MxuyafQ
H37FLRc8h0eSw1jo7ifsKJs1cy5gdKtZ601HNhVCpa3xIss6DGTwMsKbKv3qYb3IuPXRkpCyVc1Z
yTDgQVdaLovmC++d8nPCk66Vm2P13MJg+T78rp2p2wtN2uscw2qPe/4cHRFWRgdn0yjcinPIngG7
pd5Ubub24ot0LXlmtKqcXs6FpNkyLf4L8fyjEf0GIszucWuiD8kfBQ/jeezNf56h12szl+6tax1w
HhXZODqfMrRmorsRxTDKmjgkOc/wrabV76ZjBkfshiClDlGeaiGZmap/HN4zjE63JB5MhbtceUnn
A0MhtkQ7NqlxB/HEJ0yh1u1rLca/fKkIVPOkv+s99UA3jgK4sGUL+S6g3mGuzbAMyacHzdc/ENam
XLKRLT2nxr3hlUAM0Lg4gI/+goGKlCg0/fsDJZTTHjZ6sLYZfZHAUsT7SGV2F3bujl9B5vrNXhze
eYOl3ZunDLTOfJKr3F9JqG+AefaRR4dsLdIKfITvmAnZjmWTA2yak5lf3HYROqM6RLkdCd0Jlk5L
fJhSIri9KAzT/EnlzDJ57qgaCYUEFHo3A4znjef65YCml+CveqgdbLIqyay4WqCuizuxmHjF2r73
aREm7Vpa9lYdCbEdIAyiBIzvaa06VgTwy3PIMa3s0YIpbDCzkSKtNq8gEJfmBwNOpcDu+uZdj9S9
xPCeeZtsgnl5TH66DKBOsYRE71Kqv94KF6cJk9wLndgsp4VUdjmlAEZm7CNiy9Q39895j4hT4ylC
MANqNBINGcjtfl5oJu8irUcTXQ+sUwFwPB19+klxeLrfuUJJLypYnIYBkfbpJSHpOklcsruhUBg4
KLRoMTsNJxMyIQBFicgtlbmZCUuLnw5/MK0b+IoIULul541LkTanHU8tx6678jRaNfnByMMLfzEk
/RnTyRiLKKNJfGu1zkI/ybVY4Qu4MIu79Xzm+Id2NheZU1w0b5Ro061MZrfz5TOFnkq2/E2FhMA/
U8pSqBJFKQS08HxG8VKCy6Zo7ssfDI77iA+2W/6dlkM/6Eha2RxKCRXbr88fMabRbog4ezdr41xc
yU0MsIBERlXo8wSnaBaYbzocOKKhxIYRVRR5aVAHUp8eTmgVvJiqdK31dP45tWnaF+uCDx16SNvt
dM1lHIIlRE2uqEWqqYQsumt3jrZB7wg0FOrcKF3s2ukKVOrRyBgjKsMQOy9Wi35p/tpH0fYtBhb3
ZMA+DRnL49OSZg6Oq5aNCFN8gDzn89rio8tzVoTguxOqn8hfq0dMlN8fD9y5FGFTXlSyQaWmD/b0
Cr5IQ5RNxueqeKRXACahNNQT5xsYQcX4fCt6VcL1M3P9QM4FHZ6PiahPXjqXwsjnPhFWgUuCOEbm
mvLKUaXmOHXNZrNfAltvMsE5rgQ4dc0bY8e1SbklyDsXF7hx0uenjxTRGwxB2KKAwJexgTXn+jkI
GHxDCGnH3D3M+X1D2ns7oyPToKJv8/9j6XNvgxrZrdwwp9/1TKd2gXchkRMchaBW5nXzc5wWkf/0
5dPgpEpUWt42NM3tGlmi8HkpdvSN4PIadmEeF/t9IVgWAJj5iXwlsMpy0NpnavFkDV8XRtxXqlQj
oGNvMLycg/UUc9/XPwSfKD95xKXC4i/kCsTvmLXND+uqtQdGMN3EfxnLkTAJeJNdcROP53Sp+Q/L
MXdMMvVdl7gJXfe+8bXklQN4KnaKgo/SmLEm0GE8UvUyue/us/cAUaTcnC/eaihJT42TfhkUOnWp
C42DB0VDqK52ndT12hbSCZ35X2iYJryufC0s0KChGUW0Kho3h0gkJSS00zltPcOeBrnjb2o9hBY2
GX4aosKZEJJPL168JyggrCWAx8hJ0OfAAdb7qiJ2iAXDLZb700NesDQ21NtK7KO6a0Sm0wx+E7fU
9BDd2/BWox7M9P3p16sKhAG3LodjI96xkHYotMSXflAFeIWkiHq++QF4+096NGHbLkCJTaZb/1YC
aefdpgnM/2ePckuPPsoRUxEdhv4cBX+nDYhXa1qUBs+pRHQt8mW8pHPsMx/PSHP+cSBHOACyvFdf
WN1ZvFCRe4VmWK9CzBSmRDyQ3HierH2VhXG4rNC2wdIiiaAKAjU1ya5OFHBEVg4r/o6Q8sH26nMQ
Ypuetl8J0AxOrEdbfQLFKeafSUKx0hgYJ7tIH9AvzFS7ZshBt1++V92VmFN/oSiocqWR22e1dI66
S1gPyqHpu0Toomf5c0A3Vba6LktKCaYruc9ja8+/BkxNJws0MMDuy916sZhvrDo9uCyOfpsVwY60
0Y5CImySstR6paFI5hzmbS9WUt3kuNwtLjMvqtaBMiOZFc75PLwo0xP8PJJRlMbcybRz69O1xOvh
oSxgBfU6OrK/kCkkTsaJuXb01l4TTbClqny242al9+rOrFPIXR7tibODJgInMkkiV7c2yO4g7u71
jt5ZTulNb3ohH8bWaRjvZYNy6Mnufba9nc+yAQWOSlYWzLjEwpbuAWcdyh8ryRH4y/6eCnDhulKF
LCitYChmgy94O3pWtIU6ykbe9xhyBFvIFsMIvJLf7x+u2ka/RKUQ3UtUMMvqf7kD1ASeONowd5y8
S8/N+gufITFXW4U9YFO9W/x/ZEpNZGO/lN+we3md/i7DvbaAg8Hck7zcdHg73hBSiQdjWuiwsOnV
nkr7bss2ZRPlIcUsAfJ5AvJZZAhwTAYpwgp6CMvcmhDqIG6TseUMIYsgYRUlZnAVI4huql4fsFxz
9a8Fucf6hhiBi/29vGa1UQm78d0C/00nXf0hwZn2ELd8fbgAqdWXy1ubY+VgN7BrZwPiVlf2QbA5
kxxMWmiTTaLt22an4kQiKGV4qPv/kAJ7ZBE3PLHErd2whWAxpN3Vj9f2u89HG1Zhw46u5mdc3mxo
BrTdnOMMy56RP2pDupHAX8xNS6C7da8jqUYhrX38vQAyiiWUsL/34t/gvUNJQ9NL7q1+KsxZVv8R
oN4Korefim7+lCYXsGSi4/KJ+Y5wrwxHU2kgOr4CH/5SVLLrwyfMotHgOteK0WTfk8RiMDbIUvlz
oloBaeoqBuTjIF3NI2HKIjxKNSOlfXv4SCFPJLYaicnL+KH9ybJgxRTCki7cU2NHAuzZv8yycAI9
KaxEa1OmfcnVlBlaK8ImCHuTpByVLBSWezpiGclv8onzvrhwYUWN9uqmQ0bWRETomMGpF7tDKDKD
sFqXz9Tsb//CDX8hwDOWiLYNsH7Fhb00IPjNmrutykZVW5MyGDAQB30nowhkxiAz6vdOCFUu6cK1
Xy8twGq/V0ZlH1lLDx3uONnxk/gOMSXkKHfw/MS1qKoiDGSrlFUkZAGlny4Gc/+yYjfGI7LQZlri
skx3AuUsPZcBbk3C6mv99yVBMWdjJBagWAeKDOaSoyJWV+oMr6kp+A8IXTPsvqLj2idRdl0gNfSc
WREr4efAdUVk2c+PsAOVKOd59Y68ZVwmcjG/hgZj70h2GaMueoHXlwDzFDN+3QMmJmFUXIU/KkDL
DifoCmecKfCUq8e/wijS6Vyk1+AO/qErzS2d0AAjlxkNMLyZ8PXVDtdDH8hoFXue19y4ijZkwJFV
pbsIofv8OvSG0OyMYl0r9gA02xtImGrgVZcwILUbGbPdhFXECGxwe8Vhd5cgjQok+7bpd+O8P3s+
KkGyjGJNU3FFsMnWUQ091phxQnk+PtTlfESfTO7foDPtD24N2KRwghfLaOHIyAyNw5IDk97RVmWd
oQSVTWYuXm5DwqvAiVUiF+M5SoDkwiHAsHEbYNjh5/E6OThv0VxwJ+hJb8Ogcu7QXy6fra/9VY3P
XHDyqidvI1GT9XEK11nTb5Bt9h2NldtKJk3357SxRdMCus3Rv04vyY1Uzd0xBFiMy4YJKeXfksGX
d2uJXPJ1upX3cN+MEBVhCx/iPWYwb+qm//zfyFC6cELRkha8i4TpShONAZwSN0upgVDUbEBs1hOa
TWrw3lSa39neKEX87+kPs2iURzlzDBDGrqvArMdgOUBRD/zriCZx2b8h2+xvD4bh41wHvwA9a15p
Kz1hl+ixkyhkey2S9dmVi+l7DmtsOyO6JKOK0ezRetxSLihiq0CjKemCCe7inxHDOKDhGmdjZ+KA
HtEj5N105H+pP07EZlI1zwvZ858QqkleMPGvoFVflm+Ata7EJIzvaPI/iUdHo5+QXgl5nK6OlEt5
sI1CItJevttGOC8kWSca/bdWj/YTTzcOxPlieKdHq7XdMcfAfkK65tYeJD3xJFrDb5XeFiSUVPWt
zWwxs6ga3/gcTWI4cbDnODQV8UtuzJ4xea+8CVrQTNv+eKVD6MfeLO4CUEv/cXuhJ/OXm94sQaPM
4d1anVDKad4SG8WFbSoYViIyl8+xd/G09VrEYJtRjY2AEjcJpp70jIhmbcC4znT9Do1in+sWCai5
4r0S6S7gmdQC5ObBfcgsIKykDIuUSpqX+W3oRo33cFCM8c+mCV2lVrJivR/kRpnL4cXWOF0FwZTU
X74subWbQnX+GqbYQHfJhCRYL2P4qPhp4CaWFCpSZf5cprBoEomLPJhzo+9fYsgv8GMwBUjVcbje
2nlJPUymMwodajIRcQrvY+nArBVXwz7319A9dPuPbMkyygqG8hO1zlcSskUrs6mTwCYeytEVWtes
MSisLw2DEVOmHqutUGYnqCapLqTERWDSN7KJHmQj7uil27oZWBGpabn5ICk+L/glyfdTni1GTAEE
KEVYCHANvGKGXKI6+VzE9m3M2CEragdxafjm9xigsB6qcuB0QI4+5yK+gt2xDXRvywkBq141v2LB
R4k5Z1GFzlq5sNxPLsPOWLoUods2D0y1sLZiWS1jV0jgrtj1Ty0xB2XxzpK7olhdwG22EGA5EpTh
R8TYmDgKu6FlWq4DSISzY3TgcNHcJTr+z+BnsYkuHkLcXcY5/JIag4nmQLvoxbZYJeDkEo4dQ+ce
GHKw1CIu70+c6MyJPgvNQeDDkdfGraddknZWkNjI7kh3jvpuS6ssnyW28kRQsiYLlGSDxKaev2hK
6JysAUes187Kls7QwlkiVmiQYt1R+aILI5O1MbYVAxxIbwsxhkzTJKpD+kXVSTqkZoP/q94VW+/i
0EzCQtYJPxxZle9CGJgkYtzzI4N8GRrvEmRn76Ss7b43FqAvTsdTMnu1G5CJS+hDGyRFzN0cGRtR
UL4mK/IUDuVqEWjVvGVesLsP22TTVUWVR1P22qE0e2znmcxVEnoSXuiI+9T859BnVafXIvyiORap
9uL5Q+gA1y7hYkKSvlOQbGhSl06tnpjNon9PSsJzvE3Izz24GjW9UfW79x4oTrM0xWONUzhhLSV6
kJ4dLJS50+N5uYdmNJ85NohovmF5e/svQfOhgTjFd5BcDC3fGxmnb6gbdVK7QFRFyg+GlEUlGqgq
LjAmsRVfWclMKoBJPXKfRkk614mD+eaqdvt2QVpbnQdNyoQVirSoj66tXEHntoNNiu2B9ZtS60xW
betP9uhjPwSjWbRDrSupPSPaOwVNfHkAJOSSTA4LKqNXkf9KYwMD3RnovI1SWUH9AgpDTTbtDYyG
jk3JONgR4rhgdvJsLCBPE4HuRl4wnpW8QHU1TuIY8NTCn25nRETeZOZBFrA7TPhtWu7ymI8wg3mk
vZ6x+fVwqcbcl1vl0UlSHAex6t0ASIXK56Mrpf0kOH6XBk9H3sSEQ2wnbvGfa8mzj8GQvVzRMCzE
qubPQ8G3Flqd0IXCKVynanBTz/YAptJhOSTD27wJNX5RT/IB4B6gOLw9kemI4Ic8xK+5kPI2yxtH
BG+Otu3BZ8IW8rZBNw9v1hhC2vhn6ypYqhxrbcWQ3e65Dsbs9Tjt/0EFZjZHEAFsCK8iWFJBrvVV
tJvdJ5D4OmjWdp9L7EWUKG0St4ggdVkqrNum4Lsxr1R8hA0COqQOhSpTkIxJRHy+M//SHRAuYq23
OAsqKSUN2a7m8CIWlCWCeBEmhPU/qXc94H2esgAIsHws/qpOHyPTUWmVqpw62zT6DBD8b4vRdSlB
DdhdAcWHypsfSSMxfcTYcUTXBvQiUY5y+HMonPqZsqvsNJozP5rL9efIlVn8fEpH3ZK4jw0jQKUq
KVwuGw8QYThJ/qGES5m0KOfPuF+VKL7GP2Mm/QNFBYwEJ1QBa+RSRW8vSq571EHQ/GnBZwLb20dr
OEm8/dgpwtze5BLhdPnBnyjxIhJZ0PjNLpWWma+f9KXgp1m/WQibQCi1jO8w4gTDsCVhfX6qOn+7
hr7J6U0lqMW6XAb6KF3WU3pW5pKxs9vFcLVo7uhEls0iOXd+6qUtOX9A5wduUoR6Aibw0iH0R2rU
jnIf8vaRkBcB+kLRHzqYWvQjJ1GlithW+/xN7dMkpNBXP0T5R6MYRsuPfATQVAgpjkpaG4D4ylnh
iN9L3m4kiBEbuUoxglron2+0UkCqzw+kyT+Y+nx7QU3ZtSvSlOPe+YILgJX4FTWqr4CkuGmrkX3v
XphdKoZiCIfk94+VD4QT5cJkRbLEJZoPAF6xcvokysmIJ6CkeFCwkwZzUMpL+QBIOcB1zE59eFpq
kqxFD6swviLOlSLN9XW+s+H5MiMTLrcihQI68PjvvzCe5TZKklk0QFq1BxOpBDNpehkalqAJfWrE
0B1O6dq790G+5dWyB+B/QmWKbOm4DB2pbwaBJ95e5BAQmzG3CmjB1NqWf8QeGMrUjyYiknZcBigA
m6tehvW75IgFdewc8AAala3VsnfOaZ+3UZ9XgJgzIFudHuhNQFeoRBTou+45S6gFlB8QCeftDN25
b9NYMjYDBtNcNWitJQvfd8rP9CP1Yfug5tmlvD1ilmB5kkb3HQgHjm+53OB53W6hUE6PA+YhM+P/
IQhpeeVopwcF9sZg+sqYVTJwldnIDx/c26Y3XfnReZBBKyY0UofIgHix6Gdlft/N93RZWh7EgSan
ZG6pjgzE0TU92G8wWRTvKuGYnV4VOatRp57rvwDleEkrnU66OgQKjjEsIpjAAbrMDkOXbzO209/u
HaeDwKDtp8PElEDaAPrFuH3xkGKBVjNh2GPabVKrvd+yqoVH2IuFTyfha8ksf95ChzqPEBK+UKml
XheMKGIAythqXpd10cDUxMbuLM/MxkmPA5bJ/0R5X9WWF7cq1pZmXGZAcAVxgHBpSX0nmHCHiGVO
qoQtyyQPNqywfBVthecyVcxSY+6pc2Up6xTpsmHDKDCu6vxACQ/tMWCv/KumoM9Mh6mUlsAIMyKs
3XHPhQUlVPsToHTVSUZ7ieSziE9Ju4Qw8CWucrOGWR0JXhR5w0R2KatQnfGk8vdAltEX9A4/RXGl
RM9zfQOwgiodMGys8CESAJ7YROrX5mmhjd1vrM05EDiexIN7lxY9eVrSNd6voVqirAsQHMZzsA8T
Xbq7u1EUETMFdfkrCJQQ00ooufmBA3ZgHUhb4VmV9XjQylz1n6TPw1VXIjHs10Z4LGXa1q4K6t0N
KVntJsb1BuA+R1AiXrsy395G7zudscZ8nNzMnhgATKvpViBBHtLzRmhEcT38cR1he7RvRVwuPpD8
m5LuJ254aYzDOn5JwHxjK0xX++20HiA9eY1RXEA9rSHD6N6g60STB8Mdwh6mY7lpDkeyFsfOPTte
cCq9wyHnVHTjQOkiXT6RalIkwCwV/SlR1TtNOwV1K5UlsF94PVwjEt3eVjHaj6iR2e4+TPXYZauS
LXqALMdKynUu3+zdqo8UboiHuEII/iV1S5VRIiplrxF9G8bwGTJRXzljoHbGm3O/1eoenh43S0mN
zKRG/HPmrQMSHAmNgXxaoZOcTLlJNVU3eaR8LduJpBNywEdmfYPkI3+/XkA8fhqM3GD/91NtZmE8
PlaUwXo1uq5aEafBNaxq1jXhA2sXiB8udb6TeOAUXXGkofHHHKIqsqst3yvPok9ih7Vpm8if3KlF
hkIYdApTQiDAjthTj2zfA9lsU84u/bycZSJPN8+5SkIl0OzdesjZdCIRGuwZ8qcCc0d08GpmNCtx
7feegAJYlat7CoUQTN+xx7UPifIS2r0EUvaMkPPeW3Ely7abSR9HDNEK/gw1w0CrrhXpyW5iCMuB
toHVRn6ykfOMpbd2qG+mPkrhgCYZ1F14JqNj/aFh/oblzSj9Rbfy2yWMKerEpKfiy+wUQIK+vka1
lKpQfdQvlMdyzydU+3DalU2o4wExx+GfRefSwoD3y+hoZq3SCT0Sq25oiwyIoYuKpfHnShKCre3r
FAA4V8TVbXsD/bpRLYzr+7vLhDg8/+8TSLdrBqfbfOIg3WwWGUNZyQkbafXSbtiJ4hkZLvKAafKe
U8W1jZFm/bfX8N1YpEE3VwvM/fL4roruzeg32fVtE3+DBY0i7k6O8w0t5yNVFarFBlncbIpI9k+I
jx0gJOUghsuKeKMqUG9DBze96UfrUxmqD8gBoHza4XIbwvwMzOAYJp29HkEmilspoFtUMqO2v5fY
P8vlnUlAnBP4au2lXqz1lMQniyXhw4ReMDBZ/AtKfcQY4xeXcbFxiDTehe8LcvBVbW9KTNP2z7UV
eCK7ifVzT5cDYzBloLwDx2IxzIn8kRJM4YL/KOf+VTJt3zC6tVcHiwW+KqXz2EZUDjTwU9tVEGSQ
UbyJN+k7wBxiKHAa1V7kq7N7Ol5+C1Rub9NzdzJES1PQ0e5wt4RU9KMKETiEQKr5rwYeQdnDTRdy
dIEDSguAWrXKgYYNCl+bdNd0b56dTG9Yw5IyuXvGAE/4qGp4ZMsneimpdTiF4nG9zfSXxKKhzviU
NfRZOmiEsVIXAHocrpWUTyu+kTPnoz/tpw0Q3YBOm5OjeMUv6pS9GFY2eDwB6ZEjF9gBM0ib84cu
bA0u9phtlf38/lfv5LfdaPdrO0tBSF/wPy42cHH9XtsiL+UhRuocnCAgh5JAKDBUu1DzGV7ojvkG
uhn44JPULJy5F28FGMzCw6/5m8mfznO4xqgAPBTEg1u+G0S9F5IelMVPg9aPNnrBTT01mKelgyga
tsBJDBBjkQcTNGW1v6uvQxKBiedjSS+f1gOEbV+ImMu6Ltv/o5vs51q60mLUMi7rRQFpu/l71qLg
Iq/igMxcWHo+3ko90ec48S+Hs8TTOPj2+BEmcuKdxzGCt/2Iy6yGuoBHKQU2jQhFXxKpyWEHLsa2
xp3TO0HLX5j1ArefuBhYZ3K/Sy5knsvqt/KajnNgWtrJEzmJVmexWygx5HRCCH2QMyvtA6rX3LbQ
gr0N/v7FqfzUuBf684E5gW6/UB6Lx9lCWYFFh1N2EDuaU8/Sf5wN2L3OVfbSZzPpbg9qkAt5Lshr
GIMC4DYCFZxuTc9rYhPYVudkcZWAJ0kfNBKB7+RW/3diEQXF+X+tM7jdUbLOv3nkg61Fegi5PY/W
1P435junZ+xBiMwUwZbKdCMtmV2wziN/Vosi7CMxvKP/Dz7wHSzd7FR9i39zB0brCVjWnTtdgN7z
ciKmUO+nt3FnvG1pzHzHhHdUOlCj5W0DdAvfwUVZ07qcPKJ8xLhiX6Egsrz2+Iy4NrMXzqY1k0Sy
MbaSupFaRxKm/wybHULvo4OpGEp+kaB1wIpS3JJ2F0jixM8mQo5ZXpYwsHzps5HircJzeluX52WJ
VytJ1j148uynfVhuwXxr6qR1pnAwLzEx44f9Tqm+XqI8F0LafVsTXC+wi15mgpBFM3DWPo1u2NMg
k2lM069nxaj0JIuPM3kez4zZVwvQ0j2GDY1hsnStW7ZZ3r8rVF2Oa/YV8pKzE8w0PiIEhS/JFyC2
osqS7zV7EVbYFxz7BtGN1T/2LjCPkgAizoIweLng4g55pcLof0kqDbKJ74YqrG3+HXl5GUsr56cm
/oFmhn05EX6M/IAmuwYse2qgUWI6KY1X8UKfdTSoP88sMKEsHTC++UA3gB2Cuf9W5pvIKMIvQo9X
s6P0COHqW7EsmQbM+4MHMkqzTvlrS56UixMDfWZ9QuxD/oWGhpNkxAcQNvT7las8cBMu1/zivhtr
vwJwz7qKA8fVvtwK9vLbc64LU6bmfIJtfNk4Qd6ajkjRUQtwkhDPlKdalFXKaQCCVE48d0DefA6v
G0Zqd7VXiCE8GhDkNIe9WpU2aGEq45Gefkpa7AYXRdUpIVrh72ceqFZDAU7h/KRkTcBEfkWrDq3b
xm+0+vC0OOZD2tQl2qwTZrcSHXIqa9otA/Gvy+VgQAUBvoDCdKOL0KvKOwjtXQ2btc18JCgFzYlj
UeOM97yHNXlvb1xZzZ2TqSljWLWQnIopjmapvr4UKx1QlrIiTcGOehLOXsJ6b2A0+6i2VrFHTwEy
qGFcBTc44Uy/9mxk/iPxZoFBfLEyVgDybfS1WKscd6gsyuRjMM1gP9xN2j+CMGBC1g/XlZxelHk3
68roA87gfjgQW5rX3uWUDjecXo8XQ7jHRmOiAcColpI7cQJgZvHuheHfMcKVYq+tsNCGJY3LX2lR
Jkp1jJV0sY4JQtNI8ZaPE12Hz+nWjvB5iSNrI6st3cc9xrVpWGN24ZXTiq+JXkSNnSkX+SGwHpFJ
A6Vu6E7rdkqHw0kLWLM8ArUWZRForKQ04xTtQ9hmgoyid43IVFzl7pgO4U8YHcSJ9u8n4AFxmkSK
d705ZUmImcaiQA941AhHVcOX8+XIR1hCfegoOd6HwGwCOsBL5srpdMf0ne/LnOSZ3Fvr+5kx9pK7
+wGMyYlTX1X9AsZ1wXr+wdeeiB7NIG7l/lA+nABRwoabFOiJI1yq397J2L/PQjo82/OvptFssDJt
ldzzJ9r1xjTN4km7Zb9ghyR2mNlbkr+DVQ7yVA86n1BgXC9xeoS5B3fKBPxbVKAF8+m1gyRR3aGc
IZ+KxUr9mtm92kXp7vzRX3oks7llhMDb0MJW+c4LCOX/6j6vNMOjcsZobGzY5iQ8SI7g4y/Fi3V1
YMDRhd9ySd/V+r8hw9ubS02WsZ+wT82/WVVxAwrW56WjdvHgS/+MhXgUBBXyozGj36K16SUQut8S
6LwqjZhI+hXuatHFkuIb7W3xLz1xnytK0ny2FpHtiWLNFXrqg0RkV1Fv1pkR7mhiTKB5k1xFfUMZ
eF5CfYT8duUxGJ7kFebX8y3elTPwLmRmc+jZccFvie/9gcyMgHW/+wmpQB3hW92Q0arczdQKln4t
Rq/rX+jtpCBj+/7XklM1iRG8QlZXX9TWVqkbWip484qmr0SaBe198n927A4yQWJuIybGMIA82eEI
2i0iGILxoDW8pjTNYuCdSROkEurv2tLg36pWEOXbQvMa+rtjC6BHmlaUIEMf/iVspptdJwMRvem1
SRzccahVipszMrg1J1t5iiQk9mhGCIvIxtmn+YWYWDLY0xlBOz/IsPnw4jPfk5G5kapmqhqA0yU8
97X4rdk2IrpQOk2CYcdNrf+AeCeNCowjJdWjKRWeRP6XBRF5DPw3z3hUjovjOAuzYiZXN4BmozMT
hzXKsQAI2IpNNk0b6D6A0yzQt2fz25a3VDxLBMmZnYF25IQXwj1yDzHhvaWB4Ejx9+qHJEgmGdur
R9ii0mJzAISOBQrFDvSgBRWrNigzgo/18LXzE4FJrtEOutHKWlJpEZij9dN0tk1FNvA5RBQLjMRT
ykfRRIV1J6DNea3pU6C1LnYO/gch7K3BUEmEQxTj5YS69m5FNOyAh4Lzs46QqKUXzuO5+y+CU87r
Yd1Tk/8kx+hc4tG2jCGFRkXESeYz/YEIdRIwFQcbQU2ZQeLAH0SdFt4zndziM8WjGTHzhTUUeVUH
tyy7ylJOu/xU4dx4H7xdbRxUfvtD1kj7LjW9zYbyls2upe/wEMUZN5svqu9VKY04dPOTnaouL1io
Dm93rnwuZwBw3EHwin6Ys4yjryWplBOmHHnwtvK9olU7WVYAGWzT7iT/LmNzoE+ySGn0Y6SqHGXZ
iPZkLARl6BMtV6BQGd3EpYawdtMzdt1rHjiBPb8EveOphTidyVsmzY8kbUtzQdWGmj0yn5b+Ku+u
+jX5NBFkznhfcW5xBjWy7E66N/MGkrcTnslL/GPcJ1TTHLd0dOJ2jhVI8w/eHyHXlyxdGWVJyqlP
j9I80Z4RkrKT3ouCZwRWat6YBRD2wY8rt01a5cQvgBYgYVpUF2R84vcX2zpzRBdpymIRHPKtRGpc
WL/fIcLCSBsR4qoiC5Y5mRdOhnlDDwE16M4xEDbJmhBvnkMyNwM8PK4wjYp3CtRHL3tIQB24ikrH
t9xppvD52R4bwCzWZ0Dx0gkPM1vNKx5EDIfPnY7sWEVcWbhDV2Iuf7CbLaSIDWLJ5nErb+0SRQc0
aJ+ICjjFrgbXOpVMzPGuUbpc26afSNweDyIUQ7fkKSpRIVeyLMhklTeTBL5FNbeyifaF2BxGzaya
XEYu1AIGQ/rqQcD0LXt+u9KsyGGMoF2SjUPwWK/xZ3ZKAgMzpnuTzHPyyLLNOJTNX9iWw2X379cm
X2v3H16V4tOpqJQNqgx2A+pJzL8KH+hLQL7GioNAsY15iV5T/Y/+qGAeryHXtzoLyA+IINY9FNcC
aXvmrRiifyNR2X4LuKTk1LeJTocr0bzyHw6aY2MXwYWevwNHpBrcXlT3b+VGTRsvUTn4i3mpQk2T
b6E68BiiOBLrQyyr8Oybr7FWdrFbozQjNNuuOUApN9+GGakKE+84Bg6NrcLOcQp0p962V8o51zkC
qmCjpqCRrNpfkoGqSC0hbsYxsTAuPHIhNhDo96DwF6LuJMqYzWXTKexMLDdzzUo1hRW1ReBXpk9n
DsmbODyfcZpf83hKhFQ6dtc8WPQ5i2+mH4nzptTLCPbAE1LJrlrMF28+uWXdz+ub4hiQTTSYK4EA
Y0DmynPfVnR5Q3x2maDyzBz8SqTY5ZlRFqnYNY/HxLtF5r3RV7QZ0X+yZ59M2F5l53ywVlDp/xo+
W8Mg/5f/IEoqEiLrRCMmOQGpNMmFz4eLpbDM784N4Wvj5UbMBkkU9jwaOQZOxPOaGdE85hmzomRN
6nhVt62sXyEZQGF7WmYNCejRM1XGPhhEj2UpsmMOl7EMGLisJh56s3GiMaEuQL2u7sxjG5QAgH/B
BQPKEu1+0kqvpmTOPOeoavQdwMk6IiLzs1PeqEzC3fiC/NdZLXCvm/8rIkE6lDrJEd/UBgLSpX6v
a/H35oNVH+a3/Bj/58A8RXmGFNeub+tUATZjuMiATpjYbzUsr3lYHN34L0jElEO4wW2JedfBKjRJ
CWaNXVK1yvyP3RrXKPnk39HOtPXoLpAwbfTEDD1YNopYWR8Uozv/qg+mmpSMrVA48lO7OOWxk3lJ
FeBF++WD4OSIaVDgl2q2gxSlPAObhTnd0VbH/pTDRnRT9ZM/+QLeLwWy0ln4ohLcS6y8XHHr+XIE
EkOGeeqPac9R3R7iJiqtYSlOJi+pQthdBIUBV+rfZqp+vsrYH6NdKPWMsgSh6WCDBzADZ9dg5kYq
OW5MxObI2rwjhfYga4D8xqecjyF+LfVozlvHgSPULjqmxMHQL/lcv9VUmHBG01IIUQp2q2tNc+se
Xi06XPN6k9mh17BDUMfwysIW5eL9Kh5wsRGo2S+qRmGASPnOSHNduNgBHbVbedYGq7uadfc8vG8U
ILoda5u8HBEq+XsfuKvhEqtSlQMsPa4meNikIi1VtNZ2aUkGPV2qjh2dbOycBeSCzx6ZEUpPpIoe
CgLyafRxDQImhDpTAukmd/elvZzlM/0gWCK2QMP++pf9aUzVuRF2JWxBSMaUAmbLmvqrUTodWlgb
pc71ZRnA+zNcUcac+A07GbADo6QHdJLq2R3mfsdY71UCOvxbKFFoba+wiPXGsj3coJwzPMWBDXt8
uN110266fwOAqqZ1pPebf/2ZBdX+C6GWk6LzoMaLsJR0dToFjU5jx+LE/HqFg2Mhc1q8n68QfA9J
A/IacjzIyfrwrk2bIMc6F2MU2j7rKyJh3ixWx+dIHUigp8J3K237BlDN43CIFA+zJuXloFvduWpu
1JhSXGnWDcBgyMcfaaPbURh7ihSOOWQ7k7XkfiWUcRs4YalwrSR56lZOa0S37m2aRjSOahQPBYw/
tROrEGtqvHkaD9SDQ/19rz5awy49HEtRJiVKQY7icQlEVqGWm/EYeB7HkGlp0lLkSvrJJ9qX/b5N
vSTTe7U5SB9t1O7kVmImHiGbkvh+kIuQnM17Ig987lV0Qc2GjQ+INCnUrwTI2Nwu/R8gEC/TA7YA
O3CYgIm41h5Yw1WFx/owPrgNpZ1w75QYRw0rXGc7/M19xgKBWIkYr0b1IFpho0kPsD6tottwbTKV
8VTmn/w21IDigXQc1mLWVRY7E0nxVKxW3YyDuxS5rU0/75Uarw8Jw2nLWV8DdPBxZvnqOV9D6k+c
sjGJNTlCehDrT9+1+xFY91WBwN2U7r0r1i7NcH3RrS7T5CxB7aUtuCrCHjC18e+UuG+RHrolTBND
RyTJPI2iyTxdRnqYJu8QTR3tz1oiXy7E2e4AxM3KDyO9VW7joMqkSnUQCmN4LTvbQDXpisNDsTXD
MsldRatRlK/w2iieFlzeg3/AvJ0RX1bWkfmNKokL5ROnaXP2FvRJ+KIK1Lc5rScfZL5MxA6mltwa
pws4iu8nHP7uAmH5zkxL8VljErGHwT2aVunLK5TRBTUpPK0+fzmVatZ+yfpGuIWSjNaX2XFaqxj3
y4/AQE9wpnZKw2j4u8YMEJRlvLhTEXYyFGp5YEj2qHPlYK76zxXgskAo2doFip8BvZJElIYo8Xau
2EQoNMZlblQ9XfFQzLXj0RtrgEOV6wSCf6kP2Vsz+0ZufcHjgUiGalfQw2+Gp6T7NaFJG9wUZUnd
K4ok/DgSqpRsJXdGYkbgJQmF8OOi83NqB+V86HGg2wOexWfNvV6G+HwjYKX3E1lh05CnZkwbQnjq
VkKN6DyWqtzGhOCsIdHyHDmZYq8AyzQ7InDe4x0eLJN1J5t5HweKt8go2Ohw2gFyXoIQW1207A/t
usDLQELztuRM3+mSx7VbAKiE4UrAh0iwtP5OlbtQo8mHhEZzOqSnv6Wz57+YP1gM7bLfey6fK+bv
+qKniTZsMsvbyCHYF5P9gYs3wpaoHIGFLySbHBSZWGsLlzpA/Hmox/J/XcGZTm0dhNo+uWpQyzyV
s85c7XrMqoPuKqjDKJS9wOWxzDhzjUHKqk9p5Zd0zDZku04+H55oKa3JbKeSsurzMdbrSIMwoWR3
oIhYGKcn9fpbUqTigtIPJEtpoXcrPfbJYbmt0wc/P04tCdwbkcWDmclTpDl1GxH3frmjq8Ed2JDO
HSk1Z/0YN3TptaDCvLJ+W8cQmO9q7XVJ/KO671LL2MW5NuY7B9HJBymbdJ/4Xil3PNJRqKetcRCK
JigiHXsXsmmRfi/vxVwp0bhJ/JjMLwcHPvfoKIfvUuKInGR2uzyy6fikikuwQpqR4xIAZLwYCl06
6HQ5/rrnsN6a+/t7bhsNaIOX09dld2nI5PDVVd87D2KhR+NKdkhXGBXFxOLsVb0sn7ZJILW0iFg/
1H5hXXeEB4LdtoHi6z59muH+k0hLYWh5bBU9GLXCKlTwi5JQnAyman8zbcPt0aV8/OCrLo0vYMnj
UvrfYdLL+V+SsdY776ntKwl45llJbDf6O7ykR93ub2otVt6PJz8yj7TObUEfC0YWCKYFkOOlhB5j
UZP0UbLWImSV6uyhzkK2TTzR69ySBSFofZp8L/UWEVKCQY3JmtgZC9RK+cmKqJmR1kDy78Wf3pWq
btBynsBnndQb1wMaBpRZevwrkD44g01mE9gR/D7BeEBo2MvVMS5tLIRvbXU7ro2m38ibWIWJK5+u
XofhdnA5gIR1doIrCN3qgeUXxp+R4X18MV6/gcf7xAjStBG6SZ0p5knUUZhO7sCSHg7hZoPdWqSp
A9r54JoXmmKhIpUgw8XxVe5nAqEvAhHwTxyimd/a+25CPTriGjEnUKnh4CdJaihRNu0KBohu+vdA
vFKZvQ4hPMMs6Tr076hkDH1dYc6IvWv6R9I1FqDygm2Kg7Xzfb775dCzw8P20aCgQVqV1eSM5b9c
fGlpNfJb7IJvWNIPh4Cp8/CoisnEnQgY3x8Z5ThZWZKx3Ml11zyW3ewyR7zQj8ZVTVFOM3RhK7l1
fgBL0sm4gasqDgeKg79btVpnP+cxF8fqOvnwWVmSaQTM07S2vhltu545VC/DXofri4/QUTjSRD5T
RNHjLrzrVeTn2mWpLTWq+3dGdNbWUeAhHu3gZvlv0hLP16HzfqyKuMG6+p6ggy/XpQE15xKC45Ku
/4Z+kIRpPC2MBEgdbc7163EDbLdViMVokC7BiQz5TuFc3y6ZtKh2c8oAWkIfRKuKxe92EyTOGN2U
vnW3E0D5weZcZG53+lknVhM5jcFSYhboeNLtIPpycddF5o7n4II8LHRRP1FSXtuSfCsk3kaiKGud
ZaMeTIDQ0JTh6v/zwPPvH05x634GRprqy8aDs3F3N7QS4lxGimxgf7uI1PDOwBrsKq03yr/f0qRO
K+pPur7cIMnxp+Hv5R1WcC8jqBD8ZCHvKxAnsufzHYD1LOzbnYDJwi1i/ecBoQG1eIkfy5VPTjTY
9M1jMCfXAYtXipeO+KKfkSDYNtOf+kO1UFmtGJpf5aKvaaOFqiGLXPMyZiUmvYd4wcbAEkFvSJNg
kT/+H5INLM7FIND8SfPS1Hx0DvI3L8DwCssiLiYVDRI0ns8vlreX+DvbouVFAM/YR4n9/PDF9PO+
P4DLOOUwm54UjeLJCaOjzbxoFGi61nDCz8hzmWpgOS31issSaj6MiIzApOKiQo2JUoBLvX591EOe
0Cy7yr3MYXiRYZ2P90JXFTBIIlxnrPnpaXgQ9da/dl6np6AAls7STfmshPWkTz3f5LoMUFYGF+rl
mIAHoSJcHiJNU8JEyFn3lKxWODH95KpZbEr6IGtgfcmKhGWnXW4vihHoE35dYwPox43kQMDnGvm9
GPS6ukG0S8GBkh75DjSr/l0zoJdFLF+9UqTzbCBHqvJEy8Ul5Ux6t0Biyn7n0XGjMJaUQt9CnNux
3X0dAbV3JuFjhX2NZS+vomHzI8G1JmWjD6dE3GrM1p2bMIdWt0Z2UdH87+HQbzEP4Nxihl4ZZyU2
cEIOCAhk0nureZ8rdroyYHWuFPP+MCGBzlbISQ+/dnuOh76MhU/f2nFd/7bLuHp3kbcXNjLxWDOJ
3Xqg6qPSvp3orfLEDB+MVt7ANHOArak61ZAH9ORPTLmU4Lm9zI4el6GbuqKdaLpVgsevZV2YCxoJ
dF1PkvvvQIRKhq1aW+S5aDoxcOF2FyIhJtyXCIgxHmBKyLCpvUZar5mErmS8MOCthSskdw7g310Y
xHshvkFaghCwnicSIWFfzfFkt7AAqR43Yws2Xgx/GMahdLRBKW9Le8u8Dps7PBIXIsRwwEA6i27/
jnSjaCn2f2uyUZdshYCSeXHo1CpWEWBxDrYBCC2oPy4/MhwZZg52nd8dvBgbhjK7yvA3r5IxFg1o
MHfVwqgHvp6LqUu2wRV0yWshy0vDDe6bBI0FSSir0FpFi7ktZ6HREuFvmIHIJ4V++i2NIksgIzzj
YrX746fVy+pi9FwcY0/6zdtAtS6lhxnI7YXwBqWUrsVeaPKTjVOk80nY7QKC6Vj+D95bApi8ghv9
kjhQRII2f0ihQH5sWzavjBAomBMs3evA/G2TZpm8x6eK0neGFAKz5hxZ7bxNjzZ4jNvPrEqyL6dR
484oJcjoNcyEXYE5psgliJjpA/bybUGz2hfe5ygma1C3qC20T02SiPg9ebHKUEKgOaLuLHhCtpOI
VZhhPiSsgQhEV2Z4KKSoz2B/DFqGpIaTWS8Xn/0p0k4wlXqH1C0Hzjh8pt067hXwolIwgJaukPIN
oNBmda0anPySQE25n8SWb/0wlLd2bLjbgRK+QhUN5djzvMrZofLUixOVulKjVSoANELjTxzm3TrF
y2nsrDfULrYniAtmaGsq4vBssHtneOPlwskx3zh4qJXTDz5FUWX4Eoj/NHyE9NT0DKQ25oE6zwl6
NWxrwee0AScy9dQc8QhWpzXbi1gs3PBGACTRjHPfMOlX0yj0LLK+rgSyWN3X4BKcuuFd6bpYujlE
U3sBmb+wy8gS0jHENmj2b5Y7a2I40vXa+QLM2Ja7dwll2EmsXV9IVqfWcYd+I17aKGF5L9jjBqtd
jBvNohujBYfpo/fweWnaAyU+t/eqI42z/rSds1rFI5D7zVGuDZYgWxbYq/0ek0cQGO+1ENArjhX1
+fWMQ3Uvowctq00gv7j/42Z1b8dd5mWtjtAbTtaEuNYT+4Vf6tA/tsegUQQNIPLQnAKDa6nDtVeW
fHa/C3mElpw8g42T1oG1J5bZFke0iiRwjxeMZ01FuncPD6nwE4MunpZIJpX4fQ8xlD6QDlJHcM2G
noDtjAOAWQmG1j1iM79pP8BudtzWRO16bSjhNklwEzkr3fDOOQES7JFGwtzU+2SmnPXmpuDDn+Bt
uO2cZinYFVEJSEROY5jt3uvxgyYRDcwLG9uRkuyEPMnGIZDf9TCDLxZ5cKCmTibk/N4MKPY02hXX
cDYVw5sJ97ISmlJYEJjRTSO0svlvLjw6Fx5SnulBk4c1hePejB/KwyznSQqsrroz8Kn51tCY2Zbr
HFh9j5l/opNM9St4n7qHoQQhMPOryVN3/bLGHZ0E0/5y3W3VsDcTA/7wyuF+tfArMOMr06omTbx6
dlPZCtOBOhf0n3lliGcMd/+ROc2GTC587o/LjdzB/4ULxIrb7X6P9U3sod2Fpr2/0jmkDJlPo1/i
c8BgC6kx7Tl6j9Jz+ivQ0ictznj5su1G7FA9xBZHYG9DDhufCCijdYxUfkw6GTzSIO2qwd3IfwS7
9xgP5eu5qighL9osagqvlO8bHT9Tc3DKMMvvkLZ0rcy1AalYc7qccYl+weQzS3bJKoUpaupzc/Ow
SUzzlvyZ2lUDceZP7BL+hGQxRGyfnKm1Q5JBezeGbp0yYbU/775mteWnKKiopYldO1Er+8o97d0/
U5WcOEuQXsFnVypOYdWrNQhAjudW2XuMBu8U/TZRYUpF3RchuiZ0klehjbZQ6zsSOLaSfoR5vLol
nCQAJLyyegsDuSAhQAjVbMAuh0oIfrhRxlV5GGjxev00QXoHqgms487hNhyrarZ/elIB16qlUHEj
VO27Fe8xAZtxUWh1mXXgEFQ2wWTddEx36iyIN9mTUX0mfXNxF5pDQNF19erhbhdzKPmFWHFQcGI5
W8NbLAqvopw5db4tJUmFBoKMRloYZquKZQ93IR4P3ryQYhOjee1poq74mmWPKqOdAIWX0oghnkni
XGebD04tU9omlkW6+IIwnl6C3qmVEjoDSXknuAgt+dE+gSMcI7oBRMIQ9myTCgiPHcHoh1O4RRPU
ErUFlNWESjCYOVTsu32Q5xzHVpfGtoZnF/0+8n3sVuzSplxvBKNl9bpuFZCAoB+FR1LCjpJDf//u
+JlylPJvVgAbDiUTSQGgX9sgAQd94L8jWtxBg/FnyRnUw3AzHKE7pwL93/5QQ+byg9YQE17+no33
ykGe/EdG80Po85i6ygSSvTRcMp8d5WKuDu/4ElNJuXH6+fDXJxqPptzvPOz9vd1LMqEm2+SVCZ+M
MfpyzYT93wOda9ACY01UKW7ThU4n8HSUquwFnhkpMneFUbV9PxtazV9bA18xPZ6cJRX5CySdLJi2
oHunwjntWK9d0T9b4aJkCpnZScIOoqvmmQTq/S3M4FYdTMUPlcGJ6/6XSQ8R5yeF8y5U1FDPbcfQ
rA2Ngf0AAcKggCTrRlVCEXt6swi70E26cAZuH0feOC91PgJUJNThhQCljA8tc03x8cgQHoVRZdRn
vcstPLpvkX0+cXspHNbnW1Ycyihnlfpmlvpcq/39hQ/DeW5iCYJaoKcd0hLPQ2hzGJ6e4W9COWv4
GsxNKDikTmQ2Dy7pGzK6B/C6lSPEmknJeIc87ksfiRBdIr9DnwbT4HX3nvnHHqGv0D09n17CTCTs
dklUwngH+EkhtRVaMRztQqrQLIYmIO0dwBLDua4pGghDGhuGV3IX0PK8xoUGI4mzQX9cceqY05uK
nSgSZC2IJWappK+n+ZB8BKJlync+5ia5BifbLDnGUykcgWxIAg+vyb7W0OeZcQcKyAjgW2UyqhSi
46cv7m5C5rSLZQb24HM1/zyqV/yrpc2MSrXT2Z7IgrWWcNAu6RndWlAOx1wFMn5EW+YpAopIsQ2m
krb+9VT8Ipb0T9UPEGMLfCOnkkCwHZeK6ziUwGvIkMfJSjJLOyDsUGg7/B1x1Ld1+6TlTmQ2pp87
40CayyQcOQbdJadg1vrBevx+DvgIPCz7CtIibxZQZ/3uuZT10CgQO4TmJExOd55838Vo4IIrSAbk
ftfSvBpecdgmO0IVkEmlm2KAQfegEI2Ys1N78rEqHjvd6mWJq5Ym3TNEgxmuI+KdLiGdu9HvSp3N
uTErTKULFtV20CI6f/TABwEPwP5dW296een2HsdssYfxGtecO1ORgq0t3ApsxscyKE11mcj1/FKk
Pe/K+fa+KQTc3qUU1fpTciuAkfFehVXdQAPmTkVjRpQSqHVFUAcYe63xhE7aynFUWeU08jfP5wS+
/hwEt5ViNAWyfBAk2XZd818U3kfC47em2OoeaP5Tv1khpXvHRhroQTxHfpkNExNVZFxeTyNlCVoc
v35xU3mdGtqvIMinRlZ/0pyTkUAP564sNIs5qkY4Hey+bTfm711flG63UFIChL27WLAsg4QIcXmD
ZjJBS5Np0K6HdGl489iEEhNkm4z5NznVq3DQXmuyjGGL5K8FLwTuUeZ4ksA2Zy0tKYVtCAfYn0Sb
lU+H1rMy8NQ/j54pXzO5Lkf345nHRGZy6ZoER1EjdN1k5XpMk3f4YzJrlHNwZJsng4tGSzeXXX0k
yqiHK2bIWXZ9RJzq6kripoqABFzwNGt2o+RtlcqjsmhK/MRbPaPfjvZVAzjAWk825X7Lj+jNqRY9
CzhnePtg2UxmjOlRtfYBKi01WWOPXDz01lFgknyq7owYBlR4EoUpxhYjPSOeSpobQfeyWpwXb8Hn
ZF4I5VwszX7b5MDt9+pyHAfv4RcUG7p90v7Op8KpHmR/eLRvDYVViuXHEvQJzG3meRJRkQXDA6u6
WP8pgOi4omMUOMLaHLboQrfxlFlfog4yNsFnBdgksB1IvWdmLamQPalWz1KF0FSjVfNEszPpyKe5
akBycv0D04InWosWDKzmF2HYzMKk7U73m9l0S5HE2+V+pRA6qdGYi3gFFhyV7OZa6XdhBDF2xFq7
Njn8Sgvd4XFBqwFXN9k2WBmK44vPShDMSXm5fyjdcu09ecFMfpwQVsABuZUWGUnFma8/3Jtjo3hd
WDpxq0p7DeIVGGoO4AFF17/jkNFYJ5qQx21W11oezxZPdbIsQ2zen24QkdIbQ1W0GlvPvR46bsDP
p/I3Qa+3BM9HvTAHFTzBBPlDQK2tU/hRekJ9B++ZJjjFxlIkfqZpB0FwH2q2ScHt1NVn884m+dZZ
HqICx9jLOtQjon4AFLO3kdllW9VoZOI4zO9txf6np13ww+blW2f1QORhr5ChcQ//3Oeoby3HqW6/
UPXa46v1pw7zBOGoO1BTk7+N4nhDIoaGVrJfRACTy5Jeo88/t40t51SHLcLBDAwempJgRyuh93Eu
bdx98fBtmK187WaYeAScIHl+uALbFSEWJhByy2mKnh6TpBp5euwgxV1a7nQxGyPpar2B+sUH1doP
Q/9sL0yvqWqMfusgRJ8PKlSblcu6gNLheg1/qDSpwTg/AqAILgxT4IYVVpDjpElnpCkPUZfr7ZxC
VpySigsNijSGil0hDtHJHv6Qf9PRsE8CkItBiGnRIazXe20HCup1V0/lSusfLoIsZsHWe4noFVHx
PvjFpi1rufFu/3oddqifw9uud73yy/imYE6g8lx7Qw6qWqX+cmPSRO7RFtrcPdLwYOjJJbsiR9tQ
IGP1JabTT4NIMkTfEEP+YNSAC81p1zj0Hy7hT53VWWVxxQ6prW7CsYa9bxaus6ZvCLQrWvqlCveN
K2jqcNCqoe56tBjHCZonMA9tOFor1VZAt0STz9O9M+RQ4w5PBMoh4L+RQrhd2al6Yba3fhpnNx7G
exYYsTT9/pQy7uZs+cpqNacaeMTnnBS8NzpgUEMnR0mhg/9JuSw7x0a/ybmUsEr3fwWiiAtJcpVe
pR7PIrVMe+VasZK9LyE4IBJbDF887J7IhdZhFCdlwa2Uaw2/VoybV7/JwSq9xFvi5XH2vVEsAAiv
v/5VDMJRG2eMtvmWLwIEMZAyBdXT95FMqYzJD3Ioaj5wFZKd2yRGfEliRW3Q4IsywtWYp+lVlnTO
hSR+0YvsLPG5zt4IbN3l8kT2eMw/nOjcglOTAuxTJsHe2vxzvK+uN6g97VFsZ8NMvEsIVQGA07O4
Z6LD5PN66oCqUME4zibG6pSQ672HF1qgNYsQJX2xlIBcQKmbfeC+MCo76T9EpMPGYs0uj7NACck1
65XS9lPJ5zxzOAGw8WwEGIAAjxSR/m02nOcasN8hzM8M3m1XdCjclI8L0uPBQzNuaSmfU7tYIJK4
i12gGqXfnyPbyyA7YCYlSP+UFS6fGzXekCWPR0ctF8Uei00oSNPImkTouKr7Y3ZXnJ2oBgKwtL+W
11eEoMzvaYD6Ef0hjvT4oaBSs8eMt5dpEvQP+3oPHZQYdA5rhfGk41k605yPQ1GAok/m6c+vwRy0
pkMORHrK7ZGH9F64aI6qRjF6VJpYNqee3IvuaTBor7LE2tXQCUxCLgvrPpuQSjeyYC3NLB7oQHD2
duK17UYBJF8wUYmnEkHlvlsDUKRv0sfQ4fYxRi3ldRVU+R2+WuxsA8N1JUDRM0tmaTQSe8X7YtWu
FkL041jF5cp6086R6xF4GtpXDyf+fJe2P0LAsXBBV88eQXdaFvlJS3oMCwegKwyrE8dVqfbiH1cq
WM1O+aQQ58meuX5FtGtadux5vDjbyFolv7sCcFOyBTnML1DQa+NWnS1IoOH+H7XcuIQdcj3R7OCH
3/8qEADGSgbbXu0NShUcJI6KgaaDr1/H/m4Ql8Z2Shv4xWHSRSnUmpfUAXb8TRmhRW+KuuAs7KX4
rPBQpQOJSSIMIh0xUl4DgEAkgrs1BSPS1ZLRnvnQP374xVm6J9J9rxnx5RO6oymmfHtPuH5npEet
5e1dpldqOFxDJ8Ixw6iJZl3Mgg+2t13oxT9jZ2P++9ZGwM0vpZfg2SvVlzsxDcGQPgU2bJ/8Xnhc
fRrQIYWqGpawGHhF8+a22CC/cBgkwMbC7BWtX9BNAh+fUNWy+ZX6d820rSYUkbnw1q/vUqktVFrT
fyvDm7l5JlCUH8MLhJ30HRG85IG8+Co5xYFfAPzb9kahVyuPHrG5tHlk8Kg/9ztYpLAGSqLI2B/8
Xdoukpqer3TA+ugRLmO7wb1PYL71uDvf9IU329hqpvZqMBvJerc+6ExpYm1iU5ZG8G2Ld5t6lPIo
3ZCoT0Phv1NgMDkVDT1uNbGJWfF5bD3GSkT18w3CfTsBx04pDMPvtpvyEDY8u549owucik2akxJd
uVVEcD+yX0M95Pk48t31sh+E+JUeOZc/E6FKHQmyLZadxKCKw4aAHgimeZZnFCVpmu8z8lRWnW1V
Z78Vw4ierQ+OKknoa37xgiwQ26qVUwT8nquQhHeT8L46yYCOwbpH7LrlqfBwDoAdRcgo7D7vND9B
qPhc3b7GxGRHAimXVl769fjRS7P1PXggWlYuwfbVktyeD43kqienZPGv5Qhs5C2pkrYHVPON5PBe
2zWQ8hk9/PViDPutRrzGSkGIsWt/Eq5xhnPnN9iziX6/WndyTzjUo7QrJ9waA2sXDvglElbDvTMb
rHDBuwVQAMNeS3HN9ymPPLO6DQNhMlxXnBZVMeUuAELicLOzFJga7WuH7p6hlSjSjck7yjJGem78
/LvrHyo2wsebgpXV4WJyow706eRgkLutx+CxIYVSrcjLGRQCjsJyk6P45F26y99wNfX/kfJBcCAP
Pb+iIMF/huxSaRT3c/cP3DrrBWxXwt414Clpv8RxstXl/1fiMxs2TmGqfALR6NyK79SU0l9hP9vR
VI8TADUj0XzqL9Zi4CsgsPLhMUQI1VdX8uZJPLBqED8aaO3lle6ozFatNqqgusE+bOKomD1BbYj6
1rEt3HYfsQhh604B5A2AVdx/AxiM9a0VeG4iV2t5KrlKIwcKhOzvinPYaKMdE757JEyTkKoyW0cY
igI1fHt90qEIu+gDhMq3iZvnHQ4iOrkA7PTURc4A/vV5wFKs7YWomrI5RXcF40YnBZM5GJVgY0Lb
gDgqc0zB0vffHLvyzF4OJt1ZCaE4ALaMpFuhjJTND4uqK4j3Z4xIKoe2NrMIm63JkXePgTxyuakX
82wwoimj8/IN75rt0UUoCSocqj4GRyk2TfxIpmTnkqd2Rh7rq8VLzJA8685sxvov/gPRfTAqv4QY
haBxT3eSSXNEaySAwDl0jUQLFKO9lchWujiSGlmPgu+OZCAjAzQ4gFFd9rDbmsghMp6HGGaVvkAm
MBd0pxrcgfEOVzIjUuglxjaQSlDqVusP4uihx3QsDes9Bkx/yncEcc0JLWGL7gieiF2q+cTqJ15B
ey8EC2QVzPM+MyTZ3FUnpFKk7F7f0QrgKjNMms9967CVWkhzMbU4CVvZpLdOxPo8DR6aUbKqpy7J
eCrWE2L2p1GockHyRhZpyhep+XNpR1u1hZaK3iY/Bg6aHRrU004u3YKEriijvcrreP2Lc2kc7R08
PY3t957zxXG8yoxl1JVm8pVKkkLucEWC0Ggzu/AJ2CFrGDIIBwQNmX1EPTfTE+kw3sVvRoqOVtxZ
tQfSxy9WLO2IPPcZRQamgX6cjLOEgWxGNnKr2lUs3205HdxnuWBgYnnVYpFCBy8gWt7PSBhybw0f
7Cd28m6DMSAhKYz1N5UmqR94iNePfo2Kgq1ccKpArI74SbfbBbO0ngJ6T+LfBNxmyNEGZLf2zGoe
jKbYx/x5l2hlwcBhheK9mh7Vdbw6pHNVDK1QqTx+XdfdtAVfCxJ+Is8cE9TJpvN6ios08vDp1ldS
btAI3v5cdHhQJZi0ifhDxaqsrz2Hw7Ae9k0/lUjeoWNhks3PNsBJg9CAMLm3f/xreFeHi38pEGtz
8Qu9uNBTUCoMLlCiZLHAAE90T6GX/IWp7yhrf7I+LYgXQwzgugqqM4eESmbaZmqrWXKudSM8mpXa
CDq/tQzWynOgbyl/wMfwEZ9qUf60THNd4mFYjbi4hh4hZnip+wxEwM3OzWUC59GkFNdi85Z5z/Z/
i5cI8T+W60g/Dh01bKAOB6hG8+nJa/VsaOQbb3+0S+r1JNupapZq75nOA5DHl9aZrG/oZyCA3ume
3KHDYqkfIbQW3kVXe0V3OFktYKX0fzXX7lyFwXnEq5BjEExZjdvzOfLmy2pLIwduzNO3iAEGMTrH
LrN1SW+48VOHpl+56fySL13fhcedYHZL9P7nxvCBRy6xYpNE/3ybFRMbhJO9eADII8FmClR2UT3l
x8euIN2AGLY2rcVjPkWVDvw5zABphRZq/nZwyu/josns/ZnwHTrtds87yDwwOxreQn/ZC4jtp7zU
jQtdhXkbs601vSQiSNvan4IHhSzt0/WGxt1Lvd1HjHjQ4uK08QeZoG5Bs1qA/yiOJi9urH0aKijw
DKrjUqGrBNq2/YMHMDshXh2QjCCMrBtOGwvs+QaJAM2sQhuoaN78pua+1xdf2HplITI4aQi+PH5c
cyhMlxMqwYO34BYf39iS7Whh/Ek3yQsdBN+co6LygvYNjSAoGOT/5qz8jl3u2BKX8WgOOeL73En+
gfa56trrpKDRE+svAdAyNDNMrDlNdRJ9SBm4S/1NUIMi032Ue357mgjEUEer3LD6y2LWOMsMN1fv
ugCS9BT08DKRdqypMAa3qf31JOqCT0OcufZXDgSvCYYKVArQ2e/P837thTt7sZPQP4C3p4alO5Ot
/SZyevzjk0EfkxvZt6TCtzvI7Xr0YGdq01V9t3I6XmCH21Ulz/5YGI29PRW/AptJnm6hfXjWkpQJ
PIHaQ+f4p47qF5rMg5fPF0J1hDvZ8X1XSwNQn6sMZAiDN6+AtDXda4okllIPqqnj/PiOVgiU/cgq
U7DY0Q8j7NMxIIlridl7BXmUPqsqCUSk9f2pMGSkcLkhwOuxwXF5Bm6QUaTcqqBD4I/B4dht2N/j
Pu19i5o/HBqrOAHaUT+l7TX5QpX/TRIyOy4LCgyPOfJft1gn46y5PC1e3I3mJYmjsMmxM3w7Tqb0
p1NHQabDNrqBYQRU2x3P3m4q9vhgHWAeHMArNDbXwOLQvInFtN/YsXKyxIpKLAlpT9c3yJzP4kyQ
6Wj71p7LsT3hI217ZUYlgmkh32cb7PMRIPEtdfWL7bJ7XonsyMnhDZF0LO99P6wp1PzQjkbwpsff
NWX7Lj2sDO/YIh6OyxsXmF/6Kr7Zr7UtySttmGECmwv7L/YFwmFn35mW+t28PaAuAwjXy2I3Z3JC
XwhGu7LsycIGdZuqjRlW279hSE7lVTiuUZEcpEGzV9G3grROK3tGuTpXRZPx/cFRfA6+u2L/HhCL
7VHXgYLISKSOjU6cvp03zpuHvTDBIRPo9zdSDH1+h/CXK5dvWnRGfLmMmmk0YBIDySDQ1+nakBTF
4zRVUW7c8hR603rKmM33MD5DYhr+V8P0ZHsC4775gGYdwsDfHm9EruI4/yVh3Cy+z8bJW8a9io3R
Yjv3XCq5rHQZfmlf9V8J+zphjxxkJb++4kYCoOIInzlzEsRF5kElQlS9+l+9w3Hb3+jEGxfnyOyg
p45fHfnV39ycnwDqKwm4UfEBwzHwojEOE3Lde7vFs1jeblCB4WgW65m/2q7cicW7eCXo/dLs+03d
xvpv5YNVeUiLV+GZ/eXzf1ctLE4peNxzOU5AuPUucf6yqh+NfRrvzfbFo+3Ta813R2WaKdkMnkly
7suj9P3Gx55BMw/skhUYK+nGV24wLid4afyYxFOhxR+yc/hmitLJzqDlf1Y/JFIFQRuJwSf7A96y
/cn5aYu8QLqjvP4odvwe9K0PJ9X0qMS7BA5dwd2UdynVxVGx49LuufdSsl8Lh0Z3S9UBjfSA/2mh
SvUnLTHrf4XZufFBIYgVOFbCakrGQynEl2A5QwOvmvrxiH1T9iNKBLMg+qKO0rBGyX0k3Q76wx54
3V3wjvDouPUci9Z5LUkDCu0OqX0QpUWZ/5Wkb/xyn6mJXywBddqhXlmIYkbgGcmFtjMkgF4Wp7qM
klZBcf6F/e25Gbp+sbzV2hIRb2o2xb+ZdwG0HfRDJMqxGjGsXddKLbot9jdz2mkZXr2OK5p9XwJb
DeLR81GmnNINVLKdGDmGH/9lAqfzUIdGnp++uAAhburGAWxFHbKTnaC/oV6bzEeLgxwnuGuOzvsx
qAQU8OY61+8qhDieiJL8sLspJ7awLWRFfttCUg9JZuvR8HxnQoBRI0dtJU7JL46oP+DAYqETJ9F5
sDEGPW6NR6mqecMlRwp+Q6tE/DEleLe2xK/VH4qtIqCRVRqfMCAwm0IojxHDOJII7OGgK1273HLZ
Jr1P5kLOCLouBjv8f2VcN6m5Iq0HnItNAPc8SaeTAWKZz3PRvDirU/cv/xYpXlN7DcZhC6zwSrfb
uWqPcbz6v0XFTQYcQ8sIyICuuINxxQifjiVkV+Zw3kqwj9o4PFaMrx2h5KWo7Yvl62vlOCVMyDL/
AZkKjxMbN501FPkWV43WaQR8qdDLXOytFgBPhjvpQ3DV/O66+hFrX1qOx9JTtAJWC32LRkC47My0
hfZ4QC7wShuVN9HLSWhJEctBOjZwC+uKzSX0TIo58UFqt0axGWJsB5067+ru50BxcQsPPSg3QKCN
Iyqv81SssSc+9ZleIGCr5u28gYPskMtGxZPGyue1NV0X1unW5z+e/5yTwUZNI0QdL5WPbJeNmHW8
0HYSyl2Wvbytoj3cK2CoDgo3imRR7Qy2HybtpI16XshfEtqlA8ryoSPubxpFzqoabsOWpxHYVW2S
lCJZjvOFnkTQRpOW88wUhbJXHLEScEuJxmaGkjnSHB6NtRdttmEuu1jOi/10LykO+Gixpb+oxQ/n
3bbqCsjvG5dKeTPTAr0RN+bUW7ijr+eDlRJBRbF/Kb3QZTGpGN/HH7fOmJxexJXhnaQd/9A5ohdO
dvEVMGxG2WUcile8B58fV3xyrJ55LEjP6ToBhRrLAtasD0ErNOy7UutIe4rxnjMncTPgoxUvi0mu
AV+KNoeuZLSB95gWOTYhmrb3oP0fh5ab901TH0U0KPBKI5fh3aE4f62qRWhf7RWn0iwXGdHbNcBC
6WvCdsy8e0ggK5JEoZoCK9yYyHQwNHgVzRzL1BECHp/p8f694CO41hvWpEjsOC5Qz0uRa1gNBX8O
mfvKK0OaAX3Z2m+RCmPYFtAcOYYaMqVR0xcom9eYaNW4wZB8uUuE4dDLyDXYHtrylePWuvPsfWPJ
+YZNUwan79wMeaER+GxBk+yG21aetiv2Id7K6WGxhICHtOTwclizjcftk10dRNvC/07aXxF5ccrC
7CQHj93JY+kZa58+1lomMBQ4vpNI65U8NnPCrlPoN+pN/3ZaKtuKULZBa+NLqilahrW54oHv7ust
4lzU+4xTT8nN5Oei4qHHC6xmXaa3KR/4R7V4etJJC2l+ShZwVYOEFL6A11woxBTTAZgqWKyxh8vz
biW51ZnbqZBIswghVwgDqBzLL1oV9vrpkvYtzaXhUq/mxqv0VpTYNhTdcC4iLpLjX5zzqL7nk5Nq
Fwck/VCSAFuOEWCXTB44TYMxGYnR2H4RDCDu41qt0z6X4wlSYTwdrcRNY4Sbqxtnf3Qo8WZpxVSB
BjKMvn1y5PQlGBkFNGjdW4fAAjVw3yOfyviLbesgWkoBYjZp9QJEEdFErYLohKgf/RXEKc9KjfY7
2tNnOaZGJoZyETdAU13LRT8sXlpMtHU9AN/IgORXE3G4XU5YsaSrnqzFHELQvl2B19FXjTSifNzw
uVnornpRmSN4CTm2b0vYc41OcQtX9MM570yPhBRLJ4qol/1kxWti3FkNq3/yUNoVbqFgzFdF1+OJ
r7obK+PeHghbMTWyEChEk7CdV+oa87RnzKNyhe46XSz0dv3Pc3vLOD7n4swPW3nrk2+M129IarLB
B9PFsfe7lQnpdgFkttx3y1a6M/gvWqyvLJ9ONy43dfK5yJzliWmd0BXQ4wSEZrGllwcQ39mlAYBp
Z+C/YPzevrpiXldAbSB+EagZXF2tFC4XYDzXI/hB1+JmQfU+9px6Ykr0RQHdZyvbze6jvmufJf0P
nG0QIlUrsD2fhKD5jsVP3GIdv4jbOvTMAJjKoOUXHcN+/IUvEF2T4/jx/q6kyJQtSX6stqvaRarY
z3ttRawwIrQaIBvG9bQYXzgq4VE2v7HpKUsFTnJg9c9w6509yx8WUAmy4tsJLJnK/GrKZ824G9jf
cFcAKlZpQqwwISkYYO112KsYPCJ2OMMGK0IK9L5a1HaGcfR/K60c6cjCsqJSiBAtfdZFe/qKZF3x
Ch6wrIq4V96rJsIpCCi2/k34wy+CDI/DM0EAKyoZ1i3nMtujVZ6mFdsTSyUm6WLlY/jZxfbVcRR0
uNlCkBcup/uSn7x3JcF6VOL1eoRql5oVDZeVf4zCc4nYD9EltyoprK8lJdunYxuxZqr907U/hprc
d78Rws3jw3nNm/NFIwn3wBA21qspkMnTk+sGCdF+jyy+itfTYQrXkIj+FtQXqqCly2B1WP64g4j+
Q45kcFQrdHyzYIiWOKwutPLJSwLs0c7p6k9JE4DR1uZ29Qy7yT6btvrvkW4qd0aUoVjvbNrv1ei2
hnYCMa6CdFlFk49vMM5WiJnSbdWfgBx7Cdrrxs/szVlQSBnpirL/WCsp35NAbjUG8DvK2LLf0sQv
gEX9KGAxJt9zDC7T0PEfY1kHbJ7iA2/P5BiOR1uF/USymha9P4RtPDR+KjYUBIHvdPCYyE/ZqZC4
b6maFLII9vNUuMgJ6T0kVxUWceBw3mLDfP7Mb2F7uFCWFn8s7YUaSkTGmdbP3MiYw++/CecMeegv
tbs+10fRd5YG+dzgBgk4Qv5CBXO5KTCIJ9K4b9VQtA1s6TSIA0nvKvCfsdN2J8Ylmz3DJrOaAn7T
QtNr6vJJBpqzUKELiQIvQ+azQYKbJpbu1HaEPuui/iQXgVsmkrjx/eg/7xzNsZZZTKRIZ9y3b2IV
uFs1po7h6tEpURSuVee5PYd0DSj7qB9XE/BHXWzAyFHyImzhgn6koFpB1Jwlldt4OU/MKzNJsv30
nxsJ5RTLPIFyDDqFb97eUMZW/+DvCtGkbZySE9u9iH5oStbabW0e33OBv5jd+MyLRUFSd5YPgQSV
BFvh7ChXfxuFXHj6dwLhj39Z0xlmj7DLFxdl/3eUoyz3s7pbY9PgX3Q9d6dlZMLTEv9ZCaCRn3dJ
YQjPyrUfv4QzYAIDoncZJWnBJgIGEZpmV2AGaqPYPDG9lPsWdNaidXSplwiVKyL1kqZxI9L9a0pd
89FicRHPOhUsIIw4DM704MQZ8Nec3gbCNfh+pTovXC56myqHRv5KzSHofKRTzFo2glxcBvmsXouJ
DzdAIMkV/CtzwlqNfkjGjUyKKx204OFTd4aBrK41SQfcSj1TdcGla4h/Fl7RTKTbjhnuR6xrqXj5
VP93kftWdtM5L3IDdJHJngPmQ2UoqwSpj+k+CvWcxVrq4doJntDGcCKZ3gYBS6c8IswsjpMf7kAj
QEqnnFP99tUtfQl1yBVj74UuMfulcUKWvLSwcx0iOUsctawySnhsGBXOwQxH4mpXGlw4V91oHePB
3JJ9IEWnsSYlV3DGQQfp2ZjGSgdBXSLG1BOaYbFlB/j2iAs3k69ZD1prrYuri+te+kw2ltxDySrz
Ijk39acGXZBBS2pKgM8fUoAGIGQn+W7WvYIfgCxoryqtVovghnDp0PWy6RwTs9MSl4PftkXkxS3A
PPa/VcuXmMTT0uZoJx7PwCRW1Uq7FNG2mUjPvEza6sTTTYrj6/wZkeqY55rkQLobin+KDRR8bLpm
VYBnOuzkf7Z54a9ynzevTRYIqG9Y/C4piusY8uEPi3dbkAc+V963slpjCcvspz4xzfFVO1Ui/eKe
IFsqSrQysO9FkMh0Ivs8z2RxJ2OTwG3lrZswTW/0R7szeZpMOnlwqBMoR+MQ+fNYK7hw8XapzwoF
aYqq7ceJWEU7z4QkGEnRUVHsyvKxv/2DTZ8YBwETj/dvRyv2CHBrXZxDanbpa3GtP8JUSvpBAGuu
qeHTpqzRDB6XXr7HRLVFwcIsP6jzwwrszpSGe2h4M4gOpt5wb4DsmZKTuLZfNtyws64M8ixrYJB5
Fx+6wqHgC02mTeW5ZAZRoF2Z9hyL/A9/VdDFaF+7jbLvhA2asGbhQp2v58NOwyn6nUvw5vTvA7P5
j9lVmL4yzy9IIe5NXRb/yXcwanUOiVjY5/2u+KE9PuLgLa0hl7Osum0RsX9YImoeB78g1dkBY+qX
nVo14Q53XhXLIYdN2tEyrv4jyufX/hmfxswLvq4NbPLHD4wSUwjxpMj7i4k9sWNIy6T+n6K00f9P
xIZClBT2cyGPu6GKesE0tAWgnp4Ac5O0WFRME28/SXnRQzbS5sVDMfTSsANAF113k4fXJvmIhFmB
XPeNdAEkHEcr2jg/lwsmPDaZrDrPzeO7z8ogzg442DJQ9eNtZAcsS6j8EVuOrWfuz+zpuSJBm7M7
V36mX0O83dIhA8aCTKk33RR+CU8aA8FdqpVEsG4Cqnb5Tx1gxMQPTWVcoO9650bWJ0IjtHi4i/es
CnElGwhn1KeEleh6j9au0hWkROoH28xF78YIt9Vdt9GlePfGz98O5oW2VJggw5kuDj8/gJyLpK4g
QH1pQefincWWyMrOMzzYX0caVxkJLsi1GBYKt6hmePE7M9b2flMVf/8YzvmJ6Qj/a+u/9s5y1ifW
x2I76Av+F3I1xt6IgTxDRjHP3hHcAkszS4IISKC60NEonlJERdq9lPtEZIMBF4P9SiJjKFYJTEAK
zWhtraM233v/dsYUWHcL9+/TG6VQX1cCw4q4Cm9B+0jXhxqrtcYKP+Mw3IPnVDUxK0GXrXCPgNFx
FOiirGj2CiA42JSUixTMNUNqVRuEjWXJ1Be2n0Lr/YGSDbBPly+KjVek26cv+VpdIPawxm4OsGLE
+9RszAJYpBSYSptpyIX0h8niOU5rDwX9+x3ne3NErXZ5IP3Lj2t9M2N1MMfpt7yzFXN29+xrvobc
I69CAaNXqTp/+qyYrxvh4VnO7ksMyIGlThxZoz0uOlyQifZTpRkdRFT2qQlu9aGVHPXoA3jTft7v
GxHAxVPej+sxBeF4XhjrlAZY5Zaguim/rKRtIGPgMJpb1epxM3uXXBM5I9M2lCHv/hSiHww4dOG7
wOd9Q4bRlTJn8ruZ/xn54pMjSYX76qbRPJ5VlfrsPPkUJUbON4FPSGmyKL29z16YDcqRIInK41ax
XvqXkZX1+Uw9yTG9MHexfKyKlSAgZilAy9umg/OdD7jNfEUvkn441EsDG2ageGqQ/YqheMzZt0NN
EgMQ8sCbKkN9KffeCHwscmCiYfFPfY46BFVlxmqCtYc8OPmW5v4mSRmdixFmCOdHCSX6gWTFdKR+
BOx78p45vHCEfKkV44OOTlW360t8GdFzzrhn40OiKbZsPjjtipp+LMEDj8x6KExJnWji2+yXhiYs
JxfdFefTKMcxMwsSOiqLegjlSu0mpz6O5nONBj2mAQhXnWpTbOvgvi6D4i2NXRGDJv0v2yliHhik
5VPBIWTQ+r6swKZTh/4ZPzZVRwRC27UWcEMW+A+mGhYRSVt75eWrlIgDhGxqvltjg0asfHu0gXH0
C9DldNQGHTeDf4zx38PvjbLmdHn+BM+HJcBXRuGwZE8F5Ru0OpYZkfOmSLWARuw+6ByIwgPbiC7C
szx2DRCfoalqeTx4Zg+bFdE7wUPk5g7gokF32Fn/xHpMh8vXEIYmfVfFrv6latnind+Gc7dn0ZQV
PGM8HEYGlvbRcaZzJZbXZMTONqFYb64N62mhKvykUtJ4E74WEIhF7q7oepKJa7eBu6ElGsat11Om
OwP/GKPgjNhSPmDRLTR1jdNki8JMfVt4c0L8LfKv0PNn1mZYd1mYmj2LZAOmz/4lJum/41B0ra33
ipbaXEggy8GKPvfOS6tar6Y3LL4LkOkyBjhqadBR+0nywX0OrEKOyjf/pBwLJxMIvcppyYLbvExb
sv6BmUZ0g9qeD3h+RUoqj41eFnCcKIjdw1WsLbFca3SYA2gxPRNwWTAFHbhJ5lXmhSw9CUu1oret
VLo3qU4v4dZmIc6kqblkDEokdfY4Pz38fwChXXgVgbpIDL/1D3Oyn54EtkxX8AyFsnpIy///9kQX
jbM2UlN1lvASWN33JKlQJJQARmO9jZUtC6c4NN0GTSwUhBNpZ4vB1PrKRZnvCbamxWGc51SHSAt1
Y4tPQbL1uz5hrPn/dEAOMnxu80GQmBCN6ItHerBWJ/oHgEMh4nw+vtPRYhB13WOHyF2TRoSekDGe
azdMWcLjlDkno1nXgIB2rBZFaXXU9rMqutjejVNPOdOGFHA3hnOOVOI3keawQROP+bl/pL5JZ5OH
Nw9tlzPFEqG8wDYza+Kqmkp5Gg/zoKVzIl6gwkDIPjowtxN4qNw6KYb+pChmpAcBQ+7o199pGAh2
tx7TUlxOtcvmhgEDtbA0ax9HhzshZdyFd+sCDYOyDfyzecKLUJJ7XJ80kLJaOaXCAcxmS28dmsc2
foObO2EAKB7ZF7hzrru2WSfgY1m/nm94wyX1NF1VcVpP7OF+rSBzMjxEN/M086cvodbf9A5xiskY
Te+ulA5746huvK0O0QRvw3tvwB88XGMUEu3PnoqS/1GmBT/hpuffe18rpvoCvV7T3NspVuiGxE/C
74/ozRqjZf/yn7FcGLjFLc4Vqa4wOr2x1IbqnHoHknONPvQjwGZ5lUT+t9YnjKRfrZP73CPlk+cV
VTiSiEzdus6VN02ZpsI3PFbh2qeL3JXcDM1/8sTrcQwZ+RNhkylYw/cI7y2OOq8sa6l6rKWOSEfL
T1N73eTvUc7zAQ6OyXnHoimJoXMNIaNQMMelJ/g2OelecGNnGh/b+tFCdbVUvUt3rqKURX3ynZOT
Fb+JddThKfnWBQ9b/UswlgzGNRTqfu9cImwkbElQi48U+mLtgj6JPSORea47R1nW/0yGqkTL2WsB
Luwx9Wfvuv9zv/s/8mxk7fZt5P7BXstiMrEa05GlAyebqPKPX22po16rMOBnbkJ3Feb4t+NVnL/N
BeBrD5vH+Rv6rgxMIV6/8gS76P8heYxEZS6MpJ1BboIFCubaBN6v+2sv9XxnGfKZtIVcR9GYTvwK
ZwhFOesOynQj0GwhAPPKCBKhlM8yjNXuvie7x8NTZHFrKfTSMbOIOn3jLVEiJwDx1Doka1fIWi7F
DcTkEi9sAv85qwnxVPXNCZwiZYPod45UE9x5zjebyYLIASw88dhLU2epUcYoQ8kLSZUc0cxpVKcZ
HapjC8C3fR+HnSMK+SvYkGEXotCnOd2L4JfzETIQOaUOknLKLfaoMJPgnwa6BSZmpSqwDPfR1Uek
/KFJr8KxRu6Q2D6kBsNjGzCx1WbtABoUth2lc/LD0qfy9gBNYISnhHK0CCiwlxlTVaKUiScALX48
SvdX3NM8/pw5Ogy1+HpNbywnEl0x9piYl8uEWC+oGwpwD2iqn8L/RdJH7uGifo6yjsNXqHpPTJRi
vRHUNik3JGR9aySuNi41egHn3E9i+nxwZxAIdKd9UXFIEBBCydONO4H1aKtn0IBAjNllJ7rO+wrD
xJPTeS6v2z7eQnmDYygEOtBipohr8Xq4O46/uSbxpxxqAYOPIOFVbCkJAeBnE1Qpf+ymdTUbcTfC
UAT0uf7CwYrbLsDR3WDE2nflc7PzNKumRfXazKNsCpfnhB0QTMddvEt96rMFa63l+I3r6pOrZYh/
vpb1oumZNHYYNxHGCS6KXfPVWezLMeTdERuf+dTa9nP1EsPvRxHOjd1vjSex7KnLoQjST34Nvk5N
l80vZopKrH3AfVIj+X7x1y1qRQ/i9nX4VL+CsS1/Yj/MiazL3IF6VrDR6c1hbAfDZ0xllAzcmV9K
qNGNoPAQFngr6YaTWp7pawyC8cyF+tDfirEwkVkO5jgPD3vqiupDJFDSt58TeuMOi/yL0n0JtRkC
doItrOcmMfl3ufvSDpU7Uum50yLreNfRj8CMo9hUSqs3yh/m8a8SSEiL+/jt2bhAbW5FvFE2qpgp
Xi+qTZC8C/bo9x7jz5FjgzRaylhsJHMkUcVO13lITzFjgFWEkUb3nwx2HI4DaBV5MbSIFWvG9K9z
KTETVZLWufir85vV1sWwXrdRFZE0FAd5Ghx65M+8DnJVpCsL9vR/KXjaAdmR7j9dg2Ihhj23zjjT
vdspz7BaoVROxa6qtn8c1NWHRc0jRqTZChqiF1citCH+CdcTnMzUzmXTpnmx8uf1WBUdDuiWo4Vk
zKa8sPZR3PUSwMMD/JOrHIlNk84UNVZ/aS0vkj7wA1y+eIORSJz5JkI7eh0Od4qPmW1c0oF03GLc
IJGlhLCoN2nLmnk7Hpo0foI7n1901ctwya1xtGb3faC97Iw5pRZSt80OLN3PChdS++ENd3lnMQzk
2dHjS7RO/v2fgQW03q02Q0XvG4HrLsi7+DTx34qaRxdP2A8IJnN5G2aasUvC22HYf1lz5VnbJC4G
pQXne9/jTBWahJ8F7d1fgs2rveSIeQ8Eer8Cii4vXMwqfj45eIHXwbenmpGAmyzWGLozM/hAtRMU
206yxGI6GGci6YPGfdWCM2G+eTBa8wNLR1ZG3nmZPJv8E0/ZRQgQxJVCBpnZ//7sA/csRu9V9z62
w2f6dSjNfn0I3zh1vDsox70s2mUYcMkHJ8rhJYQ8pcJi5rf9Tmaea88Anml7aBxvpwYtkMQLeGRk
v0gXaxMjXVLmKvKUAvQ0s3zqJbpT9UCQFVMUs9WiEPZP24nkqkYkvRH5FkDK17aCN60Y6/PStJaq
NjNKuRzf1jN0yXAKCstII/VbRgHpsQhHSq/NorQmI2Q7i0/5Dmb74d4DH60T+k+aCV2sTGbAfnKr
5+NR+0D1+9QKovcv4fWdyfetJN4eiQ2poylhENjlNidAI1xNpdczPvlJJtFQDJf+XSiTJ1Ug0zLC
en/oYABr7h/jSHHPEXjV9BZ4Je5QDEDb7uTrJFgL22Fgj7YX3TkJJ7S0xKgPXH9p0HjxTRkGeuLu
frQk0AZQgFYz0l1u+ymr8GFz9okLQwQ7M7kaghhpqtBgeRQ3pdPcu4pmDR2rn+U0uxrWHqq5nX7y
IB6nFke3k1mU1PfwIyVtEuG3acCorkWEd8wPpfgVx4+osgfqQAG5Vo05XH/HMhONQHk/aAcaAJ2k
CdKKPqBjVHEa82om4ATQgnSuBmdJGcnzPIXgVMvGivBltwQNL627dSColVfiIqLwgF6XBik4vAZ3
sY6+eR8DnTi095sL27nEVYEZJHRoEzF3RmFMkEJxAJbfcoyrunlGsho88olW/binw6zWuDNIw8WX
4Jc7mCP/xSgGp82dUCPHlTQwXg8N+376zyWP4sBrH27LwYVAqGirpwekl9qaQeZQWThi5aVzDIXn
L/skB0YN73T48q0K5nujl1zAHyBjarRnOzzZCrKdsLnjKsYyOtHkvgj+ymdIZAU9fWDcoOwaZETb
CDiaHIWXgrpMGjxTRLqaigvDY0VYh05W/JIpATHoLkJT9w7tR/LbohFI37lxzBEC5aJqorPabBEL
Y1iGeGRPxKMB/VMHSYLzQDCJ7VWAH5lgfGGOBt8CIM/Smq6xA1aT4jLydTdh59CrvpjnjpYYm2+L
DdMWPJSlHtMquHt8XtTRirl2IMitikYxnJJrAqqilnzJRNA/+9JKdiN8mfOwt8O3FNCX4lsz4R/4
12LqXNzx0Ez1rIFh5gofW/VMbnsOqKxvzeE/wcnrtPQZoevLJsnCpNhyZiBW7p9Uz2Z6yucaUf6p
/O8kxGRQJrJRqDE6Fsm2nzIkUSLsk8HTeDllmWmYrjG+QPjGYOXo0ydbggh8XJHtHYD4IR2px6pe
aotNYZTdQiLmGw8N4pQc+fRCZNUSq1XnrTHMIrNKc/E02cYJpQiScVIu87El6vtgUGySEYKxLWUW
DrgzaEuQaL7Km4BEeCzKzytIqLYzUAYSxzWWuENGiurLhEHrwXd5IxTIxDeThTXqutCkTBYSY43W
ruR5yVmpo152tGF8O+sTzoiufORRD9u/varUAmj7JxB3CcBEnd4NxDv1QI95wWDqp5NtX28sw/O8
V4RjfG/BTdYIyA+nMOZTVM7InV0/qfp8RxYLhZVaFh4pkdcSoGlmeJKbEHbUmlVE4CJbOsCPnn6C
3aDDAdNnwMMpg/1XlD5YNe7Qoz6NtQ+49OOosB4p/iZjJ9eW3khKVEaPCAFy/kAhnMyBo1+44+mL
08cj91HIsFDMEHSU1qFgvYYvMRZN7ljrF3nbQc/gLJJOwL/kM8FbI35ms0IABnTWSqUFHUZ1QIpb
1X1kclspWgTrb6ungFQ1A/VM0HUHDnk4BPxRT6CGVW05xAkFq9fozQ0+bOCK1jg4zouWUZ6gUGlh
kt9ILSUoV6zI5cauAZz4LHOHrKrC/FM5gqZtwBCxkiI6F/4QRCzNHduZE2JHcJ4X8VlbILrlXs1s
c+ytb5rtbLWZkhlZXq4Aa2sq5DgVPT92eCaQqz9peT1y3u39yAp90ZcqbcvuKT09ICRlZKJVv09g
P6SmzNbQckjRLSENjWIm4GRR/n3SxgbEuxzGp5im8IXlK7bd+1LEDlrQfW/+Ues6Ttd0CXl7/p+5
2laQ5wJ8K4jreehlktFuwKZuZrm57HypMsfYxN0MpKACUf1k1LKpmqf0VL0weUQF89l1T0EyPT0o
rwz39jf0pbrjtMxRKbM1zwsTsAmlvTLuuH8xkn2Rc9vSwhT1FuhSqlj22vdPYRAiV/DrhJIInqTO
q+i2MVUvbd2ygXPXGE05zwPKfbT4IW0kPPjztmWTfM6yb+uRGTXu3ZzcBGSOZl77nbtmFcEPWD91
w7d2l8Qg1WbavnQsMr5k0MiJNzCIJZKfM4SIAqUkcvfQstXbQGTVkT49oEub6WQ8MzYBjQbJgQqX
ztCVWTsHzGA7J9/RKmwG3tU2V+kymVI6pju1xAizvER+EHsiGdGYxNxi2s5TOa1u5OnS+LgMRd+t
k1RguEe0ZEcJrah5VixwBLGZTyFtvzDZWZ0pay4KEO6ntUli2H31OcGA9BANNna0vVCanSpMgn6G
uyGkq1MlQIAe5E01pPSBLv+IyT3ttGl7f12rFQrTKgoPQ+qRKTWJTZiVTjD1lOLfCnyHmavfgMwI
0pdmLG3nj4IDGF+icubzzLq7cbXGDu5oOKn2awPtDtpjhhwPxZkv8m4WvF7SLp972dJcJ13jozrv
y7ZE46qGixZWUV7IZMlzAIdqUkr2kz9FRp1rVJBxjzp+qslyymAxxdeUGDqMxivGiACPl/nnMjoV
NpSHzQYj0mvbXYo0Ji5lb3jlVuDf7Oku+rxD9QFrHm+iX4+CLBIpkR0fx2pPB7R005pmLydQPonT
OF6hz9SkaSPcLrTwRgEEedxIm7XXSvexVUf6aGpcJLydQ/Yusj7mrh5b2HiXhV83+sLPEkKMvrQS
5Uh64oJtqAXMIT5NijTbwr6jR6Hf8bMCb4pBPV0hAm43pU3lUG0e956A+Hs4mc6W9tzJlsudDw+o
i8W4cFP5zjSICPHgrcNOAgV3i1COsoJsVoPQ+6xdwU88hOtyB77CYEShmwKBjsNfhQMhpMro82Ki
DsX9twB8rO3EsPkgRJHF36YTtwIFCsYMNJMQxtLca69uOAJ5ZVvuY4s2WMkdToo7poy/vsE9779O
cFrfJIBT6KIvqHjHdivM7uINmXmNlZ9BRiVF1HN2bNfMnXygcmNgnCf9vHLe/FbXiv9RXDaJjF5v
/G0ctxOOeCpkqrOuNxWfK6PYTY8Rz32bEo7EQJZyazc5idfL7mNZ1AquWOQXDAQ2zCk2QF62zYA9
aP4+gKIvowS27O9b+ziPddvzt6LwfBjpZFWEQrdJARQ88WGaDcYQLC8ixLBa35EQR0IFwBBFFkeZ
EAW3Cx5042/UxxKEJvYdSlzYwreINI0OOePEAnc+7fUKBuoa2afDlnGEmFiIEMBA9SNG3S7GDb4C
5nQd+mjyPtlM/tfWPPQLu+ddhDKXLexIJ7veFgD3UU/EH3QO7F0aKkk/NO3OSjcL6sEFAh/WhnsZ
85EXy+R0j8BaiOGrNkPk1x6QYcUmnSMm27jwyTytA+ASKj7IF+Xf4jssJr9gFNsC5Gnq/ADDW9Z+
VWjfucdhfGdYYlX2mx3Pq3/bqZtpzXELrsIa7yKkSbee5P0VJ+0y97m20wC26KmVvxXZc4L/B/u1
W6Kz3X9PRvX28xb2zHlEsnzpNugJGDbSHfIO/jlqKrwbRDyWkigfEUq5pbea4FEdkugA2esFF4RJ
MZ/BeMhYY/QodDsuSVTE9Yk4uF88oqnTeaNsM3xfXMebL/pG3XXC+2Wfsz1WFSa3L8nFELmVH1za
EBofR9Z7Fj+KoPOpjbRuFJ5Tb1stOH1VAnXCy2/o/QUcEAtZv9AJ+Z7irb++Hc7qUaqDbJIbPnBj
2VifJT7ClAhPVIeo/jzOmj6HI0HwUmOstyCR9D/v9DrHFribEkhwntYnj8Jch47zMGG81ygWhsPk
fOLGXR8ufuvt0cHchWMYE8oDmVhHY1J5rzaoZQYTz5otw3zGBjWxfB9HVRv0tMWV3l0qoNmTgu0j
NSrlSjKOR2nIYgpankV8cAWIHadGY/dOkt/wa9Fca0sB3mftuRMOlJTcFD0Y9K35QXHDvwLBPZBV
W0da+y8NiT+vRGfJ2Ciu3khgjt2qCtsdjuHS8ZX6IZwdntVUDZlElbd/4sDbsP2/lHW0ka8cIvfu
gK45CE7i6zTsRg7HfAx3XfKtt+lGobw2CXRrEI0yoGm863d2T8U8zhWRImXahFDr0QmGyFMKvaxs
oC6RykmsDGU+Cw3VGwpy1l8dn63QHUjlZXJONpVfEaxGyan3C5tdHPtGR/ck2OhPJXS2GAsG2amV
XSQXkgPKvJwPO2k3vPMDGnrcNGOp0rFZKK2U3Oe+qOLi0Z3FghD1Q77rAtYOj/16akYj0zAuDcaJ
2VC/fFapNmCVDLrEXnSgfNb7BwFmpneMPAIPlUBds4Q/dGYO9GdK/vwZXvsedROHjrMqNZIX9nkM
YKlogy+Y/MHAodO43t6ANZnxcBHmyC+bhTVDT+T79O1XQBLlxAjVnHx3ku4/7MApPbgr2JDQNGSR
Xb/o1G/S3aZHPThzjnYTDKLaJVKE9jgk+MLOGIumdj0qJgQxG5nHcSQyrTrrUDulYpHoRTq0GHbU
dvx/+Kdsw7Rbf9LThM6jz0Nwe3rf7TPNDvwEQndqxKttYdkT3P94OAJCTBeZSZ0kItFZcxcvXDqz
qKtKEtb10etTzRsEqT+FZirXcfUoPBIcYyKmBpAb7khpLZfh3wGlCHm879/JXSuJcAC1HVsfUV/C
17CiHfkBPBzU/xg3alwiHeqd+P3F4znxxvX1qHNeqhZH2iZIfYZltdloMavTIeLj0ibB1ZzxqW+K
/0xx7XheFMPEWTR9+HvKbcZ+61YQOEOMyQrh7WHzPRBRTxwIbeWVXQvDqLSk9elRMifssZ1UUeO0
bXzs2v6FABWcGv7HBlfc9FGWA7duLqBAz8bcWlFstJelBKi68mmUcArb3ipWpwosNHCtyyiCNiUt
seOGvfOZ5IV9OZQF/7A76ZJDVsvMz76Cu2ZZMaz6ttjluh05JQU+87Y/C+Hv1u75LoWoXaHMCl+P
YZG0Y8fB1u8waJwibimOQXGS/vWbrwZnxZeLXhdFLaVlomASUN/ON0+sMcNE+kb4e7VcIVlANSkN
893skBLkQkY8jR5JDPr7AX5D64dK0UWS8P44SYMLoAWaseQ3aV6p3o8Fpoqu4Q3+QdCuIwngC4Of
Bgj+4cWRoD5sKwTmeP/iWYh37qM+WrE3KUua9jrA+41CrDmYRFBIs225uL31FtZ8jxRX585wXXep
4mMSBBHh7ggs9IjW+Cx003WJtftpUKnbzx/urW7+eR4T1VqbmMk6EBi1GS86V9RG+gqdPipKkFnN
eBcnHJoUk+jZAptbpxR9rzbBCSH+bjoOhcmtVMFhWGf63ZfT1oCbu31TNOmIYqftxQhX2Dp8k49z
Ygk1gqOLWl9wpOBGuVyI1dt2pPNKiBi14zA7nMXJFEEdPApHFV6Rtzt2BpchDN3KHZLG+eu3bOKn
0iyp+ygnrqfSp0BmxorvYfvAgsX+i1s6aCdPadYtxjlU3IB2PlTyGAZ/7f7Gyls4s2qrpSNw43Kc
aOKVFdshPMBMbH5/zHQ9WROin1QIRtH5iYPDdQbJzseG+hAqhXgkp3T8T3EbLWLxkQ8nkGzYdH0l
GgyKMq9nBLDv2yyuoBr+hSI/1JxWnZ2Vl/G2F9jeWsw7p0b8xvJXcOdIz23t5+/fVju9snWJnUH8
RIdQYKfegc2KEToA/ILMPPQnA3dOqA6g4El/EUnXqk3sOtPLljrbpaN0mBDzdP+j6JjgEBsoBeQD
hoVn6pBtaYnxVLNz8jAFEvQbwhQYLBa7N/BRMWrpq5jpb4Di5c6XooFLtLHJUTnG9E77/UOhkgyn
TSgcrG3n1odkOjT7aTcJQ3JEnJwhv/vnsLED1fYRG+liKdyvtqYpLs2c/ZuENiMTQcDWU0AbAO0o
LbGbbW4FdZNniT6gjbOkJSJVpdgZLQAPtYCgTnT/rJ57j2j6ILAPQcrVpfC0S9h3pcQpGKa9YukQ
Wt4AToANX1r66CyCMZKUXthBkYLSQC6zKeFl+KJr9XomK9QajXl0GMf01aMFeqSrna71wZBhhOPG
GXixdsMBlYANo9TlMut58ku6nVbNPQxB7aaSNOY+K04JxUHawUwUNqlzTTw7XUGpKKh68XD6JaVL
7q3m+xCza6OScJtR8id8rSiTk99rtYEE8j+Vic0ilXNZpBD4SWQmx7IxROtssQZhxM7hmGQiZveV
tEGESm0z3arWcTste6H73zksGURRBblAxyIWQVpzkFepmFhgn82Bix+u3Lg3mW6AkrcaqgMOsULL
Ohm3uKvOArpvk9OObgcRkn8FqBryom0Vyq7tcOJ9e/5OnJ0V0Z03E3Y7iDgPYWPpapOHLh2GgQS6
tdLhkAv+uMjgX4ppc0fm6fIlBkNRli3GpONCmCUa6MsYTKHakNU1yubureB8oJsbLyTT5dV132s1
mW8VsF4ddOHZMSnw304bE3LPnLbzDyFakKXcyXrlgtQ4knug0jaioqni2b5scXetTu8qVhwQFncG
zQ16DG+9oiKl0ll6EwdkqbN2NglYE1kQVVYzAqxmO3cUExydVocsfu0gViGG2DmTfL4pHx3Q/41E
9b6N9m7ZUBXwjBouNlqPERNDB4QmTf4pRGDTfAXSfBPFqVwKJ34v3MqDfB5/VY9pg3NZV0mlnJB9
KU4x4aMdiNrmUH7CW/N2uSM0nP/Agr5XRj0bGO5b5wIIxzLtmNGgyL6ptq/OifUM4I9o+BYvBcMh
Qag4Vu1dS+eySs0XJjsXNPKSkSdzmg4j7adzLq4hQMhPnyXE0OZSXhiMaF69AWJXnLAUfS5AWLy2
xFuiyM82nLmRckwTJsceTqHFUnBuM7v3EOd1kuxEAFpbkZHbLZDYk0tgeSv3HmkQr31g59jvF3wc
H3hEkWXbNtCI6VEMxuyNNiDIGAaEZzmgeXhzTrCLSp72YhWndbHI2CJ3PhC7ORL1LFDNCZqZJJzr
d30rVLZN9clzk1/+nx3hdF0MSaUSl3AUGc2XB/Xkl1PlORo+6/tdQATMpPk3NknL7IX1wrUcnKdm
kqEnrAHZTuxgbUTg3zUR4xtlyOfGDxZ+urTy+XkyS4miRRK6dyT6wwTRod0tD3FODOIMiG6mptAx
Me9zBED2Y87KOUcZmeBE9pKhAww3phSSclZD3kjnn9AGq0I5++NcVxjPO00Dz445ovG83SHmgwEF
nWAXqzxRg58vY5jBtSrBcU75h8NVuLBL147F2K0CYR2k0cIfGWPQjldEXtd46d1cOf4CrPXlX4YB
txWkMpW4q2UMPDBqk1z5LvZC5lhEnloPL1s3ZZ7k+7X5zeRaGzqUMLyoetgw8ShyLlRKo4TarqCD
oUF3D4AIkSjnsJSrTpzn2D4yCuaDnH1zG2l9CWcPISTIbZS++JVpKybAljg5zRV7sJi2q50qhrek
PuVo+yxqwcWbSII67YyiMIA/24F6CP8/b2mO6pgummM9UjkLhVWnIXcgg56CBtDQj00grudXWT9d
jrhrSAZkg0sMW1uT8RCgEGukQmu2xbFGGKEubvZb64iVuu5r3TPJh9LxYyvyIp2HU9yxQG+3FmNx
mfuhzp33f6gp6fPN4Axka1mchRbQ4WzcUgHvoIypimPPrmY1JE/KCwHx8qjo/u23saWRjv0j62yg
xY/M8vCQDYD13x6KB6mxXavhB11viB+3mcfVVYtJGJn3jixpVOqMQ7dkhKh6nYbfA7m1TX72jYAE
t3Pb8tGDFOtW4Q3EvI0XM+Y2aMfNqzcoCDHoWBaS3dD695iAPmd/Hz6WJpwl35GdmRWbYLuwisgx
//Oob6H1qetaXbUi+amrBs6SbdgMUjQqNHEkJeElcad6KpiYkc3mdZ2N4V0rKyiJbI0DOk409MPB
Crziuf/5f5tZKPTIUJsEXR6LxzDZtnWwfx/LPBKl/KFVJUimlEQZ7DvoDMsRCEYVfQcKOSQhmv4j
eVi1DxfRl7rwrsHwkAWxgMIEPR/FMOxOSkSDvWGHQRocCEjNLGoPVE0kdoKcR099WBz946icZAjY
inmmumaFNkJxR9X0T2Ai1V4u4P3Rki4IaNLYWGHy7ONP9cyBf7K5lEr4qIdzDehhlDIDcorurhu5
GHFuus+PkzEwnts9ww8DEXSwF3kkMx6YxhMN5DGKzbF0pUjO/nx3N+QuTDHkAKObr0I+kbtxMxDL
e9wvjVuNsRjBJFfjTwL2CaOKvUOP+oyr1wh28Q6jl/Tc4CU74QPj0uu7JJX6RdFPM6Ru1T0+N9vV
/JQDiYNK7coHVxx9/5XhJXixqGgjHvlBAts4Y9qWVUo0qsiSiBa1VRgeopJWEPb2E/XW34vyF4kk
lfXeJOY1cY9nIIuIGetaZqjOxnVEIc6kpDSweqln/AQyWfZOvnpb9jWfIGUwvbQQ6DQnAaj4WWQ5
a7a118fP5uhE7cTNnT4l9HdYBEH9cv+cDiMtgUQjZG3HzbluEWhapoPqiX4LcSisLE6p03N/cg7T
ZbzwqmoZUcm8WmZOvGMlK1bjircL+bDQRkWMpdU6MuRaY7HzK20VA0USpKYbzWownDw0xN4TPeUs
jfM1b0qPDx7IY6UIet3G/qjldi9lUODMLtlXJ3UuG9jdY0A3TX7mCra7r7eUIeHYxV/0TlTpbh7U
aZ1HPgAN7nyudQnbablnFCFlP8m6LSUuqwnpu1DabqA0gTLjiyYUmVLKdydlAE4LJyvna2YSRTRd
B+M6lGUJ97xFGY2ONwUqhr9co9sC0XMLHj92zcM+gX3C5EZRTFppF7OLGyzzEIIjaoFZMGRyK/De
8wpDmMLAgMbBQbsPQj377R2VoWJK0eVR5jxC+2DPd+icj9lKJDOVqLzsP48A+Tp378oa0mXEgsuu
4Vdc2DJ/1FBByxa2KSwhS0UWSgvskiD1k/7T97+vlk7OoLwhXgXtjj+77NeI/niI8Qz4v0eIFfa6
6UzCZjZtm6RU5sHjWi6p7fGmbiN2rleCW7YCO4LagZcoa7B1IKW2dU7Lk+jiO+SYY8RV3EKyL8Bi
Ss1UtkB7hccvr9EJtwGZeDfSxAM28uZsmZMHZvxkl+Hu46017C3SRhw2PnvQ/yC4bmPgA8Kp+Fd6
ehSMuCzK8+sLzABSidpfNG8lQJCR7LnMoPCs7ShVFX+Zy5attpdjsz5rbUkeVJYu9d8QBtt17IGY
xzhtFUI3/A9gP3BZ/nuzAC/FVIAsYCvHcvMONH4rZiYxV4qmjdX0nCgXrul/kbIsRNrxH7U3zR8i
la9UFGTiq03SZrk7dO0yA4MspyYOuS2o4YvpUA3M+clAsvAlRiHS7CvNooXBhDzFGjSd6i9USNgu
UF2iVNEAf4aliQs89mNNosRQ41eFQsYQeJm2NRnmegWRpHKGy3AkXGknAsIOUvJt0F/s3oDSAVbi
kfrZF/koXbUppKeNg4OuuzCwhYPQboCYg6tRnScH93w45n1s7E1KqcQXXj9G5AOC3e81FkIsy9QU
1Bkv8rZ6q14h6e+7b2YNwPEHWbOXG5V7boMAxLczEloLHUL6206D+gjFdIgDCZuQrgre+cL9TSGS
AX+p8Pw6giwWwLiiqoJs8SM2Kp65MYOZDi9JkOV+FvRS1odKXAe4BiL9HynOfnHQBmFRrlOoapMg
d4X1VSuysVcL1wlmFPBrd/r0gjyfmQajv3g4bI7Ip2fvlSXLy5YBrPrTwX0fOz0KeDy/qeJLFNZG
g8Blu7TostPvHTo75RIjArTeIm4IZ1FI5J7WkCjaszZDnokOD6/fM/Ec7YhRRY3aBsUPeFVnoTFo
zGjYKzhgpV1FJFzDWmzziWpHO6Bb8jormi+ztL7T4CcXLh7ug0jcu/pUi7r39pB6tb12zmSpOKew
EiFXWnsq/G83oiAo6TFV5h2D39LUoavZ6vmxxMyufhZZ/x+z5nKFmlwQKQRvfDYS8KW3wN+eKqYZ
yhrxTgD6YiJ5mYztz7ZIy8jlKHIQ2KoLFhOhCDNrADYI3DdqrWhlP/zAUG9p3R7DSPiHj212EgAF
JYIu7PhcMj6fzixicAEoz4Y0QqDgzgjmzrkxPXQZTauLxt1EcsE95MeerBgqfNlKruIRu1rrpJvo
oIskCiYlhSc0LgGLBJW0cZmZ4fS1emkEplWF3IpBJfbPJ7m7XN69JFjgCbdzt3nOnHYjm4n7kOZ2
PG37WUSNK3Jn8n5mG3bKBog6SNg3vLg8t5D7hH5mIxZ9nG3+nO1Zb9UiFpO163jg3y3w9jxribvl
SXdeTgn/18+tW/9Ndpkqmg+DNNbOud3x4hVlEaKfpeB0eBRcivNrzcHkg9jv9qQsNAwdlYWybZkt
Nk558nnM4lkBFgTjNk8+9s1QGigj4A+XOw6U4SfXrawqeTfhAbnfrMGhiVuiq6Czw+2DNGvcd/6W
4wvPSMFejTn9Bvvavzn3eSwiCuFIS8b0aDID9umnCfZrzAly4ovmk7uErwg+YYCexuz6eohxOM76
ML+Pshkm+Y5VneEZuu2h0qwr4boZIgXFKDAp4h7X+mCr90gOAOvAbmWZx3xlQigbFQc35cgkuevN
pG54RO5YVbJZ8z0Ar0pxQt/Z7mq3ReY0pofqsUH8apnjeC2IZEis3R635LJLJasWG2nFsAZgOrC0
e4LT5hMxXxs3hqaE2YAFNtgaYR5fW+EKVC3rtdb3ICSuJfXCchN3vXIrU4505Dn/AFIQEobb6OvE
gsgqekjY1FxYXUDykDYE+FDnAbHAy8kSwfpKnsn+UIFS8dhLj7M8G1v0k9MlFBST/bb3cLt/BAup
72ZLNWrMpQqn9BLL+mfBVlHaurlRTwtegs6ieJXjLkXrRIIdBppgqvf9Ct5HQMXrIoB0o9j3D1wC
zJU65o+r3/hTET2P+ydGJiRHATsUeyNzidqSaEkQj1MzndD/KZ07TssAubDw2cKx1YcMBJq1CxfD
BQrRr0r1U1mVkA7w1ALblu/6HlQ1AEwOjMqO/qLGPzl4pyZxHr5IwMRJk3QawCpnJ0D1XrB4UGTu
hOPLoLLUUUBUi4Qnd8k7sSBikvVvor/EiGWfF8bzOv063drbjGyta1pKFCjM3LnFEYbnmfLTYeA9
n0vVgM0seLC127q5zRQy2haAv87oGkwRA2bXBOHMhrTLOLpnkWgTwXHVObNnZv8pWbsfH9CNTFme
ctSVqlZkyZhssVBXrDzyVTKA0bMUh3o0K7GKAyVklPlGgt+tbsm2OLR9AZ53PDO1P0xSkLo/Ou7a
Fn9rLUO5rOHw0ZkBGAYggazT2HUbF2HPFc7pAi2V+qAMRCdjPYqNPQxZKfR27X+iFtcuHMycQVDl
eHBcU7CXc7+9crQS1XpOhjy+Xqf84DcERFXM1ULdu0tB269l9st1bfvwvDRN5V96QWAUcCS4LxM/
13FwSe7GMtwUeGNbG3HBqzgg706CUGJX2BMm8KHwKUf9j7zxr8vAhAV5j2jsQfGh2DrTgeAAdfAO
+zryQcB41dwtPChyiOgn5vkw17um58LlcpfOeK/kIpAKk35BKP0p/qy1IEsbrzwSd8AJBlmOEIO0
pDmbVddwyAQI0QAoVEaN2L4a/4JDqXQz+Pk/eOtoGPD/jNEF/5e0CsHJz55g7+5CqqcTVYx/NVfQ
MD+wZ5yJ55p9YLJEnEG7RUWyy5yeeG4W98Xx55UpBnoccDk9ifR6p20EJqAglzwVhqYkRCyz4mAe
8xbbR4KuwjVCtU/gpZwmGzUMsNOgzLgwQBJEx4FRqnLGWXqS/A9uhvbBJ0gVVAXTUN+P4tZboy6y
xg3WvYkR3+lhsZUnd9JBgl/D88XJ23P7DSANbg4yGAzC0Em7cbasOn7JIDPZFgD49St7XmXgj32d
xQZRZ1zCZ2CiofAY6Sh3Cab44o+5L0Bf28GQP0WsSnNzVhvXa4mTMz1CeQ+AlLjmrE3+Dc9OYSzR
YUYhZc6k1CMZl02oU2hujPtFjTrErRALY+aZOlr6PtUs2d/rs0n4pO/2SdgcwJ8sPHpW9+cDiv/k
j9yRf/znuyAldGHhaBWjEF4+/qxY6W01AD4RS5Rfup10KAYq0FnzY8qSAO2auS6soevTw3WI2lq9
wvBACvUS292+I0/4nFGvME+uQeyImgdYZvwWfCWp9/LAnPjI5waY6zXIS0YmMiJUwcmgEyKJG6b0
XTceSrqMURoWRyZSkdJluLXESSo2R0/TMVE2xErnZGgtvezLnDkthr+lDxkjs8LU49nCBKbHAEJN
DWuRbNRyBdNPRveCPdTdmFGdlEug1GiYAwT+hCvGrsrHORvgyx0kW+ek10R1aREFwCA1s23y4mBg
IkMlrBheXezivGnTnuCqe6Slp1ngnzB+sTx/KXWrRkYxOPI78ZEWGsTZveYB3Zgdok7X6ig4f/X+
eeX7PqiEz8nWQEpi6plAIxFl+uuUqNpzXOoQVU97zS17fBJwT64OCAEVwXzcHuOeVTR+T/mVRv3l
gIDDTXhK/IhQIwk/69PE7miMc7LLAwoesH8Mw3q+F7bKUdg9CnAv0rwt1DCyLaLMBL3ABc1SPCTI
CDm28I0iUOWDoK8qGBaDdw/Y4bYrb7UgX77S6eRubcHsJjZX0tAdioC6NFIs1vx/lE/3k0FskIrM
kNxIyDPbuWo/ZQQgSZT+qBBXS4WN7feExOm5YELTc4GpoEquceGTOomDwS1VDaaeQ0Ayh6U5Sx5z
v50IFJmfIcThS2fy2iOAoKz6WvBAuFrvGvNgIxWeyhQhmup57lq3w7MWLA0PjwSApd1nBpzfsnrZ
v3YeuBnAXWORsFNhUopR0Zspa5fs1UzzqlICs9vehbUh9wH9wzeaTiFeeg+cz4EDvuvtLrlbq/lP
ixyr9TL8LAAW1aXJr/WjuyimjQQAMUcDjWz9SF84kPPHqeE/zZFminb6P3SR6pGZ5qMu8xbC7bRY
7q8U12w0+bblsiDUajejR27H5czV0n6cjqTVN5mNNO56O32MUYl7L0hHJ6dNpcjP8E/WmBhRdfIv
iVUcSdKhxSvGDU201NbHqobhS9ZDVSk6jcPuDX0u2E+8GjfTHZDgrOSsRKDpbJAQQtn9uZxbcP8a
Y9FNzdla/ja+mgT26uVtdjFIdvO2hnfwmtgzYvCFJwsaE2woaYS88/EgZx+lN3cJ50Yp+ITUrsY3
Hm/hLAzcRg1Tj3Cj3gSDDL+wUvFwWvNC64kydLvvHE9tKaspsVTf45pxYgcb3csufrxrxI3mv5yj
nGIVRmHDY8Nd6Fxf9Jj8b9u1lHXvw/3YmA50GuzPw/TPqS7tK7ZFNMu3XirAv5DYKRqyi9/ogy2t
g/gj5CcTkwH2Cu1ze+nZTEygMyKBOf6d6QvZtCZufSET13nTuekn5hxL014rYccfOxiBSdqwFic9
gxPizijMgIpJ+3z5lVhZeUFPpwy+mTPLKozMNUA6MvaHhaDhgBbwO/B/UelaN5y4HLMGUr4b5zZb
V0DpmCeVTBYU8fdictZZHZoOK0rPFKpUoPz2d8yAPCkYS8bf+vJaV3Ql+lC6Y8dMOk50N9mL88dR
G6pguRpBgAuCxAmrSxE+E7sqQF1dEWGFreexrrtrjsgGukP3cqxqYC4OmdQNRjGfGlk3THcz25w+
dA40+Xzt5l/WHUO5R0IUlFxULiafBwtu1kRPUt7fWchfxMohsOEyrYGVBbdJR9u6PddCqHCMUgeo
3aGSIXMohz/xmpTSqOj/O0kjoQHXmGZYIVaGB9ZE2lPY/lMakgHxdYwGnKjdlux+o2rcjdnoD0my
11xD/3Sk8SuLc9rMTZLWHcnl7VnobeH0TmsSa9QJexDIlb8cnEp37hmo1BPJ0f4dGgfJ/MuZOSW+
akh5toLKN+Cuvs5G/9r9lt/iltRdN4676y/Xnsv5I5qBexng24/xKIGsm6OJdjkHB19uZbFmaGgt
13USYVDrLbDbgM5CTMh7XUvnYtYiHXpuxCdT2MtfuXiZpCM9LYXkDfxvdWtKnSzmoIQOtX/J7etk
xKwSI+hYms2bC8coy5eEE9Nrd+SUhqxD2StxlgTM06AS5RbhQO16wAY8iID3eazCPCiCVNO05gOs
/1KL7ghuv4LmC0eEHmW/CQyOGWBS4KI7JyShWTvnGkxcCxxT+84wW1QpTOJ+l8ZOxeYOqA6WQi9x
Ju+qajq1ACcOEk3cBL8uFktrxHsDFEBS2wLqeGPe9peWWfnS+8Db+ZgXuNJyQF2YPwBjVMuLuxau
uiAf6owIveHsHexplKamnamX0fyqpB2X+09ebQmt+MZwG86MGNue+81fuckdU5LdI/I+QXWmIjWr
2AWnYp7fct9Z/ahJWQx/neST12YhG8Q2mCRSbRUvlWr95D/p3Rmc4YRGW2rTCUvPq/SPaNwO5E0F
f6fYFnuciaBGFRKUDwK0pk1CoNbw69bAe4YJKcJ0KfeBwlW7OoQk4QajCdSfSN1CvFuccomRlhh6
xhetQkrj+3gUjXn6yyl2Ekpq0XRFn2X+mKtw2+exU4KNdiSRXgEUqkk8uSTS7iVhx5ABVcKZjHD3
h10AELsExLBxaKiP1y62xQWLRNXzx8Ah8/LlebUX9wezAI6jtgZHF0HAtofC1Vxn7ZHZMwYUMW1v
EWZcn4mmb252VH56uVoo5eyixoey+EpKHBnIYCOWbLmteB0IgAqXsCiwCN+dTLJVF2hIPIhxwwYt
zrcTe5uPO4qWJrEtVZFFlRkl0Zbf2ybSw+3xDXL/kffevFIftuDRP4tWjnnWhYisvegIcQvXEw4A
sQ6Q2cnqnJl7uMhDPLr/0zwoeiChGcqS77hj4yOBLdHr0ISEb3H4Pd6CnYQHllbyEB0++379+KlH
ETZI73X0glw4JNPBsn4xEoDafClVwK9HKdtQB0YDV+CCyCVWNefsWra3hd5lif2ik9LzdZ834kRA
i0qATjKNyd2N0VcpZp1/fOY8dSzITNlMWAjTYQ0x28UdXzMry6v/H9OKTYP5COP9a4J0MM9QfJuo
+JKWN8aydzrhXmByo+8ki1G4zDXXADXbJKexSFpBcIeXynUffwovPAqp9UE/wQVdU3alFfPPR5qr
8aN658eQ9lt2hdUcj80UxSuUl2NjiCWGy5p7VsvzlE6TRqExrgFd3kcL0b74twKrnLx1/yeO6CTb
575E9DylketQ+bIP+SRKwAbKNaEexvoAFCjursIbqVhJlbefvtae7fVSyoa9hjSOikA5RcAJoCFV
X8wN77iym/bh6AvjUGIXxG9TwjtBBWUTCl5oSuZ3sLZnGMTTkwvI2X1dPJJbI1So/9sRFDS4oRgK
nt5ZKecqwcNr4EAuT3RcAquR82aQbtWzH2K0WYzqNoqXVbougpXVDRtpe0ZJa5YMBmFVIHL2/VBM
/MLjWjObaH6dTx3p80nLzJL48dxFS2N9MuyS8VGRzorfymyMms2b766PkohaskaBZm9+jY05dZLw
p5IeGSP6NujVBB9asnZcPFCpt2mdv0KXDIU1uRH9lp0nqQ70MN3/9C9DzXP3HQNwlFk2tjYtEfzS
lxMfbR2Al+m5f+rXpFFohzjYbuCMupkU4CaWRFRdw5ZOvsMuhsyGCpa9ztxR5u7EMH0OSPhmhL6b
Q96W6pktmILmIbfmb8fKrXccS6Ae3XuNBrvCMcocYjGixlPBfn5Fj0x3ixnEj2fETIUy77HR4Yf3
J3HdSTT7BB3PdU/3OqwP3OG2c415zCBwpTHTkA+vXCX/JnhVYPbrnngKxAfK26wX3ifynNZYfPDY
6yCLqh1vkiGGH1OVaydGs8Tg854vTTzPrdmWw6KnqnjTAEZS3WSyRVSEuqtFf7YulBG3xT4K/uM3
8GKmuvSzP57PPuAvZHjB86iDHHRqKXDQ/6l5WfzPDxZwD0Ky/V79O675ngK0ltAt3h8/t2ijOV99
j/slRNCJNbZB9HfIldg4AFJy5vJcmJL4hp4ObzxmqaCyzZ5pgT1wT3TXxrZe/CS8ZxEPuHYZh8vJ
mEkuUffcx7834RNEtBDrd0GQBFyqANRW6jno4hRq95zJhosftdokkocXqAJKPFiqJzxjK/yaKZP3
4R/GfhKwr2IYz37nmCETLPMZh4iR0fptQxkfDU/89td59Tci2nSVzKBsGfJOZIkJNjXhmsTICr7w
8Uu7P8eAWbkdfhxpaY8Nyj9dknpUbZBLSMfVKxGP41xryl2B7x48TCOD6qq137e5AnNFbiNC89YT
pJUeBpYnjcSmUrxraB1K6VuN46cDWDUvrlJngNG/IvmEt5xj5PLAr2m5jzo3uI5nEkdfut10hDQW
6bvkppJYeGZbc/5KoL5ssA+PAW6l25O28gh4KqsBO51qCe92s66WH7OoC6CgPcg/st12fpxMxr84
8apYZxVfycZm+1WiDUzMVuhaJPBv6XmMo//heIQbkS1gZbOIowcSMBaSvAK0JWFDFgae++SpNI84
PYsnWOABjDzSzgXbZ9cUo2Y5NB94UkK1hiu0q0+GxB/ECrZOH4ZG9Qn1BzVFwXB6JGsFkCEBtt/o
i71JWVMy/E6fUXmMs7P4HmD8PDsqrkhmsdQvxvl/c193XBH5seRVtBJrDigkekxfsSrDBUfknLeA
F0ZpKZ3eBakEH7XShQJkmtVDtOlPrkfAr9kGOEU/F6SwdDvP9+OGehH0w9Gj6wNX84SbSGCc7Dx6
149qvfD1WoHCampg829hVzZEXFW7H5unX4znQ/Vpc94eZ0mbiP7BgUJsO/kcBbHo44g8DWZNkH98
c+qkjehEyLuSiAH0/h5U+YHFqvkb3ZXmJ/l3SlcIdPf0+CQsNXICpHWHGvQ6+El2V2rvpFeIsY2p
aiFBuJaBtXB3rbHO3xbgr61G18iyBjp6kuo4ClU+VZFxv+vmhHdWUziQiGKzQNxK7PqdGTaRuvBH
TaHkaCYp4tFCsXUrtRr892fOS5vqAt5odKSa22i8KHi3S6vZuR4PUAuKk+d7EG4vjl+BR6EYQgDx
ElIGGU6QiF9QszeuYXS4mGFJ8IjHmy/pJtjZ/vk9l8O2jgRmj9XM0W7/QuHpwmk3W2Ig2GLDm+pm
uIdZkdmDCac+FLLoLoKZGkXeg8mmgwyefz6HkT6iq2b+I0NAfIac9Dg3QkwV+tVhx2u7VFMFw1tA
BLBtGrElhmmll2sTO55G9jm4ZqAc+Tm+JseRoeqAQM5hR8KhxAMgIwWzU7XGnYVNQIDJLw5apNXQ
Z+g/n54o+8ILclW3Cc5nO2rDGKKwQHYzvkDViyp5PEu4JqyRg6tuzI32/rpU3Lm1i1zj1GEOW5Ll
cDfpylR1x85xo/gYyjhOasBSoODB4h8byEkQdsihHTe7L0d4PszxF39UKMqs1sWRuDjvwg0diVZl
PcB2gZXKbUSp4qmkEfJksWZI0IMGFwQnK+e/Pc5t82oqPlO8IvcEA4YCnzVpOB17qQS6QrvHF0D+
SukZgck3E6O/rpIvjFDHbEt3LXkDQB7DjJNP8Mlz7A3I2H7NACebL9fsKPMYiyTHmnCZJFldMAdE
NXltcYRHzf/gzg1QYJfnZFuwerLLR9FF9tQ6UA2IZ3ho2F3UXoQkSA3Pzpf6/hawx93EFyiPwMav
3/kcMm8qZXFXBWOQD9J7mnrNJ3EmU/HIo12uqmkf23slMr33OwjxLUaZseNTmhklRbITAXg6SMP5
mKLpnVZf163x7pcufjuUsLnJuYwB+kMcVf9eTPIuX2WhkY7ckk5tGuAegIbF/G0WkzWBW7dDXJXI
dy7sZu7MnjApy1d452BjchvKk7oFOP8v9mCmLlBBJ8dH6bOZZ+4Mg6pct80M+FKcgKhBFsJHOjet
FdL/w85dK8e7h+ATOf5Gd5AEfoH4fWT/IAq5HKS//FRnje/1aQkEHTLYaGcLpUPNRTq7ShDAvfyi
hL3ELQJyN/L3h2ksJdJRorj57ANRXwnubJrGGklYSjT2oS4OQ2kFzzrTfQtLWpZFai3p0LmKoxK2
hLniQ49/yUnPKtMV9gT9MeR+2QWODOFjvcG1uOXCNTnCILHPfTojlNlVJPeTakxnY7eM3/3JaZGM
+jhUqmsuZWiamZdrhPwhH2Cb2l11qKWWTZMFaaSbEPAcidZYFT5Rz7ilfM1p3kM7J0Bq58QbxDG4
tt9XQID4jMKOTyNJqRfQ6GLij2R+pNVj9a6kuboeCwnYLjltrZW6igiCPMdNP8t8Sk8xyeeqXcOB
1YHQ4pbeysjgn64MoQxg/AlphLpgJZ5tmwvrOc3SeErdXbAYPy4Ede/q5EKFAlWKog6k6jWr8Ol5
pgCRXewhQu8E6rwT2NMcTHOWpot1i4ldZf4OXGeeYNr4DgUQzhMcA9FhxxOPzARfHIuoRQ7HXDb2
sVUGmUyJyje9fnYbgsBryvjFjw9IBo68gUkLItZhgCD4iW3bpd5ixyg5ItdXEBQRNVF13Zezu+sE
ZtyCeoKbWQNm0P6pVDxBNXYbJC0T41RYzuiwVxsPL2EzXcXZcwOKvCJL85tjj/J1DkrhICYDZ9VC
XpCzZIL1Tya7JwFTkqlyEye794M3za/WFduXCUMk+n3bBIl7zKQ2o/cwLbWftBdYzRJq9/SAUCYb
SrHyF+oXOEhjr0L3K1nqych5sieOQZf+ye8U2Ejjty5WMIO3vlfw9Ue4//vN8IQtQn0LC/GvsJHg
DU0MMmruArX8GiIDPVo8NYVwhen882CRckgKuHXMSsRWsiwwSlxa9KkHUBbQVP0f2kUeOFU9cpnK
ipOmmJfNXatjd0KRLPSfOz5R0K/E6XJjjQHbEmfkWgqkHE9R/GLxTmXlmD8namcfN86aFthe97f8
5f9gpIrfdaQz9lsTkGGsqAncRNxViJMOxHsynoRYOekzUYtvj1naBD7DCdSS4/eptXV1dLMH47so
lOOA4qGrrBLqR2cGCkacCQUzblaYgFtGITkNSYUJcm3Ft/sUpYKj1M73YGIVeg9zuZm40M5XFfBq
Rw/5bR4R7pWixIIvWMkUA+/x2Vdka41USMBwpfelB7vAlVZdB3IX1D5KIldygIce8EMjC1h0N2W6
fYEx8D4rQWZB0koH0gz7RQfHdv2Dq26lps5oOmgiKvDtBzidJimR2wj1TUoV7NtWg57RqgzYTjB8
aK2llp5xDDCJNe7QtuEB7zzfZQVT4pWzqQFnH+O/IRh4bAiQ8cJQAYHmxnynFByu2OZtacPLMDUh
0z5oupBTyJE6pvCdjfxBo4E4RBftztePCZpZrKbbG9gWkUQmyQUHMVpjQbf4RLlgz0pd/YcGKccb
fJLnyM4eDM+OTNSz5xrWo+6kqlpcZJ/rLBQSWDdjk7OoCud3XyBysSe1o01GI4ooFjbFjFaxx4X4
Z8afXElmCsL9GgzomVwTFMMkDbvK+YSNYAsPwjY4dyFrWrNynsqv+GDWtHdSrwklM7URU+qpPLA7
9o3diea+c3Nq24HEYtUws7I5nrVU/3GWnCOMfMP9inwSSmCMVCZoDrGH238U6Ku5nWiKOQLI6tdc
+tL1+pnoBHKqwHyLSRLTxtpMOQMqlInxBVbllc4+pMPAyImTz4EjO9MhFXJp+1pHZOk8C4+atqgh
z0qtYZEAcGsHyEJIxhjRwtf5NvNcwgxnftxyTaWgRVcQZx7JRfVT2hBqZrXqBb9z2woYuAMCBhbG
DY8+wZ1Jn5sLUMRdteN8zzYivQsszJFX6Lo4bJnorOtCR6bliZNnE+R5L+5cin7LaqX9+zqTfSgO
rJLOhARekJWrMR04K1lgqkzuZjR9oR6HYGMGjmpMGxoeq+84mAJktyimRvxObTD/yg6LL5c0Ny5R
ohPAS3Po81cnvMf+1KRTr/WKe9T4Ji4SASUKv4MBhSVyXsgoPeGkTZnITeH12Lpa28TkKUhbHwd8
qeS0oPovhXjLNRp8uruhxLB1DBnW2K1moh/MhjQR1WsiOf/2T6o21SsPticRV5R1Xdo9ngUv+XC5
veFLoJbbUKzBsapixJhTkOQ7m621SBHbo9nV5h9dfCGWkk6XXhX2oTN2mcowBqa2DklETI12Hys9
RzOwxF2CkPWfpM/B+qkMeKGq55d8/DsdHbRh+Jn1DlsDdomaHB221mCj05rTTr+HvAkbTij+dzf9
aFjnvEhFfcf4EWTur9CVDQABHHoes3AK127mojrq7HZJ2Y8sAY6w0z7cH9iMVn1rK00MKdfyNy9n
aW+FUXtLnRLKAO0SlljRTDi2MYIZ9WuCpPljcs+lY5qosz5p8RAWium5qxxKvL8Jau4ZjLYkORfv
jA7GA5cFEsjiOaqvAy8KGI8ZVx2n1iBm1zg+epmmQvuodW3CK5Cajp1y87Acs9A/ysHMI/tXxQKg
mRCg0+ZpmOM9cxndGKvTIb8aJaGMSKH03NjGhhEJGBeeBLvpyDutRcPMwupw5KCDazMAztnqusDr
dRUcHmmfTccBa4b99oFVrf2oH6s3+5QPS2/KqiWzZas0hunm56Oz+UmfwzNCiLRwODK06vEug40f
S0KvG7ntiucMS20CI7zv5LNKiiqnc1sgW9GkcgHYq2l1JFh2UU2Z5ghPsrXvRKgETs9LDqCnGHod
1iZ33e6gFLEqvI4vYc2zys524WvWT+hoasjw+Bja2RdFS85r8XKz4n/LE63/oZpSyvlDMGI/NBY/
kY3LzF/BJ20WrS5LbkWi+2BC8DloXQ/kvcXDUTJTl5Na9nfMKUA1KUhgtfS45hIcY5VhNUZOa3vx
DwWoqPyq92cD7KknnCdX8iiUgk/Xv0oTLHfzpsURZTThPW+tSZc2k3j1xfLPaWLOkKW1pwbWYk63
VTvDDc+/d+sPVIxBZnueeMXWTjdHSz1ekHHw05hweQbau+xRFSHkGyHiVgdEQgNKRI/8+DRPGnJ/
DfMFF05Qqj+WZRjg33QZbcIbzM+QGpNzMOWpvvZ8u2yQuO9lsF6t9piFEbHQZyZFNaFp6oCEZpAB
71/f2UPDlFJGgqIlMjC8eG3wxICqrNpm8xDc8wWfM4dxj3whBJqOfsR2t81nRExzk1JzittH2I6G
0xw8jCp5p2TicSgkyN28wY7kubby6Bei4bgMhHJMfGtZj0q8NCDrUvR3kowUOyFqfVRS5CU6zarH
g2DXi83DugR+GTWt0c6A7zNLclQnSVSAJC1YwBfutihm2boIKBllrj98R2X4HA/cK2vLvcGwf3J6
r2oZa8FgvhVtQOJ06U8AtBj+UV0hAN1oLCK4pWwTv1/3GAR6HW7gDC215GgFkGfDyTMomrUT4jpC
0GN0rgKnGNTV/wY7WWmj/w2vN6kAOCM3cajoRAAz4Oyxfm4gHNjo1apOa4FMWItprqab+NqlPJQm
fF5dmS2XMGluw2KOecMZk3kYejscU/vpxMBdczmAbvPeQo1LkiqG/3NJRI0ORaEdjOTXD3J0wuVo
le1L0Wfl8Y5Iguu3RXSlfRf40Zc4mzhLQithcQLjOCMqBB0Sx5Qj3VSqoiJpm7/qZMAQLJRqhlTe
7XkzCbirfw1jd60bxzRGsnHIa3Ay48wEcI+9/YIFGolgVcLqBNNZYYXSeQ7gC98akB5SIgm9GB5r
9wUkdeGozDn3FcSMwwD7KHF6V5sScUTm9zEJzxH7OXd1hN/S4oo73M6I9+DKylQIg8smeYjU31Fi
0LFqRs+53IJvvvc5grJ3dk/vmfA76wm9jw70WiC5Rg/oGwJbPdPGZ9Eo4CQ8zoHL9hD2uBUEFtu9
FeUkRJUTKzTypoo/2Ih1uhjsHAmIC8ewszJ4DixD4klllLtbmTzMBf32rP5YXEL6dGoA/fiiLN4v
d4rsFKGJFd7BRudzWIkpx2t3H5Sbh655Qlq+kNkN6867+Rrnk5jolPbXITSyVJUdDvVvavfIO9Oh
bTRZvE2ebFfzK0YPLgmN9q1HzluZm1xVyGlI0/I3uGFH4dBuBT9Thd9q7BkcKu/lbIrt0hGC6KdQ
e72i9wp1SLhqmWR9OSF9Ft2exswTlGlnBr38z3E5p6L+HT4W9M3YOXbusUxCjdxstsc65SG2eFIN
PNE7bKNIi2xrjwVRR4OG16aZlK2NXHHeBWlbhZSx6QLvurfrPC30RmgzeHFXkOVKwtGg1T5Sg+NU
ohk2tdnK4DsDC8QO+sgouOVg9eQ7YJzXOIQPgwy9u0tVoYRafI5eZbugEGAG0nZ2kQFeyuj86Vqa
aj1GaHrDo6MYwWsP6E3G+mf34eIIlJzNcJyauDiL6ixGxcYihbI5vgjIn+mcUsIKfpd4Ss5GIHnF
heO9iQLtT/spAR7ul/Cn1WSgMWzsIXcReRUYOixZrAory++eEoJ9cnhvmiNGmS8bvkE/2XjBt3Ht
kj30FRQ5UMkTIdQdGFj03LLM63ZAg8u15frLX9QZjgUp8dQZjSNG/3WSDc1u88reo5v91HlOM3Mw
JmJTjnzHTKEhvA7lcx4LHZZNQfscJeeNO3tkP/6kwM6XvJ7+8MH4gSqIsV6YaFU1ngyDs4YLWyqs
Hfomq3j/H6m25zSKJorKs++8qn5VA9q6Vg27ZjVEeFO7fXSJL9guUYarzMGrT+rhmvGcM8ci4RIm
4b2EFY58rrwR1PYgO8QkZxqBCFZTN86D0QxFZHnf89c2O6xl7DTpOHRiF468lWYWgXIceOnj5od0
IvZaw68zGAeFWdDqCV6Q+/2Uw/wtCs2x9DxC39kMCK10pf1j5V7s/fV27m50wuYCHMK1stEkdekn
xD1ZgX7pyEj+fIPNsCsby03djIk6X14Red3WJwk9suVY3VDzpUF+uiq/FVwqsnsFkHFGyHFQh09O
+MMrznzXNuK+KMlmmzsmANV3UcVmvZUIbUaKuTaij9GHSuTK5P+VeO/W6cEUXoUhf331ziLPL3/k
1iVUqtL1AV8U4Br+s8em4btpWNiKrvFl4ILbFVsrUxijaqsgwBipzqquAk1kXsu71Weh9PU0MgNf
ekHWgKTVsiRK4gt7NftexglnfB9gFEGyYsPV9/VXQsxEogomvHiP5dT439Zmr34uPG9H2NZ+S9Jb
1zbYLq9SkHpHzauwqArXcWlmZlp3+JZTgeqjBYxs+GXn5eBjk+8MtHYwytUKiaEy3Ni0+DozkDYB
84dlyrSGvErNOsgB9Itbfx3Ld4y/uKHmp8wDn2fzwfz7aJxQas5AboBMc/5sdjXtSL45BP0PQ5YM
sLi6uXjYEQ6vva6bXcQb9P79ZDE3xcb2Vo/VpjF1bqGW7dPw3cr3s+jSm1SDWYUaYBUnPhV9GgZS
R2+xUMAIBbuMChPAcq1cSEItmd6j2fMTvaMM/u6aFRsid9P5K7WR57RJ6QqWYD6deA7w2F2rK6Se
a8EkGFQgo4OP0RukWPk7XSCCDe0Ns4RsRXb3MvyzMuNN/Xbvg2JWvY5c9Qc88mDjRy9DNrEaDXPD
FC6/KhM+mbs9VWjFSxhm12anBiPekasNEllEuHZH2wXppI5CMpbxGuml3DJ3Hj9B9ar0Z9Xt5mtw
rl0WUN/yGdzdD30BdC36V3mArsrx+GPzBPZ92+se2VN1NmTzkHVy+292+qj3If4B1zMEWyB7VySr
inKA7ylIi2CudWksrCVeaCk/oo7zdhVW/NTkg2jO2JTMDcUaGa0XnR9Pp6cVM9MF6i05Hx3hh9We
U19BWrlfpfV+krnmtSLUChxOrjreBuILsvmczmn+8x94qMStO+NCxxeSzjm8AA4eV0wURlWvDwbg
Q7uTDAVNQVZDfWqnLNqCL6w5o7/1QqAYxlxZoaS4fd8WrEX+8a1TXWq/wPPw9pq2IbpMrNn97vxC
BeKG0NZ56z3FJmG/BWPVeO1EMnrluQUFBmsatEA5bjPKvPFX/tlmb6gDv2H3tZx2/BA0eM/yb5Dm
8A60jChaoZHoxO3DM7Nrcad5VggehXJhzUP3op6RYlbTaRd+vnXTk5lmqv4e6NS+HbkCey7nwE0O
3PWmalTSEQM3kwU2VqFffex9ANWkE2SZRosMdkVtEXh3hQ9Lawp3PrJBgUyjQjDZYZOvyAwx1vVh
NEYUQf1R6n6TpNwFqolbcgFmsUFs8lMr/kYK4D0wAc+KCq4/dnm3Yf2CAF5I2Fbk7/vNLX/N7O9e
G5fvm3auoikHBtqQZ/XW5ySw7vTiIxS6e2S63gOxB81pzb3jEKSYa9JYor5FQCK7kOG8fB4xo+7u
d+nPyvuhLVX0V++ukuR4QY1GC9olRA3iqCMiy/2+XlDtghKReg2y+uF10Qn+tHwo//FQEpXWS3FT
HgmBPE0VZvqrcl9sle0MNLcQpRZg8NIsmcexCvJHcrgTz+V4hjr7blV07wSD4YB/6c/GKVpx6PD/
KmKKKepN8Bcuo3mI8iZQkyEngBUW24R9iy2nnjq+cbCsxDYF7+0KQQSCN8VpHwAll9EjfiqueV5u
sYwvZyMIGtENcNV/3cfLavNXX+8o+DkqHtIjST/aeIOBj860OxScpHn2SJ+e+b5bi1g6ANqfZpxj
80CjrGOK6QgZCxi8ys/2S/r6ZV5Se3Lk1tfKrOPLUw8ALKy7X0TQoFmZCMZCjWM2X3b8hC4QBhAU
uc4OjtpxmvbIMHwY05BnXdnvUX6oU17HL18EjC/K2G+dBh+T9Tutbsj3I3lxSncu3gOPzL165oVg
RZeZhwsibjo8Bo5ifRqFzzaqWuybVbVOAl2Bgc+j4u+jDfr/um6/KkEtw/DCu4LuREzkIFhOBmZX
09fD/lU3mVrZw/HC03L4+6byN/tOBvwrHorq/Z42EGK96uKsIJ7Tk9sInAW0MmhjWcJq6ouZ1VBT
dyOcc0du3VUrrRXNubFsTT75BZcriAd9ur708YwERIviqrmwt5Bp4J150khDPxSk8VAvt9zUICeR
+FzTIjG28aSvL49q5Vf6LeT2XJY/uldy2jJeNdV1CoZ+amN9+f3GHK/fXkn9H3lP61f6mExwIE8V
aebiaS4o34cz7pHTDc91RCLTlHoE3CtrSgAMH+TdXEhRQ4c/R6GBaoToBc9gzRerzeOUKP5cvHfq
X+aL55fn2b4cdMjBiDGA4AtTL9ZIQ/cQXWdSjEVviMkdNAxZTCRYvxwwuClkf5vh2EHoYVgNjwNV
f0MFz5OrBocw056CruyYOAeW0Q2+jEiJiBRGrL5h9G4yl5WEA10h1M22pZG7w3N38S5EGNtsrMi4
9xPDZgP4s2MR2SVtApw+4K0VnTQJTOE6ahbuhqrviDyfbhOdtlQQIZmXVTSlSZFSzI38BB3FgyOo
KtvJrzk86PCLtxhkb28aoaOSFOT1rRDib1HG59TrbIotuI/fpJ/qcpYhgBwW7gFLfdyipIRdfQvn
1tOl8RbIlQzdO+Omq+3Y/LQTvifh1qBIbjCTBT3+VjefZlfafQk9CexabLodK5iTQDS8b5BTLXgn
QfxFcS4c8wANSmWra025vsoAqAq56FIxvGD1nZsvn6eS447omVTbz30PAxFDpey4FXg8hNTPuV3G
eeU0H87MdSZPRWH/WQSbwIdCsEwj/wuIoJeoQ7w7MbK+QBa3PLbRKzO6xgZE4DiVDlDVZEYvW91H
TwXYi8TZapaD/yH7PD2Q83zuAD6X62L145WYQ9XKsSKQFTQBOScveqx4vSZzAj4xvdCrRh1o1IL2
vsO9ShpoE9GUyf4Q+4bJSFFAGFmUX04T3y+RNrcn5hh9bB7HDH/Pxn/Ou9B5viilkC0R7HtWlLRL
R7neZtwMN8cTIzfjQ5g+NkXfWjY8BjgzAM8Z0HyeRjpuJT2x0qwYnKEemD+xasr7xSb3w4mVR56V
BAUiPHRE86jkGWC6EP/RveSfWQanq/TgbgtmTjk2CqI7GcWRFJNDag8aPCVZHkthylbZV2QD8P8n
AIBRo1UYticSGYshh7Kl+WpHaf0oZpkp/vhIkNlNcVmWsFf62LUwDfIryhQibrt4viLLWdD5Oji7
bz8Ee0Y3YZbuFIJvXMrrGMBEC0PxDzbVsRJv1ieK+hTArF8c89YK3YwimtUmU1/vlFu1FlPofW1V
771hxkbqJ29ndF0n/o/3rxrfaXEWOEmL5cGdz5/oIBtPatHumNYvJ0eZxI4+V8KuJyiXx5fxR5Dw
0pztijFGS2/0TOyrmnISD/dIDH0M6Isl0zY/H2sbYMH09b1sbFmYp3U1fojyOmqZ+WGioFkAuBYD
aNPU6Z/LooBh3AqbkMoQ5IACL7SK0BcpRSQT5PiLX/Fnbb+L8sqTGJA20LCC56fUoqQp5mFfZBtW
z6vNu9G4BrJmMeYdbvLEqRjIbbJ/F1+6IfDGZenMr+yQv6mcM+6tIzDycH3Log6U5b7vpp5b53z7
JjELZjUds7SVUz6kFlpkb7hEE9AWSjVBH1oyY+mhoHByXInlQGIIF6hUEy0d4iXOQEjO2WXJR4pU
zXkO6MfCvgGxNRu52pRVxB2sUvSTGTwLfirPalrEIKOdgglCCqddLZpIzdq6bnwZGRTP9J7YAxD+
gokHkOIHhZDfFg9NeJslz5ytE1RwxPIAQcDVjjT6FKBYjSGF7qkAhhEImnbJfSerMf/rJtC4zJtG
9JHpDdspCvsyb+u9HqIajEX/ALSdIClHAijyeaLtbLAKm+yB6dYL5TiyKIGbTCvEdAeqVbTwzpp8
QxIvHTwL9i/zTkwD/sUySOfVuM/zwyGS0X4xdgwX4mwWZ9JVa5Fht1+gVZcuSO0cNUUw9EZXT1t/
E/4C9daJIuA0qIWah2q/fU2OyBctNhHjegq3Z32s4F+SHVznVJcFdqEDwoqhRo2//eOOq6i9NfZx
ezYiup+sVQEcWw8mq18xpDeBquBOYUAAyXh6z2nP/CdvQ6P44HV3n98sGHDVYOC/JAKQq0/mfXie
p6pV+KN6NEhpeYH3w9Q5hF5OovpsNKLQm/Wm0nhjooykexGs026T4u3iaMgzK2MgGnjHC6rSwDwB
BD2JY/ECSn/cxngXt/6tPiuKcaGp7DBmCKkoGFjdehOv6Ii3daBiZSD1w4v2Xsrqm4YrPc8A5Pct
9OHsMkCvg7+ZoIx9hCQwZbF/OxGEEKmbOXVxRQil5eqXCQY8q+GO/D0sPbBnZX0jA8pVTehht+Yc
z203TUXiYavKXzAtCUxKLRV1Jp63u8lxm8KWR/XabKTxENd6+utgP62sl1uhoWtT4NrUrgjoZcwu
TBTGynvCVsk94u6a5VyaxnDc4QAwhnGocwFKuQ3DnWrP6bOVlq7PlwimPID1jsJxS6mx3utF4Mnl
nY2rUnoJe4JZrpqdHiGa1uA2rv1xZOUltZ+fpvWZK4IbN34kN+6ZeTqrRq56rXfLrdkZ0JkNNw3t
kuRdRwYvkvnXFoXXYBOHxNE8cCf1D+lfNrmI14sFnKUHqz/E6Al7kgfA8cLhp5WlBBFz7xlBLgPa
GX3gC/plfKKMdobhcC4xyv6b8G90Mze6QfUDrEtsAR9O8O/2e83wLQ3H0lH+Snn3ZAGKB/bBEnMU
v1xvBs3soOxHzwTQ/ZBlFlR5xhp6vNDQA9JWdFuTblK/mFLRHlqXFdz2ZuViXdi+3ELWcCX3P/Vd
nyJqGzg0B+XDxfCO19wNd6Sm7Q62q3Cv7XKhCzod8S+fZQfB9V7ahq/OMsm/0nt9lFcT+TUGjhF7
s37ELzn5X8sBb7GxtqMnS57RN/3WJFh3S7sQcFIESwAYp05ikPIxaBpoICGqeUdrzcPTf0e0XW7K
UES8XUUfQCWt5ieV/AbZX7AkjfMbbUYPNUozuDIq77LZzbMY3MMyeqkZ55F/x0mEGbTFGX+VdXyo
FStry2JpOcr3wOZa3oFVibvmrkQOPLpj3h3jURSQ9gkWexusvm0d4S+suQSKig8etFou4rR1xIFg
NQI49/Ia/RRPIRsurJb2GQiihSzMJCCJzZXTDu3x8PV7hVWSahYWHJV1CYe69e9X2pqfG8NIk2Wo
LkWVsEB5rcgkkboLOQS8udK/G3QXwvPfithUsNtNIMqgi3Uqaompn08RCE24GEqMCR2/I/dkGYE2
G6gcjOY9AnCcQ27di8orhvvAB3bgndj/Ku9aH+ObyDlz9QaW5VbrZBWheDVVDmsltmDYU7ttMB6M
dkFrwxGAgVZGWvU64WtLw3Piai9p06ry/3AeQsL3U229jSAKIJ4g7io7aArv5mKvXoIDmNDi9dSA
eGycsUc9nxCahuAmXHTVDMv7W7p1qgBLQataDcuxYWOcZCDEghzrEeo67Tv1gwbGWQIuXw1cA8vZ
WT7MGZwO1BY52Nx02UWCAadCsul9Dztvdr8+msZGLGDEQxAeNKEw9vCRc+qQCYUfN++DYyN12r/a
nH5IDIMILBbzJta00gkQlRNVTB150yYOM/cVL+HYQQP4rFQwekB4ek2slZgy8SEIsywSagL8bTRt
ZcZCqwzPXmUclW7DxlEbcW6Qjov4V7YrkvztVLxPdWYZdhTQOuCOwLQgHbNq4zTDJL/MUd26lXc0
Ul+QQznBqeEZydwFOtSd7SZjNjgBi1y4E8pdVN9GlnuO3SxL2EPGr/zHXomNg/t6p3mIOrKwS37d
0TM+IFbRMWTEhvelhdALGzp+mGoek342IiVN7N6coaHKBLaRPvj17HZwwGaT67KMroLEQIcNxS9o
coYxDdvBPUeZO4ol7n2OdGuIin6NgMUXrbluWZuQykvGOKNeyXaAsRURbFvLsi8jC7zJ4h0Ya6f1
DV/fm7uQfQ7kP+yC3v2gqDq6UXplNhQnosl8lsdVuyZY6ItPPXZk2TconmqzjegC2MRwNHzfz3zZ
IZc4oklrH3tPCFc4o5g3f0IegALykMzfTPxaSwovQUMrcuP0QAin8WGtzBxbf86z5Kq3o7Ci+462
TJGBYWhbsULmkNNi4DLVWH91zsfkYYEX+t8/69OkVS/NV3iedQaqm51yvDRYMpjTKm0E9htAYPhq
IlwW8nCnauWf+lu61i7uyofEmJPPq5jyJb4m4+oEMPgjR0NJtUA5fPGn7czsSrrIy4HfvDl7nxSS
yTX7KmY7/I5ni1bOH7/y00Z8Q7JwKj9JYyvpEDzH7lDy/02L6biL16fmvlnopoa5snezteiWT2q9
NKiDc4UFcTpVqQf9sFbMnkKcxMX+RIJ+5Lil6j+nQ3EyLAc5mUgJFZ5UJNRB9zEY7tuf4791bLdf
FOsqMHO5hUkgakD2N+nA4hh8pXy4hsfX5Jx7DlnQUasc8INMUNJULoYgZckEXnX/Yc/XOqQ4cJ4A
zIa068usyZZO4EyjG+xWW+mVMt9+BZU/Fyz7mR8deGMzEc4f/gv78MdTpCU7OmQuZzOTbptWVq7L
AIAjZ4ezYv1ttRjeet8niENMkWJj6MlhibFe6FR5UaehgdvlbM50M2/8xlNRq2x3gE0QidtNGpRt
LRAmgceSzAP26wVuBctouSuncEBMEIOd6LoN+oKpsShn3ZJ46hcpqbIyJtvekFxiHa9VDxM0Yt8i
wDtyMSvOwEe8ZyGoz3rO5J+4FvLI3v5M2isvq6kvoGhkHbsz1Nupk2M6itJ4Mg7qjmWlUrqgkOZ7
8MNfEGwfTy2BcJO3X4YAkgzmtob3af8dWnXvB85Pt3ZRhE+VTsodSi+hKIpgXkEYyppy7UdYMZxz
hm+HPb33OQWQsRNctLg8hW9uCH3tHx3gOs5fxNw9hLvpGvBzkHRZWofGra9BazbJLJFcgCI/+SyL
3PAslhdYuEk9Ufe4hjiEGF5nZjo5MBDoh4kAAHvUr9PSPOcCUuRbOIOy6JOcahWa7QfGHBnluEOH
U4aLLN1y7XgG+L9zSwguwoHDgzofGCjek4W/NLhcsFARXfiiAbNQNltDvVzKiEYnHo9LLVlbMMGK
l92romRl7LxBE3ABy+RfxjhLuO6oMpXV0zKiwCUUCBsrBMg1iO7QAgoMJi3t0P2kh7JiZpBwVLQy
KZEMhW/0IYlls+QXBbIcH+S5EZexbJ80au5kIS75bAtcxXM7u/w1PHTw3SFkR+oQj1whHf+ns1D5
crd16bw2c0xjanpSzFIj6F2ifjkqh4WhqFguB5HpaYwaIFvPLrxqunYwFI5CQka6/Cdc1kiFXhxY
0yf8N6lLFWfXCh2Y+tNot+P8nWdSaKcPaBp67jfoBQG5Z/I4grkPY5jLvi0GGuZxIlEnxD0LjvrL
7FtuaCAlWBaW9MnWiMBwdWMGVzOEkZDdDJ0lOAZtK+fiWn/PR1iy5xbJegwiHS8uFevKwPWxcQ/E
kw4jl2b8ZF00mwsHFSumC5S+hQDaWnkApUM8tllCIi34Sy+7RsLGKG40851itBgga1Kz/SnB+uFT
5SJNf+llki/BR4xCusL9eE2JnmkfEFpmu8NwZwMlcsVG8e86Lik9gHHdhy98Or+5WisI86D8ziwr
cIPy4D7MmysSKaZ7ZeGqMTSwGxoWOs02u3WjlekdpLeARwTjrIRdVyBPURNHTdYDu8kzyIuKhKlI
SfVJsn32W+U4KmKk6JnQgYvHT4hXyHrhDF3Z1ZepvfRaHiwxXNpZGoIPlzA8xbDXcI9O+TPXTNNj
+9OAs3OSCZhEQelmxxuYqa5Ywkt6Rotf+1CkjDpQcT0h6gF9tIfopZCnvogc/K/H/pbdTbyNDVXS
Vz3vFQ9/KaYAR7Njy8IsrVI5+OEyVKZZXG156kdqqst8Hn0ACcIh27j9dClY5wbS+gJHBj58fSGz
zsFPELUEvNCj1te5fe1t6FH5TI3tRTlIPyp6kp53C84y+IBTs+2fJomY0QafZrfBy/Rg+B+72nmq
LxlQJkjR6No6WzANcrDkG3A0qcD+D0cq1lD8SV3FnnE2cWyXuhJs2cNVfJL6ly28zMMPAXFt5meq
2VSn8bKVPo9gU9qPPw/2Yyc8c0KVdwUgKPsXNc5Ws+hTEU92Q7lIectMtM6tYTJqnxl2Crg7GGct
ROWPUWtnicDO/KVhKCFcx3DQGyXi20Bk4br0o7atCja/67srrKGiE5XLi/5wCwJfy+7znqIkSQ5O
EQEhWeLg6ZcPcM4SNMjdpxadNQNL7ELjq6jzfBAfS/4k1d/mu2k+xY4ujZTND+9t57YeNkCL3yMN
f/9HXtmQxMVoSUxv7N7G1EjhdL1nZO7u4/tdGirm//I2FQWaoAdEV/egNa00kdFmVN16BVKMuupF
+jRtm2JGfQlZfzQb0zve4nJHGrRTjEdz2npgUk0nYWhzHx90BwnfOINybP/z9i2iBzRLSyPsc3PA
sK8wA9h1WDTQ2WPIczpK2hM25hp/UDTFPfnTgbtXzlGYzABOCIsAKB1FS3t+RbIjpgRh1TtFZcrI
WYsCTXfctpdAPY9NMvzvuwrIthhMzXI0cDHk5x8k2hadqHRqvHPBZk7Idw4MLL8QV5jopz53XPnS
YU2FUOoKH2YZlWiAj7hFoV2tuslt+os9zbc1/wfZOmEsfgmTbZOwDeBVYHNc7CnGUyHdxpB5hF8Z
QhUmVp+ngSqg8eSBuhvTmreegMgEheGBJfEmae/OZIXu0gGNeT9HJUBPx7RQ+Bz5tx+xQYSxmMib
Kqso4A5imqeg7aX8XylFC6rkQ8B89wZWoPzF/lpY5lx9AXwrOlpNRJwmHGbtIwHUbG766r3AmU6i
En9s1YMAI3TohLLqze6LLzfcFAN2KDuHZe/sZ8G9TKJl0qb3zgjq5m96cSpi6R4WTA+WrIrndo98
28zLFGRpQ9Uyuc+oZcMEsQqFUfk/OEdpA84zPhtVXdTt+bYs3N8XjFAybwVbzFvCjv+C6V1/zJae
lARzt3UpmNY3+0cFDfQtupejBuU6yRL4IFH5VhXVSX04B2n5OyqjYKPay2kVp9V71rpLpKAR7MTe
b5IEaOc7qwbfR+hYBM1hkoU4WWvgxtn0IJOdyX+1BnjXIMpfrUiWlxHnanJhmlbpJxslB6Pb8P9s
Jbz/w7xu/WRW4ceRCW11p3POP0wpK0nLrSvQHIHWwvTX8unV5cK5h5iPn9z9FIsqZJup2wvxpfSe
m0c/Dhj1CRjAZ+PJyGms+wME72ag+QAvJ2AEUFSwtkqtjq2x7BTttaYCzT3yv29tMCIKo4ViH5km
8G1ZJAVgNg9hirEg51m00Zr9Y0PBaXm4EHgjTevq8H9P9m9sQur4UsHD/z7uZn8VHKx8aZV3z+Y8
/p754xJWhM/AeXT6oFf4ODifv5DnFaN2QAHbcnYUlJWdjfd1Or3s5xXyCwQauSAQaQtWLi0xYJuz
JjLpGmb3BPeeCafADoUcdHSqKZBZrS8+F2gWKwuWrRQ/CnzAAUKHUaUYTRhwb4h+LDz4t7xJc+rq
wMW6cS54YqEaXWVg7i6UUBPy+fvJKifY0vmxkNW6k9SHoxiWKj3nxfH9e/b9oqQ+zDq/AQfeNzqJ
29jvXwg8/C1CyZ9Cey4blPQyFbmrVvZYNQ6LSNY4Eu0FF+oZikh6leoxXaZuM2RmPkigJBu/M8Nt
if5GUvm/WXNZURTV0HRluA4nuqU6dBZiJHlo8AGtf2RBaJEOSWOeFvNep7/AbzLXkAjshU5fuf+j
qfqYlYGbVo6mp69eip+G9P/aj46zCnyMmEvJJIAHXtCSgl9GKN0iGe6k6HYvIVn3w/VmFL4aJFHx
w27HveKw+DXTxoQI4gxJBPaj7j04QlIlgK5hJKb/EauSNT8YyDWFm/9GixpJoBJWhNSfwH8JEmd9
FHwTtlOFzJbBvfjDuahPdTXnkIJZNoGBs1f1zREgop+qzBBgcYB796HaVMKzp80AsZBGH0c/eMdn
Dr4HLZBPlFn0/hVFq46JVGsCKm0pZjoZDbpshvGkC6eTF82wXE1yjHj+XX1Q91PNgaBwslt3fAkj
7pqTEFyTwPENoOqctL/943iurwE/cwj4Mt05rP7fD9vMCjVUbpV1tx4Liz4/lcbv71pxG/1V3KGF
Z7BocgxpYSHUHsnvwAVXn4r7bLp+R1FJ5d1CJIUBmj+we6vEj9TZXNmaDLRkPxqqI+Zx+mekqrFf
pCbDIgzYm2fdGunc6ArD2RIfyWcnA5QXn/sp2BPmrOMHx4NmFrDSTKAX15Feldhp1ybJuqvJEqLy
yCDJXM8EC163Z6TX4jXx5zpoBbcEvJJeZuP9Z8zmlrp9bvEHHaGmIFR1bhi3UD/vCWVaYH+Y191M
qS7mPadWJrcjH/kcFBBcfBdWP8PynS3hyID6F7F/dLk85lW8kEbj05DRJ3zt9nbXxSRb/Zof/b2r
rP3wuh9haJ3YsXinG8f5EbJ4KACLqlQ2dhj3hWovECy05fuq2jfwGbzW4srlSWgbinSVQjUJiTGN
HVRXiXTYxAilKGEB8L3BZjsnNMmQODigVOARs8+CF+sOairUvinCa+mtRRISeeTX/kEM/hlFp2Dz
VzuNqtz1uuaFC9SWF+DJncMBBz0n9VNHjRiyTn8rEyaBhxo1C01a6EsIV1ioybWZSBR8HQ2U1fwW
B5u5X/Pn58d7GM/9AzCL8KgkSu62nve5gk/4bBx53r7I8IzZ8BH1clFpwj+VV+9tyoJ1IfxD3IhB
3zuRbYec7kh/T29FOlKUncb3lmlfG5eBQjcAQ8K8ptqtbJOWNnGElAublWNEAHT48IcS20D+nPeO
YnPP0CkRN05C3QGgwPf5ZrhIV/ZzmsO0HKBXfvWqEU4ELmrPYBfj+miWrRm808PorNa+C2rffwd9
HQkJz2EHyP+gaX/V76wenMZ25N14XjYA08qH+mdUmMllbbRwvB0kdOeOrxokLHdjoxeVYwRqGzlT
aQl5oK/uwrkTnjGO8JThwLEbgb6xxy+2iCD0x3CE3kFV9t3W/pBgGRIVqUCErTzNOi2KjnAU6OY3
VMGwqxH2LBhAR0lms26gB+hK1Uvr7nR3vZSFqKosY3z+MfeaY4tUEhDwEVuUYHAsWXHhA5SLyjII
WHvClrhJj54GotrL50Q2BhcQHjvKOZkrokDtdCxYagXFLrTTjVMEgDcuSLNyPnFhoLr8TZG+MeOb
zj75Nw0rcyBOEuozNKO9yS/YUyCOpBF3gzw/yjrlxLzLK0ynfqRge6Mh8EXyvuzSpJ6byouJA0t7
8RTxv6pr4zp7PwhEZqJ3A5HB6nkjmUbIOGOsK01X2FBiT2mWhrM4bP0H8VxfOwUk3DaN36e2ohWv
yi3gIoe82jLHHxHGDLNh4bzKkSDMxoizUS914P7I7K+gD2xvmM/Nn9DL6ui0Zb3HL80DpssJ3eog
NwMrue/83MRGF+e8WjNFDW3Gfn7IyVmtJaEy6mJDT/LcpvUsY34j9af+ESbSxqQNMLilgk8dOv5h
1haiJOnaTOPI5wBxY1BmkNht4yfSR9o7D9/LLYxy9Zwz3EanvP3a+duNk6EKe1J0sJO+1Xi3NfMB
Wb4+plIR/e6JapiWLoNuR1iQXe3Ch3MTjKrK11x3my0kaTJc3tX4YhXnWtAtORuvTUYjAfnd/2Be
3AHxntNlW/v5W39DamCMHOpvmJ8NPAtcnUqbPGcef7hZzIF93N4nB1MFLgkLryo4aS4utYp0AvXi
1MtN4QjvBN0u5poNY6D/icqxSDNZD8bHKGUE4ypXKwzQ+KzWPy8iWrrf4XMMjytrAlhPace7Kxl3
8PFDLYeUZnozKyDljT5u5gcvqelmN12QoD9u0fUlD+qFgFVC2QA/ocHfS5HqYTf4tm35/bJdUXzI
+mW/E9a/HuKQip0hQFWxNBvTzCADJrhngqBCgqFvPNhFOuc8Doa6NnRv8n+es/AwhGmEEYJdF0TN
nFSQLZR4Pgnkwa+Faw8Y1nU31QdQVHPBvxz5CgDQ3g5Oz/t4OE2OafyVpxeXNFvdsFbAVGYwt6xb
KTdEReTlz8y3uV90dRLbjKYZl/Q8ybhTu46EYoavbYmd3tZ5gECtY9EdR7WxRMC0ecjKdB73lAFp
fXIRg7EGhqIio1GnnotVBM2/yw4RIRUeGv5Aj2ARkXhogLlDEUPuap9zr89Lytl6sgrQZevA89Kk
wh+U+xjsEQnuqhNRIeAjzGLKSB/pV8MEspgfaY1uHGbPqFpmmBCbg8G9azTzt9RiLSv7vUWFAOx8
cX8r/lno/stRrFl+yZwg0qRkpvMBSWMEoCAZsfriiJOqUhGoQl6/mDFLRVSunhtG6Z3i8BIGCCIN
tkGcFOauG6rWpwhttpUItYRUQ8AU3ZsgNS429ZKGf3lzO3nWXaBeR9b2VCa4K0jAdNPSr0gCX6kM
79WNeOA7Je9BiPBNVg+PnuuE51OqG+hJn66co5AooajdHEJmUgkE5OrlBxglC07UArlegNBOx23n
ZWRZ0FSkfJyX004f09BGU/yIQGTwMGMJYDWJ+IcultmB57HJEUbH6u9u/l0tru3L0vZ8WCRxpI5w
oGG0S7+Rs095+dWcck1Dr/Brcoh+IVh/KwbtfaYceWdVuzVCdXA5whtJ5EGcMts0A9BysfYBN2Dl
f/PX+wl862eU12mRUfHXQzXAdXbd27jbi+F51Pa6Uocz/P9m2dD+zdavc1CzghkFmwq/OKVuCwUO
FFBlDPr3a9H8ecUczPqPr3i/Vxgy8P/U3RmW8NuaV+/6i/JiZuF+V98v16n0fJOGg9MA3eO6AVvC
MjT718E1HeLP50rr9H8diGsUbzX+2wI60el5m6NsJBBk3lxGQsD7GtYZ0w5T9dHr4MsIpM3vsQ2W
jaRnjAgLeUyS5U6b+u6DVi6eVRj1Tbg/Ob0oJFS+fcoAnHotDnmnOuwNnD3/mq2W74kJ/bHlkvRE
RYAMWlG7qeDYRXehDMLH069kNaZCpelCbkoaykL2cM8uS2f+v1QM3/MhPU7AakrqeANGCNi7U+S3
ookM2TALdfh2SI3bSM2UBjSeSLby3v6XdSaU5YI6KjtBg2POPDxLnJBLJHI6fZ5YWzbLAHtKLqQY
yWYbK+cD3WUOHfhj1+P1qVJa5rTrlz8dT6HmMEI5wi+o7AOGCZoaqx1KnK5D4Y0EGkueK4HK2HPS
qK+gneEtC/XpDg9HVt71pb86rS4vK/mjj6I103jnC+8SfCMIZR5jNEXSoL3bEACThZAQ693Bd0Mb
G5tDkJDeWXWUBEmvgvDeInoHh1XJA+9xoSErPYjjFKvULJe4MGIKM46KAFX5H0TEoH4jx2D/1GdY
q3hSnB948Sm/ST2RAckOHjfamM6cdHqJqoYEuwAXkyN3nzy58U5gFAvLGV4nwwO2vA8bXWzdFFVW
ai32WERl/b3hFTbc8OcEal3G+7JsHC4BKYIVUWrxJSZVN2CENKJi0LkSeIPIsQSPIlt0l1EAi5qA
krqLWXkmo5LuYJ+3onYyxeIe6v96IN8AyYcdTto69mx8Z0uQLuLAjgVZJ/EgQJLE65i2xDoNjV8l
iaRwzj06D959Z7J+WlgDbY8pBKIMSAQHKk1hHCmmcMpnnZ8McfDZpZbQR/ukr2kwx8nwSvwkpxuu
PGO3r7ljRue7iPSiG80ahAP2GUHpIJaSivRL3V9kLQHc1HMQICd/ZFz8Aa9IGLt5XeE95rS8IqN5
yUA9Wf51Nn5RqfJQ9gYyOAA+MPlPpf3tuPQbxWI3ZJjOHD5l6iWJgxDqrfTOrmebeMluI1Ez1nOW
V2jjjE8aYx95zTRm6tcnO+T6GyvIijZ5TXf8MaVioNQE+r/f1DPgXeB5KtT5QxrygZSp5BRFQzvm
5qCx508NQcawA8bJkW8PaZxmeoRJuw3Ti6k6xUdy8fLcwOdHdrtAuwO+beujUzzsj9MTzLotimkk
Oe5hFPW5teaG16fq8Ofc3rHXtsowHNss5wHuqCGNuTzV/mZDUM5mTq47v23Uo7MuozTpuO88+jop
LqKmw2JpLP4z0s8CYX5XLmz09MYG5ItQzgGj9Gf+zrh1EBHxz1dwSA1nZxiqpfZD9uFbL/bI3sXt
Fn9he3EA+WNRJA41b09qhE00090RftH71l0zQq1aV6o1idvHM30vVljc2y+l019sARJRMqPhosyj
E94dMadja9HlPdEMtSRgFOh28b8H8TP3QJ1TQr5UgP+5CCwcGpt3qimpaFyJ/9RYHOWVUA1P/gTc
Qtk/DZKjEYFvUn92rtByBg7bulrYhyEyW3p44bfQM3w2ZotCwv55b8XYsg/KKCvlLdqY6cfydnBL
aNIfjN0fi6vcQNNLCGAdx3WcL7L5iv3x3br5qxPRPak7PB8AU1VHbuBBpWnGdRLN6dEuLkoIcUMh
b/lRJh1d/xbSTAmq4/2UTL1ezzl8sXyfLxuURnn9sMvmkS6mdEtVcJCXiJ5vD9hIqqidDmioc3GY
4SfdAhDIiV/QBYFxqUuA7soMJtAF1Rl6xkzTIUffN0Tf1ouJfedruBpCBJ6XHQ59iufZ2Y6K+Luc
s1PXSj8tWHyssbaeKkWkLw5TO/v4xV3yC1BhWMtLCfM/vEnXLt/ZXrMEBPuBwLJeaJZdwV5+DyMH
0TLfHIJ+wf4LRiFI533D/GUydX6TRWQ+k6vLbos2WEqYQ7JIXzPs5OJvSHFie52OeltpHLXGz/9L
9CC8YBE9qkjNg1G9J27CiZASFh/P3+/3+4ti5APhvUvNvBhB7avzkY4z1AXN1zvQvQBXLWd7S6sn
7SMt1QEhfCQLAgARsqU5wdeH9cpoXK+rMc5H55w+S9OL6yhbd4Ndxlfsj4p0JDu8L696MWio86rX
w/IbIO3exTRj5FEA6cfjZUaCqf5GXQdlFjoZheK2jSQHnQbNeJrYBOFYyI3MGJJsae3beAmlad0r
X5Niwd1OMtaU84E9T8vYfkM7z7D5MgxOYdmFESPnHB0BJJ1y9SoEBhJlrzr00ua01vYN0o8NANZF
SIVEp/Dllv1uHd3VA2aJ6SWG63J3oBBEOBSjSgvg+VInK+SONkrh8qcHTmIFtjmi0rQBz4ZVALUC
X0WO5cz0BjgaWczKSTkkxgluNP+MCUS6yY0LKsycibshGPu29jtPSbVH+6sq7tbNCban54cqSIqS
BAUStHqDBpBaXGh7hYtD7taC9/l2WlXL0ORr9jK50r18vKVdpwo+5zDvDuYglI4E/CDtzKERzv/5
bIess6KbzQoDlZ19et9DyqDngB4A6rGdLY3KVH08Kr/oQXbU3s4/AsUB0qRhbqHgbUAUUVFlwUZ/
G9RZ26YMr6FgnPcGbet6Y9jiSzMG5B/fJrw+V4Dv+kVvDQFW5nY8fSBKPoQNLcTePw/DOsZVnUwl
HqGZ0yMwtv/20jlL2DZgWt9ZFqtYWdgxCUMl+6eoD7D2pW4o0ayOyRmGEA6oKFXFXiYjZMj3Q4cp
HTowHLt0UisrihO84rKxiq0eYh4EC9yml0DiLgyshJjGrouDmosv2D9eSEsUhX18Bm8BQvnQ9k+h
2X1Uua/SYZhJMjgi7slRH7HsclBC4hbDi+LRpi30EYh28pEgliRa/4MN/UvaZcu8x6BlbJHNOzp1
sK9dt6STB63PNgb9r1JyPVK1yyxilEhh1AZ7ZlAJfBa+U8npBrxgScNVaI8pO+fj0/YDSMT4SW41
8F7uhQeu638/PfF9XQFcA605l3JBlkfzTie9lNfAHgB7+KxY+XSzqb6hGI0PSHriBdO5MyvvF69w
v7ZQZpfCg568YmmyqIQDokMR4OqsngdUBz03RbD1XBpnWZE2UpZcolEykhUqaOp/Nk8FHKDSFPay
PA5LtfFpod6xAWMb0Fb/A6Xo+M4cPM+0nJ/fKdxibad+32uHVkbgd2V8P5ulwqdJ+8bOuszhqBLm
iXFnbZumBDTsNDQ8gFpQp+un0puYp82cttY5Vbzxwoq3rPn3zt8G7848O+4+lfNxRONhA1AAUyl0
Gh40xTke3O0ShOtA2OEoAQZtaTECRY3hbX9eNlwHehLKM5NeseroE6lQtx9MFFSmHVvGINOyVJvL
swm3mNRMskYkdDF1uVWA0YtFXZ0tRFm7mX6U9e4p8Hf8fxhGsJoCtnpqt3wRdgXB+qo8tVZd1CZ4
JxoTmn1J2LjWL5H7Y+8GIPw+oIrn+TLo9Dyq95p8yfqlSVXXb6vlSPAA9Gy5uIQHbA+tjJtKC9RZ
x/9lq6K2ngXR+vJK3sKoEARBXprFeUOWMHzvA7bT8LlVhgKlQagm4jBDokxxvYJbepOye0qbEegU
xIXuIddwb9MgCSTY5KHe5IP9eo6Wv21fZeLcVXVYcV1hJDznSbi/947/f2hmu9g/d14f1/sUPbCV
EaZkG87IbPuvUyUGcB+fiw8kSw/wjjv82Hjr2spCT/et0J1srpo2acROxuVrHI9mN6l5eoEhnXrC
/MwuFlPbi9wEVzFDRzZcOaLqv/VlV/KJ4iY5IgAaaUYjdb/1LrBETQfi/R5bnCOF1thbRFygwCOe
rbi9gmsrYYILEet1R7e9w+WBBDyRi40ikeV41iq25AJB39nJzniZfWsrXBHxfXpblBaD+5sxCTDn
oBt2ZzbjiSCcsf4GAuv0WU39y453G1vNuETFtf57oAdtrIQ4rxlhBpVMncVLL1LtdN49w2YfZ9Xy
1UfX6vCKRzgk+1Z2479Bt9OvjqTeAbdQ5DcldESu4rnbRRMFXPejKIXR5UOQixti3yrA0cA70XNL
a3fYI7JI9N+RB95XNg155350J1gVRGJihyU9D9UfHRlLAMvMru4mshwEsFgqlDEBaR+HY50MYbqL
adiwD+GcE1nF6rnRHN+fr1egANQdrzJMEcVvvBCwejMDLnusS5fosKArKkY+ULSmh8Jo/YknaaIx
rtn1inEld4C3dccw9APMMJPqfTrc/UeUFnodi4JHV9BNOXgVt8J03bFWrCsxa4FbW3lLYBUoBw8Q
wxrads9MvYx/XBKvoqA2ww/Zuk1I+Iz8fsPBz/WRjPpHu7IENxZixjnnvpFyMQjpdIFmoMPhMet6
BJIzNwkapVa3QBKK0ijXb4D6EJAQPQQLiBTYz1Z8CurS86VSEDSP7Hf+sjunX2K9YO60OfdlgJHI
WS8s2Xf69CDQtbqxYoFu9cAZA3ikCx12rjw5Y5eL1wB8y0q+qPr53Jv7VUiC3CNgk0rgZVCS4VrV
FogrMOY6nNixLjk10SbALyhMAh0BA9ooUk9bhZaBHNq04ACtQqo4OJKu2khO0OMAsKUeIT76dA46
y1U+1J0EhUQHl+zPLpkVpmSmQTo+gQTxSPlglosOy+7C7loQISkfPPVuP9ntD1RxVPOCzlPhhxE4
EsafMFWM0Idd5ersE1yuJqmgHwWBk/WGURrxV24TSeev+9DIyz/nW/H8LJiDe5EMK3jVzLi8WgMG
x2BlgcqS1UzutIojwTjnqO4D2Fbf2wifNcfzSdcxyilaM2Ue/I8uMDx+93B8NzyWvIs8G9UQWzvY
Vq9WzVA3rPyP4gfom9kpffYMQPUEqk2wZpqFxLBw1igQZGCw6UZBNX7rCJqkWl8bIxjNsZchVkSK
8JD1EdkM8RNgv0b0CanopO3MvfFiQGkyJGbkBCPkBAhlS0bgMl/PP1zma2bmRKOSKsTyuNpiQ+rt
GvWWBxVjRN9K9Q/ZmU6/RzSlWR03uzMuuMPK++sA+ldgoEE6tQ6aiy262uI62jcMh8+rU1Q+L97X
mF/ikWa/Rljcy1TxV4Lp/VbGui6XF8Si1qbyO+WpXDQdJz8vplOt611tqRO2usf5HrzjImDjTpwI
NLnNobWpDSbvkvvLIQr1P8eHExr3HRZ1hzSLVapSDjlcvh/pSNWiQ+51N6QeA9zAZt7vJTTZs6uT
NB7sehETdzmnJvn3jBa/H0Dc2rzACaiorSJ7m8exKoDXIUL88lNwE9BJW+6gXZQIz3uUFi85nRA+
vqSpX993KP5CkEG/SaEd7FrzszZ7vS+6LCxglm2B2ehY2BFuSZEpc5wSZB21+CAk/J1/iq1hdwVM
B+wyB0C1lB5lMkCosIcBYJUckq5YJQ5F6uCMjG7Pgs3KaGIUUfx4tRAIkXghtii0l6+HYWIa8Qwr
nLopywcpG8KI2qQ5Clv6VSlxDwJpNzk5jLKgVoaID7qCbrg2uGyTs5/eIWkMl49Vmu3HhDcoB3v5
/rtMK0rifPnf4eEtngpifK/gwL4tYR2/ZS9Htmm8V0fTULRlfK9ATlQCh+vmkfpF9wBXkW3mV8bO
oECCZtKy8TJzXa9yqZvzg2D+JQaBG0/0mX3CfwgFvUx68wXLPHqw0zLEYFqtzigpqOmqo0HiREf7
JQqukJjSYLOvdZPbU7zR6xn7Ewsnpb19FINpUbMAifNHjRkllbZIDzjLbUDyzq4zZeqt9aprr2zY
Vt09VLPN+ihycgRDpxOSzsDRoYNivilyWgxIDIhyH0g2EaIBuoK4i8Use6krKWEpVbRwPu8eLrzT
vICwHoIJDmQtX+b4bA+sGhl/CedsKq4Sh7uWb9NSf/ZagD1sHqmIN7wJylNRcM01K0hc958bLVPA
LsVLh6k8hVZMU+FabOBJaQJxqcjfYFfgONk4hAMGNLI6xpuE8LBMbrdbMkHHLy9iMba6AVVC5N+f
T0vn38C8+fGWDpk1ovStfYhC2diAVh/9yrlZyMazWLyANfiAIf2v5ZHxFzyYrqKgcL64UfWROuYa
SjcOl/tMrHX70sJnC3eg05Bh4Xl2uOq5IYmwYVVDcHoMeRhd4flSPw1VJPZMwkNeYbPAuGjy20Ax
JZpZJnnY7oNDTOW0rIOkOaP4duvsLb9UPJuPkwkj2zq9x4tWVRM+ZvkisKj3qf0G30cjLuUH6gWJ
bAW685sd1eC6xpfrHD+vsuNJjPv8r9zvffy9tM/+gt+5IBeHlh1oMZm+r2DKhV9eMz1Pedb2WQvJ
nZsrWiVtE+zTn24NqMS3H3Q5J6Bev6poP/rruPz2/D+TNwl0+VZwPe/5ItTMYK7P1gR5Oy/THfc5
psAPGX9Y1M9beqX+6BzHIyjEOddApQIar0fyYTMD8s4HIavTW9hSHU4qbXMixvb2SMPddDugjoGQ
f7YtXZVnkQdRqBiIHW7nWeWtOKShhG9ypFjrz/BjAtWk0z9sTCySzn9QuXmK0bRMkEhB0rHT0Faq
rsS6XxIRGNnMob7dwwMyTreyZHzizY2ud05FQN3WTtnk1sH98Xo3DTRGnnwkFM9dG1BmOyMg55Ad
5je7VycmQP7P2dDZCgQz9EcB8n+aXK98vvVKxyHZpr+WuMbwNKy/PnjtzQMPHDynAThCpU8x9v0h
ctMt8GdLGLGN4Q1V9l9OY3aVF2YOcBo6Kt0lNi4kuuz6grMmNiz+aJhjLRDp6JgiFSS9sw3eT6MO
TrpePWa8wHXXYYaOtshxm/i0SSLi9j/V3MWtO6/3jXzNwf8u1m/eItlBaHfRfBQ7OL242pEYXgFL
i1+W5HdWvjC5Ix1NdOLUgz/Eje72pN68YMLb9BpyMUdt4uQ2IYbqDORbkZ9p+sRc5SrdYukZG1o+
6jgslEwP0jelG8jEBkRdOHnr0lw5ja7qcpLbl2g1xVeg5e2IJEYdCUwZVYZLd2lSBcKMVdbWJ15T
w2zeV9dllTPA+sj//g8Ack5wPH+YwVuCNUrLurnmqvj14PlvW5lK/heFUdnk9EROzjxAeZ0JHLUj
9wd5VUknCDvLmeNPbtT8IE+bR06eOzo9wdBQeGeHmEHNasf85a/cgkGkbOf7mrZPLMg/HK/mWbfu
4lgNdlFRMQN51j3KLoO6okDbYKDi0wB7PuLExPZA/I55GLXwWGMK8jkHgoGOQpg0U32HgrogxDqD
WCSI3Tn8/IofZt4hQbRRwEUMsdsnrHQ1xlsnNC28+EfLLit85kMaix2keXJmqCGoQI2UD6OnN0S4
iYqQOutpfgOXJGiIELiALJgl0o0mfggEHyeJaHlvRERqRFMEj1euSQ0K+gAt+nEcQXEIZnsAIS1T
5kVpr1opKxpHh68ChhwC2mNomAyjHHXQ5pAtlxUr1HmtlpHELB8uxUVUchxDKFBweCvN6cIDPjJF
8YlSiwMwMBZScgWCljcDzUEsyu6tk4VeCqvgDEHpQjTpjGJo7EmPB+/K9DqKbK/oWwJTpbwm40oV
OloCdW+0i1EiV6ZtnhIc2vCkWmgTXorhtrSlNsmQ2tp+nVEO9isyhsNvDIOiru7Da+tuT7Yy7p3Z
mzCtvuEev8CmEv+kezh2zCfOEKaLtDurY9HDV0WI76hMpBtqTv9oeEodziswIj1jjJIrMa0qA2HE
8pmbUjo5yAnONSOfpejinXDwui7XqjBC9foyRDHsNYVAFbcz3KAYjZn5Y212sRORbtXps8MRu/aP
m9Z8SZTCawzlaqSEoS6/kH13ttXUHaMmxYAb9FsQGJo8sLNBG8VJPO/4dJlhZ2dnajm4HvbzHLlG
ODAy6anHVAsB+pD38V2FO6n2lInPVLVNEkQwmwMIEetP5NpNElflD+f28n1heSsgJcV3/LvyssGe
w+BrQBOtRWl0lULUAjgFZfEu+E2etJwmNNmjbJGfaLNT8oMsVgzkScwE6RC8sYoO3Ih1wqd9yTIp
ESZBvDZ9DyXuD6bwduSed6wcJeyk4lt7a5EVc+2OyJPOIQxURR4CMEH2XbTkP/uWlauecX00xI8z
APyvfg5VhE1BRNUWii6h8LVBNAYDK0quJOXzz5c5JEPD+bhPI6+MzaihwIuGjksDrHbR+OCIB+J7
15/xSopCpBTI9iWX7m+0YgkObZDalnZeIwiHfkHnk/DGu8TwT9jAJD0YI1e7VIgkI+u2XGoMkhy2
4nU/Isq4vBzrc7ot1H3wuqid29s+/T+cQeHX0mp544v/qnMyQAm/GPRnILE7i4pwlVCNY5b1JsiM
QpHe9drWuqDR7RUb5Sm/cqzTuk2Dx4PuSvNIJyElrfw0DqXjE0GwF/ET3ohLyPsXjllcetSnHvn2
kviHv05HJUIG8r/jDdzV3panFClbxcHR4XxknibpIj52dwB6HCG+y0MisSBQgrKPduS7f1aVS0D7
J1LaCF0w7th4DYLBAcXlY4Kw/N0QrM8YseeqUlowCTECbbuizP/ruurWFJUFWN/ncrJsYJBQ3u+d
fYzZFU+MHPSmPCy54N4jZHHD9QDdRXd5fy6/JgG7RZ9QzgDjygSukOziyp31OB+MZ2s3b3l3sQOD
gfKb3KCCzHNxFg+kPubruZOSLAkCdCQ6PfPi1bYYEbeQ/Y0vttdNr1WoJQi9XRCYZ36QgukCmZ8Y
en527DvHPB85MZHZiF73OwRypUAPqHiJmeIqQC4wemORy8w0DtiLL1yhN6SRDQoDCEp18xM1tKPT
MbrT9Mf1+ZL88g3NKEDGSlBcxb1gT/C2oL2O9W8hDttv/FVYuiHjWlxbolok8rYdrkAqwY1AdEHH
SUY7ftIJ9/ALvhYG+LOR4GK1NYLayaOP3Ypi7pKJQCJ0OwXgvA5Hzzz0YRkgLNOrBgrgNG6ciHpK
562jZUwkquVPRYUhb55Ay+iiOaCRo3FhDptczkVDNPrH6oMea2Nc0bBOw+QS6PSqJl6B4nDHrw8I
l9hfK/LxUlW6dlw7yJ5XJac/KIwrtMX1nW0Ky5kPfaubNyIfzBzwu8b4BQPDLzhgNQDu9GeyIOxZ
AgqY5ne2xobc0+40mbi9VxfDAuRTKIoN6Xa0FWUC1X6tcDAXZXlRfr6ITZpVrp76InPGP5LCV1f5
RH5ks/bzSifjPY0v/TuCz56A8gFhJ062/bLE2/DX7Z/vMLMj1zBvyDbliuyokoP9FnzLWYE2Fq0Y
HJ1H9I0iUDCm8ln2mBnxDKPw7NDLUT8S+k2OANrFftHZQS84nzbx0RxkpGiJCcqj3NxYyb0w3jsV
6BSPF7qFQmAsbfxjhPE1mtaydu5+ukRweeLUipz66MolVbX/QFW3IZEPjoWtaeRib4CII8/Z8HYL
NoHsbjIDJVW3KSCrevcULV04jlQ6BF+FXKQQLvZ3MjOBUIOQax9sO9S+xi6a/HNxknvKj058zCNH
DkH6ZH+ma2zE28ZkdAe20FezlDFN0yu+uZ4626Zmu2RngtVWcxtNXioFdFTaV+8JWE3W6jiiUS7L
astqRdiyd+Yu/ZC/Qs4dGCLYb0cspZ6NeFIrtikyhthIdRJp7LbPF4iR44d1ooQxlY4H0NbNMahV
LwW69sZy3n4UN/6OpsxlI4ahWlvS0q3gjNLucafjAc9bPRhRR4/YZUe7CGjISU6/GU1KzQCxKq3H
aWquOt9yMQ/XU8evmEH6FzxwJ9eZLAZw/NbK0UQoDObcDN848YTFFn9sKvrv6Qml+p9p0xJL8gGG
82+eOf2SZN5Oe5kLecQJnkabnrI8RnGz1KsV/iZoxpL+4RvAgDW8e4TKTPUcu2LZGeSah5HxTY46
0dONVRjs39kNmr68UWlq+Um3kVwZv0/jsBFerBk+y1JITcjJ9OOKtaS5NABbEiqiJaXksEXJnANW
7vE0J7KXsnslBMAdQ4AFVb7NHcclT1mbAFDWkGM0xFT5EpN8A1Kv9Ne9Yk0D6MwDy/Hl4ACAgSHI
NTiu4kPYPLNVq7hg6nlUSWvomYvcTXvQh3DUbtgdPcL2OB7eV+wukyJN0+Z75MTT6w8dfdh3dFKu
/kssZCuTw+puusgIZ90lF0wAS4v+oD9DUcNbc4nx1QhrGA01E0vDacNMMheLdclpYiCs8slh+Gig
xTWDKcW1+HMzd58wZBjM5AJgm882NEMdbqPpI0CfykUGAi0+6AYwDXgmXAYpjS3/YfI7VKuXqMMX
j8l9NBxz9n5ZkIwWIXSM7J8Bjxwv+1oIXPtpbPTAnre1vamC2z8n5FKBsrarBNcvYYdYZ+BaSOnf
3bL1wCDFF+bcm4nnO4vAaf/cEdp+YFXwwBSxN+jGFE3zQvhvdOsC9HQ7w7MgNq1jAf85JmPgvAV4
r+LQtsduuTuXfN5QSqamZ80OOaaHR6X/2s7w6HKCLsws4BxJ+7QoJU2gJ2r6Z8+Cr5EzLHEhjosb
vtx1XGM/BarVBcjk1fJnWRwo6dIrzyYj3yrtk+EP8Ggz2ct6xtFvgCB1VvleJEdc/vKft2hClS55
wfLCwgMPdCYB9ma66jWJN6kI78n8JSpWRh8vkyhczsWdqUH4ylwZMAmd1pI6v0QDMJxF3L6t2rLX
L3FyAMJgULt6v650aZpPlMVyKT6BKynLONRz+bdCQ2+8wYhbce439LXOCzWEsd5+obIefxDdnQZQ
/eTxtjowbNL5Onol1JHGLpn1UbOObAeONyj4NVYYzwG07IZRld6Pr2yt78HkAcGUQTV6yTh9BoWm
33/On/uo5S+px3/r+u0p9iBQFU5+N3I0QR5B2vpmmlQG67mc0tQhGPDuFWAXWGXn4/Ms0tCQi4Nh
b1ONF4PHoTIiRpErSsyLgqZ2dpRGSYuyf39hhoP7F8YX5pMArOYEesCFM2pb4TW5LgF2++3uOQuG
oEi2hp997zpg4AUpiQmxk3l6sVa94FTe6rZC9aJza+fECNJWJOzUCjmDrNaZegRgiu7F01gKadXx
WMceWOAor5fOXMpfK2IDgf7n4ksZlRAuteDxE8ZbOk5QhCWzonfBB/7neN49NKI7w4zAfScOePml
I7nRpUX0GOIRmExZaBfAZMAVFWV/ggHacFvkdD6/joTi/0WIHHuAxAhtrBfOxyg33roAq/7Dpje4
JOKwtGWM/wHzGaIGPDhFUe6H5EryKUtboHgwjGg2LLCcpBYRzLYYk3gTYdc02CDDs6Nwmce18R75
Hi2p+0pFRXHUQqffMCu9wjSlSX3NRxDIr3cUrCWWRhbsnOdJTvn2pAW1m1gzO68EED9R0B1KNZNk
qbaEmSrHlIh7uBfPr6MhnZ1sg7jLL67oDrlCoLNGEuEm8ShAKtXDnFPAR0btl7yqC+MsqpXj4meF
q4lVTmGaC6Fr4qTIzyGPqEM+3pjPJaNCWyLS5rY4AcnYaj2W3vQJdtrSRPY6XzWytecSJ5BtvNd4
sHbieCd7FDgmBUB5eLRq+fAvZt9ThnLjtRE4eIffvmnWVIK13XGCGE1wqzMvo54X4vJgrT2ba2Or
7j9P4LnbsfHyNHFiVmoHJSqJYToSaubC+vf/5Ce0pdNiNssqoqUa1vMx9duEbOK0wMR+NDGhZQ3W
MDBvag8RGO+ABc9JhXVbAwrTfzBkcLkmNbf11dwKiGCzYX5aR4DiYboRznkLDRdDkHpF1aABBvW1
oRLMBckhTSdproJYO3Wa3hUforZWS1xsmqLCay6fyIrTlBrlDDMcaL0z7ZTwfDAueVH33VUO+VBT
eD/2/0DoY458yNGKdU2Horri4sl0fFNIgrBxVoehqaIttAZoISfSevC4UEh1BqGHny0KhdJNA7Ww
2f/OatYD+AkBf0ngDuvdSdBgvK+Vy/kLGTuVXoaoZPvbt+78dJb2fPMNwYXi0wgNH6nLEj74AGtB
LWBhGDoUf3cstC5litk36hyVFQTrQlgunGqNphF7mvo51T+T7SUVBt5hOTEbSOR+ius6jG8vwI0V
WAwlJK6oJJAcJA774DS0GlzQH95c8QAOAJ/lnWigSHJMjjdvs7zOu6ua/4pnU2j3ZYqVqi1Xd2Ca
wlP2MkyE3cVAaSJfYqTaoHwfqPHujJhxBxFOdRN+DzKuv9KOE3lCkHcm5FjvcAv+Q2p2IHHiiwMZ
1q0+LFzeZP1t+7LsDerByc090SHVK6kgUEY5NPSKmlBzkCPSusa51KVkMk/jWfSmzri3ndRPrfz7
MhULgc9OTAdK1QuAnKU07bWsykRbbrvIwBH2/32QKGuCot4fasLLhX+AtxfvJRbzQW4J5cP8bz0l
lTrLXCSLJwUDtELGzIOrVYJmxgNQJHNZHE713/A1u/TzoVJJnHOR1eck3AjZ+0QGotu0ziouqCUY
1gcn0efqqIOhXTH2Xc4EQ0RunopH3DfPMQJB67oA7yK+1Z19DGaHymxSNruJeuLvDs+WghBsKp/h
JyEM6aQmv2Muka/WoUri1ABRnF44T80LbCHkSKmRsJIQX2hIdkDhG8IM9gGizj3YxjhipAFFg+KC
UGc/hcJucBH1tsDhTP7S0nGTFDf8HfMq+E9/JEzuZQ04zOtVWYjmy7wnjhTS9Xe8qkSyppGUefm+
tRYYpOjk64zMu1P8uoRH7mieTUEeUyM7MsY7eClA6d6RH9aJ/P2L/m8SF2o7L/SURZqiRzy05GuC
968+0qr4QjRESma8J1f9gO5S4PtKHiagLbPx+9Okf5CDJyP4ZzZK7uDB5p6S00aJDG3XXzZDMLVu
TmSldOSMckQ52oQzy/o9Ig/CQcLIFFsNjRJDobieBRm7jFbBS7pZ9qzXH7Q5NFnQPdVda7ji7wCO
Cw1ccibM351R83OdgvxXvVhNCt4Vb0hpy4aa+e9LlHEsR/YStwvcZ4D1J6tuL5gmYQFE1421JIUy
PH0y0BQpOTOOvHXYM7Ex48FwNYXkAemJMLUwpjY1hkXjhMtG5alnDs5ErCRoRkYkGxw/6TDCxSFR
5n5Ge9Z7MshWl4jFY1SYOw/XvPU/BZhoreNLkoznL7VoBRI3paU0G7oeU8ncbGF0B/7IayZoJ2Qd
PIejnHg0imMLaoxwvuxVzvHOsej2YzPYwl6MVdXD+9oCAbIobvN6khZ6SM3jdj1JjCYL7ZpX3UHI
if80MQj0U+0h5IkMzTr0/XKA2J+7yaECkWr7unMNwmip28RBQAMkZatMT3k2LJTY6vAsF8guvxPt
m9rVnlkOVesIMcdPEx5jGE85BZuH9GWKBv9V9/9K7ZYFv5891O20DJEpyji5yyZPNIKB1FeeLgeo
PMi4W+Vew92Aia2NVKNf8TiT7ee4J/EDN2D8LU/0oRzggEybpZ0kd+In/JQHQ45D65z8rQbGBvcb
Jbi86fuAbsuD1ZS8jNFGCRmGJ5vAbR0gxsnlXKQ91Re0Qiq3mVgFcYqJT2ZmdDgZpesRYdD6wBO0
2U3tmmHnz2JGK+9klMcxu1aE0JGtiOTT6b52LbQkLPvisnfhqC9DtGX56FcqS8wvp6zDKwUy6KZK
f7mIZo/aH7wSUanAn3vMQDaxCvgbPTwQDQEmfjErE/D+NXJ5LF5CPzhCMy3fcDQYxQ9CcwrW3kKV
eOmWa/EbOGeg0Qv+peLFLbIVQ/LKJGKwJxy12cBM4Vn309FbWMRJZIDOweo04w4UDGJVZWfUw01k
qooOlAVPj7xwiYoA7osxvikV5FkKTLeSvPUnUHWKQs7sKjV5p5U7fb3rlVfTFnF1mMkg2Dzi9kIi
7yy7LfKjKIWJU5A50fFv0CqhY7vT+DOR4PMIuI+dOO/hrZguPJAVcPLgE4QDTpolyFxIKLD/cp+u
yROgbZe0NeekPCg5L98MlHcEB6T17yzrWTrkvhg6FHUlTOI8i81pFns56ppZOZfShVeBaO27pfjJ
gbGNkTQ97XSnundqqhHKyCahalHxe49iry6/9J/UUdHvltYApYirwoI1KH/m3BQ06CuEhvsEIDbx
8myk6Jki4qWtRu3xGW+keNGkLrlBe6IT/ZBb9HJbh4g9uejfK82eVOGZAsEwuKH7cJ3Mo8Aopszs
gK8ssNYwi0gl5Lp6zAjpuCE7QlpdX9XPOAQZBPHWBnJfqBXpDtUjSxZ4928S9Vcr4Yea0uY5P2CH
v94Dqcg6ixvI/G6fR/98kyAvy2dhTcxmGYyu3ebuASccQlDuzb9EP9URxPGhvE9Keac030dMepfQ
uiNPyGzJw7LFFAqeHsixxG/35FDdtayMHBCFbH3+aiRFXYGIQe8JW7KXsiewkulrtiuGZ+UUFqrN
xO4YX1WpsPtCc4u7+hAVgsSkkMPT2xAyG8W227pZ1sNpl6nyzT9G59Lh0T1l8ALmpdt6WtwYahUT
5BNcTnKGCIp/a8tIy/lXSimhppsuunubCMSohTCeE1jDXGeipmq75rExvq/cTgI6aN3bnhcqs0nl
mwuQQ1urTR3q467mhWl5X2JW1uEDHRe83h6Ezx86/E9Fl5o3ji2fLbceRj49UEOFRfqdjmosm939
DlQQ+kOTmzfksqFa8Uw03K66Xvn6ieT+P9L5FQkg0YYZUPQnUQ7HJVdGQosvhUvS2H0MuK4awHy8
Wpo9lfdJ/FuU1axRKEiry2TScQHkU7ir5LbyWEoosJq1P/Q9qHAaI3bcwC/bQ7Wck6Vco1yR1pNj
xmarMHWDWci3CWPUDOdjZmDtv6HsPvzZXhxGwZkI4dMQJrpmqY1AkgYR+7X3LnKu1EiJm6rPdzL+
eVn/1fbdwbMqJZeCrrNi/mEduQwcZkhjNSHZG4LPrQcxByw2fNlr1XQlL7KO6Y9ildWcfyxLFJN1
x4D8I9pVz7VNLyy/+NMLjJhmrKjkt5R/HrEHisJv8aj0cW+jjNjIuPNxGSZJEQbeAm94L2fl5wvT
hQ/XyhFkRk3wF7y4Q4BG5YUYoLoV0ZeqOEGDuq9tQw1Y27+Y0itQzaTSzw7BOrAfbPZt+xbHJKnl
zd7Qc5k6XgtkTAlWqIzdwOzqFc9NXWp5ubrn7mwSazOSZaFlrL87uiQkKXUmpNskxwuYUCim8YN1
zo0CAWxzXzFA2yeKOGIYCE+82mV+o18/45idYxkvaHo9bw7CXaNXVnE8xYfPcP7ij2duAjzwEczM
xVR0yNHNQ0uaY1W7KZiTJXmpQaPJAyisAurM7tFrpbmtSdSCUblKZq2ZrhcEMOgFdb9Xp7EyiqzH
ri6eGHlLG4/LKD1/OXKnArCTY7h92lvQ/OzefmhVweHLW9YGA0MD3SNDVg/yQl17eFViLqGXupct
B7UoNGtVtNDEkLUul2oZw2PhwcmcTA9ggNzOY0zxlbITrgMSxL1HV++4S/yfb+6aXvSzsZv7HTpl
zzmRUMwt8uH4tgFEgz/08wbKSWL4EJkiLmppKBWPbDqOvW7CGiREy5rm7N18PL3mK0Ejg9gcT119
G/mn8qx4lAstKUK9UaOPQiezQRBiY/BpGAjyN77EtNmK5PdpCWBmx4jfpzhApEO0YOlSItNZfiw1
mXpuSWjb3i/yD3UXFxhWHfS6aozXX7vlIpQCFqPSFkpHLJfZoXc5ITRF/0Tvs05mnnb8mog4nzdW
T+sF4ou7aZFk6gVcmrFiSwXbeuDIWX75nPcFdXIm5cKsNLnjCcYrHyIls3AHZptfjvurdQ7YyQvt
lbQeHTNBZYrMo+GHFx9OIy9TsYjALmL/MuebCwOHVlluOVYqQTATrUpPMmqbksHM/ViMhYJhcY9e
QK1fc1e5sfyiUyYsJK+RQUU3zCdRWDHmTzdecb9odLBCltKO7siEClxZnK62IoR/KSEMKbwopg5X
2bNRjydUYmtAiJXLDm4FDQ73EDPCocVIajdgQ9Xk4ZQNCk1VBfOKlrDmsWRYa3Rvv3DvWNpOitYe
h98YkcrPj3Krex62dPZ3mp4HE8CCVgROWQX1qIQUjHK/o/YdyBq3sz7NpoABgzxIK9Z6PEFI+8C2
ABAdKwoE5/5E1MNVmOmdfMVqv1wRpcIBCSFqaNskm6LDDvKJ092nk2mYSJsVr9yFndqetkjM5tF/
O9MpgMuXiHIJ/bh/xdEi94yER/4CM+WuzDlqwfyvM3CASKYQMeWkNL2FmDUxlFsfQqZ951uWo3Vl
R17IKEt1y5eNaxFJbi20o8yfbvEwIG5/ITOpCz2Vtl82GVFi/dm1ZWeXzgJ5T4Ee/TqrBjKIgBfp
mHkWBJ1cuAAnof/TOsUyTiQ1fEg6enwbZqBmdJD0bW6icRIHFA72RryMk3IgeZNpmX1ui6LrGJLD
v62/vijPOPY5bFMilWm5E3AoAO5DowoOJ4vRP1Jkag8rG4813KC3oREkfSi7nrZ8zkDdXVC8+jmi
czea0CaMQdd3oIHLBpsALe8IUW7mOxQbtnY7zTaXxmzCDjEe1sS+5BH2T1af52EJBmljhpq3wqL9
zphKtv5yUfYnzWVFeCNV0erDJd8Tf8gRSQD0fEtIjKERlPV/4igQu7IqQ/wNAlOB+ZgTwFhShEXl
RXK4hxReIIIWYCp2r6t7/gwZe5rAxaC3OZ1XcNLkBNA86j1aAmfrj+TKeSp2VkdkeBinpEtviYAd
A4aBgH97p/etv62HSy/7KRXEFBTWMAC/cHUQA5Y1yxY102eSLSrHOo4wtDKIE/Q7+Yk0FUFPfQDr
yshppaGLT0BYVrGhLlbubHS4fQrd+gie88jwFa4U3TrCRrzCq8QMKg95wp8KPAH0Dhr43stBZZWx
Bnb6WBmr53Kd+gK6J9tYWm3MC8DgCjMfQkoSxDJ3Zp8HN9K5rm0g8kGCwgVLDfP7WbWAcuwmZlS6
o3pWHbg2sY1GZmWf3ZQjT3XK8CNeBXRnjaSn04NN0ALytu1tvPN+NSyE4OMeXPtJJ2034Mx8LU8K
8/ZV3X5VHlsT+u0p6UCY7BiIM/yUBvcpOc1TJdd8/JgHPDoL+Kjr5rlIgiYRCWnxKCHhlspjWph7
PtN6GL1yYu6m8fNYMiANxO8xw26TXpbWFSsxgHyupkLNu8ETiDtwUparyCri453AlFE6KdZhPHHq
TJwmCJzJv0Tgdy+u8EHIuOyc5QjSELr/sZ2S0EMhZc9iOzJYRdmLf3EW8ymLcSTGeRYRpPfTSjXD
mQpsbLSReGbasMwk6ilybRqBhU1zQa6fKD9JiNHLeNQliyW6//JLvpzboaQcT9yZZXKgyK8shdfU
0DGt/Idm503ARfCmKi1e4gFJSxwXiC4znEdMb4OMCk4WwVrkEUtKO9TgItpPCLuBfsk7rNHR+Jas
nhLVPHBIaEM824MqYTLe2HFnLUlRGqbt9PvcWBU9Cfm9M30ysqXnnYj0MvXpbdkmzFC5nmm7s0AG
I+P0rW9F21C/+aA/olfhdaipfpsENNgSlHtvTxuUTiaF/KMC4Bl45L+wqGn24koLriktB3PPg5KX
VyYcP/q29klfu4coBUigP4yZEI2s1d2u2jR7AB99B2ecGA+gpwE1kWb9oV2mHvXpT3SoW7kPrOC5
q08BlfNczEzJ1tSoC0i7toz9gXwluWc6lseGtZsDpoYRWpkAuCscMl+JBI0cinAi1CtkykAOVtYQ
OR3Fn6Sjsx8W4+N592TEPuD/uj5BEz9bHAD2WcjZS1qVEhBjWfbMTTE573av4ES7aeiOIAn461mK
VTteA+Dgkd0Qdb0uvBf1qvdTjA7Ang9qc0FJetgHTn4deudeV1QHtuoDw13sPDLJLW6Jq9mF4u+j
0coZOn81WTtd604z+bPnU8bCgjbH+mdY/JuhyNcIPA6XiuQfxxbNR8+JHojOaDpJDNQIJlO84zrB
lAK2J5Ute8Jqt4uLdh9XWeesWHUppDfLSSfo6udtYwgTHP+eptAEIjkpnulo2cpgLd/bh3MyNa02
mEuSA49kARj/8PrqnCqgCr7KBdjeYpxU9fkfcDkVKJfLB88G9aLefTo9fo1LoLD8gJPI+fAZW6Nm
jenE9yhwh0iY7Sc4tTOJ8QSmSu/XD6D60F64OpGbDeJPd85pnnOQzQ4seOMF6sroG2LzwHYY7qjU
yCpL3IpUT+DnAswCM4xENMeNEa025n+HhVBR6OkwZBucw3FOXigNnFgaWJfOtvKFq81hbY/4FjvS
2WSr8f3DfOh6pJksmmrTTQW0mOep+kx4wiyDLnRvtOtQQauwXdbEAYQWFZg5L6Da+WQfcoL/Rgcx
ttvRa21M+9H5i1LvnUT1GlhZvtK1xUVKUYQigA0fbEnkm+q/K6pQdmqf/YNr5uvJpEc3FfOwFaTx
GHPOAoSibpp38ebpLEOTlCYxyvXsfXt2YrhJcm+q9XlRu3Fgv7EyTUB62ni6oYFdnKZcKpjAKhlE
bzeQ12zfA2nR1rEGzcGMdib+0UtGYKzneEK9/3k+1S+uLJz+8cTx7WjvK/ee5XZ7GqV6vdZzpedI
3p1FaWQteQa9vu2sOonRzbHn0AkLGG2G1fzdiEsuvBicaKY5Yo24hNtZGIzJDl1q0BQHsxb2BKC/
nh15TUkojnvQl+tHZsHz94OjSSlKyaEqhn/OSAVZgWf2cyIS5i8bUaRMa6QD2U2yQs1JaZMxavQs
s5doc2DqewZj0VMfVLkkPiiRr775GPpFYa2w1zHPZlo5brM6aNsG5BxAlDTRzL3+r2tlMuIkL8rx
NFeucCUt+p/hkhV98sc6F7WW837RZ7NHnOPtZmceJuyT2+UuDJI1MehcfKHO8IIMW/1KCSwmR7oC
NWacBWMwKvyzE7qcSRCKe6SqNlT/KaTqz9oXhfBgpOQZGRyB2pQPcUnK0TmPY/q9RrxNtJkZJEWb
FI0AXmUaIS8xU5cjNXetcjMBfTZs0qj0k0NQzZFgxYWd9LnsuQXFTEwo1WfDjdmEwtSzHd46CgL7
au2KyXtG4wUBINMoYgzp4RzodIFMwNE6jlk0UN5N969ThwEwgmhzANHzZyb3G4gsCks3d7qNWcdc
7K2kTx0TNhfJmGGcyVXKWTVeY9rNdSGwgem20k3OZforSFc0dt8SZ+bxByGaLoQ04r0It+4Xt40I
nE1by0P4EJiXlvHWCQ306dmuS9OrDFuxrGfinb0RMdR2aIkfKKSVt5jcPMt/ciBft4HVN2VG3B36
cADLA4gZr2etAruc6z5huMaqglH26agKo+LAo9cxmxcSW46YJGZ29mF4Sb0SjFVtMpwIdIYoXgiQ
mwDs88x4yT+7AFAsxks5hpFHCTHqUvz4tSEwiQ8JHPxdTUesW6wM8WreCaovyazgpFiA0za2drxO
pLQqJd9TdeMZLhlW5UNgkDRRWbdQ//itIEMrEpXINSweOM4vdT/9sS9qZO7uAlIDc/nmDVuRvGID
8EGYyuic6cXJj5lCctHDtHzWXXlT42uK32bpvh3RBBuNmNyFgn3brZqSu8GEUr5p8d1+84/MaX51
QoInfZ9DZEZ6pIhfPNp1sbM1QYwaJKxjecEHi03tF13KrmoRWtQTNNvTNm9yYGwa5J/uvjwlxtYQ
lYJiYTRwysajHS0wtNh0xqkT2g0m7unMktmXCSgrgFImGBHhzb+P8yGFSfDf2MPlizDvSwBeAE0i
MJCv2vOp3GP4jm3f74TbMiAfs1GXCuF0mDaPtVRbrhTgK6zaBxYz7F6ma1hzfM+ZTQjFTnX6gDKm
6GUNk20FC10+RK0vLdO/UOY5xM0+ro6gCGFdCXa8xEtnhBwnvS1shLphafj6yy9F3o8iCy94dh7w
TXSuU1fkjYyeiDNnhwsBrlz4B3FFk4PIeC0pbYJ9gGbEWuuZeWlsjYHEGDfL/+G4N3HcthrxfAQG
FmSxrhcm9RAZEMWtr1rsDjKXeqgAWt8H5IgJqHCo9lem7IehgpFNoJlzz58s0oGMlAnGMprX6pMD
dvQvtHqieyRWGp+ca0RwipEfZitp68VZyinVHKMeDF8de10hpE2o3J42LrzaJiExLvEQeT6j8dM1
LGf1/MOLVpWKJit8FhKmDSpHKkQDvrcQW05iMNG7BY9wyZf6MOcHQDO4jaZWO8Vnl47gfgJTTDue
nd3l/470Kif4nVrKsbvToq9doLfo1jAWhgI23o8V/B3lMvZWesv7YKWv7pj0uTVF7rTt6ihFJOfw
povZxGAjMUmt99SUCTkrLRFUiQ0GIM072XY2+iwY3Ndsxlc9sXi+GpQTxXVI7JR71znjUYKid2Iy
OnVOGXjCowz3zQ9jXniSg9XyDLEgJc2hSWlPWGmL6/eno8nDuVi68i0HtmEoPf9iBmmA48E7SX5P
z8xQg2tZu1YY6FxLPrMYjof5aYnURDN+K+p9cHr2tw7FPrJhroq2fmYHMyBhPfmBT7ve7MXPZSin
XxDHPit5dgz9IDMK6TGruYqSFkPvmp70oMp3tI778C3Nnxph0/pOVR3z52I98/0vSFt0C0RcBmKW
6eXW4XmoE5b8OAfdyikT83NjyIPkNHk7zrCGm1fPJqjWaITXY/0KVt1VPnn1IgDKPTod7z8NV3fg
EoVurJjZ8k5QMdWmCE9SF/c3tIjJrrS0taLar2nUpi+SIW0FSEdPZZFI7kUU1rGkuQtB0IRsApGP
tgM1oMQmvuaZJ01u/NTVZCsme9MxApdewcJBo41tUMv9+GDx6q6i1lzO+jJtgP4JBZzFxHBD7/CZ
rrCj7hW3TTHXVR2e1CDKB7dY7+hbsFKdgBrbCv38QUDIbiIoYB5ZBf0Ccje/mNlh/EFb6bguqdWT
W2MYAGyI6vdr6ZKJc1QizuIwo5sYI2zxCkytDzdX64sapNA3zhHBuXeGTWcLxil3smd//sYCKq4N
Kj0oXMZou9uEIaoJu3GySZhML+4pRkNzjGKfa8xjp+uKuGNRera38sZT5dVt4RcbIEuSJoPy+LEW
AZRDnnM1cLq7XR3YNwbLG77RWP+jmzYo8SJSBaabshX3ofuz6HSryPi3G68qA2CEp44J56t/0E2q
LxR08hmnEdk+Bc0iwLyd2bUm+kUWqsFVdUjU2ayn4xxUuzJKMLQOCavV66TN9yU5GeCWaTo9RCza
ncHZ/6QIh1IzFyzSrmIDaIQ5tNTjO1VlOK5TEWtIygwr4K8UD8PRZHz6FUihQCsk8m7eV2p+ScEh
hrO/fB+ZZs6zLCyDevVuzrTCdiZP0Qh5vL3qTtRZlEV71lWz+MRzQe4YSwdPNyK0s0ygK9uMTKOi
8LY0C7QsbfjLvVCMAxZj1m0j2dGeyO6EmcMu1dUvs29EuDlQsTgxoCKs5O6eXGzn+WwRECxSQuGF
A5ULBYdNh8xWvZ7h2awa7cAfb6/rU35a17GOC2sjnvjo/5Gtt7q9cnOieLh3vysthRf0olmvi758
rjMOjrKDntcNYIYvzzg6jUPH8btL3I+uyo5XAkjyrvTat/Vdgw7vSgkAq2+j/Bj975J6KRXcp1pS
RieMLEydsKFbSQrxi9lDXnACRAT6gVhHiNV8RMyyq+Y3ns8bOzSfD9uPO2PzegdjFo97V9TjNDd4
7Oas+0ZZlmI2rtIOokWqVwR0pvUQR1VyEbQVM1QR41JTUunopG+qCe7akv/bWEZhiL8lr0d7hj1l
YJveX5IFFcZwsEDpgRPtY061nOrNE2Ly02ZqjrHTPt9FfywsbnTS55tJBFBg4q9zfOUwQlECGn5F
iPZ8D6pItIuJYq/9hdTJQvalEEjq8cNEZgr0k/YXNQvEPXZX+ZIghO13mNtz0IuRoHWDudi7EjQd
YUjtsqAzhMvryYu3XXbZkK80/Bd6TSv1w231n4KN191XLulhnOFZOySJGGVRWgeEQFpWNMDhCgnz
Oer+J+l5mRYbSQfqghuawgI/2im1Wf5sUnPMoWuBON0si2hV97a1mFQaxsdoyG4urZ1sSojazBBF
uOZwBnEJgkSa72gLIYX8EveGtBWRHT0QHGGCwkriXv8yaiuzH/gHg2/gNW9yJfD1jnuUz49DKPSV
WMDLsumXDLM/Cs2fJMrQK9FNM/M0uNCrBwCAPBlSFvxwZhlM8dBlj9X9Oy9M7MVc/4JB2uavqDx0
auwr1Lvphvp3qFXw4+GzRIGewgOZqcnUKDJm76M/B3OYyEVSj3FRcIyjdxzIEOmoqvgTvXvNDq0Z
Jv179RXh8b9nakvlmslSQd/1ztBuDHD7zSeqLsQGmcmXSmhqAOCahQeLoXxudmPc7YKjBmyWC2Bk
irb6gCu1kplayu9bTxJWurOXhGdcYxxl+M9PM8SV+DjkQIPzmmiuKRx/qnd6NZ5Aw4655LFycFt/
xZ2aGWki2eB9LBOWlbkDoKY9nYXeVPN/rl/dZIP531uv3tAKmTWfIPlrKzykFKP8/8vMy7oD1tZK
38SZfU4isazVoJrPl3ZE0gvtvsq7yZ4iMNcyf1wWZU5H/Sf5aMIRrt04CISuApVovm8ddeL51ZYy
fT/uMgQW1EHzu8HgbyG8LXsotEku5bD1gLotZx1/Cgk9HiudmHZIsUNDVyHoKxv8TusaiqCfj0im
R6hs7azqSojEien5VQwyjKhLP4/oLDUiRk/wdBYoBlqAMeCHmyTlp/NV2Qegiru/7L/rnqOtB5IA
yFe1poWx4vI5kn7ZOGDks27huMNwYLONQux0OQd8i7QBgYuvAX7lyctH0sGRT83sa8qxClINcWAi
3Yso/maOi25+Ppyd8k9H83MrqLTcxNBDZIIIssrZU4+t5oZu62cqOZmbKpWb/AKuLkUBizOB8aUl
i7tB39TCvuwJcKIIx2KIZf0mPWkuHXtuGbu+Fss9zDCzCwOtONdqB2tIrY+cFDpD1+P9TyaDANje
HxCxEgJKoMc2wNLcyC+l2Qm6jYQUU4H17bmPdRBX3tTwpKVccNPEFz5H9jE97sOU8PVeIS3+A7zQ
1UfPeL0iAzc6LHL/iEmi39Q1Zffr28bv9L4P9zMPocArwISjNDXv/8VtN7lIqCHuOKVUq4DkmUAh
RO9NV4IlHuXMXKXoKHIYKuYfYP5bsEZrXXjRoUbbSphRSr3YzDBfooCCHOi5L7JSi+WQqG0R5tMX
1anl6Y5p4la7KdLdPL8yoE2hBPkmvJbRGwYUq0fCDz66eXMU15sd9qhNCaqIia8BLuNQkzB3zNvF
dxFWfpHRyHIqVKKrTRG6mnkIZfgwIiovsQOV6z1mwoWoDXa2o1n78HvWh0LAYt/A61Om9VeIuul7
ovE1P53oYx7OAv8FIDyLwD7VDGbcgiJtMAwbxD5vTrQj8F+7VJPdN2z3sxyBVG9DPFFeGrw7laWr
pFJwttgT9flVVKV10KkvZ8nvprhti8nSFJfJta5lr9FGV4dIrpbz4NHpRKHM8yV76+IuUUzADhzm
lZJolUKyAJ+eCegQByKf8uKX8TzXScMd8bmiwPzPF+np+zfVMVBljGrOhYSimSdZn66zGwWNIy9w
ae/QKyhgSbFQkGGyFTAjF3h6XjPIlmkP5xxBBtlpN4mg0aOkIaJflqtEtEvZBG4cMWTN30K7eRCY
EVtIY24kfvwYu4JEYOUuyjmz80/VA4WjEmBUV3FwZ6xGbgmbM09EXoj5lzXE7+YUDLtUvcUBCojy
wIcrc3xqFtCLpPoYQoLQbHeLzZ9fnTT8F8MzX6D1JtNFREyePJgeHLXqfQFLcg3oUR+exjkI976N
09619cChsf5BZBcHaeQ/iDsbThxUwPvu9HDU3T4revQQgrCTR7pNrnWR6fUbFRn+ItkWNJ3Uvg9t
Q9fKqyYkJn+1Dfq6h/hj0xFGGtX7RNtDE9hclrmmHJ9U+0wW0wKJEdGhpx7yBabTZKLSZUrescoA
VKI16NEivKEaAVQdjm+dFIHjNhQ+9Lss83ILReVrDuIf3dob1tKYWBD9qCpFrvDhO1MoAVuANcD8
zvR7XhdnhOD5ynYRIGi7iAOaChAGE/MvYeoo9gdrNbjj8FPzV2ejzypnGlcsj0I4pI8KTFV6JIU2
ZTAmm633QrnKiFgOJcHZPjuPbWnmI5gRWgXltMN2dzKWwLaB6oMgtAosSOlDK6CZcpb+Ww86tuXx
uWA00Fyn+lrXqSCwpBllp3svC1vXlExFX8I0txtf+3TCTFJWja+juyMCPHnjkci3OZxZRuLnGQU0
+gPU5odEbrFXwuiD7SS+YuKpHERqTD+qi6I1hhbFdpQl0oB0gocVE97uW8p9FCDuQ2J0h9Z2zd9J
dpqW+ZqDoXsuR5CPQS7g4s14aSEYpYWPWG4zcepbK6Z3krVBNUXshtwgCdjaGn9L4KLS/xfWR8/L
P2UyJ0ZLSX121ZNxNe1Ql8wNLvo1dhQwuTqQlAY9ynG0ZXbKYNOC0MU9tc9C+K8CzOdGF+lmLopH
08V/O9xx605VJt7GUXplAIk12Zr9IPwePiaEnDloykvGyRt6xX9C4dz0zzCN6FQSpI7jYyx0CKQI
Kxwopk0Of8KXHC2bymGf06ymy+Jb1e3OKPLM2Tlcmb7RVsWGcbVH212rv/9g3nRkCzwK0vmOzlKG
b41CfZzqirF6weMDKSzVF+061F7+xeQb4U4SG5JlrXWZ9LonbVAth1R/Vd2k9MF0wSLBpMWVrV7f
d/PEtp8+jsSpGLCSMCTzfWp4tIR/OP2x3TXfgLoPspoJxeKaY+atYy1sLHnLQ2R654xSVCKdMCA3
bHErnqRYbt5VHwnyc+rfU+C617fSDJsU+NzdPlDrdz7FxrFFDVyuEDW78Dg3qOOoLt4KxnCrphTp
TgI2jKF6tSFoxO57JhgZzCthUtJUYXfor8wwDp//wd5wFKCoHzJgCUzu8Nz5FWYx9TYxKZmS3trT
yQ9Xjr6gdQdH2mecTdqHpD/JIkqkC2tRgwfYDQpaegCfgLVEJnjPGYZARD8OowGz9syViT8sER2q
x3l3rmtS09vCmk9vKds4YoZxa8idqU4mlmplbS8wYuQlFvNkRwhNKe9K7DUS6rHHLctCMnPRAqKq
vVcb2u+HjnVq5Ha2QIrUWZN4b9XvYsnvoBKGJIK0MWz0s/CV6Yf10yE679zyxks0r7cK2Ks7W8BP
CY0J27yEprkcuuPyErwALTQHH5nyrjonWbzdbrmwvD0t/bxQUvtaUPZ59ks5nDQ0icP4Qv7F1hVu
F3V/WUabjb1gulWDAd87TU8wk2hMqo5ggGgZHSMJ0w/RpNXQn1xyXVkQx1XfuZvAOS2mqznVEgpa
HPG8uLxfvYbrEhIJ0+pnhy0iDnP/qcIK9/Pw1rLUoLKkk1oiLh5pmzxmsTpt/UomDAA9XfPNnPLp
hDRv7G+xCb525utyv1uIjBK2T3NTqgU4w0txBTUa/LBHpvpfXQjYBxrzYKZ/VMPIod3moq3jy/tN
nQCzAOLYfIiNscKOQPYGu0nBEKjprC/wA7LY34dSv9OcABMpGAh52DsV87oaWHs/gmETOoFsbK/o
PuhIEF8ZYYhSMA2HAMnhi0MN1vncflLHQwIx2GJvKwvXYa2B4JMsjkfM6qYfypHMsnuydKlXAWvQ
BrwwbQzs6NQGNKN9xeJO743fwwcMcM52vahnRkLWTa3powfDa+9juNStwqAUohsHVq7j/qPk8z6T
9Tb5zeuy0O6B4DtunCVMdiJzqTWREDvlk4ti9qmJvOFdkP8u9Ju+EHOXT8IS6Z4k/eLWl2Q2s8qv
gtKtjSSoULQH9w0yOVccFBRcy8ad6u7cvMORV0t5QNSF37LldCwvLvGXhRrZMi6Yqj+ldbWR9ImV
RdBL8sdXvAm4/LyeXA00aNaTIG/eiKXyF+ZXZuNzB3eDHDIsOPci8jjZARPr9m1N0zQbgBkQoAAT
3u9u+DqZK3kgTqzhF21hCeqatdWZq182qhB07HFE3HOWc9/S0lJ+ocXdwqIDQHSZF7f7pm7lOgPc
dxi7g8VvnoS7+mJWQiyVkspXEEqxV7dNHKLW1vhFG+v6Dubh9UkrlcnTOpAVXHDfk80p3EE7D/pZ
xlkqoqEoaGJxP9d79xebenoT8owqyBaTFj97Bi9lJ9QN2xuoPeGBnSP2HLZGw6ehDm1zzxA3I5wv
XynPs4br/qOg3N8F4J+6HiT3AV4HW/z+zzHYHpOXXXasiaM0/d/C0wlZe9ujpActpwp245NilbdW
Nj3+8Ti/3AUieC1oixAP1lA0xeguFw2hKQtZnCkvaKi2C8+QckL8CsBuloMQ6ZKF+rKlQeAv9tCX
ecclrB40zpYKn5vwcvF9ItytUzSr+nXvwxopLRVSylIVDNh6hIO6P9JZq5shYzhHlaiIM+VheQh9
wVjSVOmttu+cojUIjlC7+l8b5fhKXbF1gK/+i3IhdKOJlGBd1BnPgndpk6qsVFI2ElfWUzAe7oeo
YHvui9Ucadw2HSpRm+8eKQFgrsE0TU+JglxYA05F/zqdXpyhSSSFMThjd1ZAmK751Ujx4VvUuOgH
fHtHYk3Rv4wskoyYKHkgMgQWyyt3H2xT/PH+FZdhZQSgd7Q38wAxILsSJ/MJTUdN09H+w2+9WFVZ
G7Nh7un/KWBvXa9C9Hm3MuJOiwXy2LmYeW3+oHSui2aXU33Wy7cB7uQApdYG95tlfEwpUzwpziXn
rSad9YwKn86SYCdwnm9TgiznR+44l8/QPR1jDaHHHxLGTf6P9ECAG7l4eHkubicaTe5xAVlfbvFn
DdSf92omF7nvwlEZu3Wm+ZABNkvm8yiEm7ZnXOqpdNe8GSQaKReK/A55wiBeVojjj1y9GzijgCYs
CnLAWZk/9a7p96Bq8UAPU0sLHVX9MGgO2kgjzCY2LOdvLoV4/LpNjIunPg3uTYwdScwXnVgjhPBj
dJo3A1dp1zuPl1k1MhuNAmyMOu/ko+esp/6h/rhCqxN7C5pAXFkl4t1qnG8YqODaxO9dquFi4x+N
0e1tS1y2iS9NGBAZeGG9bsUYuF3MwQlp4PfmHXBKAbhhwCJUgdeX4rVYZw4eYPA9nOUb963uSlT5
xSdp20H4+VrGTjYWT34KuHtG1alqr6mRZ0mkJ+EGbsosW6weeBQk7fQHcIOP7XGn8gpAZpYECZwA
Y2f1+Y+WICrGIJFKG7247ZJ6g1zDXbf3ujTBNwz2tAd7wNTUQwS2hr/YW4zRTmCvuQqx1l5BdkBI
VozMw04E/eQxELUiscKi7+cxK9v02q0dkTo/sVp52qIqOIDtiqPOlp1N1Ol1tilXjmLpSFD0SKer
UmOHg1wl/z7Cafdrc0y5uI+cI/2fHkRx7Eluon35SJaRoBpweroACqgnWxK/5qCIf5TDvFmnD59I
8guWLGO/6VSfAkzd2lRqs/hFuVY8lHASPAeZgQkkJs8IxkjgSLtMVyn3EB8o+93EkqKejXk454+F
Ag+eQJf3RZ8nSEcbIwK0na6dYUnPIUDRxhifwVybf45jSRgZEUynRchG70JmQeJwdUhGz3DkLzp3
5s7u5eQNhrBojwWYgCmTfgxqGxxP0seCgr9p1lsN7uqjnRZSWtv4T19li+mxcLCnHGCcCRi5osXU
41LB8FXByOTHf7ed7udA0Q8KH+0aDrLcPtPm4zw1C9Arkb43mkVLR3WUeP52Fvqpg6yJZGxPDVAW
8UXyaCKmtuj39wFh+GBsVC+rQZ1OgGcfwm7/eQ0QImfo79Nh0YBsHOjFesSEpYIUQzMU2AQXyuIR
E2k2b3Ui8+YTKoFG8lNWG71ABFoLmIl/wjYrnrjB03tc5mCL+4V6GhDCdo4MeQpQMbT/fRi1ZR2r
Z9Q/8NF1XqvADUKC8ipffaECe8L84sWi5qPye6c39Xtj4I6gp/ps173fQ6CXFWF9bYRzXI0jCNNt
KduaLP7bVdlIlqwFL+g7jplZCMV8cldM95pAlURHH/xcmtCAs2FfXOdYP3bUY0ER75F7elEj1AfR
pIgHNibrqRV1p59fmSK899rpf6R9hE8N4QhuocRUA+W3YLLks69iqoqLRFTpLqbpClnDcWznDQNQ
Asoff7M/RCPRkXoeqEhr/CIeIDQEI2ZI2KDNlqn99SP+jAVR4imJIwDxBbnbF9Z/fn6N40gYXuq9
NzZa1MioIM5HmAoELzCL1RjiFYr8Twj4MTfULqiGaTVY2Er9GPF/N3jFHGb5W/d1K8DU5Z0cEY+Z
2lz5yqUBsp6h4kZdz5biphee9knkckNh4Xzg1X7WkMn6JjRqnXI2+gx6tuxkW97omhYjW8TiVoDu
6Jo4CTi0dMWtXQEobEAH+Ddg3nTgd0/CG+05LX60myM4Zrj42ndJsfNH2oLpMKMs9LwWvvdjL340
GyCC28+6K21DcotE30G5SVslRB0X+6YRwfYTl3EQTtSrKfWq53jC1fNRLGhRU4WXRqXmbsyp6jlt
VxwxFr2HTx9pEWWYwcAD9/TPFny3LQeqaxjuE4U3LS8eA6+Ghsq2cjgxSjFGEH199bQCyHVEN8tD
Ltrf6gYT8EmMCPIlW7II8UFN/ktM5HihADL2imsXYmX/5m/nvWmsS4G7zxadJYkLLH3mIlf3xMVG
XeFVv0fjIyfCzWBvMXgDvK2dULkyWA7nrksSyCw+kPDr6fnB7KOXa5NcUf59Vmj5V4bg/ev+IH4l
gJCNhrGUYtuaoxEfpgfB96/xf5aRr7Iao3/+SJORCBY20LyMQjxyqDZ4LaaGZuDSpJNyamKLBbf4
/3HfYDhNJBejxXjC9MjGIzn87aacp/o1HDwbT0o49Hl3YTU3SkZtiF4SShLUSYE2oqsS6tSF4VF5
A3xv5pGrFVs2xcL5+0zHdBFrQruAJukZifeoqiTq5Ra6ODLvS+K0GXxvjKsIqPHimWgWnOQfo4Of
UvK/gMod1ilYYDSTzjPDyhj+e8lF4GmVgbwsOQO8eQQURlyllj7c5X6JROiXUwrZgNCQ+2PS7XyQ
Z64PCOOQN9GeWAXf3vYQkxQbUB62Yu3yemccbfXsr3LckBzaSO31UCdw8QNYXQwCyHqdBCPaMsGw
n4okctoUp9QhzAknp5CTPe3T9T1xtSNaHY5dWBYbFONSphqOW3bB18OtQXrkZbPaYCYMY8zDbxYY
05CLnIPgCF5WRIa6+e4WJvf0D3xgyHhaoFql/WHDPpViU7CnCS1GcpfN4RJYrWAhk8WTh6EURqYw
uwX6x2Sf77vGDKiUMxhYS8qRRQ9a4xvvdiBtnDyKgnn/u7lLE6iiN4zEC6GWbI09UoxtA7n4gAfj
bae9WDo6foAwuCsKMTV8h/0VX+j5tvBUAC6edFlNHySTqtlzetcT0IIruWN/awvaiFP5eA6jPX3m
PEEVaQNjOC6F/sw/exxbHR9c3te0iXZMDg3AWbqM+Fivcztn8i4ItxvYRIo+bsotR9CF2IrGoqfQ
KXTn00ejkXtE0VZ0qoeYi8pjwetersVV7X4YjPOIaZXBCMMVHe/E6NqF7MZox+poXUdo+Wr+zjRV
EAFj4qL+bTC3ZoKuWkAaiC9+S0fmi/+VobcQ/r0VBQyIq7gPuO1DicpQkLn3f7CjdOz1qz7tBpBP
hgewnQr7MZLTIRystgMyjPU9In+YqeMErR3xZnKQOxZOyfqSR4LHMhn2RMSyOYlC9IfdWBwx+mBt
is/b2d9Noms8vtsl7y0x8AxZSbZaS1z3qVU5CLBfQ25HY8ambJjOQ+DkgQH9Xae5plQlx25wVODP
Ue46PN2ZbiMnSNlSe9mBvZu6shSlBOoIitKzqRrst32DAZyjHyMmII5JAB5ymXAUy3tNUf9FWsR2
DcfkurQwY1R0sVzuFQ9yuCzZfApCkFJsWK7bwQd5/Yh4fl2PYxP+bnbrceSrT2WzE09xjstV10Fj
TS9ifhAJueAvm4snggGZrItYDj3QQhdDIMK9ZSidq7PZkYlqtUeJRmS5cniTmamiud1eV7+ghoWw
aY5ZbBmGLO4Xy3mzn7KMU9SzHq7ymC/e3LDnHd6TzwLOwq1T/wES0Wb9u/9swbAWaVYx9E6GhXfm
TT9W5uHn/OgIjdqQpd9P7Fwbiv5oQhml0hJ6PtvB9SdjjyDdev/fmRepzzz1Zp5yFj7aZ3YVNEMq
nnyipy4dap6xNdLzvpEBMK+BsN8Dix+JfmEeC/mTn4CBR0h77ZoIlzphLALWpLBR7At9mwUt8Nib
eDScAmHOX3pTdggNXKyFqQP+QtXh5b++pclHYigfj3z2GcWWNhnEmrjeLw/2yewVBhxvHfMjRV6F
zGcqIaKiut5repbhrjaAZly1PrUOKJlU37muCyp8egrHnGe47fiGhP4S/XWf5N7AgD1xEEc1FTjC
jUJxadV+6HOA3f7pFPh2CjGfQWPYt03hqRG2SnI1cbIDcaj+Iea5Ycu4oY65gjwcCsCR0RAKQHIU
pPdO95zLlMlTBppKlid4LZ4FMkjtp9Sbkyi1SX9XXTirSn0KiU7sU+4fmVJi4IGoGED7z1KvLPX/
QMSlmKK+dfG3bHTpsaPKYrpdXDfxLQS98ROrKBr7gOW7YiX5XmgC0/gaSFdV8lPl4JGe4QeFqLVi
rR0+8O7sIynlegQXsync3g7uXPVg9aLIIjaW14cRyCXnBbnRZLnrf2vxc3fFpTDdSmHce8pHtV8q
nV+g/oajVmHjAcJ+NuI3OMiBtwIHhqYkj6HKlvYQE4KqCuf9fW6ZjNFEfuXnT0dFrLt64uC0NWJf
/JR9UToDFEpU5/YXxgdfj6kXYfbbSm3cCyGPyfez4Kys/rlOxgSD4ucCOWMdJAhBX90unZd09+i5
dEMpFQfLY2zbwlzci/Xz/eiReM1hxX7na2WZp6vvHW80Bfk1xYA9OBHGr16o8qavDEFBKzo1C0T6
4fr35p5rzpJ9Yxwo7LweN/+yzJGgccw3QA7HFETNP4JiDjrkPyf+4NqiDyZKm2HNW/ykJtEfEtK+
kzSzAUFF5Lit6XPjUusQiUflDnTgIVHE4NIoGcAwuDWJgFt9vKpqdFAymy0vGpBQ5BCmGf4VKlYd
xfXmmFt6SMpR4kkNnQ9S0S/Ji7TCmjhrhjku4yq9gwT6DTFVEQ5+6k9menm3hbYGuKdUlEibZG/L
/8yn7Kev8vzeyjNgR/NsBZdMvaMAa5aY8JGqhkb7XQvdpxig4qodbmZLGk8una/UeWfb5L+vESoE
V5DsQWOIlwP2cSPNKA8mO94+ABK4ZaGFyaUK9nWLitv8LDWhsxhr8lvrrZCPIZIxcNJ28csi/HRl
sv0v7PboVHvib7nYyWq5IEcmUkjDznd3VZw9tc5Bxr0XZ27wprEqD8W8fd9ygBk1wmo1ODVjdxbx
AMYAEGH72LIvMoBs6g6AMfnc4VRGw/1WCe4XUfGWeMb5Qplr3nztGIVvE8Q+6ipzWDOfrF+GT1gL
mGpm6GCGXq3SyLQv6L1nQ2cR/nivL01ZbcPxvHRvVZzKyCfkZk5ymRaZk4NDjdpiEAP8QznCwDtF
VOkKehU5pOJLbxdbboYj8qwiB4Gi0poYYRNdLKXIobbQbk7EnQUHEtgP9U2M6vIVlBLWEgrrr9B4
Bf6ylHl1ZMPJDTadXAL8ltGKD9idHWXcCTh3/6CoIAJpyf5sATkjKT9JOGm3RD0s42KrMzLw10+9
bbe1h1MKU2T0nvK0hiyaEQBIEJWISAz8uVpuSTp+/T+Lxzr1z6joRkPdF2QPDDtf3jDgDR/TXr2T
IuovslhQrsiVVitM+RLen28Kn3QOq7vw8ap4oZIfef2JhbpLeY1cWRbXAbn4j6EY3SsyBFEgtElf
Te0RwXtcW1kBb36m/WmCAHcJ8lQWzBY02EeHAj+FF4YUp2Oyv/09yneMwz7OY/XqkQYsqIR1UJdq
x223FIqvmw6yTXMJT/PdX1jKEt3KZdbKWSfh161x1HuGyOIH9sp+OyF0ltvTykC6YVzc5sihEOlN
4P77RZD+RBo9ssPcTnuTMXNf9fM62zJyprFe4BA7W9E0xkVawi4rXumkZYp1DkckN0krje6lWTWe
/SszMzFKxtkD8wpY2wQ/Vk3ZHDUlbChiqU8nsj0UsfvDGq/sHaFlewBHvYPvWxHCJPNHuzGg+LhT
2qfY68YjmyOcX8sbi5eKbSVybw5BUwPh6DrYYhAeWx7eOB8EzNrM80/flhJ1vgSIe9Zq+M0Ku1zI
VTna1EbiMgio8RRdzMdk67xvkgKlkci8C5TbinEAANPbcPr16zvL2Dvrgynd28B+vI5reGNtkP9g
i0wwphrEwIJMEB7HYRcFSl2AonjUgF8HEXQdaygRuuqxzElyO55Tzq1y6EGrdTBuNKcnugzmv4WJ
HVEwo4RO4rmjgZaO+bBOg/ahEBomGTb1RUhf7AnUHuuhX4OuWE2VNqPwibZJ2w+noO3BdBQuLA2e
V/hswycWB7sXmA89cmiS8NXCSg5WZl6y4z2JlUF+RuWHwzoy0CApk0Wp7phvOUo0MhecI7Vc8rz/
k+6/yo/OcDEIbVY/VFmWAUK2fN/bfUsdUyU1lsqp5Zif2JY7yjmpcktnJWIqKKoysCeXyyhygPgz
uFHrWEVqGz4SRqE4k/eUthVX1BBmXtmBabUq79DxMOtn0GmGTxb8nzhTIFetsRvLMQZz0tNTzTHq
n/iiZ8xe1et9yt2WLWloEHVUOgWKXGJ+eTzzaiaxjXkmEhN0JIKkbOLxMYvQ3d/H7+xF3CmG9PaO
2GVrNOW6mBA2isxE6jYN6OYD3DTSANWsJycTJs8LD8+V1Fs/xSLxusYdBjFf2CTePMEANVko693q
szIK7LcxEiQXbZhhpT/g27sQVpj2x5uS2mWUmdwhdlPU0C59xm7T4/PPKqwMD/ezIDVNQm92p5wf
Wys085FTwaWdARGBaRDnP0Cso7YRzsqtctC3qNutijSNL7wts6ddj2kr8K9ZgA5hmhazRDhJpOz9
dGnxNkPlstxKBBaPbvfv6UMjL70hJJP3w3ODDshjhJJ82xIpFfj5qbES/5S9w8bTN6g+JCx4+eSf
5lCFSqnY8twoeqtThauIKCcr/2Izb/p17+YgfU2ilsbEfyzYDcvriM5TDFnPPeJXUHvH+9x7TG8T
oOqfet57kawqKpwstVS6y4qd3g2SOC5CkB2FMcbrSEMNGpguWwKXEqczgSvfwV0dmk9ujDFP8An/
+sk1zt8TeSUpDdG9y254olMlGn2qP708/LTcIo+me6BWmIVHy92/2hUunjlQePoYLYRZ/kGPhIAv
Wcf12X0X60cnoixToVn29n+3u5jao/t92pw+VeWiS9BuGzsAouAERgYqsoTmRIw5QQ3l9WilnPKY
gIsNmzZVD0uzddm7eYbgFkW0p/OmtphbN8H/9cmCl5z464aOEJ7oPweEyNCmDM0KRf+5B/+rDoYN
Il6boMnAzt5OkGyynZsEr+5zAYiFXWtcD/B2Y4mOVBbug4E9aAicaK3przVTuJbRrqMdDgjU5/+F
XJjbKje0xTSVaDUaeWVQbFeEXpcEG2AqWjih/6OPjAJAwKWy4nzHOGQgcoKvLm+nbVUKvzWshSYA
sWTHAVA9vjx9Sg7ocyjAiGz9Evv6EhXy2xsCcFHvqY0Bnu9IaWcufEsjN20M6GyPISb72jEYmqPq
0j8ah2pPLnnREh4SjT15wANBHPL5q31g7wpGBASMgeJRj5YxYkpXZJGhl9UKL/aJpiKZcWCzqYVu
pT6/OUXOkP51T0zJBjOLo47UDxz7z7DeyrZHa7vjOd/VULBBYWjvcBND/3etyMRkLI9vpalV4XWF
SXAhH9rnCGXFTktFR4MkZ0Y9sW2rqNBrxrblnMGDe4NOnnjT1DUq12pSJqtEZ1Z/Gp3L/2mWN8IS
s9dUmepZs1dO+ng3RwN5S/SJ2hBBQh8b4KPDpzV8WOZ88FckMsUud6mndOlwI3jKNSEDrHu1v1Uo
ZkWPlOCLLKzHE3xodsC/QAe/Ofms35jco2NTOc0hiqHcF4qPnqr9mp83UdSfJCWllOJxwQsq8LfL
IHMJdlkLGRwjrTIX/+o31lNgQyIYQEdX3oBDkci9ZtjDsb5IxQ6d/XPLbORfA65dYBvYZqsy9y5l
DUwfcRv4BuO9Tz1nHScHFIsGAemLwCsc1GLMKsBAOZ7te01uK+bpoSCovn3qGq6CruRc/tGMj3sB
hPiGnOpjS9MY2zVH40DuLTiM6w4Ff3GzkrXiLRSulNkdxizMq8+jVn0JlkjczvrlZzkvxFhYlZdw
VHZaC9B90Ej5N1cPWLtNcCg67Qlm5ciEuj9pxUpuFn/8ILW0N7Dm0bCEEBSYFisL7ZaDy+j8Aa5x
oc9g8wR+BlRBnQhbGwrjCplHM2GUoHpMzTLmMClbwTlB/VmOzHTPNRZA+I5/4FlDgXK8Sikmc7BC
uGfaofhZDXX1liDN3HP9vErdMW4mJ3h13skCqwMxFDUz14KrUWEwifRu85pCCGrWEH+GbzxlmXm2
MuGm2CiMApIFKwFvrEp7sDR3nwDKroqh2cL1AV6iKKUsO+CgqSwki+FoU8q0Weius/niLJW4WIZC
jWaVD2xVuBFyhOH1o3OZgJxdN0SbWAPWCUZUJiHMix6MYgtZrIowu1x3+CVAhP9y1sdeF0JOuKqm
BLqAzPz1HVLtvSeP1HksiVMwRfvGCnf4iOdO09c5KlXdLwTR96k6oH8KGPoJS4/3R9p7d3nhyJNI
TNtI1TsYy3eLZYBjMIyFJePcr7vhU+O+sJ7cvLu+jStdzq+TIxSm4yCw02FbS4ADODlWGwtsVOXk
j2XNOc9nmUOb02rq8ZY2wTPaHGXnL4WnZLEwzDLrn7KwsTVU7wizpNeNx9bQ4WyS8P0WNMJZGG58
vBTmzZCqOkO5LzqGIwvj6PNY/q4HomxQrUTkCi1ffi7QYaQNHQkivrg6OInDR4Nz2wuB+TQ9WgzR
e4edbg2R5HPlQkhPQsjotuWbF/tDx3BJCLCTh1WOnBnYt+a8egL6yvpPjGTRIl+5Jy2uSs4ZyzSG
R9sGxpH92q/hyg6bvFdx6Lb0QBOHOLifdbj0kg58g7si8Ul81iOVxas/9Zh+gtUOJ/pdECyta3e3
hT6/1aXYFZJwrc3//j0TAd1pC2EIsk6PfEyBVHQNnMym52RBrn2z03cq/FvVhxbyuDKU3aDYfskl
y2ui1fLTemrIvPGkqTKPJWOBRyeSxE+oT9rocd0cbP/XWDmfsMlD6s0LuMNDMDltLu6xZ9ihhoe5
Z4M8rMFfmxXMU08/BxjSMf14v9ULnYH8cTPVJ1ycHAY0GgPM7U/AHWESqL31UKvEvlWGcG52WWFJ
x1wWzeFVc4ojpJyAjDmSHpzvql5d4tCMYmMROU9g6J89+Xa1UrsaGRzcU0k+gKU6pJotVIPf3uNx
+kQ1H4YNHYBZ+SO6IcLLO1HdRqYGYSWMi4Ra0zY/DmF1e1yIxLt+6vi7oTzZrqQOT4lG5XyX2Z6Y
t5AAgtNburx1MzD4/42UDV8QBI469jAS4Wmy7Pc2e+0EsZgznmYTBoANBMb8Cu5cx1bhzMU8WPyx
+2GzbbJBEcN8Y9qFyhn6sO9L1a3k2OEno5tM6Eq09JEe4Ac8qnqUvr3QknokPGoCjMgSExprydcd
WYJHm9lNroZPwiqFXCi6zs3qvqYW5mxkt38L+O9JR2HJYpjaH/JQmrg4ybm243Ca91knn6/wX3Gm
XoGQZmXkSJsuz58veRBKvBbYem+ZNjHcXFdFjs598hVh4y+/gNHt+x2Dqt52nk7vZUki1BqCgH+N
oYbM/ybj9iIz9tNzYB8UJr6CWvgTOgq6PBvYqbkeED+HrgmHrT6NymZhKMfO7Y33E8zCLUDFfFez
9MBq4gGDbNzGd1RIDBq4ywVIkAXSoX/hRAeosP6MGV/GOjbDbHQ/2UZGF2K8YZj1ScsrksPlKPhn
wotvC6KHbu9a4vV3QZm68PRXk/6p2MFAF07zoXDJElCKw2VgI6cODfe0kfri/DUIUXV6atAImOrX
WjWgQ3Ycd0W1WkM1cCKvkuan6+99sxgfj+82FYdbvrWOgREXb4m3tHkExjvzh1tUDMIesTygSCeo
joRlRf9IyQWFa0dDfk5OQbyJBunIjm8O0MTEH1u6/SgHLDfyTnZGOSM7XNX+RJLR2x5Ublopbp3x
3o4PznpQFQfULYhpNwMulQSKg4L7xaHJHATmfuBNdpjwCb299lzMYNQm5wbRODtk6KYa3lWZ4BgM
K1A428XlXKxlcHiILXkW682NO4/zZ/9Jvu3WbutZkyT5jqqeXtURSwxafHs3Vd68PuimASAY3Rzy
alViIIMt60acmOSkH85wr1chSBhGTNdTw6nMt91gVwvxSJF55RuIVQMkEVflDr/YP53Cf9vTmRof
yIgYZYLhO+dVzSf7mn0O6uU/I9xQizLLkUNqCp0HlQ4kuczE9HlePDUh32/HVkxY0zqX3HpnL1Vl
l2W6e8eBoOGyjLjcLqb7vCipfm958YFI0OrFVW8VQ2d1Ix0c8yEx3VIZW3UaIW36sRZxvpUJoWgj
sXieZghblOY7DAsv3iTgPrTOaT0SVsj6t05qnRk7QlOdXt6QFly+E8LlOKEBLBniudRqWjidAHqx
jnqL+HBOeEFywy1NxHoJOBHhvR8N/daJ7HhbU3XeTZs+vmhew/DQ5ZqOq4BpB0A3kjvB1ug81cRz
mUGcGthr24oVxaWUZOMKzCHrlARCIbjajgsbEg2F8F6wruOclKCOVf2Y+dFXAnUUBjpXNEk7q7K/
COW8AUf8jSw5cEcgdwFKJKtxaWwILyEGVRErjqyD4u0ckvfpQ2yFrXWZ+184NICyrlk8OzsrJRRN
bCSRzOygp/u3hDkSjS4McW74+lPKBBqaJWDd8QQX1mGsV59SJhIdSDs4O/dXoLJ1dlElftsuxHbY
oH+XZumTNumTkbZTfu19ipecQV7ZlBXnHf3+yi5QVN/RIe0S4uwN7/BLi+kmztXDtdE+eUKjgHQt
LIw3pec2HcBjyTs0R3cvQm4WZfwyIVck9g9PhuAniCtc2aOSqw5/QdXddINnx4y7Fjt+y7T7LbJS
M0jAM560hnmIM+N2q1tng9P8oKzZoXWSZZCrOszLXyUVLGEhxy5C51JcamNy2y8v5PfpEM1+g3hN
SgCb9YGyeqBkop+1AoYKIbaE3DRDnQMUdnVC04jXGBf6E69pQbclp/buC2DNmXU8W+V061B27rPu
v6Ua8XIPjDLHQOPagB8loCO1F/1QGJSALJi9B4zLVtwtTBhXRXjETvpWjtJ35MEM7yWyh3cMiSeK
dBqw18bVmjpXDpRajEDCUUnayYV811T+PTlia1DGFAInVToLx88hV1LMtxz9v/+HhPeitycuJlxM
xURtLYf48bOWPGd0PfHQmuq+kaPIWvSxyUbiosY+iVBA5K/nYE4rww1NiTafs0stTrxCVoTdEsyu
w63CjcNDfj1EePqyAiqUU1wEAqshjBluGeYXPVgodn4M9dJM012a1Trdvv8n0Jf/5QyDjyPMOJ7l
m1dlXL0vKzRsrAJgBhvgzrDPdlRhSEnNa7H8ga04QEofG/A3N67SEpTufzqHNxSDSOxMHTdO6X0q
KnqFyueQLI0owsGBXUyPxnGNmSUJBwckSWTmamz1Na/+T2zGeNb4tEdS8AU2SQ7H2iqJhOSvW/4p
Obp8JvRWNCMWcTHTHdu/fenKCmF61ZjmAd2u89k2tl1dE+eP9uLeZ6prJZfz7Cy4/Iq+nmL0tvwJ
rFyAsdbAXA35vZ+A0AQFmZUoGWfymyj5mlEITcIH4xgGP0dCejqOfwjNNs9zANFtTtSoXVZlQKHt
3Sc6e6yGtzHcLlcor6c6IsV0mtFVw3ZNkgxXK7kXU7sdovP0JqKcyjC9zR7wAVSJ/3rJOOlbIRbY
NzVvkQJYAS3oJMoeThIm5Mi+Cziz/vMr/KSKVPvKMSJTUKiXprI20s2znssOpNkZ1VnkTc4O7bR7
eSGe+9HC83xJlCEoUKFjXmBVTWioboKlEk0P3SC35QnfOZNyfltfP53aHEgDodjAFv5PcIQ3YFxH
NMtQ+dY5WXQe6emkCbstKR4ALqsC5UhCYiEmTRsPk5HeTa+sodqQ5myeVAxPYIvMpUw9XaFZyMlM
0CLv6NlDrs7wTBOzHPzGrvaCzZSWVMY1eVqFcbW0O9/URHLPMWPNtUrzZsDBzf0U3eUUzpMXyr62
YG0H2vf2TxETkHjieTM2cjsfibS7w8cjqxnUfqQG3PvJwhrtoiUoJ1WpwOa/SCvpOqdKO88FI+iY
PDSADL01IK9Gs4y0fcmbgYal7Zl24c8FoHLN5K1lmvYOX5B50DttwQDP24jyurPD20QtQKXeX6nl
cyosKZ9fyZcb7gjIqI2NWHrWW8nSdoW9ytBG6W3lB8cR3mqP6N9F0DS3oHkHISIbbS3U+nLJ7LJw
jAeGU0OiudBT9jDp2wwTLxMajr9/GZrbR32WHR5evO6lfqusi78lubToX0Tw/EmzUo2r2AiS6Msv
tiN39OQs8QlqTSEKawEA+L8hFA2NBYYQenrtEzsGL/Gh8wa3RF0Lm2HnRW/MRed+2OwylHicX/Cw
lWTm+mM5xR+GK4/MISoHJo37guMEHkOtrZuQuwyw3+bbVcuIhyZiZPt+5vDFAfF8jX487Zfk9L//
FMxKev4+ngshIWULpyPB5RpSiGM+lSe01Fv2WdnlMtloEl4Z/VxsYWdIiavhf5X5AKFvHi9B44ni
g+ch+gvr1lhdsRs/s0dfbDGlq5TJRQrFVHOl246lVJWn9f40v5AbehXoSKn5CpPE5Yk7YNlRaoJq
DCV0bS+Jd2EL32ZhOsUzwPO0a8aFjv+bfM636G6HK3bqKl6y4TarqxHDTbvkumACbxnGs1FPmdFZ
jUIxWoPQp7opgNprbrsr2UyoGXdgymZf11fyRyt0GrJA878bbn+3zBtnDw6B9BkU+OfEr8c8ff0l
MjaMVTK7jv2K6WqMFnPrrhkcKAXzw0r1UQ4wnxAWxD1v3Biaz3uXt9+UO++PLkbk+zTz6eS3zemy
UGbRQVXS/8YSmK2kLouxzMO6PN3rYQwQ3Vakf2tCyYq5ohDBj4dBfKJFoFC7e8MtAou6GcUvkGqY
SgUIF+ESv89jQWix/Z7fgQzZCUnFxKXxaBqbZXwIzGV+AP+s+nEdQQI6pNMZs6xTCU/hjDGRv/f4
DAgT8qQc0aMZdSeJ+jiMyJYrX47I5rkfEvs3n6lJhGRqL+1+mqgAS6WzXCO5sw/GPMDvdMYamh9g
UO0UMz2bf1Lasua1C4SKlcEJjILHDxtn7cdW6ujbkqfPBkEpqvM2fEd5MEWA/5JWILsqjpvFRQxn
q3UYy3yE1G/DXPtyf1MqL0n6ug8nfxxtILcnCL7VFeFqunTbyi4OOx5XRFfQOIgfhHStPTAyH3z0
Sc7OHJcaJ9dZCtStckpNsF/0jWhp+0uh/6+ehQaDLO65GyZi0CPFJ9gnckn058sSX3pN9Q26UorV
zbd6MMjgjaXFipwA19w24TsaHGhpHHHJvJuTX/iD2v8gGUY0X0eCWM3PEa8483oBPsOyRi1Ziqbo
NTIvJqLNUSDjZ+FpOzk2ny8kLgIrhgCWWMGqHYNTrQ1roSuQUO8nU30xny3qlSZQK2S0xeHiwYgC
RQB+IIaUS1aYYQhZ1uwMyUaOf5OJ30+mTppJsW5jHm5p1mlSkr9c19zE7nPLNz9Coej58utxYiAL
9uOJQGWxXzRTfAUd4XyOR4vF2QaumlZqWI4M4h7L/agsVmvp2oK18NVxeNtMJ273skR4KW219nyN
CF0fxhOKtnzjoxYHfIxISrYyMH/Oap97yBqEIA0/zdgMzZOzVX13/jM3oOvotF8PU1huB/8H8nUp
IcOQFQDe+6D0XLVEsmkI0Wb9wTFklSxsJxhM5bf3xhvnhvCDdO3mRC/jfhvXmsivx5LTN9E7XFhG
ksUunt+71jcglcSO7MQ7sRH5WB6jx88D8JhPQzQkzi7naSWJ0ybJVs0c1I5UHYeJ8un9ZzpDAU5p
pjOp2GUkEo0UbSoRzACh60SyLmZLb/rmCluo3QpS2amS4NZVN9g1bbUMeGeoNVKpRBdNtRKs8ZRI
g1iSQExQnTKcQw6G7nMX3CB1OEVqnUQBJohU7rsr9Uh3GIqOPd07el427T5o48u5b8zotecc5FU3
liDbDn4A4MJTlO70C67hIp6ftQDq6R+UEg6VGrBdmGa71XFBkIlu2gA5bVZ+pJ+vs0D/jGf7Kv+2
JiiNx969pdmRi/5m1yT6/+qEsWEfq37g6VEAcuH9rTADjXjf9LGpcBNDS7lX1OBq7ELW97dfvRGA
dkGEUaUD3K8sb8NGtlCfSHI7SCaqfupEWNpuenZ/G8a0W6yIK3w0A3CtkAWxS4F37YsatPZd11aY
xwWvOFy+e4pGqu/VqwiGMu6AdGyq26OnnsfHDk3bpk6u4bZg+/zV0ZpJQk1Buvgxn+RVcl+CBXKc
7CgzPK/WyX7WdirYyyYm2BjhE1vrOQ6POohkjU4BD+9zaBp9m63S4c8kr9w5qm7QMRRcHkEFjS9x
NneT3iMAzT7gP9GL2lQwCoy4TYvKMPY5yUZ0rRzSrWrxuTrRlR2FUgs19OA39qS9by7rb/4e7RTc
LP8SHeBEjCkIUo7rNH3opSSMKVaVPKkgyU8M191F8KtCBieCYW7X6ZlsxuMDmEhfYaOAzu7W50DO
204LqHFXMUm2ZHrUQNp0J5Mm7sGeIUrdVnP0iJLPUV4zlRu6JgO50ZxMJuXr2GkmrIRXGqVg2EA4
cWV26N+1pew2EEHOyMZSiON9dMz74wbAxGY6P0i6UmDGmSn8OwMp51hvIFRatD4HJNDyCBNxCGp7
Y4D03Wbk1VqlrDByTjulKfhbm6JwDhjeinTJdqxVSaDlWPARqqkX3mI7/5+T2KYqZt+yAlk4YixQ
KJKIhvIQjlHGKvheTUMCLMISmBQ2Dsis+N+nltISUSD3Q9bHoRsHSiwQf5DOL1Mh1FrelWSrcFwX
OI/pwXS6/ap5uWlVlunigCQD1X+Ir7fz/CAO2DVl8GlvviSHCoiy2dO0rOr6xdvKoV816qNlvoyG
lm8MA/Og5ETxyPSP8FzN6QTmtHA1/DKuy9CtNWD2huIo2rOyRmyc15YsauDRImjwKA62p4nR7jZm
V7HFVzTsqACkuaacJh/4mrcPsVuL8y8xn7DZ0D/c3UT2W+de5KeyDAkFqG1L3JBvGUfpwUV6YClz
EN2lOFInXTc9UYDS/kO8bfHe83E0JJcwDFhY85osMsKVSHuz7tyeIEoHRy5wzXbdkP98o1BW5hXG
bK43O2KOIFeHA9ZZuvlSGnZlDn5YS73LadjuNtQ30sff9c97FgxC+Fj/gbEJZE380iB3NHMwWXfO
itTbXnNmvmTLsxoPQJbmVqYtFWNp0PYCnQZ0NPPXOCulpeNgCPUKsSAn5Apv9ynxMf8spAD11Q+v
CGLMWv77TacK9NO1ct6VxWzypYcumecWRmVU4FdsjpZstS8opj7nBhjIVDl8Sjqtzvgd7YhWHEdx
AU3jz1p7aqbFJBhSVcxJwQYByBnPmUi3IXFYX9E7cQcX2QQxgvbqb4txgddHqUGSN81WMf+eVpD1
qpDRedaHs3ycPPnsE2wLC0zFrAn0kGwmwaDibYssCdU10XpY3HfwQfZewj4nmqYYG5RYxZbjY4wt
MoZXuG9K0uUkRy016VamU0gwu5bt5e1Uqah6eRGIkedNVW4OauBp+mrBcGdi97ZaYMQLc53mHPvh
mDWymx5ueQW8OCbOvaUTUrhPndIaUXpAdCvOqHG36AX9qYgnbYP6kklfZeE/jB78yd0e7Bbi2GT1
N7+GQwUyzPBKmmPri2dRzeJqC7RWtQpXFJDPbD98u2vKQUvTX8fX4VHj1EhGkodd1OJU2A+EDt/m
YhOfYJopU2lU+0tdvKRqjmoYG1/N5D6PSwIkf7KePNrSLIUidZ/INaqTAhluvmPm1AOeuXoQpUNh
M44xeR8Rfawkoz3jYbpkBXx4rU163bL8ol7bgiJwoR0Ih9wyfEurUWYu9WjpQKxcUHGgzd+zOqZx
of2KolThq5giScLRlWj9pVLTy1OP4gz9s01CJIUqHPWa3bOOUaMFCZuLawV7y8AIZdR4c2QJG4qs
LxEchJEpfz3jPN5Sznb2qcPvG0/S7o3p+JYKJINCbcVzerX4IDV6Dqj5fAMtCmWvNEWQ3r9LhoBN
Xe409ECn9cHo1TJwPVOUc2QVm/MEcmKeeNR4+5JVbEg+GJ4SGqMbllkziEymL8uOEVCxAnRQfBJC
IgXlcwySocaFUR4dX5sAd3muci5Rtad1DBpiIzwS84rPVTixE3v9bR3ClxDiY+Wfbc2+2L6WV0/I
VNjFGPwjAAFnjOlj7Lo1qx22DLI5RAtlhbDKP6JD+/E8V7WSOZkO7EO5S9KFLXG+AdsfmfJXFZ3B
wJcrUXq5tahtVBs4D6ogSYmZWS6bNli4tVYc83YlCr5EWivRS0FsD/XdR4K5HU+I75sFRG3sIvBf
EbsU16XLPp2Gw7qLKo9vaC/dVLjzdn1xDghfn0zHU38YWAiRX+G0Befcu7DvWQ2IdtC6cf5vm09f
ux5hGIp2kKRE9ls2W0pFhXtwHXmPyIWVQJL+6Re0l1iKODTBAKes8oDduX5PKwGGim+ruEVfxDOH
rOf88ZRTpM/SE9LtmgfB81868PWlIEBpbxp1RmibaStaMBzAK28igs+tJckq6qbmtYL50F2oEOd6
+zo6F+Ib1giGvqqskaQyIeDJfWa1P26IJezWMR54xfryxlR0UmkhMXdKyBAny+q8FlLrveHhus6I
pT3rYCnp3R0nyKed6Ga7tK1paD4IN21ymHkanUzq1tAaImX67DkZC5yKacDHXUH4VXD1Iz/OP+AL
ZO8COHfXLeAoGIU0IGwxdEOXAs8b36sKycu0PEI1GReZyIbSNV6jw9lnrg7y5MjUaqUNdW6iiD1q
RFuHXKzMwfH5Dw6/KVl+901UIHqridwfnLzPfmbXUdiH5w295PloQ49RLKCiGhIo7nXH/RotSHnf
PQJByN7cxUl3VZrso3zgqfwMHeYROWviwlIdvbZHdcZkee7y1DpnYXEJ6prpTALN0dcyBJeqi1Hf
LSjP11u/WhqmuXUNnCaVvVMHiES+0NQW4ordeOul4bNGi/QNTKiEu5qcLmB3oCZF6MBFJ1rPic+b
VIzcJVSEXcSp5+K6Tidt/eR5p4EWxi9pH+JnckCPqSrRWqyLoeiEo6z2a9pU443wUccg/vORhndn
43W52jxHI4md+6XsDc7xZXJOT/Pi3QJHX0pcN+y0hKjvm7i2Vi8AnevXXK1/wtnrHZnzK9xgjiPi
SmHJJae/z9BgR+H35nBQ7u7gLeaxSCUkfj5BZSSqY0rhONZbdYvEMNVM8U0AeYQcV1AE+Vaoo9c4
QzOoadR5fTViKLaXZ29UxmqWlQN+6ECAc19jkf3+th0JZyiGSwHkkj56QMr5BCfgkjO1vb/kLpfX
83/ttPuCFmYw/0g5V/K0z+VAslrj/3v4TPR+RG7EFWqiTYsPMjy/uHyHgUG2y64dgbhjva65Mi9y
ll/89fWZNRPoyBpE+lV3GrzPFCbZosR21rT0mjGwJwWdWOoqgksHflfiLi50vQTTNPE4oMfcAUsr
pdspae2yFdYDjDYQFKQNVB4SFLPzjczlUA40Q/03XiM2nHHQ/iRDqBetBskOpwmd2Yr180DDoGbO
EEUcXCNx3Qwr7oiGDdfSTGzekGWSRjO3ae1cuRZg05Ep06hBZF91UNUprHReU59A3EaB6DM8xplu
7KNajZvhwixPUeVlryvBc8D2HZDGxrx1QdXAZ9pCcfTAoc/kG1f28a5G5tv3GVFshhSOt0WNl+ii
EWuXbSZrct+2J7ivtD8pmsU7Ul/QwdQsef4tQi+04WzNvqRzUo+mQ0jVGP5EXbdb4tk+M+Z+B6dR
cu61R7KHZnj5qaKpDfvWrsYJteo3sJyaHYstp+SOwZii5nHbAjQl4Z6GJ4uht1m/l3Im7AQy683K
H4kEViiI1GBhCMoMmNqLZOzEXdILIalRjfZ8jEpJ/kWw2x89NJ5YJO2ow23GoGGEgR/LXemZ3bb+
Bvt9XESMXe2KUQKV29MBk6RnLWRVdN5aS5gzs8CjqBr9hIHwlay1ORRZTP4/tAarKQNrVP2SxxAz
PbEDWyOCCGjtEa3dxFXrKXgVTRPXmnvNJRfygML0e84jhkE62SmGmhnTtFjWxRXXx2q/v3l9hk/w
8x0wLnVBlvbxqkuyKiU4R48L7uk0AsKmgzTQW/kD6Cq04MfgBDmn7jNLkdwyOGw8inTDi1nxitgA
+TGEiK0ksYuHTQFSL/pA7gbcMufDudhARSZ9Bo6SPjfNoiUifsAI8jhxwIu/HE68AtfDi041VlEA
UtU3z0z9k2IxF8EDwOTkvZ1KPo2zy1OwisNtfaP127z4vGi0K7FfgZGW2Y1j6OhrdDm1Eu6iRH/V
puqcDEZ9MUjdMbYH1DCQ6IK57TVVlBnyBFf4jfCtzWzdj7wtjy4qAoX1DiKmLKmvhd10nk8HGYfD
BHeOiYZ4xhR5pU0KdSey/BLptFB4qIKqQxsnVdQ8w9LNT7AWGqPGAvWQLBTEQw6rmoPirv2FzHxq
pSLI3Oj3hpF1qvqTORCA8SWl2XwkjO52CkHtUXvLXEPOhXR7QsjvRGC631PVoXkJCH8wwVgoII3i
eCB6vnNHpyuOY0M71fVQGjIUxnvoatk1IMRw9ot92YJtnvDEdLLMJ7SbRcrjq71eQF68wRVXtMjR
a8cNEGMG1D49JJSym2OKTi1TGUTFRNtB9JycXjSOL5fE3JsoUQuoJ/EN0i2Hzxcyy7UzswsYMmRm
/Va67jXfYXl7VafSHyYUJJjhM5GsUKcnoiv3Bn4Dkf8AeR5/2ta5IgAk6ANK+MR5bAGnI/YYpmZN
uQ/xf3J6d2u7jgabNjUf5jRIOJZsLx89a4F1Hudgl0LErsSjwmi3fgEctXMieoGv4vr0MsLi75Ax
Mnzri5K5N3CyZb+LjPq281WM+YDy5YGyQ/CRENWM+82Jowyd3mU8VbI7VFPn9aHBXOIEialafAtk
ppO8ZPS1Fj5g4X3GElWWdIHP/1vSE4NOvB5pADxIa8o7rrO8K6RlNrEiOzmmwEEZoXSRCtf/3P99
fxilmxLigELWdvmLj6GNwN6r/rBLo6K1+MxMnRTiPtabgOibcK92Vb/rClybk2SGfgILflzhcq0A
EHbw1/HUTt0Rna6D97Y1cZJMOS395KQ0WkhZQqDZEPSR8ANq0vC15exXbb2Bwift5koxnL4te32y
4FH0BG+cx2/Le69lTRFeIZ23B2YSn80Kl6je25EULbZGes3wrAg9Op7dAbdomeYcnnVimn48apnq
JDY9xe0oH5iI+2ELcHvq+Sc7IU+7Co0mzCrz57ZZUMn0QXNigJUAcftnroo/ZnO956J58QH2xZds
cEaCXTdmCizmeVAOphlZ9bnNuDP9zCoH18IZGZVr6Njt2Ecq8GGsZZzcWvN/zhYuEIQmdxmpgWP6
O9lgaNXhSMGX3Boni0Mg+7ZxLQGDLl8fLnDhPev+2aYAeiBA52LZWHMOY5LzDaY5SXDK3dBLmg1j
lJNaB430OF75Xu2uXrqMuGBMTDaRsjyr+wuBuvJg/YJI3oanGp86f76d5qkTtWjR8L7XaxH8a872
ubF2cU6szKqmLeE7qfix8EkmIx1uqDVneGolPuogMtAqJ7sIM3PuTOCmnfH7hK+3JffOa0oefKvm
9hBpaNoCkABYbbk+E7EaCRsIGFbPwMX5O4qB67uReOwbOmETzdkgsOo4B10ay81iDynNBMjoWvae
jTqXK6GDQ7cOAWhPOTf8zcEXzppk9WOa13xj/5u+TiCUISknhZ5/R5MnsETNBxbcICIXcpMjcG+W
iGNXCS8if2Na5HJ+s+w8cxL6yuyWOj1D6mIz0y3mnrPANn852gQQdmhlCPWc9DXIc40CxNm/l/OA
RSwFWNLI0Z6E92egWTnk3APAGPPvnwnBkprvfB0hJ9rOs+AHHy3ZeJNkspU7Fg6wKG9R2kpRFm1j
nPMJA1jnzWak5EMEfDWjTvStbC68x4H9VullF8wrZD3xXAEWepe++PZMhC5QJEORuteQij69BYcB
+XWlGxrE4tsbD37EvVgTIu73lq2dlTu5u0rUt+tl7qq5MsLDPeuKsIFpc1suXBjfCfVwv73v6fQn
Ne+vSL+0Jso6qRMBNOFo8rCdywr49Yh/Vuk6XcvefXZDPiLUY8B3dGRTKTBh1RkgnDrvFha8H/O/
XPLrKwB8+Zu2KvZwibn7akS8YP0uIzUed4tvHOTOnO+C4fuuOqq9Sk0LmAakeL0WoExnxu+sVWfC
EZJ1FLqsamTA/WcMX+c0rf4hqQp0Sz6t+CbMZliFOkaYsIsw/4QhewU9+zMd8i35xCst7g62WBZI
M2t+va0a0qyx/boVXvWI6MtH2xJ0NmAAYrVDgH90bu0loi/Msp6akkWUlU1CYHotFgnC+vG7pC4I
/c17SbTHhFlPAEEyK/9D62RnY0D0VbxRU7MBpAoHME9GWGcCSZH6z8tXtnm2J6LxWoKWXXWiBgL7
UqCcM09ee4CZG2dwHSa4uuxsClCenVwO+6bAU06z9/EoXJCyWSp7b1u43m52JsguiI+ZszojNq8H
+PLRvv31GWxWyfrb8BEPUfwCGQQHLzanPdmfLf9xubbiRGQEBO95mAhqAHY5NyCOdwj9GRHSuV9K
nxjOm+sAFa3xRhwXb+1WnxnadbR9TirbLZqwA/zA1bj/o7pMTUdFRqONX85QyhsxT3FhX1xic/zi
3rZNzmn+86zQ9GJjK4srhKppcZXIw5WB2soZWOUeNe/sVCDz+ouQqxkVcryJm6KjRFQu/IUfbedb
VjoxS6S4YO0WQmklJcGdGVC9vYcLkgCb34Ca1vZNgwRMypnmkxlTrxP6olj0/j+DHvkpDbvl1Uaq
JeT/v1Y6s0AOBlJcxd7cldbo2vq46hxSIaWNcWb8sMl8FlXetJVzxpS0vJWXYeZMJZIdfjCc1M/y
DL9MoDMmwGzVUhz2/+jGdWSYJuHZRAwSRdELVnwNtBo4IHp3gyTnW/oU0jW640KSgGlYKmBENUOr
ehb69q1sYAAlXO/EIIz6jROJ1PjVuXBqCLoB0HsL/koyeL5b7W4h4+JRM31c2eT+5p86JkD+rgkC
OaD68rYam+CAy+wNb9t+RjP/Hx5qB0SKVYR0Rbkbj2cmo69dk59lBqYdYCMWFKjul3m10c8W7zL6
0eDVeJqQB+iJNileYrm2Tx439LtK4QrErQo/ZYEdDvzWMXyKyumZhLk6QPPJvU+itBRLmBLDmX21
hwrzAejRdgd4zQgPglswtnnYFyZ521kU0q8ROHxc+JM5oSsN5qfmaCIvz5xPc16w/ftG0L9Se4oQ
R8ottWJyPVlhKM3cnB8h1JzcpYz37siHRa4OtmW0iZmf4zqZoVcsOAL6yqrpiWA/WfhY8oUUzH1i
LgJYpKfrBkWLMvIUdzCkVLY4nv0BX8IR0I8ZZb3IeATCcyMsAOXuunAoZ5AkFn9P/FSXSoROz5j2
BLhGeqng4zXLHgS1dvau7BlDxaY5ZBkD5OGanR8rkbSZCU/hOqpX62T+Qg8naB9b+iO3SEGTZy+e
DzV5tBkcI8gnZzA+Ooue4h+COcIdhbZlUGD7xk9vvPf3eNsJy8G0xS+9i8bN7Bpb0k+Ftgo2c1hY
O5jqLMv3aK7EGX8Y5L8hO9ib0atbd1RVXSANpP3+9YtPwq/loBc8T4CcWFJdbuUz2cvMqIXM7Vxo
WdEUwbc8No3IRizQeq/LREel+/fMR6HEWmb2eDuCHx7r7NM23ndqtKubdE6j08sK3Zr7yWsxuLpp
J1ch7jMJ+KLHHox9qR4NO3kBn9tJLJpW3CslIWCqJOAY+SG74tZKUTvNVzEmOFDtTQVuBfqBLbfF
3rCpGwtgyhp7n5JPWEMHcAyvtXF9QPbponjiwXsS79bkhtOaAQXJYjEa9GTUJUZ8hPfJb1zJVQfE
DqnZoLyZl3AMUef//zjAkQ+TaDjTK2zR6a0eV/81h0tJ9kgygW0yCUBQf/cqF2YfrTPuhlvvkbPk
/DD4CHHqCxQGYx7PRsDt6MWrkYiVRRLn6Lk6b6DPCeKTAWda/vzVFMfSwyHdNCRmDFlSzTjauXye
HNETx3KefLkkDvYuHU5FpfyYU862fmvKUwzdY7nKbV/V64+3dR/ejSLS3DIuZXrHRkDgt2fitPBH
1pM5hfFwlbBgi47yKbz3yJo4QsPdmyTDIqIWKb7FWLOaP3rXFxFQNwthp4PukMRXhhBgwH+U6A/s
L5aJSoNZbqOq7c7gD6/dTtn5q89EcJF1uOAcOflJBtlPhvJNXw4Boi1fVUZ6KlwIsHJ6w6rQu4zM
rmhYOGxU9id09P0/dc9s1YLHwdFMH1CpJ3gM9+qIBJXSFdykd2C8GamCI8bb0FDTxIZfPBB4+zpa
oHgOJ0bZxyVbnhrDP08UH9/tl6PaEKoYwx1q1ZReS2zQkwm1ArF2tkcsM0sl5oBjMoIMOaSK+sUy
j8AXv0amJgAdbhAmRhYBQKRQzqlF7pmAWzyXq5Sh+1ksvM3BJfArExqg8OIMYiF/DaARnSDEYoEC
qsgqotKgS/md8Fb/kia+ry177vJQbuOqUt5012f8AQpVVW9FbbQodzg9dZydaAwcqwhi8E2bHF5U
cHN2CQda8SAMvn9pDDh4jEAxjThXceyVPirUg1uATT9iBA2MSRHDf98gPGCRul/DnNKtwRWnEOf6
0QyavZvmea+pwSq0c1zqerb/PAQgv6wBZ5HNB+FA6TcxtnWfjf3aJuYE2cVScX4GkaCPR0wJTtEI
u2IKaOcvbpSHUZrokItODApsNXyh2Smg/epi70ArcZ5VIHK4EBE+6QtvMimiXTPM1oNU1MLiK0vx
oDOwlEXsfXDqVTJCAlqJNlUOgNLfVlWD7VsxglN60AjXstP+O9LO2/bSNPUAc2rvcOiyTY3SC8Cj
Qy4PJzMlQXY8ZyMii0tSApBeSxJdCV6dzuGZwCrOtJOiHTSaVVIrB4XmmRRiF0VmjFoOPA64VyLk
qjD2kMHpEMM16yTGpwMNXpg7XAqWGX3BhdAWl0L9NKLp+8HRDLUXZ1dnrQRsfZduNbYvZ2dcSLRK
AiF9BiXWqyJLBYKcPx+1fSY/w+STk4MQpwKBUI1TJK00k97p/zb6oLUbR3hGpP/fmDoTwkF+JnB+
dyU+Fh70DbU5BaqeSamI3pH/fMxeC+oDHBpKERX05bTMu7sqfD3N9ibsjUDyO2HFgyPBOO1f+FpI
xLYF9rWQjGwMtKGaROvqGKCW9R/UH1/q9vg4Q9+xKTOrOPYLgKEqrUZVsRNdSU1IsuQ1O1iM8gaP
UWOqI8vA3zwEqKR3bfywSvnIz57EiayO7JCKFf7xm+4QhfgXen/GT3vwZU6NnylvE03Gh4N1bAXV
27hRLTGw4YXJVxSyhmIO1R2wsfJJVjoDK3GcbbfaPLpnJjyQm4MBa2bER2m8FPd5o3tjFfJ2HW9U
pgS+Z++m+/nhKPgiq9fwikTVMk4qumqCHfvhBPmYOKfM7Td4n2WTV9L08JZNe3FS5G0zmDnDwMmK
Pz3EpRvPkp6z6rCgp1QNEewzfxE2WeWxDY/HSRrxe4Clbm58m3X6DqozheKIr7ssgY6vL4thQJu+
tq3exbhtcM3rHPJhpmMe23eCsK8xo/QfXN11gU/KIXgCgN3dsYL/5Bm/CZRfIU847ALyRaEsOLNp
8uuwOo2ImW90y5VUUrcMtx+yBSz4lYT6WxTMpIYutNoLjSE+knoWpF6IUSOU2tjAfCbTCtDSiNZD
BNmToJjIrI1sq7y9pO+MFKkrXL1qbdZe2ExjcvlbTlbabh9wUW+NNU4ZQX383rL/Vj7c105gM1H3
SIZ7JhjKKXLirIknNaEXFkA0eeMinsNdbPbFuoO8XTEOOkv1lJIkasxXNCkydpwSd9eUHg48jXXw
TNl2GowIJ//S1f/iX2qmwKaAl69z1SVXG0fGvIGeuWc2kapljvCuwaKPBk98SS+sehrkf1/EY5Gr
G8r40lkcGG4YRLHOaxUvUTXJgRcriMYo+HSWsVeZUUuFCqpzkGFb+3gvAtwgwj8DOBucdImcVBgd
NrKFnNYbcQiLRlIuNoncvuzokgOBvOeQ3YmBzC7P8+V4ePAw7PEcPNe70WdrfZnCNbvJMwYkvkjx
xmBwG9+4EqzgJqPDh9U+KK8fXqXng4zPPrmtDzmSCfY3lUn91wQqVelwR1uRPH+S/vo1msg/uGEA
yUP5+Qc4spqYSep6CWXqHXHbGd407NoBtu3nrewFH+Q9gAmpBvAcHJvEmpYfOO1OLIwEUB2ZfHSl
2TuPs/Ct60QoIUJAxEp1ntzL32zOqPnnHSS1KTOOIft5WzoOqkYDbmjV3tED9kZMOqYC21nA4nkU
G88EL62cmLCsmY4gTLaMIH3ZWw0gqPdGNT5S3E9uqdxM6VB4QH7FDmmp+B8biq99e75mUJ5xrPnR
2YHFHOPdOvOJhQQAVgjNIAK8mSn87+YYwkE2MaJhNqP+esJUds2u3p24di0IMw7BwhD0higXAgTr
Zst/ECDyx9i85i9G0o40PS06ctWjB/cUxS/uCBcIVhX0K62nmzc3VczH3EupoqBPl3ta/NdGCqi9
ZhHPWhx0hWwrmXGyBNEBz5bvygNzZk8JNBOAzYS3m4v4DT2BJTg3Pr4S56tBMCF2OHr7MAna8RQk
bMWhg+fkh577Stz045u32tyF4VFhM+kaX/ezrfrBDc0LQVOHVeQd/JTY48bNrAqSsWMBLd4IkA8Y
VmFBMP+BQJbhampu1LjFQCJ4z2atbGNRCFTmVJSgv9x2W/7eHImN6TAS1yD6Dj9ZnvqD92bljvgf
ANeRrFYobzM+lldczfMCWXAvfrVOjz43IPelKZwXKq8Z1cYtLr9P34QWc9fqmkMJr8av+zqLN8Ss
od3Lwx0l1qHurGvUciV0koKPecajwTtCTEaDjzWufuqtZ5RagKs5iwypXCVjcHZjDVKIjA90G8fN
sghRa3OjtZH6DHxct+txCRSp7PMjdjcnSLzUS9PU7F9Z+KFGgZeX2u6jprssWD6LNMgk13AaEt2R
m7LD1Mm1ERaAC1UDdnCT3SXEU2iAoDISDDH7kWPQDPCAkw8c7t58aO5nVsk5pMC9KNL+o3Bh8zBp
9Lrps8URrtsEtWh9ep10p+b8wZdWdo3Pv4O3L4AmtCrmUCtc12AFC0msl3lqFEqxE42e8OEfT5iW
JiZ7k6iyW/kbDC3dAUdpBOEj9gNW92kCvCciM/jbrXyl1f+NtC86th4UN8fv9Wp955PM5BGcEHP5
Kl/QSTkGUbQsET3HVVFa3EKOdeYFLq6Pd31D1goulGp2PdByM5xP3IumRtB30xZfeP83Fqad+/9N
K5QbQ3q/xqiEhMlRnN5K5T/b3Bjm619oUBgf/BVZV+Y4z0f9k8llHK5Gi0yLQPsY+vnJh2Logl+i
McCwArGUJNMDTbLN+GgrGsDpyqycqWo9J2NuIF+s1JSesuH7AjjnFHwfOPcbWPPSF8ZdvdcNiblA
3LAvrSiJZcTeb72JnjxMH+QKVgWsLhzm25EUn12+p3gmfsww6UrZjxZXXltf9BouAwGaPyFF89ZC
7ZvnRhLJAyFdpyv2X9gRJA/qpIN8B1388VhJ4n1zgVs8Fy4oLuo2pqLtQLyQZe3plpIqB5rE2MLP
utjjvLXf+JTCY2qx3Fl1pDAxh5veqyak37nMtax4QrvysiSKtgj1M3TdezXQzmP2W8ur/n/a8opZ
TBWWkneBj7XP2FojY22M1NgPFEceuvR2JXDeOAULCcriZ73862YlvbolF2n0pamUVzsnA2wPQCch
4b4XWh/fNk7HzSR9yh0QkbPByLdSg5S/OtXewUpFY9mh8qIClDy6SYa0GyAi0nX+Brtryweb00Ej
ssaJ+WXfQ85a+GC4Oefh8tY7DlwC65t7TLO+GiWRv7L4Ulz9A01iqWHv8b/eYyVJpqpGCO2y6bB7
/zNR9w/5Ki0Ors28xxT7lQ88nnRyIoNcj3DA+yA7EAKw2hAjcCnxD9Id0YPmknlX0G11yt7Q3lns
zwZ7gozt7IXdL3G1ho9I5ov2k3fLzs3LYZ78BYOLo0YM9/GgkfZn/1E30c48LHVDoZDum8+k0MmH
3sbSm/fHGIE7DwGzDWZE+8GQ5vUDfVdrpVAqg0sUH1R2N8JRelKTziKGvQVkfcU8+PzbQz/fm2n4
BVEv/vBAQ838XT1Pq0ojEykOH/+C6hsh2Vi/xFp5PZpMBKTjuWm4qY3FfWzpr3JPTZIgRtMMpxiL
25IJ1Iy06eGz9HAIp6gNvfNMuuYHi3fcEhOYHBtf+9EOrnmBkuFv/xuqYTJ8cN3PYRDP1cfwOslW
lrWCgsNoYi1bCyvvuD7paEyCGDAMprzDC9jRxOxpyGnPKHypwCScfa20vHs3zo9MVxxJYsGC69tv
psq97wP2F0AjihbedjhyROZ6H+nX9GlRyuEL2aukNvNA1ogO6NjuOC9xWx/ZpeM8wB3Z2LpRiwnq
zSRDOXpcDk9+XkhhyU7ljC5DzZ+dYO/b9eS0oe7e/I/g1HYnsZnvVjF6vtWgcZK2UEXsJF+00gK0
m8o1BoZDsfXKGHP44zt/LtsEd4oJY2mPb5EB02daKToCHwpTLcPBrmopeD1bLA1k6TY5UQENLsZU
nC/eoOhqaYYmPuiIvrV4akf3+6z4f4259CdJ7a+oS0TLITnYIEzXFnaolemV5cXEl2YrNKoWjTXr
B/S/QIa2sF3BZZPXZ5GF3LjitFlPt1UG6+7JBZCG5xyDppHrTMN5Ahir3Qka/qzFpx8ShWn6uPNO
UIVwVYUZnunwfSUk3AkYnjoEApUzZR9K+g3GMuKvNZE4PfwaYwWblZRff5H+FNNC7xAYTfKR5Ovp
OW4ju8azF6WPHJAMR853SzlNHZ5fJNlEMf5y3pwjgs6gIX+wvjGTgWNTa8zx1kXIMUi7Nw5KnLLs
fnRPNdJP+r3ZUG93LskYF6+51AavDYGAlIAHoZPz/Z6Gvay6oRp1QaPY20O9P9hTgegK7/FnFPSg
Wg3Ah/VaASILWwHPQEWjasksT6/XD1m2v+xp7HV6lL4UdaUeA32bujwnpSHB9y3pvhvUuhGryZ6Q
bsbuBJcNTcwE7EQJEIPZ82auT5JHWH9QqCCVLICv6ihjC5f/6HghdRE3QtZnGF9y25yRYLYAaF6n
8PFtHYKlP6S8AMjI0v8KYfMR1W80penXmWiktUPlRvNMN7G4er7FINaMQyH7MwcAisYstbyrGwO1
NZHrW8MJaXOXTysdlR8iQK8dkJIPRKiff9l1gGblNhfE5+gzCYAwdtyVqB0r6mSOaHgShAoLW6dv
fIrVMv5WsAeA5MWAGWP1oXkXFXMQSP24sS78OJSfmjH8VTI/3xrvzgZbeqErArfx9H7edumnxw0Y
OI03CAkhdPJEXE8W48VRstnAzvGVmykUwnQBG1ltyivpbAPoxz13b+Z0X6dq7QxZKWtVipFwemA0
fK0cLPEukwkGaZreBfbX220ZGElSgdBIp+kZqm/1VDLp+Nf/Etj3Fbwlcl1tqHLI8Fa9Q3yOQQKx
mpR0od2u2Av7h7Fiykuo3ny9Zjg89YNNi4j1HkDTqQEbDzWthZylV4OiRLf4REgs3WLSyEeRR6bX
gsMaSsuPIB6uwG0wi9V9eutAf/imi4cbI4gFOI/EqWnC9JwCwW9TMg7I9hZn4LRL9pzTddThvaxn
ltAWaDYEAovQ0ZJ04FHFE0TvxnEVKLuZDH0KH7PtBP6D1gtFQFKfxPuNfkJ0Hdr7ErsFFdO2En9o
JRPJSXm8b2f8ZJCRWlAxeBk9HDRzkHlEpDUhZ21gAd77/bL/YgbBh3UN+LJmI80SwuysNPOx8PV0
lGXTDbD+2nneUP1bzIJgsQ1I5pKpuQT6z55wMg2KhM14I0+KhSI3WUOgbEiGp+4CKVeluCve/nzL
BY90UAxKbraQTpbDMQ0x/a536Dng5NBnE9CkxgdcIyOq7UIpluMPVUAfKKsChaFo3Fqy7Ouz17MV
pJXzNpXHR9AtfHs77dLSq2lhrcTvKppWpR0xMUEZ/EJ6we8+rCY+2d1MMvgFRdgfmuljTe7jwO9d
m9PMu7D3nbHXuUAk3c+aEZHlKSTdpxUUtlYHeSW+k4AXwV3W7tBggi65b9sNEywSXU4BJ2hqIHlg
CFi7oUkgMkEoVKine5t7AkmROH7a9dfbu1oJ5rxzcKVoQ8TKd8FmWLqcJd+ipvPtZW9WJyc+PNUR
m3uLcXb58PbniUZn0ddZPJERW6AnkmleZnB3tHYolf1R69Q4sFASmmnCnabDd0aG2VLPE8qN5La4
8syNlmrAXQfpaFuyVjxKAC8vxiW9OEj48za2AQ30+gmEWIf8K5I1EO2mAXV6vkFEvmATiRP+2o60
vmVhZu+be45+vQL/0l03FqWUT1tS41vfpQJ4+6IANgiUUkR9l6Ijj0hvYytrCMA6BI3eRaRSQVeG
q+YrLpdxRLT84ykzEc75UgBlPOLao4xY04Oj05njEfXKcrYVdGUuIMSx/C1BNrzkSZ75/jaIe88C
03j1jTYPqw/pTo3n/OPwXYVu4wAVOeIKvLlCuZZT/T3LXgN41A4+8fo2jSJ5Shqu55Ofhp+HXyTc
MlrnBPF+JDrSBA76lcHyIl4UAOFFK/S9RXx7Vo8u+MJrD7V0XPjjPybAV4wO1ANQVi0EWT45nDo6
3wJhU2eRr3TtZD0QqTYIJqagJ8ve7aK7R3x3LZyjEs22MTxT8iziRQpdFYUhTavnxMdf325kmmBX
rBrQtN8JtP+RqpOQ9VuqPnW3hI29j2Vu1tbs859nW2HfhqcgBKilPOp8D/umz1NSOJhFwKRKLVuK
/CGFDyyfoW9HAcCnapFk7U+34D/dvg602VxOMkbpI06bqe5C/gL5molyHLkY5iR13uWEAWgs8Qsw
dM+daXtPHkLA+9077eLBLnXMJ4cnn+CdKnUj4d3SRsohCDpV0lNXWuZcijVEdfWX+WxpzXzcommf
gsxFegm2MiZImDe+pq//hBsrSxM9rClQz55VEQMqfNnmHPm+xZalSpYC5MfsWZ9K0PThLOYgNe6U
Un//x3C7sMIHHmELSGQQdWIfl0QwMfGqjrX47u/esTNoTgNP6gjjzGBn8bENqGFVoNUdti84VC36
0mNXyR/0kffNQUZMnfELHLiFlZnumUldKn/HG3fyqBO6fvKZ+zrfuNELK5sZHzyXKWc96R5g4+Fa
nAuQYThcLmHGddxL4hnd4h5D2kUh9KjRVyp2V8voaQtE2zGtQgIYUDoxxzaLm8QKoOpVlv72k0/3
24Ex+E4en4fDe66OGI5Zfe+AhBkL6amhK+Om5qQDcy484i+yGmD7O8WkUhCLkInEnfP1+HxLsVZJ
lov0u2ftOrJKL24PNMGJKj6NOlEBomfiAlUpX5iog+LXSlNS7w98IlbjUl68sk7tVsAQBGI1MG6G
XEv/Nw10AlLQTrw1EvsGUU7VI0i1T7Jin6sZdYuOXnr0IfsVLTLp2YuyIaYodXX1q2Ny6bj69hqE
277+oeC9m5UYYMHJs7/hEZW9Wm/c+qFcDY1yScdcs2YOomFtMNYCtdTOGyW249Cwbf0hZfO7ruWh
KJ8UKH6RPDQBJeIBZcbCbo+ldgfqsmJA/I5nzPLmxGXvzK0YPWU1gBoUFKZjk+XPGkHdzzUroDia
BEdjqIJ1/WuEBqif18WJPeeDHoRX0KdxPJVJ40Fjqu9SpGBy/mWv+ZYqISbbnoagR1H0U+JQf45m
OXkJh/WM70gE4PY1LcpLXWLf/5qXCYS9gnq8L7tpvJItfujfQWFBXqvaj6RWtnCDOkHOxnTiICyQ
KGBODaCcjuwYb5mHTWbt5ncheEzZlrCusFEsxuHKWhikkQxnepcev+9YCoH/Rz5pQRmSVu/flkYo
YMNVqdbasLDCar/ii7IaxVJB2OHQGCz51zsex+3olsL78VXDqVaGNs/DyO91omW40iXfPRdTNQMC
kMfiloZMW7a0IzPfDwNTRZiC9Fv5Yi5yY4sTRTGvIelJ11D6IObhGIK8c4jFwlFLTenKy//CB9Zm
rOshIjk++oXTfgM90gFVMfNm49rvvn1pfMfeLdLgDePqJj9+1mw5zDf1ICUW/gBPxYzeTNfp+/Pq
A8RSaL8BZKST3YBrsoHEYWfuk7G7xutTUmFQ7tZ7rMmdNNLvvnB93dsJYpbkVJgFp6I+PXowwGN9
9gcpWvK8lDqUcgXcAjuzN4JBPzDGBPvZwX9iPxTQu+YEDKaLDFldYMx/6AYNoytq1LVQQUpyvNZn
lZps3U4PFkO8clWAd/ZStHKO4Nckunjz0VP07FPtY3942J1JgFiXCSAzA5TqrB9S7Pe+Q9bKcN1j
HtaaGZZCX5dbPHnv1HEfli/we9sdEdPUnaJcdaLOY3HMwGHrlVm1wx6x4oORjnwhLBUTLAObWm3a
InT0kIDtR24ivZJ4cvtL2G+ooF/FHpzjQOY8V5PVw6ywAtaizqVvEkjpkM03zs66OrnhVP9r/xgg
tkqtKGuxug38E2SDqSe2D8CH5nDipsEgJKdbgOgMhiz9Zl7dWX6KMauwioegVUlXyLPTWa6c8bTE
Cs93L/YppeDrESPAA6FLrOZ5TYVCH/STkbpBxtw6PsZo3FvIRTqX5tZHqgvlBZnm61zTnR1oIy+a
u/oDMY9n4ZeZJurMVE3nM9QcYM1hTkWSNsJAWdc3C++mw6hjKiOY0fTyU/ff/uT7dPF7Vk3xVSQk
cYVLFPOzntQxrA4hVqYa3vOokSWnOP7IfPCPEWcNEeaWmuV+pwdf7dLuOgBX48DBY5+0zI8JHcVi
n3xmnLouOIT4bPaES78s7wku8jsVl6T5TWsw7/86ba2kCrkImp3xWLWm8lOnkFzMVsKFASWa3C5p
/YTSJyebZQGpOABD09BnHH5d/dSU63kDdQzXshOl0pdg0qqk937g7NYulSEvzUSHW++ICugYPGW2
+eyqyI0iYUaEy16t++1MvsfaUhNrhMOHHrDypKvd34DvFyxkSffXvsspMJWLMLdO3LdZhr2cGfS/
qfNGEEbJnAPxgP1WPTgvQzKTLPiHu/LGEqdk7RBgWBWnesAjBEmPEMk6VZF8Ipiq/nDXKsBswyIu
DVUPIl37N2TfMJhXgIc6XHVgxXJ8ZrKUxWs9554xtkHhNWVaSPmA3PYE5pTDNGF9X2mox3gMPdIZ
DQtc/lDxPVYoAU+mTTesScVXQV9jVkXc59Rp0J2eLbDt2jVdsSIHTFbwGohqmRlBuu0GtVA8l8oh
8EznWzfEB/xYn6tY4UD7xG97zYlJcR/KY9yR5bGvfSCEbMBHO61zxGn6zni6O19JJQA4rMk5+XDO
4ugbB2TRD3g0yiLo4eJwHia9hjvnuJnm5e/BIwc5/b3ZYLODF9RnVbOgN0749xWGQztNMG3RFe/e
jDAmdfWkvjrnqKt5/da3DDJwAIJz4fEokWwTgJ2E5tbDnR8tB5R+kMNd/W+oKxQYiQU367z+y22s
H2NXcFllC/ykkeVPkuY7dfR0HValbKUPXiymsDTq3Mbg2dBkL3zgUDVD3ZfWUvt3qedEem1zy6Mz
Q9gYoz1ASgQVpTG/2H/VTLyscLwHxX9hYtMl/Ps9u1b/oTsuPyOuVoJCDX/A0tvNl0CnX/XiEIEP
8kcyFfqs94Std6HezYpjkFbsm9doB20VK8AaO0flEMlqo9tDc2qSelO5k8gcSuchWXiwsVRdK5Lv
au7Jt/daFP/AM4uYcUWjr68uz98jbGFqNfoEov10jF5vxj0jvh839D+py5pt9vMIJHIaXZyVnB7C
nS7VIF91dJde5vqsbKsHVA0GTk+vbOWwhDUT6uqGD1rC06n9QS2G4CALDDNHpNDhNA+YDyxlMMbk
SFHmpHp8MtMiAfbui0EqXLzc9Y3Mxw+pb+jP/Hrnzdvgd0c+byt/YM2gj2MDcSHAcdUOtBRZ5CQK
E8W3Bvq1beLGxsjruFzIrUG1XLtC7UixRNjWXIE0kTMihDqPRKNpY5Pr6qqOic3muot9H93iL6x4
Shdh0FCzIT3aQchyFXabqHVvHdIIc5L7B+lTkl7ZG1h30n3KEAb9wi6+UvOrKf7SNU97/b4l5UhI
JwSDZ5IU8FdiMrEb5wG9ql3CxrRfyJPTzl23TJ1eKEFwQIQDo6hM1F05rylRKeCwAK6acX5wed5M
alMSBJXl5N7QSjAx3sgILCpQ0ikAuI3yvsLglAYukRGkq6Bccdq87jsgR6xWqggWSyTZ5chfhUUw
YJyWKMjc8XdOueIfICFK/wA33UfX69AM98rf8VY6xgklUFFnIxdHOstw0a5Kh/kygJ/1d5jjmKqx
5ajOqPhzghuVJNtJQWb8+fs5Zf2z8CjNgsqXti+GogdMjjcs/F2IugPDG3IchuBC0BES2sOYFVwH
h4mjlNBq3XVhbWgXUZHAiZW4HYAFcJYj9A2X4WwadwJkRAahLy063CFpP8VvwACGZ7aVhouuCPI+
WjWkVy+zrwFiUsuvh7k7YvLoCyQDo6biF2CBeqnEBoen2co97ZQWBWjZXIL+4EDse0mdALDdpyID
ZePwPFYaveV/JtvHSunIbXXdxJdoiBSpCB2cfhKzkULX5kyUKQXH6E2iD4NTIN5hkovddg1KM7lY
Sud1Lp4S0izGB4pKTO4iHKEE63f5hygPwlJS2l2yoyA+xcMjGmlV15xoY/GaLdJllQXyC117cKX4
LExdoN37VrsxAS5u0EFvbuS8fqJFKpNIwsRH4FnOLPJTQ6l1GaboDTCmmDA1ADUWZ90doiWi12LA
ih4QyjXGPfiRJMc36kY80G6m2tCDmqTrdqFogmKjrBFZOOLCXHHaK0/xdsK7+plRxbQk2DFrFCo0
ibg1cfT34IIRJgc0yyvV7HGPH3KjkSOAqUhRhUH170kty26wp8huvDHkwHFz9yeKBQ/kW25udQOf
Oy5kOPcXCbDzz1a9yQ0wOwgEWOP6LngMAYpQfVpoK5aUB+46eiCbtU8G472cOVbWeFi5ijJbiy6l
RgYmpGfRSc/JN4c8BR58U2mA2N/YbCHo+Y0EglxesMdVZzNg5jRtDnUlBj4OJIFKA7Gk0G3RaufE
PvbZcEfPtmXirBoybJdsDwuSoBCjC6kCILGr4ZoSesMdgQnAh0YbN3AYKag2glEd3uqr2XFt0r3r
5Jjikit5535fMSefH71WhBivRXKBylWj6QDxRDIJnI5xZAr73Y/Q/lmE/yopU6tJJ2g6RLN1+n2A
yzkbNRBvmf/+qkA2tDDR5QFE3IiGQI9uxMgF8PaBYg9mB4r32i7JoV++h2mLAjNV+J/FDu7AaUoS
8r38tl1Z0D42EsUofqrAmI3jGzlzDpRP/eHqSJycUuRANDvLXAQgh21lnslhOdJ6W2XKX+MQGE9y
whrYs3ylc/jQ3+xlhhP7yn6tu5JriFo8Sd5uylHjK8nC2NeXsoMiuxDzj0R/8hLQ+IpDHwKODiq4
pRBSLo0Hp8utmgwYkavJZJCW1+au/m3+sKmdW10LEIcNnterRvIKrAybiNHtptEJ3mwMdiQxx8Ol
XJxRjutZSuhw3H2iwwSL81FBMlnWVZBwDtSycERqXo6O5j6cyYzscYe8RvCVmqZYMuXgKDnhtu7K
91+652HDlQwK3hynFLn6OXpdoIk+rzvZ2GsRvhBCE8Mtmn1bM+Vbxex/QIrZPJ6/hn930KqTZDgY
20jtjYKhts+zAKHpdG+VrmSqvib4YMrMp9xstCmndCKKtNzxSPm92cSCcjOwt25QeDuUhsjxldkz
dN9EKjaKJ0SotVVgg7k8dE55x8fjkPfX9pFUOyUOVVfhJMbgiAE5viVMa1VE/T9Xa6RqzBPjz/Wr
1kc99V9/MwuVXrGOKQ5qML/KfdSpKVDbP3a5bpYW2TxcwBtaHHy65XwQ8k0aE20+f8s9UV7SHl6x
v6mweM54GKe6jKGc6k22s4fiVxLTSLpegrGSxCQKm8RT0XpWhUyiHTOST+O2C/2lH9Y/4aB6qZE6
06jrh2LrmHqwc5f7iKagRGqnvY6vA4W6veC3acy1fe0VRLBveyAVVP2HOlH09/MV8iRGbjp18zUs
REEMYSJD7N6o422XTIfowraVfPBFsB4mnQ5pjjQHQfVie+mupLgLzNd/m9ynktTE+9EwSrtXAwOQ
MLizKuL3eGXnhZ3eWipJF/NGNezkVwPBFjH4VbJRW7vzg+SR4RjfI1ZAh8/XFNuP/ZcMI7vYMqBT
5nCSW5CKsvmpNGJImNfHfAUmpYDrTVG3EOzBhHXOSXMUdWwSEsbDqgsldkv2MahvMlZsQhoVpCLI
3FbkUwoJg+7HVXGVLXTqNNzs2cd0Q79Uow+V5gyUn2ctHX4zO9E8gs4OzA+gC1y59j28Ro5A/0gb
NdgyD1s7TSSzVwRgEDHFzoMxVpMDEvoSvLz8KABgKwyZWtLwv3RPID22+hfUZd+gS9vuhe6i3DVN
qvSvvrDAFkuUDlS9O2jE/WHscpwnuWRbw96fM9i8coJC38sAnX+K2+DlVFjks3H8fy6j2CVqVUJA
SPYGmX6u8mWjh5RRgEAaP2JkSQcqw5A58Jrxywbo8y1rjnMXFTAfMv1MadaDffOgUQQ/TFpoPz5b
XBuo211XlOTngc8xJmZ1nHjwpmD7CSHQTcueokkI2B3KXmxavfRnOz5r00ug2CnUlgwB06tdnOxx
3C0scili6IIwdxNxRHYzGC3QG7aTsiZxLXc9ogmrjIsQbsksgYEhZlZgX1PzkBlDTr1VH9Igitbi
blDBCyf0uVQ57g1/dteD2pvTsaTohy5YD9lscOH50VQgyrdLDRblRGR9HvfkYjqT76q5X5d59H2P
uCMcOE9WfcnsK2hcoR3maBprV0xjb6qgjZdG9WU7MZWQ6M4EYNT/RpE5EHbXbgtd8Q5vBvxugAmV
wuuT1dzgFIFT0Xs1EWNOrjBDgqJ8Fykz71J8nayMvwJttmSzxO1Fy5LQlkpvNIBYYf5swv+1DXIk
FHFlHOGkjm3hg2kW4r6PVpkQLXXFpNDQjqrATGie4ECpBQg3XeBD9ToD2xwI1K18hTKNuwk7kL3s
1eBruhYBMFwUyx0APGTFvkk0rizffaWkbXn22GdMPsxan5kg2hn08koh45xDvnmfFYsYJjQT/MMg
0L/YVAxNS2FN7up8mtnAPpvI19ITLMFC8nx1UClc3hDy8MRs3tBrJQs3PfQWFuUDUmiFHY/ZTksG
iqEkxTKRoLGbgBg/UAuP6LzExv1gm0qI7aW5RlLptziIQBHOtfFiYBt1W4rl3k62pZLwsG/OdDZO
2N6vlRsh4asbyP9FAKYJ5jdYKRGSTCkwlyK+n9viE7eQcrRTRaMR9YFg49hFdUZ/DaYPWfVV6oLL
Wdabjjmx1Ui/2+rp271UAoz+wfPs60BJQhFMu3qm+dg+7pyha7HTe/k+fZQ5X9ML0g6G4CKi5Eal
DaaV5Jatq8SYQHfNm+Av7pNlZN/5VLUhYuPHD7CV8viZQp/WsKDHoSYk5rhuPndJUNkETDbUC4hp
D/tBat4iX+vvgz4sc5PBiaJPp2AErpuLZ4CpmeseJQjAS8lutRjNes63SrkAs3WP1SIzW/qHb/Tx
3S6yJ8OwUT7/Yc+sOgEiq2iBH1uAUQ0TLnfcVM+tpdnHVqZN4V+mugPMNp2/c9DNcZ630cc/iDxc
q0HbARPYfAwsHMPdHFWH3EtMNG2AJ7r2BR8od96bgx3BqmpuSSTDUqA6w60YZv9NxmtJIyIq0ryU
nu2k0vMD8JoB8uBykuXDBgpegNgmVtn6ITesftWR/n/pZCUfCd6HGf6TcAfjiLcDE9HfKke4nRNL
7BOM307608Ctw7Q0VjqicLTnORXe9dbky4EAkUTR2x8UhOeg9TM2lI4oeYUALDFMwuk/exmmMDmI
jOEfkdzbPYUzR1VO/dnMjtFQ7gwM5mMzVr3dhyCFDNzKe7muWdG3itJ1STAQkEd+/IcGxeoCqDDs
O01PcZlnnkfTq3kwCTKPHYXkgCCK2OQ+BRmxVKC5R5iZDmVQfLBJ5WqNne8PUuGdapkYoGAzZ3QL
p40ii0z9JUVsScv1tHuoC/jRwFUQbvYE/dwTZfOazpLqdWxtoC4uexcxN6dU6RgHQis6ZK9HtrLJ
MNj5mqmoMH1snXV8g5aa6sNehNxrEpwliB6ve46JbYWUXtmJ8yCpdbL0XmgIKI0vCxReiojNfTBN
KCyUMwYvBV9qKBF3eCYOzON0tTO0aQhnOK/TavJB8YVaTWM8dDCBR0otYOdp/epfhs+QnBpr9IXD
nq//cMAoBoHfhuPfKpD6yKYfw9SPTKroFrpEoIRrTg8jl7q2vSj8HKsJ8x+wvYqAHB48/eJK4izS
uYv6ouyEEIY/AUD5DpiOd0H4cE4fP+FHM2XaaZN1hgWFsfu/hFFsEI6SJDsmmmkIFM6Bmt2dE6/m
YD1ProAY7/3SxzYhpdy0r7VHGLAaR4goxI+L3Bti3uqT0Ru9oyh2qraXBk77iet3bJcIX4xsf7mU
Yq8tYfaOtH9lIz48iX8Np2hpcw/iyrt1/XL+Po6Wx++iSCbs2+8XbXyQzSKrxW1166lkpyxl5wez
GTuGXsdIvn9ZztIsfJYvP/DAfUq+PIJ7bL0Nff082jhaM9FjAqANZxFdL1akufxF/VDF1o3gRnxb
vjDCjvYh3AnjS5KAZZv5ex1a+gsOuFXa93ED4Q7pbdE6MPDvjRAT3OBlu2o7htHjYjhVr5JP5Eca
4yTeZsnTx8tyATpxPqgSKZRhJz4DkziXbEIQnNYEpfl1AZxMsQhk1f/0pjNOdqhkLejpRSng31X6
afsm+/jM6edCRLc3eJAoQDHDsvfxwKwn7rARuSAEaIA2B58d3D154tPHdAXKpyRXiAOT8v9taNY8
Qhx2+9x69ZWiLdvZkZVCKAEvjypM6V+kwJutp0HwLiyNfzNJWkr4Pr9RhN17yyfY9OmSPsgGYNrz
buYJmW2QNbYvKvYPtbu0a1Acb21Ky0vD2v47BAKoLekNWg1yQOrovsjC8AwUEdmv1WhosTwaKeHh
zTobrKpvysHEVVlqpzqfSpK6nj0INE0sTPd2roqgUqAiq5/Fzed8rcW0c55lg8OqBLxog7odJtr3
qUpw8Zu3rnJ5cBYFPeeccBJImzLbCGRN3Vmhmd43DXplDlPbNcBD99sInagbImrxLvbfvQWAMk39
3xnFhy1Z8WB4gYoNhNNo9UggS6V0HFaLGy+74bslspoCmSST+QOSbIGXrrPebYv6KU+A643K2FUI
ossgygI8glsT0SicN1/61FU+hsgXY6YR7emxMlX0QXPBkuvhcIyb28SCynj/dL3BTlvVKsgRuSt5
Co9apBykKvPt43/Zz5LTr66XqxwHom4ZS0cN4UqaEqy0eCAE1HBaYE3gCgaWRvK+CvC3ny+S91WO
WpPl4ljrLqROdczT6v32EtIb6qYv5Y6IMp19ZtI6lSIZqDDlLcOZw6DT9XIKNgm0pFnYxYAnPYGt
Uvx3njMlgyzrpaKAdB3m4vBEQgZrua1UA9nkNfIRiiJAC1sZxvpTJ5QKKrKvyyHSHlx+z7GI4AB5
LAmTa4YHT6rSttl3Ui0UQYcuZ0JiwzVZsJFKW9LnvL2w3rJydqYemswvnTitk3p377XHJGA/f7Ve
75g6vE34yxVTQlUSngIld/tlw7kuGsAGArqOfqj8iPwtdam2R0WzEe0Z9+F43P0xBu2mw+9Y/rvU
t/cmefUWWOu+Ic3jc82r9KG4Kedu5nCjjx+UoDWggFUXtgFVljm9n23PSUtBkt1eligUXbVpoXcC
JTyvPOpBucKJVWvluQKKaiBo2C/RsW2Gx/zJ0yWzFXR6KppXUykhkFrP+ZIGiiz7UjTqlqp+rB8A
hFNQU+qtNIVeor/sOr+vo4KCz+lVWxCFr/h8G8GkirVfyO8w+X9yzFA3tkDgIqv7AqgeyQ4Yh2in
QFHX0LqfZv9It2hfyCvZKcpiKfFKVe9Lyh2FQ8x9I9QpY4jIPW9pO8vzJ5FtrmGNhgddZjHcG10/
LoNWj/X+iSE8cjGjc0jfcdT0cdVn997AhtPZl9GfPhy3RS/DSsgDneGJCJ9RhJmsMR/lxwp7cIgr
zbeciFA4viNfIboTez2aezvywL8j2iSQqFNcFXDK9S0bRp3B/ljmgkY1BTJsJjdOm27Gob0U/I29
g+QUZqCEnRgtLAmAalndHh6EU1+wPAkWPf6eahucxHLkZ5ZhbGA1mj5wTN8qAMmNYy7mgj5hdk0w
TZdZPGzdrsrN9ZdyN3HexXiPFAWclKTg7FJThdfQdlLWdeUIHHd+vpidwQpwcdjUs9132QKZAKqz
G8y77f8+jKGtRdQi8PLgFoxI/dA9PGlsBZXpX6QFCuDQOqxlcRggAFA+Ev/cTdNXADvTy3ZvI6Yn
ecqH14n2JFJJflbt+SgZ2REK0F0s1r0TOdINe4R9IeN4WqmB/KQbtk/WvsZKYrywOxvaeOcLeedA
RKewfxM2nmjY0VEzzZPoKndq+KbRIHJz0/iLREjOIA6oEl0LqGBHjK064gUOlxEAsMRBjY+zkf3P
yBLgOAQL6IQsAzbqtkCFbydyHOP5x1yts62lLtog7Fbmx/dKJFSHTDXKHEoN+1EhqBd2FX/K7Die
+uG+1uEiyxVKM9kpftUPLqyuBIdGgpsd9xbJar35+ZAHfLSG9xatfRHRok2faGnxsQFU/E4sZbJf
YslUNHyntjDNKRjk/lshDP3HwGNu6n641NeJsTNIQBgZUy/aL+5NPMPdfEgUUz63OejjkQDElIXq
ZXdyuHdVrgtL/C04bg1A/Z4QV2jQM/PyLOhV/15c5QcNffeO+3ZNmZcVUUbWH3rENYlib2c2ezoX
E07WvNg7Igami3yHQYftb51Ftz60TTFihIZa6blwZaCxgZqPyNkd5J8wP8/rRVLbWc9hgPSsBqYQ
Zzwuy2R0S8Vmvv5H9LRuuUZEKUJPTR0MGGErSbACcFsboL9oWIsHMGiLn5vqVHcmSc3Qe6zX/9Ii
emzSbXj1Kq8O60lY+Ag9H6uK2ahJNfaV2iHYt5PV5EgMlmkp/t5EtWZC1dNfaYGhQ60hNqeHxiv3
W3Yx6C2Y/kWvXrvtD8pdTkuOS8BBUOOfe6QRo5O9HNUk+GYqTd7MEaLxoRX9XNROqPjdlPOAD/WF
P4aPljWRMYRDVglqosWp6P4MnymPLosxRHIw7iTQ6xnlNaO4ubVPA5jDtsRBGlTlkfeUUJdqQxht
rIodSIrxt/drziz3uCkINjLgIOk0doajVP8UfPu6ShS51oRQ1O1GOkzz4CYsjN/61ucoW2cJxdmP
5Ebhejuo9Vks4kZ7UBrtVWZEVzfGtxKQD3nwVQdq57TuhvkMIoJBi1rYIsMIpYVH6K4cdst0dVDm
hHz8iPU6uyWms4+tzG65oxM5NkyjJmeUuWOmlcOqrWpZ8SOZc2BlR7fGb9tCrAo6Rozj/NBy7oqQ
6D3mkFKGzxOdXMSqz0zi9PNX49E4rrHYnWycnpQoVoeBRTgBFADTbHo3+6HIWl6P9NqI2ku+WP4v
5v69fkCs1qFFeq3L0eTu0ieivjGLtYz40fRB8+S32vH5qJCzGo9q96CLASVZjBQ918pZUtjcMtrs
ugasveTvlmsekmGa3/qm50vvysGgIoRJC3m0dGmuL8kNlmdRJdcIfT8SVfa5f+HqYumfNzFH9KtF
T4FsjUMJeFuMZDym1i0Mtq2hJtyASLeiEgequQpcDM4qNzJ00cWLvsKTcUYIDaFOmW6bXfp8Kx4k
HKZSLGCUlcOQSg6BoN0t5VZJwQp8njRqXcJRWZaIv1AwoJVwL0fo1IW/zYx5mGJvwFCQho2PswVr
dsAQ7uSHfqLbtF8aInKxllCC/q9T4mfh6mr+DVNMFcASsTubQeqvecPDmDN743ylQwLCMe+r6+jI
Rdq664DVnIVZVIg41rSuhvZLNjMHllrwCAi1/wig40yp8noCmqpO1Y19airNm6XGNOeLtLcv8dIk
DFmkPVdAGL6CrBrePtavxJdq8nN/+/ctJvmSBf/nIMKobPyMu9Of8asAYLL86i6phsV+pFmorSCX
ViVAMfLPcfQu1GZY++G5ms4y3tYHBFQP5jTWt7K+ZeABbV2BJ3fu2LhDkJxLoD89O/aV8CLEj70s
xNfWOSb7gDcSILGIIiBGm6Egn09gj8g8n7kytZ16eq2vSDps21pnNq+U5VUmDsbH9kCvGc/YidWT
7be2GvZ1WanxoI9XN4MAeFAoblPF/+yF+NGg9t8CRw6WBRMrAhtXilKXcrDLTBoC3vA/YPKSb+YZ
gTMNhS0le2SzTaQYC5UKc9eaPt19qtoNg+FKGP3Iw81c6gPHYX7shtcHk5X3P4BVc8cRbIV7EilN
RegN+v3Lr48sGEYR/W2Vhs3PcDsN2izuFlUPxBMAsAxiYkmOx9R9Okdb6oAXOJk62A5pq7cFTTgh
x6FLY5bfXso9/lyrQUoKU4oj9uWWEfvHo1EbNG/W2XVyeQXr3+SHEZdNYWyXOXEQv5qafTGeTMSO
6iGVgyuTq3KTKvLKk2KP5NKSNu6AywGAuqAc8PsoZ+K6Hu7z0ZFtFJz6L9t3Q8wBp4ToBTzFVklA
oaEKTVQ3I8FEFepjn5oRrK5iR6q5qID0vN90nE598V8gCKRYkriMWrRmQtPl+G+/rwmS4N6nkxzl
+DdOm6Ml19EtMgadjitIDuk0diYb4RWJOj1BfRY4TLSfFqRfFXRMhoilW5YzvyAOihA6drwkFu+b
6JJEvY5Kk2wszOEvInhrWAWGRyd0kftuT+2Pwq/SCoBtCNzoX1NsxU8WPMDbflqMuhEIXYh5ifW1
KFpCw9l1Q2dAGHySeLZe6gRAPc1PdDzXK6IxKtazIhgcO/N5zAwlZG+z43HktW3A0/E2fB7snoAT
LNlSTw1WMUvv/qBIc90vHH0RxIO9FYypo4QFJrkjPMubP7R0F7RwX7YxNgdUWYZEqHv2eTBSjVMn
OweeujkyDfKOd3TK2i7f7esXRaG5KhpL+yP53DNngMANqTaam5WlJP3Z4wiYeKKds6Bo1WuzA+UY
wNe+0PcKVp+q3G6xUeANo0JRgQrE0wNroFi8GDvbo3gMcP3nL1jVuvmuLRBUP2nOBgHWdZH8VHGG
eeEf3Cuk4iHTOpAw2d3Kh1kQWRo7rNvHS1v4VrJ4SjahFiNm7kW7TdAULwREPUkw64nrPBtlt97A
mlQEuQAu+AS6hxwhXSwoI5FK1UeItzp5AcE2KYZr6jErPBdGJ/a2TRJqiQXwJFX4N9OTewxOOxnW
mY4tg6yw+lh5cWLCzAmBh+RFr++m38MHrh9kR9cBe3jf7ujp3FoZsPHhO7pyT5ERgq4fWTdGDwk8
yZSSEd7FOpy6iEcfQJy9wTqd1xbey+55W46xpioQUFxtgBcGaJJ1aD7Zh+85qcNIw8PK0KeMiJ4u
w0aGI9QCkBnCZGczC31yWaEdORdS5TbaiZzuilJVGzS+m+MeqghUqA0oF2w02HFEKOKtXvjnHpo8
D5yvyNLLgojYHN/dmxt51rfovgi5d9LAtvzx7jOYQZbaql8pYJnTOtb/JVnrmZhGbkZJjFAwHIDQ
PSkMpYSpRBuU/MV/IB9TLmYCBclFVil77SAnBpPauenRSx3USFyTFITKxhOXlPGLC9wXmDjh13Ze
6BIE3mS0O8xRfyBvuTkMbeF0UdMXLGcZVQ+WnWjJYGoQQBs7R46bHJD9GQ2scHEWKH6YbFG1PPUb
1Fcx5Zgot7EFQYlqO8vSMC8tTxrJNXz5FfkG+7T4861xWu4b6eZlfqIHCh9M6GjdQJdqcLWVY2zw
zsQJJPx/Z8QqiVw0Qre0QDkplSGOcK5zL5ysBMhS2l8cjq0LKGPrrbRHkuOlZ1eezhp3VEbNp0pW
+IY5B4zSTaiaNXIsjwafJgHyRQV/6CLxRmGsH3J7sX13u0S73d3xTqIAWDDXJq9uAWLXaj/ca80y
tGrUsYRvl8e9kGcZmIm9cG4lcVa5Eel/DB3trOGzFfxaavllbZh4D1wKGd/UxKAo6xdmws66ECaJ
kpcEHE5UOcORg0i3IHdP8H4vaTOpnYYqLHThtknM/WcsBmFkgmFGouK3WyR57C6s/10mT7hqDJ5H
wFJoTYxtr++MngJMiWEiFwclN3d71msZhj5sf+YmjAw/s5kjlUOIQFcsyngC+Pk3bYrvFV8q9Q+Z
VJCdSnvAUDnzIUMdEUxxKodZMO+J1fnaV26miTp7gL92oDgow7KWzYzEZqjbZiblxaKyLPGW9Sn/
pcnB9V+UiTArobzzJ34yg0S5ZzmrPZvGqohtRe19KTGa4w9GTmgu228p4kZOD8tRy/7Hih3GnEcG
zzIUtG+SPf4RJrzr300+YMLFR7qtfSPybIOhQ1Dqd/2YHdK2xDc/maVaVdEGQ28PrLSuC95ifFB4
/sIj3Rw04MxkxvuuFvxVsaBHzn6EpkjDUW00zH5CTxCyCe6MMA6iy8CqHpqk3bB8u4eCULks8v9c
UMTJKPi5PFTwQh6xv3DRXZ92SKSmoPhF5SDJH5umgW9iI77ZRPHSFvhqQhOez8Nh3bt89M+f1mhc
p5R+pkmE4iz6eXpwUGDmtiwghQPYOXmu6uoM0A9gP1bJinHv4FtQS6XbId98V+B7OA1C3hYWaIqn
q/l+oIP0y4qUdbkcYafS3IFy7WCsXmz1wAdrtxtCTa2b0PHtLm6VH5spapvMLHQ36WnxM8a3L1vH
2MOnpq75tH+kXmjJT4yM5eSCxzQAWEuoWk49hVEavDI3HlCWLJ+61BQlMfiv5xmHnE5aFnIWeMQL
ayubr53V7Gyb1j7aXwkHVl+KXwkQO3n+zACnS0czCozzknv8rqjDkNDcHkyOIOZrCQZKp0zIDull
AnyvTg6rvPhagzZGRuREJAAkQaqAKMIuiQT79Pkk/COtLpDfuFs23sUXbXGVKDRaikgqtqWNU2Pt
Q4ufudaMME+Q3lIVvdPjyGqNUSUeSmicEOSYyIXE8lrQjlBjLrIHNwQNawdhg/YLchTyWj3BSdJt
5Kjjeh8gGEA8D6tEEGHbtUIBluVq0WJLw2SjAo8VFAgVdpT36MNBdLf81hp0LlxwQ97GHbiaddDv
S9S4YEnNfab0bA32t5n9Z8xACu71f+qTHrAj6G7iG8N7tMNM506Xz8LKYMjVR0H1F3EqyTp8R9BQ
SzQFZUJ51EKp2NQqILwrcjTMOx9yoJ79X7X6oHeJCnDorTliNth+shTzYa05aq9pmaueiSq1z1P3
iXCcFH+aWPCEB7kya/L1NC6PlGsAnP9W0E8YvS/NSvemzN1NscKPrWtBVWnMhfZ7UF+WSX8hIyBW
DFvDE7+0NpnIyf9KJffjMbQy0Odau8c/Wxv1PEQ0yLvdqNgw3uWcER6ebQ/SHAyog/mk5lR9G6IC
UOPwfNL/62gV5gaXILpivrJcTMafJ4p3uAxRRBd6uASNQaZGZF2cMNxBxvSUfQZgsC2/yDvGrA8P
rZxNk9oXkXcqhGE1yPAxE0umJlXH247QL478GwgXqlphw+/4H+m3+IbX0Q4zBJT+jkXl6hCyOzPG
2ptYh7L6aaMrFfVcoq+1DgbhjK1EuF7SZoq4sajP3EtdZDoSoPYlcq17+HSMMWc3XOLCBvjfCXwi
eLbIRJ9Ah4DCa7aT1CbhmrTvb6X3Y3SP7A3Qq6JrblKApsQaJ3LtYdSNGWvH6v8AlLRW0yDW0TO3
0rwagcgqP8VMypB+rcLwiQeTyNO0YHKtCEtGkHpsaDYXrVPTtCSWMtoR5g+DtCTLzbfHQe6pl9lm
dh+bI+QpO9SXkNB30i6ZI4IWcOlGYSUQsgpyFq2TGHgxGWTlm36FhrjWkwCgwlezR84Qnk4WcRyj
5K5y7EB8zzz/YDK7zVSVF2Vra+NvwERYDbgYT7CWpGPAeiZOhNzsMVh2QEgxrgJlkH5+8AEpr1hT
VYX1DM/NFGPYmNV+b6+4GOskRj0gcC/qZbPWu+QgYQ0WVrxm3ddwu9y06iXV3bKm0C9b3Kvr0DeP
G2pocsfYlczgI42t12fI36OyJzZq7HBWF4Ls8W8tw4tSPdzd8d9+wrmFKEkpRvj66hHUVeQ63law
XWXNcRQ/kW/iCV45cvh9m+f6eRIivfmGbUSJeuQHvH6c+ge9mxxBIKV+W5IbyMJ1SYkKGKk6Nbuj
TfNsR3ubJYcbBt1RXxWIWIR2ta75F+y91EJZLGypFIIqPy1xWjQad1jRQzdyIJIC3pDWh/X9Jzyi
4857v400uUybQdiNgaRCccIabxibuZIBULFup8HYQczHiGwdWsgH98zIperiunphpl6hs7oizlN9
BZ8AcciudCaDIYLkOfzeXoEjxYbQS+wK33T8+Cl9rbV94KYX/fb06ZuQD6kAqM+sQllzbFqE22GI
F62CU2lgnwskgUqJuF7Zc2P39wp1l3LNQcGhzggapZ3iSjFuZd4JNKffyCiVJUaKMJxg7YA5FcW0
WBhtrII2TpeimDibX1dL3fzohyDmocUVAqEyXUmpDmY7t9SbxOBRdGcyzqQPXx1nuGF072SE6Bzl
kDd0t0JgacRds6/cqnhZQCIR10vFre2MM++HOuVfDo3JOEJjrMVvDrfBjtHmnOkmKozC8nZkKqsd
Y7IvsWmK5tY53wEqGAuvOLxq2xSrOULoz8xKTScVoQDSH10iUTMP0Qe7ngasdLHlv7+FvHNN/bSO
ZPoTfq2iQ8NKrpPYDBGsDUSSy37v8DvYtg1lTj2e4xJbunhtEmdryOpM/zbznCKcq6gVFyITQswU
GfM0xFxjMlQY8NrrfucSCPMmAssQ1XOSVLkEynNd0IB8i+IWZTGt2t2Gx61OST+28T1uQ+brb5QJ
oU7leyiNwp7Sn8gh4O660czjaUG7XR5U1OK1ROcHC/s0daITKgM3SyNyVr88zejRN0jRJycKXHiR
Ybxf1oplnifRAVBpLG47ogQmekGASvEQTCpGj7WEUXAE1NaSosnnG176XUQgfGOFhd9h3XqYtNyS
4xQYEanFDgqIlKsD42tN40VYMhqwL/TTsGWZc9iNgC0xX6xfa9QBoobtToVgmrO7k4dsIUBNSkBw
xm/k0+LPfAgeqfEpf84XBeZsVIK3S/IcvruqP+niRSIpe4vMpe1CoiKbVXeVGz5cYM/H3S8SPV9i
YXe1GE7m/isMCJVz+9fL3mcGEQKBKrWbKhLExgBnkieq2AsBXFht6Vy7tnuWVDKk0ptZXqVHl9QV
TrZmgtv1CZsp5kLp2YtKx3OeAt6cNdK04Y6P6iq5bcn1uV3/g9X8SUND1YYJNB/BFJ/m1myL436r
O8zxnTRPFCtpeNTVHRORYpBhFxOM1dblPOMME3PnQ7SKSP+TSz7csLtHtY80uN0juxKm2xggUdUE
NlzCBrss8bjB6J6xJhhpRxiNGZlc7MimZH563UE12DBuQAp5LmtdXr2NpW9kSWTV7Akb/vpHySul
TR/JdZGTGZje2QzutBnrh3MVPLKSDEyGoMVI4WqYoZekTj6yH6KzMCKZAzGtA+zaDR9BHVCAdqVf
/ATes4dH+ngYfGPGxuZGHGPSX4hckEp8xnoi/286m123GkNJDOCBMrH1YyAgIaTeLwT9CoYl4qeH
cyhLA2IXWxA28sR1fGiTrt/4rVEbzT+QYIJ+mcaIpfyJ3FH+TVdLeaV0obbXli2Me56vZkODUcSt
CaYDliCTgdcpq++WhoNF17hCoosTrk1EZPCOX2/eg2P0mjgnnXjSpcGzIpJKP5e8nir/5fAXh8TE
tkZXeZ4m+YYuyVTQBmEhDTukrxVt0VMtKgKX7vy6bOXdd1wytP907ijDz/OvDiiENs9DeS3/yacF
m20kxi2J8zV22NKPn/cQ7L6RxLKmUhqlV4rf41eB7HqLyaG83TIEc2kZbENuvDULpxtilUwZ8KoT
6Y0+bXFe5UIryK2+p2ZlRHqxDpN58sE5gUbq28LxwMNtxAddZaTZ6NNAwxB40ET/OQQjqUW/Hab+
nv3LRVn4X2bsmrAlCLDYcU6ubGEKr0BLchiymlOkz+xt3qzsO5nt5MGC+BoQE9A89DXSf0x7FGx7
lTlY0M/lDWvBG8sgzXhrH+a7WHa+5Zt7v6783SwkfEsNTUJZazMwlsXpiWHqlT7vSPdEsJDtDGm4
1HbW8R8o7YpVls92G/N4aPqgsub5K7kHCoUMhHXdJuZMjGwO7ehwaHuyzY2muuMNGK1rjg2UY9Ps
7TB+WuPzcofnH9IFF4RzHfUCHHb2EHg8GvScHxWW/pkxOAkCPS+7WHH7K80te/euw8trZGsRYtO1
0CpT4HwqpgwGhlei0qj5OgXQv0wwsEbORbrdrZRlulNzFb4AsGfeKmEbgeEiA3CIRHWeOMFrn/1b
Au+EWZDFqqI8c21nbMBvRj5QXu0+BitXFm698JvwSN1XTxtl0OqAqfnBYluh8YkwiVX03mYWeCGT
G51sVySCxffnqQIXpVxKAJy5z93zoSyxkwhOR7Q78Qj3AqWluexjptAfw/864FHeHXxb/yojwOXn
C58fRWNSt1ls5/CSeY7fkqOs+pwO1wGaJ5APY73wwtZ2w5AvEuf/U7qc/0MytkLR102gd5CUTDnw
1jYwqZ1aGWx7O6RQmcvznSfPKKtB2Glwo4zHY9HdXI+4HpPBFrZptXHuoSv3gwSTNaj+nqj2oFAh
bi5FHxWDPR9WHfMxBvzzaGK8uote2OXkxzjX0BJFahFmbfKDA5X/0LFRg2xr55MrEU6iRdhFHmG0
fUTO490+kzTJviGP7N1o1qB25Yte42lNa7PauKO9VC+SPBYjpzWEh0n8vuWV6DLMyqcoavjzhDn3
u7ENgNl5DCLmu3njxynmQ0/mOGoQqsrkMS2Fc/KXpNfdcu9PwOHouUrckL5viuN0o/mYaDbwJMPz
wh66FMMCEGO3iHp2P8LLgzkB5ceh9GibcnVi/YuNqX2VgbSwD6ZZwIlrcxtWIoXYpc+q6T530t8u
WdR5Qhar257342kUVRxOdKPRhxMnvQLKywviaOzBT0xgSqCe+OafqDW/qfFezROdNnC7UA5MD17+
aU2rhrGxO0cK/+fHx0EOiJIRkzUr58WdwZ/R6YYqZTOk7LMwgt3F9Vc3Q3F71efq04CJ1TLh2pzi
so8AGq1jnviZ+hXyS4Kjb+IbM+Z4RbxEm7Zxuf4GX6/lcOYB3s4EZkCnjxMnJ9cPPGa+HaJhi7UT
g3hDSfrszNhqeLugC/i6XObZI+EY21eH3Ubgr0pBk+KfN34rAFvrOH0CQKyXDxnoIM0/+AbdO2+q
jI3M87VIKp9sur4uDzzeREd2Qmg9u1Vc41JCxQp7fj32kWl4tGKLB6DbVfrV8xIdMPbNqLBX0twZ
8Is8B00MRbm3nkdQB3LwEJgcKin8ZrMcgRNjuoOzqOd+6mc2Bl1HbeBmO4I5ox+/kV2JIKZTKLkL
q4VLnx22Jv1RpoDlMK2pU7dENI5ru7kG1xA9WPYbdy7VFDJVMBhn90W7QavHb2ld0vl9vL+3/XvH
RFRMwAm6vJwN8WRwCmV7HGLfgJPUXkKMxYVEn4qwE+Wyvv3SRUyptEw8/GbrC5TICJ73phG1EHtg
T+MV0jkHqMF2eS+DpIrkQseCc4IfrOIqhGBWGhcELwkAcCVtDfsR0pmgl7iLWEagX76vUwQU4aqn
wunQHPsEg7vTwE33kOmzFgW7uydGRPxeE/oFtFxf/Vp3pHbxIEjTtn6h/4I8E2KHUn7xa1e3ZijM
q6ui5o7ZiN9uwy6H6aTosQI8qLIfJdirdVvqzPRg2DZ+GApNTMmQdKw2VlWztAICE0mReg+cpjHH
L8JwfWj1Q5CyzxL4s6WIV6Uqyik7XxK9f9qtA9NVUucev3SsSGCi44mMkwTAYB+pMAGZmk+tNCQl
3F3vwgG53SbudMeU84lUHr7Ae6Yl0RptftnVPXOl17/UpC+w8hOAwF6rg8q4qZFkkhXtOhlhQNQv
pw616DOoaCsKRMAHIDfcFDEcKnk25fXD8FCCcoDN6VaELZ5mWgGUgpFoTYi46WJ8JfgW6+sWVs74
FD9inwO+8uh706nohNdh1R6pp9EG/3Nr2bBhNp+K/1cR+wAJt6EkwSC+VNyEIEcUma0GuOEyiElf
UDIdRRDu02R2zlvGxJry/nsFDrHlEu+EkO9caihyZw64/55lYvsQYd+AeVU//EqGfk7COni4QcGl
sfokScg2uKursYx9oxJFLafPWpgwG3bxUfPpMAVU38YnfMqWSOIn38Q6zGibuvVyDvfyBYqgek8c
FnYojEmDCjtk9Ps9Zcl6wkGysiOLlhL7wwNNmEhFyCXKvQRknfBft8mQplbutrcyacNYohKuaIPZ
PlXnWJ/u6TxVMQQod1/tSOhJBAQ0YiTrgfFbAgRK0sEKB0cSAUp/rP/6zw7iw3qSF7bbD1t7RSWX
Gp+9LtH5EU6I9T2erh661RMvP/jPwSrlgb4gPw1vp/cOsbChkcQt0A0ZS030vYVAMHQfvsM2jkQj
eugt3479Moy8Kh+DKzc1WTPcSZdqOqg8NUKREtSaYU0mfompSlA20VGGfJYhhJOLa0+G6KyFHXl7
GMzpoh6jbSwF+B/t25T0wzp/whstnvB0P2X7ugiIVnFKoRACvXZglaLkVUH/gxrbn4IcnDS/rLxy
jnyEntxUZsgcVMri/8FsPL+p1iCt9lsR8yVknAqTQfi/AITEkJ1nA9aNSzNeSzDnEGBmNTnuryVS
A/ZXW31mczKHkzgXoWjWNKMhGBFCqIfQA3tNMeiqWxPgPAvmO8CGQE2jKjoFqOzOR6SUJu08nXAx
N6gdAWE6aEukaCecjKZdOo+lhnCIfmdJnNq/lwc5OjcY2qPcwn+iO7Ko65lWFXsOTfmMxbDk+3Pq
Vx12yCvfhWF61Ah+Xjrh0rz1iW2kfPknXwmWGIsPgabgggvk2T/ES+JmLlqOemqhLxrsTqh98txd
j1TUyI2mOvQv4Mij+M1iZO5miQbvjqhphH2CTqjgBUNwEMuWDibb/5GFW9QgyI545y30MOCNb/NH
k1DrLIfxUpd1xhEWNUbbBhFiCtAMiLbtI/jplLJgU+6Gh1vyCHAMZYDFKyVqnspMao0nczCNdQ5X
fcliUVistDnn4K7YBWGgzOkuJk8385DJ2n0OdXgEfGI07fozPqHtOcoOgkhJbA/UFHY617jUIxz7
45MQ8YzHhE8z8V54f6NCvN4IW/PNdSNhfkrFMdSbItHzfqSaY5B7paEDgSvIfW5EpP/DQlXXOLyt
z7JEaX67jOlHHUv4MZ24dsofsgmL5Nv9wX0nSXrghXJMpgtzDQ11tdPTM7teYI5zi/qZSvjMmmhl
e5WxdaVdSqj5H0AJtGm2YjEbOAdTNH9WeF4KuTJZPmPz15SpMxFWoMgcjP1iliRT2sVZ/oInIjlc
MFrSDNLOfzPWL/1rylujcv5g7RkaZkNsoU5FhBhrCPz6SDKbyuwGWDPQmgDZPxwh+8HvsVBRkomG
vG77vptkb4ncBamauVGQd5P51VNnyj1YbZAHhQq7w91SQWECvQPlIYesAGe0zpZ2yjJlVujuU4ck
bzHgauI/XcTj0QEQvVNA7k8LzFtce3wYRwy682nGeISBEgK+eGLdfatWn1Bu9VGXfR93Hx2LODYs
qhiuszxvR0zTZxJ+uPPQUaiRA1I0kMp1OfMigpNEwqNZqAaNEuXa22RZqRxwg9yYKEqPABfCfU1l
ifH+qtwvYcgjR4gCxZh3BhZ5Cc51XfEBp98JYaFMhlQ3YhzysNWW9c//fHmpby9z8fKajIK1s/uO
bss13nnbHt6KPZjoh2JYlv9Pux/LR7UmszYVIpF6ypnyRnnIlGH60mppcNf8Mf4UBG0OdzTmUSFK
iV+Iv70oKD6IdZnlumAqzvFuKlqZwaeICE4OzJGdGUQpLDlHwrfcW9Wi2zonfJnLNh8GwhbLFWTn
CcjQwqG3voEVaGQ22kztmc74M4TMeKEltVgDUwkYjTH0egI0iGJpR8D1aTCXJiWIwf0ygRWx9+HF
hpwFe8p70fBO6MSNDwCj+5d0CD4+BbT2zM3DAxdJcIBsl4IoO2+DPXya/VdSmUAHYeMgsdgRKVub
pn6KBBdT0uQEFB9xoZE8QbO6wvRao0pnhxoauTqnw6qBkElWqBQ7vNoKhg7vPmfzJpijr0HUzFmQ
cbz1miQ74fV6Fr82Rj6kmODvpuXx7U1F6XXmbtldKXdcovvwM7prbKHhegGhcsyG8UK9IOzGGYUP
5HO6HxLTWdV6POWjwByDs30T+tfduNpW36OJQSsVxUxWmVdqiaGsj8amCA8gJ4WU2+yiJkuA/z0Y
4n9hX6mPgSnSmvUAuACSO0saxPkkJ7R3H6cbaF2Ng9Y9GyT5Y4sQXqJdNGmQL8AeJs0kVb5XxoqQ
hcjYSd+4I+KNFL2vo5Zh5ODhl0M9ZKkgKZaNptxwH/2xXzV9upIw7OyimEXaz4OJ0u3jzgm5nu4b
hMs8cTU9AVjT8SxBanB3ag8n0cpCKm/HWPPYzhEZo6SNTUKIRKg7RD24epMIiI9HOnnlpwhBs3sQ
wHZOBiqT6fh5c0t0RMf5VbHopyVLoBzr7PKAd1ljCH8TgG7YnGhg8rLVF6VkcQewKBUy6fHNJRmo
ecgfz6mhPsMg3PG5YWHW0viOnQqZLwfhwoNs+TCtg2c9Y7ytZ7Ia5bD0M04rMy6BzffHbu2KDOK+
tgUYgNV++Vm1R99fLGTjQyTkOP5LXR1luVc62ZZDI6boPdQh/TwVg3XmcnlcZuy3zskSrMM7jcb1
KDZxJuq5VkKBCcCOqezQTmxHuIN29XLSTJo74LzLzB8Z3LcgG3zZ8uucI57WHaN3Nw6wUEAQt5jJ
/kd3s6HBSq1KFOrJUjgocERJbG2Qc1xPzzh9fdS2Solw37FEDcb6Ld68CaiWr3jpD9VX4rDOo1+D
2rCjjh8JJHi0y7j8mXaSXG3IqyN7vLS3Sx76jsMNdE0rTyAXIz/EvGRmrtklSZtOTGE1r0Aaz5R5
SqZZ52P+7vAUOYNJeJuFkN2RX4KQHFcLI1f5bph5ukCBC1EaDJpPQyzzZ4NWGyRT3wrjWvoKd+Ce
Qz97+3Vcx5aMJEli4vE6dFv9zimmFZQj+W4ET48N0qGP/dDYZvZkNs7HtFxlLZiXYrJ/8UGVQJVp
cjhDPwiv96BNfI11A2uoMiC406pRL/att2Yc+M0rXW2ecxR5yP5PCdwi5DMy2oRSZcKSY+hbRWK9
qh1tWPms5riPMxj96LEFMyGLR2IFnXQjPJKLk6UAQIyeK5ePm3dvTv5SLL2rWdmywD+7hIwEEfLd
PMe7oW4m60w35s06g4wMVjCeSpQQWudZJleUWw4EWtq0sukUMvgwNXfbYuZHltrs8IZ6ETBRtpzI
ty8COxiKeFR4t9wTMG8SJ5/e9uwjfYlpAqdrj8v7nwLH6h96QWqlGaLaBKRmeCi4mqUdm1bsYsML
/QXOv6XVw5P1y3lQeEhQsoYHQ/EH4N+KndavM/I1u2IchZ3HT1eZRkCNmMrdXnhnbcApD0glTjN0
FFJZjFn0iQaoWCWcU5nG0rj/DHfs7QTs1bL6FdIdXGp26Aa21ME6ZSaQWed2Te/th1DcsuVgPfDt
qMPn4h8z1tihzRBlfxK3Qni7kjmCh3it8V1n4neBAHnxzQ8gwR6PBEzuHx6NX3ngrkXGsVqyxPuS
TfAXCh3ee3LwKTSYTxopnelytRZy5Ot0YtNgw0zXfJ+f/Qmj52wMKs5XsGduQdgvnyDFktCYZ9Dd
lrNOT5O95Iik7sWh5s9nbaPaWQWwuHrQ/x2s+MOsp+txVpW8d7o9EIDvXVZrgnFtPY5O7GF5gTCy
9+LCqXaAO8D+JTvPVQQHColYZP5rGgcSRSg/xxga/STk0Z2lCkp2zxyMKN3pO916ecT4oBk7J2BW
h01oAbzLZIqxjX7qRtasdeN7PakDBtg5ebHqPRnpfTppdPlT6aXylcda19hFwACEPeq6+KvffCdd
RA5GWKP1fUR8elShcq4Xe8wE7L/W+rUY+eNwSMu2InMqNGRywue2Iz+S5MocRX6KSc5/RUPEPo0G
oGznEa/9m3vL1tWmjAy5Ns/AhYg0/WvVLAfniiNaP0KJx5YLIDqG1C3087MZ08I17ipLdWvBGxOx
J9K7mr0D7dEBfxNGk5xvWhLQLkVdXlxJr532Pt5T8LpCEqUfmpLI9knY7G0Cf4+faJv/yzkdIvmq
YqLDAcYdzNfIjth4h22VP0Xa7qYY66aGbkfRfX888mPhmkLGBvEGFnbwKtKIKoX/0XhmE15cFUaT
ePyRrLEUj4WRa9LfgJsSJOoPunAMiqbDWvK2I3s8VssdmZql8RaTFWWUBCslM8zG+Us9W7Z7IK5l
DaZEsbwskEFHWhWM4qK90G71McnPs21Frnba06lF4/jIfRP/O42PrXZb7QuNZGYObfoyvf3mUPOL
RZe085yZ29Qz7eP6fQNmfzEN0JUXec6jPhsrSkIEFIwsjv+g0Txg6BVoCzzZGp9JQDM2Uugo6jSI
kTTV+2ny6edtXWEl0ehXFQZOzW43WXYK9nlYD0+4T5gsYZW8JpjruPM5BXOmSss2iAWb9UV3wDhJ
MpIUWU+lu3yWOpva2X87ioq4MTR20c+7BI7nw0CnatryuBV8Us5gkFiOTuJC7JfOKBOQRHI4Qq9n
tZkf+wXqn4BipVAjsgwGgzHzLlqeB4y+gkjJeeKI/qW76K1Vfg7SHtnKogODl5//gQLlavszGUUB
Opn2S+HN3xI7c/HIWr1E5oku2/PmRJyD6Bt29vuPtmgrMYLyepepL/a0U8fLItZHADqs7gFh8J0A
V5LE5NRgq88vRx90W7vcQDjoV8P4KMMhX1apFfYMt70JxHjWVthT8nyXpCbn+tA7ydIh+7Bzb5A5
ySc90KBHFocFjJd2q4SVnCM4pcmx9n3jebjUnRI2qXr4UfamI2oFTuSRPiYaMFzwq1vwGtCV8U2u
zO4WuqTgfL1TuoLmxRWfI0ygOvmerAM93OItReHTQhGyLm3gbtFv6FKMTaHDBEKbSSMCXq121Bch
HHybBgbfcIBpAg62a44+Xaq7vsiOvmxx516003Sa/Zw7Zfo6hWXpcjaP4p/Z45FapRphFwTwMNTG
WiXg6JhsTu9Woqk0J6lyiZdbzZhzIVnxBQoFaOYhSLy80vDEj/buyOKFmkIZvLFplJuVfIpYOe2A
BEBT8uTYpPg90XgVlDTrvgxJ1U8T2OgluZKmaomtFnsrcme6LEJ4mj11Fuz7DX+GFmn0m7JsCu2D
EP3jquuouKbW5zPUlTJQOX+hwCOXB5dYg8r2N8/bkGcuhKFccaTfKBqqTgy6YPRnPafPKhR5Logj
Cv0n3qAQPhUSDA+km+IBL9KYUe+mheERDswSZE8TtKl0pZK9f/Jrdneg9dm3bCWZqphKq/nH5jqR
yqXfz2Rb0WjcDW3NetjxUMXCLRNvq2+ibNgHOacg4k253KRd+S3iu2T1EspqMykVeDaR1Cqdlr/V
NYxApyS+q6aMb7QNTFqCCVRGD2dW+Zimn5Jh4Oa9ctSIhQVmBE8IzZtACG+FuM4uDi0fdKtOKKJO
wm/ar4g9Ly8ypAYSqIUVhAaaP1QP2sZk1BLpAZJMJe8j01OZTyaZa0DxAOifTPwbRaaM7NmA9Ovw
/BSw1kNHl6/BFW7xTU4U4XE4x2ZRSCWJmXMa64WYNZSkIYKrtJDqa8p2qTWfDmmwh/gMGSPMb9ng
+85nLeBF2Lm9V9m7H2x5AjEVqdJQHxjWiF9DD7Ffm7CDf5Pk8P02MAAlUGAyFPyg9kD4apMJBq4M
aVNKaon8YdNVGrGaZJNxtWc2rKIZQO+9MJnmZRzl8vkmW0hZu+zmWNGqFdqYSWu+eSDLvNhqVI0z
Uqwui9n62dGopYs60ZxJlp79o6PtK5xZx9kVPZ2HVczwNta19DbAdPp2uWcZj+TtgUNziirCvkNx
cczYeuytKZsBZ7B/gjqKaSrez74yKTu6hy1jIwxf+nj449R277cvXMt8Gt8mO0apOULiMUGoR84U
9xMv1XDeoCDxN+d4gDHysnw4B0waPBYbKPS/KUAfD51E1jKFtooAQHv/3rHa5qho1fk8dVWxe97b
tgqmXYtAAuDFRBep3wbegAFTyvJeWRuCVuf+NDa/eKaNNCOuKSr0ACiVH//7F4K1WyJWdhNx9x+Y
6FmyjA+B1zgLZDLQR+rc/HRF4RzR8GEZahhgJ0ovsmJkxLjRciqhuiCE6HKPLP++cVHQMi71iZ9s
1t8KJ59diCBma1XMSi0F9S6v8O58W8LLKxUIRMsufRgUb8pnJqMJJCrGZIV4GlxL2dICIX9F0yxX
vMB6LE6/w/kew3QZ2PZV0AHoBASlIz3pgh3ICfk7nUxqxBuNFG6nO4HNoEKWnL4hkxu+RB1B4Gmo
bHXv2Y5gj5tv7cShm0A2gCfreewuU74k+bOJqC9pqFH0zWTwUfqAXNfzyoE5EKWBjCa1N4edfvWJ
u4CT/GJI6c1VcqdDgiKMcfFcBw3ewA9Q3lrUu8+U7KHR/20I5A400MbJHDVWc+qSuhGUzmpjAhhX
52eYUt/MIBDvEu7F0NxuZ9OapIW4497vI1U9nBDLsjPH7Zi4oWF01OCPYpRMILcFw9T2sCpxOrxa
+Q9cL2ACsP7LD2WHsM7zEtrR4bq/W8kk1wr40XJvaZ6XTgsTpjiPsquxhd1hXfE0VCIw0bTUMGDi
x/djZkJNYbQ8w77LmIypqiQhgbhslDnxPoB9x3Q7/ym44QA4zs1laWTiDxBPR/Xx+Zkh9MOlx2M1
g7r4JaZCiTo/+EaImwBBndjiOsQSk+vRKL+ZjT7oc+ufgMMA94BcFlmbVQQJNvrUmyaf4XFs9BwJ
aYXe+yz+/Q+3SPkDz/N7sl1HFB6A5gqcqyrg+LVjXjCpMNPo5SU+8zCAIx+Sym9UXpkkxdrEq8/a
L2F5D2cCb/u6UzLH6zGwkIBTwb7Wq41jQD1WVJIL//pCIZI3jlyEb41orCGldx1z/faAGSG1WEZK
IVJl0AWWKEQV3TBqRx9jNWkP14UXKZUuFHB74XAp5NYR6okwQ6u+PXC0gs1dY1xiSBkFGYteqCeQ
pUd5uWEOQDiLCoxFy7q8raQgJMVEhOVCNNHPMHM5lXzXcIu33Ixa247jFOaBq2IZmuTPYTCMVMcr
877w5rUW2ubDOo8qpFyGEArN4HpMbgrj61f5Ts8UQ38lMFPY/OG5u1Ka2OlY+RsIAK6ELSro+3RQ
sahlt1H9mDVOWwqNeVU6TC3T1F3UNT7h10uyzkelqXOsOiWmfskvcMQsC0EpfCEq25lHvYr9IixK
IWXJ13xDtxBnDT86p84reRkhJp2QNJJQ4JvoTe2GZR3No3OnkB+H8kbEwwRkD0px1R7pujgRWPRZ
WmaNsuv34xqZgn9R4swTkcg9gEpawCgn3lniPzugYz4+mWCcnI5Yt48W2fGKlCrBk3aSI4wkm/zT
vMdIs0426KtyBNrcjm361XwVMjwk3hled0vyat40VhEnwBZyeMenBFGkZxkI2TAmYQOoltm8hwyE
YepmpbC1ARYXdIRDcKeogGZtL++qXu8mw53gplUqPYS+sjmtjh3LJsoVQwayTizCD3N3CaC+CNUb
AWygO+m9cUK6PfgYE0R4QnY2ilUqLHKZDHxqwdyiqGps3aorM0IQ6S7N0L98tg2Gv5iss/FT4zR8
YJOPlOCgFYjI8Ljo33sohX8C7LF3ooq/4Fi1wJd7aYpu5NbfwdH2aibQxd26PumQWeWqVxcSxjdl
JzpQZkUaG0rnpJoMB0JYEBJaRwkli987HtCmESfnNvdH8c8yD0k0Hsypj28M6C3FJ8mhCiAwhzRt
eCat7mKqOMGBZeR+W5z2QmDGSmWZKSsS8a86KYThoHZ3y76USNpb9rEK4EM4SiepuB1W8LHEtFCo
ee32nujZFYgTdLAVwQmPZ9v+1+sVZevVj+jbEHCoyGFGJtPOYGCsmgGI2LDSkaXArdBF5rMU+4t6
LtO+BVmuGSHP/vTLP3uXKZ+pdxhtEgaGHulJBlJXr3U2PouYSivUXwV9Pumr8hzf3Owpeu/rD3pi
19hYeA/+Evg+7MFZmRyZwaLZFELrEkx/p+mTYv59+b0hTL7m3yBnm08o5C/NWjkCEfku/OpRaEFz
5qQPdgtB5GtmYbETyYdRTVxZkxqN/yOsrO6uw3JATm8icyBmKXIxgpCwVTqNUotbHZG8R7heYsNn
4FywDDEyWyDrf9yZYFhyE3Ad/Awhm9fuK0KB+1n4jStL1azOlEV8KO31lnruFYpudSBpZV4DAhnD
aiVgDdrfBXZUL17aww2y2tU35XZcdFqlTASUVN2Cu1VirUrJZVGyyMErP+vU1jfzubh8GSr7yduD
2Nla+0AAqCoBQN0Dtk01rb7bIEOFnPIksS6+IKIrj/Pi1TVwxUgLSxGFJRTbp6RXiGHZ2hwbAb5U
Dzvt5wFjeJbbPkcJhqdGyQG0pu3KdV3XViu81pIymCV4FUEZQpbOMMgVE7EGnDE6CCAZ1Ae9dlL8
SxMzisxSIvg5E/6/TpxKYkd+ybff/yl+z5kXTjtix9Px9f9COlimvCTsPi0tK6wD5UCoB2JizOBB
L8wHicmoPpE8UIgTYKM8ZaFHclvCmh3aNdeT4zNeKi7qeFgXCr+68steNuUXqE5vzmc0O4u7KXEA
pBSBGdunFwSFh1HGEPuhF41btUbQrr9z6hYA4LjbWbZaSUYa6wUhNnY83OMdAqbal6oIyplEXvf3
Jx/eIG3NQSByUZ/z4ksHARRcuLprUlzeYGcqk6riz4EZtJ7q1PtTXlxaHFCJo8Q3szXzaUuc/kbw
UGVeBGkOgWc8txUAulRiOwuUIpbVx+1Zmkr4rxrvuBqrtToTW2lpU2Cr0q4fOdLxJLlxPmKibBj/
5Tfayy0f1usV8kYxvq17QypF5mn8Qjrx1SMQyGgzDrLe06PubmY88ctmZLKJapDfGCUwgpxZ6fG8
5JGV1BdoTXvjyHFJX0rZsKtK9uvUwUPwo6B3jzbBYTfWV7cKxpNYoWm5DoAlnbOXVuOQF0u1XMUH
IKW+O2aqw8Cgq29u/ltUFenhlBhk1AsUebnLYYBHvJMHw7WeYHsvXLJ3L7Uy4EauxR3YvLXWvcB+
jmtxzGcW6mIYMXIU66fafm4w9rovJMYqHsWzLOw8Ro5xTZVpjuovnjQrE5uzLbAe+635HY0l4I7f
oZrHD8YxBec1FTNDqO9AUuT400SwzyE+V2vQmJ+7Wak9gO7Ns6SgN4AI3CCBb8zF3NkWFO1w6X/O
44PJxoZjVkn6PdTkw7wn8Vl8O8VmbKokfRPUHFEgHzSS6UipGRm7gQNhF/RQCdQ3CBj0oFzIHtCL
nTXMvzVgZEC+7cILkF/LggAiGssaqAvYxuVmtV2HinOEdJPkvrQUA5leHhd2jzqB3yEtLGLmuZV5
W8Szfg12RKvM4iUKWLsQr1RZkCqQrdZ0nefqP2dZaM7FNYn8D51NX2PuUxY+Znw0o/m8mRXGIDZf
7lG+YVd9QaiHEcYkEaRkWfNcrjGVMIshXb8fTRAZKVtDaonA91yawHxs/TxKCUQE13JCX20iWJXN
c8ECfcGOSuDsdG0N54hheh4vqExyAQb1ZGyj4IGenLw1X9AwBEbKPR1Wx0HXKAlfCc6/x/tmlZlw
S4+ktkfejvAiHkg6aPlPzrFTBcjN1AwVxsYFNY9KllxjnTuU8Mpu3MEBzhbMNA2sivfdYub8OyxR
g2le0pAcLNkx5qdagN7upJT2pVUtc7z+4zBEAGZY0L7lXs87uXBTaZMbe9FHfvfvYFBeF3oC4qrX
dQnFXU0Jz1py2Jd5oae/xyEQqFPnZrBZdqABOzw+RzASfARQMRg90FwpexbMSrjSFIN4d92Xfx3j
IEmHQmXgFWj5yUOndafjVOOmMO2J8oN92XoSDDzFnsBLCOeYIs+qUZaCragbaDFY52hT4tAhDKSl
Epsw4UoMBGcQ9g7PtbQ8gqP9NtcNIXOO1KccKjOuBzl7r3MDxPMkySj3UL3GmkFNaC0d9iDvA2xS
UyEI1bkm3/fjSAzCPMdMnL9B8dRlBL+PGwBy5ipJVkR2eOH+8tySKLWpvmnxE2IYLDSoH5VUNk7X
i5pvtcMSkH0g33ymBsYID8GxoKeuj72wtumvNeJrMGl8Q8g4W3MWQIdIvIUxDMhA7Ai98I6KtrdO
LniagV/6jHt+dvQ4v/S+5U8I4JzMnLrJMMR/2eqxWr3BMmA9kPWFQy2xedCGSxibG0zVYZyjtIRZ
wIj6NCqJ1VKJleG8S0iACoAlQ0rlhcp82eQ+Ddnab6aBLAIW5s3LLw6wwoa9/U0pmklei28SvHqQ
iUxqjNNDGhslHcyH4HXOTwLQFLAPCNHJqdRsz8ug3R/qiyCBByMiaWEzJzeFJ3/wqotFkOMw9xnL
pGyyFo7a6RmaPjdHNWwMt5jnScojQ4dYCboEhVzy1tlAQkeY3KQYTBxPcVGCGsyGWFut6MpqAS0Z
gISu+MQyOTEEzf5DM4BNdemhkDSu/lsTatP+EBPeYpCtbjDoEm96xIhddp1xpcHKpgweM1tDp5WE
4v/MgG0di8okcDXeG2h7fJ4zcv7T6iJidD0wFjTneS6h70XR7gIx3p3BDDablzeHc3m8li4di6np
5UrzYFC115UldQojwhcBJk8mntgHeLpPm6f7cZqvXYEaDLeq0aJGqbP5vtrujpbWJThT6k9yrRtD
j+jZOVYmi3N/mNSqfY11qyIQPCGx89i17XQqcjxvI8HMgeAFCktLkg7oIk3Xpf4ShgmdxjIV4gj4
/PIWtd5uPe3K24oQay8Hn5TJwKOJYpFGqEKyucKU9pQ1M0gXCJG8IrY2gRvjEPq3FHIusIvvnvMG
pbNxBWi2krwLJXbj8+dj2TaVPXVN9cZoygo2U2Fp63jEj4pcemmxEVLv36Z8/rcWR0CTNhQwr1Qu
ocWPfKs7oGzBscqPdJ5ObsgXnSE9GvwyWS6VCPvg10Suf97gcEWGZe0vAancwfgwlX6+8s1hBwBF
g9Mz5NFacfp9HM5FWtS0nSK2kOOPwcaXCu9nYMm6MmEiunGL2nnBkckmpfGVxBGQo62PwjPoo7aa
YNXGXVeQT2aOrLcMWYoNU2SBhRP/SYeVPxQQvtoW70f3jKbOJjKZvfFcRmcqQrAay+vtSAsCAdE0
15TUqs/6TAElDVNTGrLZi8tWUTofdugkfYAJLSpuputXCQdcqKQ7PpIPd9n7KsLj11vSK5Mav5Zn
mLQ78Absliat50h9mLtE6Zxp0EWIuQODDg7PfKJpPKeTaSb1wGKZNvgq27tCdo/7agmTVKIq9Vlp
Ky2ZuvJnVnaDLkcsjYfswnWgpRPV9Cm1Hb7NZKZ5+vIJkoWnFheaVmr+B5d6J5dSnbybUHd7yCYo
nGk4NMPF9hfnSnGc5knAj5V5DgHnGGRX3BtpMjmcw6UtBRYNjGJCm35s1FU6YdgjVzxBus36XqUA
6oTFJp0l8QFmg+QVT8D/wNfs71iaGzsrCKt81JnKW5mXGaa4gllKesZH0j1Zhlg+dv4alVXabvEv
nm6wr8FW8qHYQ6cIfQFc3W1sNQpvHpiWbWMVi6drFfZE3MAOQhrH3iQroVx5Xad5kqI+uKsMPNSN
b2fZ0po2BKBAg4SwINIpsOhVSB2FJMZJGPtVASJpU/dRvptTM5rGMyT4ihShecshAQf8X8eyLsy4
OcXM4CPJJ1l6bV5j11/dxR8Op4cDIE920ksoxgjTNCkZOe+yn5uMl7T9eP7D8f+6RhrEyM5DByCx
AQPnIOlrNlUjaoPCN8ZF/Q8UtUoy10G+Bwt0AzKYv4GFOKTUqdJqnkONUGzb1aWq5DpAFA+60XR6
z17saGhxN9BkjLOsY05bz49Hv+mS9yqDqIgbOf1OMOFNf/5ShUU2lGlVtxb+BpkWcRCzkwlDq52m
RS5DoUY0E6ltT+1Jz2T5H7VqWY/d0slcxNwtivVAxvGgJACLBkqJ7DRCjglkjDajLnW3voM2Xugx
DEAsF0XrtkJetsL4sm62Fft/FkIbPNglHDoQPPd39t5UkrQUVjG4OP7OQn5I7mQBX79P0FfzViJI
sM523ry5KMGrsw9mbVvT6zPMFlM4ekEsfVXmXkKej4yoCESvblusv4LcOEKrzjT7KugG0W53hJvv
Zihmtl5Xfxzgbh/71PVq44GfdwALv984nA3wCm1EY34jOEAUNjrwTS0KVYxvpnlYMoOqJ0Px8uSc
LBx0AaacnLmBNAqGYmNkjsedND9KhlaPvM/p7cWU2S2MaNrOKS0ZEE7nSGfrJcbOfcoewc6/jRId
d8uRW51fyvLvY87sBPyvs/HUp8rncqeM6EjWkE4/H3Ys3jcPB6PzokeZ3Ju8rK4zr421NHlZOhFO
0k+1GfEAuuAG8wkqGKrPzj9fJ3ySO726IysvllpvYkrW0VptiOxmbCs5UswOjUjw3XbqlbzBU6m6
vfhZembWXwfLa1cnDD998kewP9dhSdduQjIKPzvGNsyQ4qFTQ4Lgs1CxWlszJeu8hPxT41aaYHCY
+99zXgZB0DnyVN5EQpQv8e07ORT0tr/NLxLWMYrP+4VbWe9alzlaKb2iXFdd7OB+ZsqBV37hRMXs
qcED1hsjuC6ps2V2Wd06prML6Fz5AWSlFZsd1icCppAPJYDD/+clHYg18xExdt95wz8GLmwUYtjK
/5+zhSXOm9lec1V2AVS0eL5Zb169mbj0jLn9L81Ti9oNRpK6Exzz6CR6foXDdsVH9XXP/vnvpZh/
Vyxi4fTQsWCgF3cykh5jyMZWOAtpG3Z2WxpPcL+UCR6DtVf2LiU2u7pZ3HLQGzxLMxKvBDWKoXiX
8neW+vHUVSQawXDtStV0hXHp5a6VAH/khjcrFlrnjH4mRR4VVjbAxpsgibSn7uaO2LSfITui72YC
Tazo5mWuH+kcqFx7oWZyR3szGHMDnY6Xnepiq1CaYDmo80HTfoanOhQdPZoUwK5d+Vteiqn2yTi3
/OhmkAdURBINvL/NJ3LxNIX1O2ifjtieyVadvLphGtb+n2/3GaDoPl9keD7AA+w15JNp1HyFm5CR
q1saB4vQg0DbnKiiF4RBHLu+ydayoJEMjU48o/Csw+BFZj+yV3qLUuS39RVsDf5lryaETC3nQAaX
DoQ8QdoNadrkCG8dniia6XLqD8QixQqnCenA0QLIKVP0hWJ0JyIw1YOF/yNoRfh44GQ7l2mtNJhQ
61OVjoGzw0FJGtn97QLZE69rdkB+fxy5y+9Qh+MpnWOLrJPtxew/ZC5H0dlTBtcWipvh5j3BIIgK
xx+WbaGeT8p7LnTBUcGKhugE5wnGqi5mSfTNbV9d/Qf8/rCr0sKQ3UwcvAPO8f5gM/jYCYUT563Y
tU8RYkPj2IR+lBuE+Ox213tQkbbfh6Xy7Q9a7VVc778Dmo7oKPoX6zMbOLuo8hkS35IjkxyZjOiR
m3F93NCYRD1T1Rx/cSrE4mlc5w2G9VGUlDv33N+Nkm0Ih0KORNr/L7FrBVWqhZavX1alEHJhbsj7
uVi6Wdt/hTOpstWgrO/5aHbJRKaIyGiZqptwFGgpN+UEzJ9AifMxQU1AzuUeSv81NYeszHn7nE3j
HJ2v1OTgWH33nzVuzqNNrDylH4Oc7ExMFSU3uaADX2uj/EmInBEzG6+QGj1qy0ro4N6yf8SzjrCc
lmTu4uzcpffk5e3nzXwtX5dr1jSaAGSDxlhD7AT+pUtxdUypvKGq2cZbe7pt/5hbQQvjGfH28GpX
l/HMAT6c5WGWIidaVbja+HweAS4JeQo8xFdN0jUaCdrGrPpGWh3efH2bPN/ElgcCV3GcQ+WPCMhk
mpSlLHN63yFn8YZRs5+vfQaAUdeuzKqSUDpkcIh3OqGpBqRd84D25Z/3X6jaezCVRLAjqezr6UGI
Ebtm2282GznWhm1WnJdoA2+5CSzWI/ZVKV6CSxNr453cKIkvuBaF685PN4qRJKRE4iIBbWIioftt
a+EOdXacmFxwioG1QE0rKN+fyeGhoOdW/STqu019ABXMWnsaOM818WVKbdXdo1n855vDIsFwU5C/
ljp0Raty1CUucVGVrL+qsg6KfjMOCNhjWD4iYU/Vz4OrijWKRjyOmnU9iusxarGTcbVoYa8IZpU6
ODCGnn7Bc2t1R/HP/97jlo2SVjKykynkQFFIUINxqcXUYvZfr1ffnxpDNqbWzfVCAlnyLPNdn85C
mMGqCD3pxApDyB8M4HaS+oZ0IgR2eoEZGbnsI7zDJCp3WNtFooJRgGpslelJKgjdyPR2yHJSls8V
Ersr7yKAtm/4PJ6NPYaxMW918/Ew7CYaL79kCZ8d8Bipm6C+TzIK/pokBwsEeErUF2K/j2GzcVcJ
tIjWiBNF5P+qSeWYAhWLV312MyxUUK8WmV1KM8vklelo48hpiNbgDSrB6xdf6OQgmyNvEnXGaxj0
VM1SztgP6z3TVAKqe8ovj9Yt2jY7xAXI/SG+ahU4XZj1zeosJzt9+UFfagjz9deF4guQmK+9zzQc
8RGePmCXMeKwTeA6OMR984uws584SYfJ+/wpaayRofHH9NsTXbZcNKYYUnLjb1qHoVMTAOEKrsj2
AgpSN1wTIb5/U15ov/pydQMyc7ZBEGi0GBVu3ws1o302O2FyO41rV6bQ5FlLXQ1Z8iWP0jDKJeJW
hirfB4V1uA4yx8k6n/MhEHNeE37EsHLGUeTPs/fP/OxRHEB1d0jvh35uKQklJLddly83RcYqpksn
uFkx3Ggv7WU2ivt+n7waOl+xba+Uxug+7PZ/+4zePnhKr9JTjU2P6cpZ4HH6xE/2ySnv9Deds70h
oxwoq8aeF46atVjJDKhDgDa4RFDcybP63HwwejqFAYrpF+MSW1A7ICxCjjGA2H5Xx4mEO8+cU/tq
1H+e0k3T3d2rjI8OlSkyZbMaWQ6vrPiWj2JQbrbmHsmOgb1hIBhMU72NUgyVzMu90OyYnOS39bYi
YJyP5Uf9YbFG2BkH5CkZ3mFMRXZXvvVsnIpYZWyYFijJ33yKsMbfn1+gK49LaRxuR17kfgEe9J0C
uxXEWPCVsKBUL3+rBU2CFCnP/6XIX5jqaXT9HpTfYsXCyFqPVMPDqwAxuM4uemoB2U2AHbotnPrg
DdvgR2NivSbcbfBk3IZt5Ze4Rj1+D/16RNLFh/uonncx359RMotOCMehAw2MLzLn9WIjMxSumDb3
TJ4vvyBVAsOJkiTv+lvC6ezsQ6lt9+weuIJU6rQMEJQZTp+y1AL78i1Ih3DQ1H8s9cvA3QFH2JaU
K6sRGeuoE18e79y6EXIPFlLv/pNxPX3FzrQ3LTsY/+hrD54rj+CIboxCSc6/O4Ger+RXMfc63iYg
8AnfBfJv1yBHA1GHArgwz1A5On3hXYmoX9hmQSV3nfi2N+FqP5Nwoxwa7pKW3qPqYZRRkYEN5hXd
3uQ8p3BBERsCupBcrdK7DsuZ4w1udfqJ2KD7RHcCQoFiNHYkmoO3wUgTU3s3WTRRunB1B6a2+n9i
zwJCy8D100CgtwwWbF+KHd71nykuIYzjOtlX4SwyeIpsnszmbZ/Us9zjgmN67EdVUQtKPTyGuFsg
UvfCDcRUM5S8V5IQHR5JqduQpiQXTDMlCEmxvKXPg+YQYrfJVt3XyLPpkJ1a4kLwh9xgE2htGWYU
VEiuQmIuT4ECBIFIyPgmAoiw19G2DVFlm/l1bfH3DxZR7fE0ZhdYhlKuw2Cw3FVb0/A/GJGTGXF3
r+q/eba3SphjB7kYgNzk8A1igA9MOqNXEkNuV9m0fnMDkJqm0ZuwKvoOEKn30+H9Y0xV7DIF5CV6
N8kmYSkQ73cq/c9s169+Z3AZ2STr9aWkK9FuFYWeEnJhYTR4btAQ+YqTYN7l9KkvpDeHbgF1sXsq
CdU+sLfar0e+xliWMFOFIG7mXoUmytEDvpehfJSXyM6F+mhW0j8qaZs4ZN96BaZGDM7YC75GyKoq
ZMTOemVgWul/Bzp91YEiaPk3m3bB6T3oAwxwKrXGKoXIeAdx+BqksPjXOKrwjDaM93qKxrDrDS+c
Wc/EPilgoIVUUGQp7zhdFh44T43meRmWHKBhXQh6Hl33Pcu974+KmxCpnQy21KuEGbbvNlv2RfBV
miHIOI0mKn5UAfhNVjrOXcby9TtqymxvHqMrVuK9EfzgrMaea1vg+mmK0xk/NTQwgBKaLd8MRQ4X
auEImWF91Sq7MSpMuN5XhNbNmmM831FdtwXpfbOwRWKYslil8rgcu1XUwlDWXmrm6tUEqwSusFn2
TC5qe578I40SPXPtiDf/TSYNniCbf8ExpHJRCco6MUQILQ/lF5RcdpsR32jL45FCmw2k2ow+GxZv
sK48QX6//Z9/YMLh4Z53sw9MxdPtc043lUk34l0YZV0OnwqlHrCdZ76Y2Yv1pk0AAH6UQuD/ZOfQ
8gUhuxbql7Izu953rmgbczauRJOa3qq0DapYq+q3anriFNT6ZnTEcUDD0smryvMz+9OS4ZDEpKuY
xh52BAoFJiUKqB8XjmNpZho22VJqzD4AtpV3O9Td6F9fLLcml6toBsRigXw8tXYfcJmkduiLKCMh
Kweti2IiEpIFjqblT23ktTjBXVy8ECciEQ1GPXQWvUP99MfS3wFE5g2d88rundH5hKOfhGxkAn9p
GKIdI4qEiLZUVI7ZYcGuENseTARpYywJ6IxJIMuT9TITi1JoBNbMP19BBQmDR0JrUhvx061j3MOF
yJ9mi7AR+GOocFmmTa1jE6clKL+M1r0nTr9dpz0YviPQf4Xte2LBazVIE1QjmLLbA/VOdmL6JQXe
Vy98ZsnXDWrqh/Sj8sKPNI9jhui7FWlO8NGimlBELLFEEGzTElBUv70kxV05y/YTCShgEL2m7bfv
cIQft1LLbZsFWGoXz8HjZPPoJtsYQCTExtnNTj+JnjlWI5SRDDmWEZ2YsBd+HblVEHUNwmjDlWZX
sDWJl5lMYQkly3sqcDw20C00tN6FBBw9oajVZYkmXXwN6n/DsUq2iPpwiGkHw5s0pOGHIclrgW+k
+2LREfEEjY43YDaRTv6Cy3/GpR3BLWP11dAyCiNO3PPJCx4PTxOyM5CBTcV/Fv6PlC44nUra/UqH
cubAG79pUdJQ7SR7epuNyLcel5Y81dl8SaiLf1Y2BU2vJ9xNyFkQmjXh7dLpcIz1JcXWGVaTKI2j
Wxwb80kCwmsP2KysXlmw+A3Xt/baFSv0RDsMTznx26ZvXJo+1wvELdhyT8TUS/Sj+gfibOB7WAPf
1dWbuYu/bBKI6TSurkmkOtDefT6T8+z3QvR3d8ZB6rKw2MjG+px/AILZ1TIhxW8Uu3JxJORSPVYi
7+RmZtnTtFngJ8o4IiJ0OTONrdIhL1DfMquMVyYSpXEg+zKmi0tIzEa16OxuX9BSP0LzSVRnJ+ct
dZoRwQAXG4uQMAjpzP92YM23BobhwMv+Re+mAYNL1y52OrVqGvolgoJ+9SMPglG5MHQe0Nwsg8Rh
hG96lGlYptm6Z2THPtM4ptJzMizYw3Aoo8DO4vwNUbRmHTAwtPIiIqvajJ/HyaGNZIC889Pawwx9
BPgaezRTI6q2EGQjKcxWXHLUjxpIqxfzTgTih3zFClVbabdfYCTOFlyIBOPsNv62LMmXKlk1RyGa
RgK/BGEYleUmHY5iQJMSM92lGYqGYd1pHCU6f9uhD5qsIMl5jnZAHtpJfcoqnVxHNdWc/GjiwYjq
yWghcDYn4JSrFIoDBRFkXbOuchADPJR3PNOAFHHm60yHprRzkt1nmKV/r83GsxXybrfLcxTX8ppx
elZ+aGo0y3yYK+9EoKrHKNQXo7BtqD9lNbTcqXyBPey2OuTSBM7O8a5mwX37mY4S0moNpv1uIQH5
piHjzACfJmYRK6syrqcnwKRR7TPaLEdsrj0aRRsL3IQTa4ZaEtbzjTijTixy+dCN5tGlhAg0jtdS
CUyDlYqhx+DesgWQ/aK31duIU+Phwf2zADdWQj4wh3ye4e4hVhPOL/JVuQONDEKsrj0y6m7bM0S2
oEI3fjx8/2bjw+PPd9Owhrsw3uRUBkijbwiWwUdGR/S32ZzAaPTdpJ6jEJOiDxsUczUO895Z8Lp9
VgWVxrYOXV1LhsxNAzm2mOdRl/YlY9A9taHlHKfPMMHjQmrbqukxUQwDS3v5Zy9KCOPGQP+66jVj
HHxG/ZGJrV6iY93lg9vhguDAYLw2evZx+hv81Cz3ZiD6

`protect end_protected
