`protect begin_protected
`protect version=1
`protect encrypt_agent="FMSH Encrypt Tool"
`protect encrypt_agent_info="FMSH Encrypt Version 1.0"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2017_05", key_method="rsa"
`protect key_block
JN+BeDXZeFwnUwxK1lG/dKY646NdbJNrTFrHA3zPWdAhl3Goo9fhS4Wc8CGQyzaBQhcSWFIgbQ+q
EKY9DLwi7XieLQeXyYheprjfp6fUpY79VPD16gCHdqp3tUGSSpl93tLPI4InzuHv5wObcBGAskP5
Dc8Y84/L2Q6hqonvIAEfIXEnMKjH2jsOPdq3URTDuAMCzcyYTc7umeLdavxyrplBYKydF4xc/zU6
6rjnJQsInKsKwuEsX9OJ8IArzkM8zu1xk6U14xUG0+jl5gpWQkgOPxJ+FW/SqnSVWcXi7hZJOqiw
WLghLyfmBOgzoMdNM7xFkN7srHC1cYD0KP9zyw==

`protect data_method="aes256-cbc"
`protect encoding=(enctype="base64", line_length=76, bytes=74224)
`protect data_block
cLni91RjmwLEUXUxc/kj3cu+m1e0WIOiFG0N1gQ3+RN/gLfjnhKcG1pg+tjumybkvHm4gjHrXYdv
u5M6g7CXecaCElHcKY/CbH0P2n6IV7JuArHLVkh4R5ACTRcmohjlMvU0lPkNDgsKvMEGc38COLnY
TESnWetPDuxw00ew0FJUAKtCiV8o6lvbOG7h+xTAFzSNdpL+30UAGCqwsFvG+VrTA0jit4ICQ3jW
sggeW55mIBUQWDtl3yzLz4y3+Bcc/AgU0VJzVmGxgk3yfyR+MSau3Mm9lMuJ9OBnDrvIA5W9hsKF
e+cd1h3aD7WSh5s/K5+Jp0rNVgvAiPjwdGlxR2sCQYrpQzIJ6neYAVtKg70H7RRbxeFv6NL7uUFt
OnoTL5p/hSkLR51fAl2Z+5lNI1biNTDTVJglNeeQ3r7MsrFPQCOOamixcX7M8w30k8HP9AAAIfEg
hZ9WBWx7VWGOe7774HYGekUD2P9HCZcXA2amqiM/9Oy7qtt3rHuqmzxmdP7tC3vUoF1Eg5uGL1qN
kamnQH3WYr2Uip1N4BNPiaXN+w5feH5C/0w8SbbQzJk7cCwcHjN4FxtDCHHC0Px2F42YLY5I8280
XaqXfg26fVSZZqEu0CcqOuW27Qq+x6a3Z9rhdRh/he805KWRJPpMnkQEIxtKMyw5FWcZJYz1+Szj
Xed06UMBXEiMfPdhB3enwi7Cx1du8y9tFlhYmgwVMylHKAoPEBFSXaFIH+aXnlCEFXCp3yBpDhmZ
DpubYtwFalQ7llTyJx/MDZsEDpNui4Ojf8w7ooAbEMxtMnzZuG2lhnT6pCuwhAGGQb2WKiTyHIC/
dyqXXR5BgxkSzMAtAMJ39gcpMPOVhh5xf1sfjElMegVeDaQrIgrNYWhxAnVG3lfqKNCeRkxKZ0wW
kR7OyqaheLTKZ2+tVM3arRqsQxhk3fOAZfcALU18ShHlmagDVfXQtB1fPl835PEjNE20Oq9Su3WJ
a+EcPygbY3sY/K6OlQD4a8kJzb7uVqrc9UK33JSfqH18uc7yN5cDLMg1K11bRBpZkE2Q6/CRlmDt
0MmA37fFVF9zp3pA4S8vtWpmk5Y1n7a6MjkDMZNzFAtM8i34k0ZhxGSxdAib7tH5l1gW3skCoxio
lJ/3YM7yxsGq5OYm5FUym6uyCkVT65okxzr1GXWbyj6zXfPodmuyFn/HV+vUHqMDhuy1XknVjB5b
1UWhxbEBbOYnDKSCnDhjhI+BlWM649r0cOApON2tQvwyD29uxYl+y8/9DDgJ2NhUnsERLJM+mp2B
22WQjRmFs2SYSCvUQ75zdC4E6PJTv1o01syi5/t0I1JKjFx7jpQim7IRU8BRql9ELTbxTJD1sQN1
ac/t0f55Vckd5mU7K8mLLw+Nfp7fWpdDdZprBBToVzWVNfq45VBQyr+CkCw6zMRyI4Okv1TWFaI5
Jhm6z7y8cUs+YkNZa4ITLxKNey+8STnKyLA3Uc7Rj1eDLVeH/Kz64Ek5spjvEkWpNYcFPr9mEEVF
rRQEJQdXVDGYiuSeLeMVzwrmd6k1ymf1PTZbODzlwBv8esaFARN9Ng3YYz7Zhw6f2XoqUkEwqMuS
Fs8A7qVSooCnHlyAF2/eLBwsZSv97IO5S0bSg+rI36Km2bgNNt+gPWAZU6TmsHfYmz3rLNmqsKzm
TNKIYjfMeiOEesfS/ejaXHvlTKWciO+04etDIoa1rLjWuF/2gJzEc8s3jOA147VsPQo5ZgMmkQrU
VHBsR4mVlUojS1h8iTQavrUol3QqhNk7A7QjCH1EdFwKEd/c5/e9I64JT0RS5OsQf4AQtuJoo7uc
xkfAlMUqZHCOjiGRBszqffRxDZ2RRGEM4SmSvBDUgsqMdZQuDWUiqX+PnvfBcyUN7nWRD5L1xDet
xZEjyQoFf3Jx7OJH7qMWRiKql8qPH+3je3VwI2gLieRoB9wVu2Y3lPWrhxJdNLp6pw3c1ioow9jw
94aHtquh6X1e6j17P0nmOyhvChnhEn8hUBGGsmqCFcDgbf/WrGIlVf6Wi1lViBGlrLlOpZhEw9YW
1SUvMIathn+OBtPUz90X4/xwwiI7lfqCIL6UtK4ymodpLwiD+yaqUlamV03Kff4wD98+ABdFZNZZ
6w0L3bdpETOZ6IIu1bT9NF5Yf1NZpOeEHsdh1iC/815WPZlMvJKPBirUe9SRnQUeLfvHi60g6VGp
OvOhl91OVoFa0LS8qCEuj8oQyCSaIvLWCg7qn5YL5GU923V29bbYz3taBTKvAoee1JZ+/sn4ofAF
r+6AMBX9Q/OqB5QRzXx97onk1Rgq76ccJ9gKIBzShJb41YFy5BClEKGaXYlSVyBpWQtQmwC/jZsM
tt1mQ8eL4jBcL4H+UWH6bwqTL2RAiw3lnMnYckzQoaP5B03QqvofGnipREHqm6Y+GZBDRkHNzt2N
o2e3DIXh6HMcXUOMgwnX05pDwM0E1eF1uWiWnq3LrdhpQYOkIUlvym+4qA2vonCrxo3XxT5yBkEw
G1uj0o1tyygfln9DjFvIH/MTETt1VkEEMhSDLtwMdKmby4CIX9+iU9BRcgf2fcLjT+Qg077dWsUX
V+WIHAh66QBk2xAyM/YBR1S1avRyZXjsdUmG6trzNSJ90TrKtu2Xd+NZibItrm40jy8AuK3jeeZW
roqQ7L3+qC5PqhVo5G0/YjnJgpg35Nezm+O9kRjhXnosGKgXv1HfkoHRkjgT2X89fK4UmXMN/pcs
yLVzMNTSZnN2rcNyG0WuYqD/1NLzhOYjDuSYHZwcEgz5n2TxzUXSfJUSQeqTVlZFo7av8E1Nk7pO
FlNjJRlUTNJAlz0flN8l6mPCHazxiVm4CJQ3I3dtbMB5BqbJ+Kzp9L6MS5ITstyat9Wwus4xqrrk
gI/5XQ/1e9N/2mLpQBHPrkCzlGmQKbeZO+zoR9AF8EeD4V6vKQHzS1n8p6WQIPMDkfNGzDXNUCBq
aK/dR8DJaZZ16Z00fEbOdBWAPkaJJBBcNSrTvBwwgp9tCFuzVeXNXLNQkwf5s8KkMr0e1mcvGTDS
vhnPfJi6jitWTVfhuep0fN9U9h4ffN9/kNfAz898QTUYvdn12Z5b/S5Uy3fF10Yt/fjiMUGvZFZc
dmgzWS71LaQ0+AzM7tJtjOD826klbr6g993BMeVVodYZfAtBj+cOQhFco6/7teKSJvaJkcDKqut2
pcZ7eZnYQJYtJceXpTFfpxUNmB6+M1JxCRcf0iLcktLDu+GJFinLEgz+HaCk+h6hA/1Bl5tkyzRB
3ogryAFuBtwkwdyO3OgtD56zhNoNiT9LB3OPRzcMBBmMkT472i7xOp9KkIZKu7dD0/pYSQqAPUX6
P7wFU9x+r1eFENRq4VlnqZfhRVtTor6mi8oJmxzfUk5c13tDdA5Rg7sq9f3XTzSKuHba3B5DNZXN
0WUNBCNjOKuPu9NTxECd6Sfapiz9NAwmjxIgZQh7+M/vFAIuVIRrdhOcc7BRh/DLpgurTD+Aj2RC
+mHvA4vr+xk0yPhuhjp12XbraEclwV+6AdumESHQj1fVnPhMznQuNC1KtKiQkeB1YLyLqwzlVCQQ
lHJPTVoOvaOgYniVUWfQo958vWeSNL+vMyWMO+J4TTzOOhnhv/zq0zRCdSaCG/egzy0HufEYd87E
o4kyD3cWcfzPoQrl6sq1HJwqELEc7nxlRd2c5kxBQjl0v2lT/mMcHR8PNXZYkdqzcGUeP+pGXDP+
kB5h31vJv26qR+8kp8fG32HaXO2809J+AR1DqTh4/ocAXLDpjDLqd3C6GP6dj4Ynab1a73OFYJWS
HJKpTZ3Zdgm7bKdojWmOHkBUB2rzWL6u6jtZ2F9/M15BK2e3D793IiX803qJ+qgSHg3Z4kkosHfO
LWlIxfUW+/hH1BHieIpHlUt4pXcLFxnDejGsXihzmwO4zfpuCyuXwn78t1tNKe0ASFkdrn9wNKn5
maYWIV0qquVjNb98jThoLnYXtK7cFghuHBKEiumYOzgSTWEoR/EgVKW0Quk5YM5uX8A8mVH2S3R/
ZRh8I2C941H85SNJKvv/1n5M0/05amFtkzlUfthbFG32NJaL6tbwbUjAm0aS655J+kLu8QMfl5KV
AnAjEASFFUXpB9jh/CoYI4+fJjZIA5rv8WaUrPHYMrbQNNI22SEI5vCwL6DV8FwFtAkPx2hVvCk7
1scP0GtCGPkHlLxSHT1DNMkb5+9DEbx6SqTBY0B6Q7EXogFiv4tiosmwqEXicI8pCWbE78TzUM9o
qrPS8cx0qgdFVTp9ZpJLwVFQ3cVHqKeforGBlwCzpGsrEcRVPns9pUZEC5vs6h9ORfAg8EXtotj5
J+/QoXIjBJ+ZRaADIKM84Gbdv91r9rpzsT9sZThKTOQWbwxoLLS3smkcetoBmgkgUgRwfkTqY42l
/KJAibKTsKwJ5TulGqtSh8CA/Db2dX8/WTHSZibPvPy0o0yDXaHLSM2A9Ubno7PrRWlaeJT+yGap
aY0NCogesnzH22UlgfQ2VuLX3ehAfsbHswZ+0sikUAh7Icc+zlOwytQkYDovfykfsBi+9dqCEGir
ru/1WS7NuTyezYhrkAzQ3k2BHIGEa2++dlWFQjrpF+YbowE9KdrfUtKDH+MV7drFRHHBVZ6lGNGV
0B8xQPBtZIaT2/TjBVs4k+a7BWPRAVvp1Z6IPZzQJrZVfgIa4W+OHbbNznWmI+AxZ1P/XKwja4BE
4swpifoGZn+Z3mEETue2/RFEijRIMyXd4KH6rh8ykbyofp0uz1gsGLZJayT02gE2ezoYxKit0TrP
jvQm1DfDkbPP9vsUB3dgznXaQ91bfQ+byjBMb/nwuMZFypPtUHrD026pij3dbc2hdQ6PFefGozax
/OcO55RGZN4xtgYorh+EnapwueqiVM3WvuT7mXo4B20a5Y/OP46tGiH/hKMv4CiCEGLzz965Vwya
LPMJl3AAcdl8g8Yhki0gvme3xlROf2+xn9hJt8ZcxwZRvROhMXYkiZoBokxQ530XOq5BiBhMpRcO
X4vim4/RStEeVK7fUVbjuR0JaUkLqZq3fOcMJLeXdPcBi+PxN///oIrt2nSD4vPEnNgtTYdhxhWO
40hJIrDGQxHkQZtsrXeV44FoYostr5YrAN1ZeVA+gMVodgBMe3H9UkJSaTACwXRYWqtdZYef4+18
gbqpEq8XBDkLq2HQ3JMgyp9olrFbF2geOwDfiBU+iPopW9Czrfku7PspJLHuO7LcMiItwB5u8ebR
ZksPCFZPiFhS62gXKrZHkuT4yjM/eoM8U5OW0yZIYH173H23YVUZUAvTpGolS/wpTsF+W2L6FA/2
0XM9aDy90ws0g/kg6o45JcFoaFtdcTQ04bzOCvmeR7DZou4RoCzF23MFAW1XpyZ82uG7oh/v9fwq
P7iFjtyVM36Z3bccLqfrCDiVzifFlQlf7rZFrqT68jhIl0ulKg/KheOX/zTZOYNpMR5DwtRc+x9B
6OPq8loKAlQQH0z7SDSeBtohYbNdwWLotdcfxdjE1hFlO+y9RMGWggVvp9vDmh7pIO3STyPoIJeS
pVqQyC4621CmBM4VvUqsB7zus9hanDHMmxJFWB0lq3scr6nDxVxbW491tFU5JY14S64IyDyYXoXN
cNJFFFft5IxSWUEAKMay2bPIOw0QQHZ8r956ZU2mvTWy0VZiUxJzWAG3A+5Y+p3uNfBrP/Nvolhi
gOnnn+TdkrxlgZ1I4yFaen1+0Y28ixegvnOag8gFINNtrJEHLaXynqIcpsM2Ge0kGWZUZ0eTU4GS
h/qqC+NCS7RRXBHsdTcl+m2sqrh8E5nyxzj4zyViWCgg7M/rFbyuqqnMFZN2ZMb8yIwWHjOmC2sz
+ibaCAwsRsxW1Xjy+/8okgvsIzxnJoljW9RXPqIurWJDoMZt48xYCALWtb3Ax9+0zhJM3EOSJ3mD
R+G/FnKi+QoLlJ4ks/XJA3YimFGE86r/0VbpUTgtzZXHTUgSKOBA63Znh9HjxeB80AuRTyD7Gof+
+iRhrZDnH9BHwnxEEqpiJ9do2zKHTvcjDH6U3cmkMlwr3qf+0Jjbun5c5/ch7YOtZD4kuPQebSta
Ak3AQkHKyFc684FbLizknEi4fNulf299mUgOtk5xqb5zvm2AYfm8KKNr+4GctaFevaMtwAQdpmuf
jOxt1Om11zF/9dxThzuE/1a4nO2mXso/8YsifF8Y4ZAIawGSKtPc4bj8ZoVP4DgEnTjOKFdmwD/q
xmOBPShMTb/8tFnSi63BQF2O+hSKQTGfnPJ+M00qVeL1UdpYWf42gAINEr479x55jc5PySFofCMS
EhtW21u5HC+bg+DUWMVhZEaqslnX7qRAB7P6U8cQKeVUrrKmp6M2ZRu9ckZnVZU1DhoBeOpfADIQ
/b9V2KbibrDpbYPcUPCovfwKgixH22nTY+aIJqGiAGinGzdMJvwcH8EimGUKN9gQUuBOFGzxCgQ6
ZP+0jT4L9bYnU8ZNSqLSTeTP5zMcSCc1YcXhrNuX4XjPOCnpLaL1yygSxkrZ1HbI1UvgmYMWeqKP
dS0eWH8hSuNDGcWo9+oA1wZTPFu92aNxc6w5MDwa9kB7+sdzAfR6nLtP/PhUs2sQBe1nuBsUHIQ5
/14mJBUvJET/5buw33E3r4/ME/BPGIElO2QMHm5KqSITiyZBDh+T4YWkKUZDPXTQWf29TucF2EQX
L8xqDTtUWeLuC16xRM4tBjVHZXAZTblZJLsWI4rF75nyZDyfWuqE1l9aiuFYItvkrAt5APeNprXl
8KSeosZTv+1jM1ZHo544a5eUvLl33DdYTxNO10V9vIT7EoljGYBIMPBZVZIQgDOBMyUqlLIpVJ+U
5Qn8ARMynH+uJmdd98FDca10BLDtBoY/P7x00tt3dctw1GUlHgUXFZl6qBaESKY/vs1RaRXgqydI
wFl5dzeBSKb/STNoOVuv/CoYPhsCuNSZaZrp0/srrqGh3KGFbh3WKaYXdoCHBVcUTQShcuNJ5hf2
YfE+PzS0TDoOwDH9IEKxRPkIEShpyMae9sv/P2i9Zk2VO4imzPoNa8Dh8CpaYQp0AyDXCocI8UsQ
22pNRi16tIzC7K/Fba8JWVhcYnwbF+jbj404A588bJPggNE2Uv5Y0b0JFkNBTZo7LbSytteoqPoC
GJI3eq2MuTwk6AIPiGuold9ajvk4gAACMTAsqT7JVuFiA9cnxBdvVD9dq/DRPnNOzK4as/3Z3MFf
9pT4O8N1Oga7K+NPF0kivUlwQZTQV7IuaN9KNffORK7jnAyrcP/JlRv1W8B+z4AF/B0TJt4bFNjD
JzG+ok/qmaqRjVGlf/yZ4n7+Zo0CfWLc1voqas/SivQWqCktIcRhnjB/gOWINJOdqzPv1mikO6WH
D8NS13el6fEVBqzU4euAyJkv0ZGwJopNw+gKTGZvpnmGnDc7pVh9IbNY71Hy6LwulXQAKn7DkcXy
kpSxu1f55v3h6LxKmlxq4vkHez5J/9Cocq6AwVRv0Nhc8xcpmzEBjpaVAD9EkZJ5D1U82OeR2OvG
orij+QG90iuFX2gg24ddjKgbJo8YY6RC1ior7RODvPQzmUWU6YpwVZP4VgLkFfezwPaqy/jQcd2A
F/9lnR8o47JsQAXu/dwK5xHRVMsfuvmtuTQSt+6BKs5TNk4Z+pokcag+Z/t8hm0973bjX+qFQFnS
GTTKcwpdvWMoV15M+MvLzm/28rAKrC0ourtc7J1qKNQF05GOLL086kBE77v5+Lk0j9SP8pYb5ALO
JTfd3mcNho9sHhdFbfyQdY1tT1+r6/ihYWHiNYUch6QXLg2WZYGTrc1h9Yz70KkVO26//kPY+Pgl
9MDyQBDHT2eTcGflA46ERiQjgihUeKD2PhYMmoSdELHLsBSFdAAl9MBYdjGcvOu3dJm7k0pnoz4I
PQ2UAuy0ozvAzcO7JM9dVqDQxda+TgNVHBdh43a8iDPpGYSwVHC6ZfzpDOBZJetJ0knyqYcE3/GM
Kv/ptUNYGDcuhzl+tFDG7Pv2/bzGLcUMWEZ5YGHwAufu1U0x8Hn1KaTnNFQf2PB0yRfEmWgjdGqo
tXlaAXmjQrihSLLSy3/u1C9qHDSp0jFJDGGWuCQI4WxhRXQBhy1H+YH1LUvQdHFieiWiHnRhnwqr
weeAgskOxkBBIVkMwTJtf+s1J2ImBhiHLsijd8Zoa54pnqTi8St2gBrofT4To5f7JJKUtYfgsLE+
AH5SD/4Vbv1lbIshKIGUSRyCclKlK4eH7d+TmYV5OAfFcQiDs1LAbdQHFkSOdepFQB2PoRVtlCXU
g2Ea+LTFTnN74bzbY9E6VblYnga5jBh4E2D67aH/mskm5daJ2nKJUOHPB1mixv/C1UrcQuwjW6pU
PO3MnQYp0oHDeW+qdqJBI6Ho0l90VzCYpOFJkJHj57dKTxtX5w3l1WhwjT3DEZJmWe0gCciO8/+l
XBJiANKet9/amaQve18B1T3hyYZqm1PP63ro4MMb91PQbgEU7l4T0sf8nlXSZAaO2qAniGzDow9o
dTEi23N9L1RCWhIS8nCQS4irKZi0SwuZn2mCF0CQIHuMCIhxCSQTn4cNX2TiD6MbZ6PB3eECEC/4
Gib1DF3fIKCIve/Bu7WNDoV+xdsK1lkhN+hcrcr9CqY7sQaYCBwRVN4+8m8TC0MYXMDAo1uED+uE
At890GgHaRchX77yf2+MCoZSgwj66wM9BQvnkgOSrDsMTL1irQUTXCec0FS8vRlCR+zpRuKQA3K2
UtKRxELzYjdRdMAruq4wmRcMldKLMn+HYV8wHEnzfdyFkDrF3wonNiYTzQnTheSMI1ZyfuTwJhJb
JgcmI4YIH2soLtx912tZrejG2tFDXAj2SmLMhWCXWAl2NJLtfCALQ5gvexOOaUWNXxuiLCuvkCIs
ZzMPv7F2m8Wloa14c9RuVy3BLrCZhOXv6GzHAWOWwtfXB7yxuDpnv2JU9Kfj9DsSzV86sO2mIh6z
oWSsw0LNtBmMPDvMxIDoIh5upyawTW6+/yGMHeKVAQ1fWzNKwUQxTXRqqDujWoi2dOOU84DeXav6
KGqcwO/PB9vUJAQUwtZ6tpen64n6zW1puzQKvete6H0bEvbPRtqL3/iLGc2taC/lcVL/3Pr3zlwR
qNwg+dGyZJlDDrceVEGIvqCcfAgByxg3qi1T0sJ+MoTOe70Sw9Di+XG/2brjtBT8nzVzWuQaR1FJ
MZ2zGUfebQ7+zvxRhRdgZSu/3glB2K8jt2fvYMCUY8IoOKDA1Fm7BDZoMkqXbByas5/BUOMrF1SA
zG8exP1J2YzWEq1QuoFc1v8/y8qnwRjFD3R/FqIxGzFCMzMuxG1Z7Mt/rqGP2g7DNc7b06c1Qby7
WskN6eD31S3Ns2LezasWX4MS5AKpROdwWqAr/G5H7ZwEVYmhfddYHijE4nO0rBR0FP2/M4hdXXRK
mWxnIPGOQxmzvKHSQ11YURmaOZRzwm8eFVNgecYHGrC5rNG21VWSnJkOzGSNhXFFmOlhuptcEA7p
xPqZlB7/tFG68xGaXxyRvKh8/APaFRh0kb4MhwcZclrh+BXO6L/Md83BLT3NbEuXT+vEZ2rgv0Fs
0/+4Ux8ENi2ER12dP0VCpHWqVOu/acnDPg+hI2jFcA4b0O2v///MyF33WrvLm+C5v6FZD9RyqMsH
eTwfYa9ZxlUsfMwitsSX3e98CezK/MNq7JVEzk8E1Cqd26nwj+LR6/YrqL/TE9/7CEzTXWqPMDHL
2/uLCDbdj/JOlkuNMCiVmjOsfPyHOAbk4ieXSP1cXLVf35mW3LPYR0Wl2moWRrfM3Cs52fr4Q65K
kinb3InC0oEixM4wVzGzxdv2CTt/JGNdSESUShrw9tCqDYlc/+JMlQ+nckUuQFhApz4oMGLrYR6F
eN0jciw8Dvrinuo1UInkZr9B5Jb03gQGAHj7XPVFuKKfmdAU7tKVH3dBAmRnlsedX+6ueON893V9
9SrTdw2CeEyRNumwMpdguPuM74BrYgF5+uPvWSKPT4Ywdin8XHI3apx5ov+co+Nxixne9rr4hsw0
24VgpLFe1eqN14BEKAY/SQ/SNnF9IvGVN3AeDkUw6E+oh8EmR5BqVMAVGxUMc0An5fV35vngKmZu
pYqRy3EFqhBM1XMeCD44trOHRr5xozrLnB5XYuflp5N+YmZ0HKXsXWh/xR6cRAp/TkvnLUpiyQY0
oSmoEfisG7xAEQVgIx8D5F+rkP/QC//3FgGO1g8ZiCPU+Azz2nvQzNvkN53LN+zwXFskJnHtmm4o
SM2F2nffMsjIx1+BcRockZHulGmGH9hfX1NRcqsSef4i5ZFP1jLLWmIQeTnCXxSiWZO7PPlj70yV
FDzjWxTBFdAo1qQD/Vk6WSyKR318TvzJ9Xk1cV9qm82yk/ta+mchQfO5s1WbKCKnBHsdwkYy2GCc
WlZvY62h1c33oPeOsZZDv8RcK4Ty/hcIufPtfp08y2u43ArTO66wTLPgWhyvvUDETYkIFuLcpDVR
6PKTv8AFSn/hJXmGICDslnXEsR1+3Y3SXNbnv/3FL6pUHADYF7aVqWZt5V4lPYPKe7l5nVAnd95i
iRLGY49Ea+QAi9zArT4kBOkOURT/TgOk4AtX6nNN7UhssdAR8fb5JC4q9EEMhSXUml9ePpk9aOxz
/6FCnXsnLa/9jxrz1gSv57qIwTv87dyiu8LeXhE7GyjbVnPA+kh4KOgz2gBx+H7hl6jOF+KOFrhc
BOUElpvuvjX2vCyYBUeNSQR7ByDcZwXCQMEX0aBQ9L832h/of80Q2Z+ibCNzHofrW9Fc2cSjmBT0
IsdPWIDausUd8Je3D+14hEX2fakXAlo3xyetHRSvC7jqzeVblwAckDhLsNjNaj4+L/wcKd1TiKzE
vW0mbOvcYeh2pf7hHio4gJOB+wi0ZjtUnxLDFj3u5R98zRWyYtw8x5DxNrmyL73t2Y3g8W3HzXBM
5ZJFzSKw4dVMfBtHqiYLrw8weduyS8cP4NwkmGs1m9gfQGMF4tTesyhApsvDRhV7xP/XPSWzuqRl
kz81qmBuLMXSJXO+SUifEy2WzpqLgvQwkR1valCp9d+7oVyqcYDx7DoakQdiyJ7BLZawJZnsfEH0
9sXNQso3cL/0UWpCBmAX2ui4OnItGF/IRnvsBa0eFVaghOObnzT8FV47LGVL5DTXRE3E5EYty9oX
flFjFCyUWr1NhCw+yyH1b2eg5JFk2yvcBAP/Yvtj0QjvrWmoZNp+INqAOdXoQaNLzMkDxx6ZCK5o
u9H7ty8h7pePN/StJhsMSBHbBGqkqH7YCnqRKQOuTdBE9o/GevKh4qA6cBvNtmBkQB5tJmNbg2Eu
dpaq3sPnVvcMnu903sy1t6Krky30KcY130jAuGPiTw0NOpgNcF6t7Rm4Ty9JmOP3TDakzE8arzKe
LtxOXdEwRdDlui+w/cHDLL96FCCnXLaQpA4cb7K/UOW9OHKDiQjnj1lgnbTi6gIazc1QIGQGayF0
RNf0fi6L9uvjKUwnHn8rkk2D/cdnNdjJ0/NKrp+H1A05a5sgZQ7SpAUWIzBGW9kWoTM6Dxosadsl
glunnPR4gD8PSKqGsvdZ2ZlNp/8KjkdRJcSxsc377KjY0BmU+wKrxTHyD48I/8iC+ObYPSOkof6W
6oNinIusNbRdT4bChNnHZPd2C0avunbJW5SCpqu+mrZYtEB3fbfj0CuU4oEc6LqYV0dXGoYmkXDN
xcGEwWJeYXgac4BNNWVS8JEUYQQpHRSVx2g14rNQWiHfzC9vWDACKbHkhai7+eBXNzJOR748T+SR
cLtx3dbq7358QfDAh4C/th/4qX/F0hH2Ngli4R+a44QtXnVIVC4AOFAtVBLwKwru9Ry4wG745xWB
bWX/NbkGY2qp3BiW2TWUyIJIW3WNr5XZqtq6LH+tPSvcS0n4D9DadNrZsbzyhTFgxy04GUCLlXIA
Ci8RZrAKzPYShNDFPI23eJ+XpX1Wr6Q2LeIJZnS18/S1ePR4ql3Du1pQIUXMOymP2RAeMUhcGejs
C7dTFSrXOFxFzXY5Nz3kOgf64oEKgZ8+8MOLgmfhB7B0OGQoBJ5Xg9D9SijzRgKvBgZtenck3+tL
Iys02WoHrvKVwyoSSV0Pvh0lZangg9iPhdlo5SYOEqXWlFjy700GwzfsHcX3Oc8PKvEuGc5YZVUx
0+sx8eZgRnfBmUm4FcVJz4TypXd9BbWnobSzJLOFmjvO1/StspRDML8hh9A5MmMslOOEJUMcsyL0
KGxOARRCTyVAO6aSFxqNfVJPK2j8vrfgpKq6l0RrKnFH9FlqfysxXvtShJ6ucK9RBw2ijrgPlBmn
qQssNZsfh7QqkcKSkq5BbvsTanDM7OqHgHgOtdD9SbjwoNn5DN4eg9vRvOMA6drMHCwR2M0f0OMf
gNpdYhHifPD01ZJ3ZlCD9xI3QtPlKT9TJuoH3CHAIrbEj9IfsAxwGsdvLuGUFs3l/4kfua3QNmNL
rgyAPrFW0dYAzqPjxa6kJd8CREx2iCXt/Uazp1G6qEs4U1V/5m8OrO82o03RJXyTIIuKgFTc8SOQ
XpN1GqeVzXt77DbRMahzMoMOGw8InKOgmssTcw8ackOpltKwAoTHCGzS9Y8ESfFZ6vWTYtwK+9Hh
CavBKCAw5QL2RZgi48ozJlB/Lf1x1NfxfCUHwV7RGpSSn1LpBAtsRTlL+S7vL5S7CYU2xC5S7rIH
ymih/JMSj0YdTxP1CHpsb12EGk4h53zAkACtScb84R26LyHHzyWxtVLinQHslwN2bl4+GAEpwk1v
PDuS3ZUMDp4D2cHLj5cvBr5AhdrC5SP632qU03idAPXigGVWcGxeS3Lnr3zWv9QezCUmVERLwS9N
yTbD35/ES8+eKWlHC/DDVc6k9GRJXnN8hGUnQwJ1zajPBvq+32yvbIDTmq0G0rUgCJ2hAiRboQnS
bmOARBP/nIWYdBXsJAw4fxVAgERNckWj3ZqQ0MqMAkw6i6xbtUjNuiTvrZoFkuDgv4UVLD5Sef6Y
tKo2UJpbQWBYO4IyycnExugtHVt9tJuRiM+y+AbhjEMDIrURvcgUN9/NDogZ5kDzsF/BoC4Sjyqg
FeGapbVUOyzlqfYmNCC8YIPkQC/AvGr9CjxSpFTbnegJRef/8Ywmky9Bd+Y39fJ1JjT/7p1GfKjP
C4BB5rVuOtfQb33XHLTvi0f2omWCrx1A6SRVQSR3u5ZMTaZPtX0XRVdIUbU+21oQF1btPo9bozvB
OFx+1GdEgxHafTRcKuMPEZXnRh38+Pijltj/PaHiz2cxO06Vnp2Q3K91mNoK5PGnxYqe8p2C/tuD
pXJtK4RgA3i0ZOTqISxks9mYekaizC/DhN3E048VoW5d40QDRPz2bPW+Hf6l8vblOC7lsJF9XIQ2
fDSSmy9h7yNr4KgxrkMKCshlLl59fkpUctpNFmcR0MnyhYp1IZeHMdoeccHhBVGLbNCZ0P03VFin
mptphAikz5IV+DJuXAuRWfVshgNsICv5WuFe6e83HwnArlhywWDGokHQYaoJa9Q2OhgnRB42bGXC
5VVWutHS0jZESJbs1OXo/iD7xP5o2e2pGXCYnTcSEofMWHViiynb6/7mwCk+DCERzGJhSHDTkbZ1
AGf0QXYXTzylG/Yw+jBb+I0gF6Ha3x0TQYzEQH5KpHtx6O+yIT2Ni/eJTkLDBiuvfKhrU8rDkGHe
+Uc+sK4rGqF28qrNe9RmS4TxZzlzP8YppDRUoIh+cEskuNLp/WQUGX0Vk8Iq76HGAdFcolmK1Clt
+WptpwM0jMNhokEUJJTugj0KQVOtZn22RfM/VOtEp2GeGw+JD7lCANCipFc2bug8qRN/EivdBBcr
k2Vb1xl1I3RPBAjGzblkeJIDLlVdyWejQe7jxwXWVuHx6NubheYHA0yp21n2WcpT/bEZ8QzJHGMA
myjfL2KAEY1V/PKHvBx4eCFB1biKWhsEWwOVjxB7aJg8PI+B68t/LcFAqHPsYMuFfmQHDTU1fXm7
MMPhRPLV84A16NWK0T/DT7ZQ4P0MAA6Q6K/p+OwnN4cSILUB1V4YFjX/hUMpS7ZiKffm4P5qlRb8
Anw80gwJ9bUmIELkAEebNlrJuFtfFyJJEmwHqmPe1wpAgd9ucItUduCqfh/HnZcIv/LjLJ8ZVwYr
2hzdn5Yn8+c1OeURJ16sYDFwESlBkONOvmVjyU4YNx6iHLzDEq0+zooFYUqM/iPD9eZmo35/o97e
rAO74FXrusonQIQ/W0qgfykNSaWWscGkWXwUL4tgYpE3DQ1f7rseDqY/wIvCbrC8qmlzKqeyJYCd
5rbUgWMhDDHNPCWMF9rPHdyveagF13BD5lanxRZDhvSICJEZCyj+rYdGLVC8JJT0H0V9K817z8Z1
wejrmgcibaOcIpXK/9koekbCZiEHUlCECSQxWLIq1zwne1cIZL4UuBEpKEmlme9BmeWWGQVFBvyG
jl4PWAA2JUVfijYazH7w+FVJ7w/GPln+99ajVaJAZvOqaZyYX5r/BJAtFY29ZFZko0psGsyUT9O2
l3MjobMBhYqO+phzjwlfGGKqEvgOBB9ooYY9q/tW5vgQF7FLwnwrcGMbNvRDHZ2Yk2ga5vIJJPa9
wbPJRb/oYcv7J6cMg+PyP3SCcJqV9jTjsNs0Elx3t6z04nPHLBPRE0I+Le1d4wbG9DEb51XXKBB3
FGTsEXgnmOEzv3Nd23PH9eZ7+bMob4xdavUek0dap1tUiDN8zZA8j0JFMD8S/dC9z16wjbGRmUfs
RmtwqrFwf6oKtsKPWjhbMQUvAloQ718ITiTgueV+q6kT9AFmcW8f7dJab1AHGSU4pzUVSJt7T1AY
1XVBezOTOzsSS5pvefbrJBHUPbJnxzayiB09R6WvmvOu8eS3akPPWSbEEdU38gLz+r7/3yE6dzzV
XpQ27YRSo3A+xRyapSfMa0dykJoHbm0JMOUFCWySpEKeaQKJZG7+BZIQ0n8iL/EUpZZPWbE4mJcb
6tEqSiSc/gHL/A6JHjeuXp4OmZpX0IVUAdOirR9M6w6DOBL6Eaau2nGTAmDNO683/TN7syS4Yoqh
fmws9qZ2BSL2DRdj5jNJctMnB6deux9kF0G0DGS74Ij2rZJpu6/Ve8rhFQ84ttQhLr/zpPh0/sU+
bbQEC2zgz2GjxQDveGpq7QSoHUy2Xe0Tl8JdvBeHzpcGDL5FyZ39wbwphFNDhvqLvHMDXhykUE3R
gX5B9nkdYLvtvCJ7hLeFJCDn/GPphegHx09/mfR2iqvEbL/Tm1KYcsKqPdzQASDI/g/w9KihPMJ/
L7jGs3t6hVyfhywCAyN/Z+sJ7v9v9iLzc9H8b0QvAFCQdHSflioC7minB8usHTziyM3Y3kUXViDX
bmCKxkSbPLKjwPQrQp+0cADVzzGc7eZZUs4TBoey2wJFe7sGPIdfw+fuxOZG3KJyPjGJhX6avHad
l+x3zv0Fx4T34QVC2Y4qBLlq3XdZx+sjsSLAq/X0tVD7iPjhZ0U4Q9kYVlo/yGOt+rnoeIm0oM5o
g3QGgkDfBGkDcg9EG1LBzpHVUvXhOMlAQLQ6hBQ0veq9SfBnrI58loRXRkQWh7cNYmrK79KAxrKg
gOFC3dTjpRvvJGNodaZXIIsct49MkJpAS84rUOXvFap6+fJYQ4odOhJhQeZnehEi8k/xP6UARaMA
yV6JLNEsIMtZcvIZg6oGbqvMRMbCWAG6vGlbUDtwlDSDW7xqckTh4OpXhW6yx8+29YWtDiQxLYpu
/jSin8z6Wf0xVVkIbPLw0t+ih5m/67Grr4/0ILhGU2W+aM3HAHnGAczStHX+I46GNL2nm8PjlYDi
0Ak/Iyf2E5m7b70MKF+JLLHesf+583BjfTUp67E2rDrMFcKOo8wgdJQoR6cQtzdhB70wQZMB+2qV
27xa9rXUKtk130/buuY6a/WL8LjcsRloY4bZ1YA1IYZ3Q8peQq4zFlEzPBTQpNAVgUBrx1vybVIR
RemyJkojOeR9WkVLkRnBcfFdNG7L4dYoGKYpCQb26Xc3m3hyVl6ZmJq6HQJ1WEWpv6OGptcZPESy
GeQu5vkWhDhDpCzGfUDUZbB9gqpdQOFLgsHXndFR+LF61hcX979Klj36RtGXWLt2VoteQDYhURSV
AEujTFZJxucC/HXC5jfUyPaeC2B6gEDIge8tI0dW2jKGYOIJBWJh0kyLkuQp5XuU660HLXGEY6/X
zF1Vx+QRWPISfb8yNrbTzzSdxml0iQK9fFRHxiD+5alPwznUTitwbyb1S+/Rga+0hGZvwQ9Lr1wt
q0+liM9gF65V3jgz2DjoVERAMFQqw4VUx6ceI4Odb5ndK36rc1VkC/34P/gBksLHD//th/HWqRIz
GsJ9botpapA2cYwFkE3wp1gWM9BQPg4lHrATC1oA3KDviFNQcplnjS37mEobym7SsF4wdpty1nfg
ovpF83Xt5HYpSfQvfPx+aAOFevQF2bFmyYse2cXx6dZoaEs3nP+2HvNTGwjV/sYxYr8mPwlumQ/8
rHx5N3tZJ+hnLS9YmxT8J8zgkB3LiTMr8Wtl2eNHiAOvS7XvUdJ70nGviEpS2U9tAjZnL7DqMOfn
Yc1+ZqDJZMO5EF3GpaCIANx2oQuMyXNfQio0TOljcj9PB/uLgB0cKQ2NAMM9neCoNcN/yhFPtwiL
2ym1/27mLRdG9brm+z5v1J3p5B6k5G93JrzTLcRNOP8l5eiL7OkfeguKnx56DIYKEMaQxuev4C/w
Te0D8QLGPg0cASeTrzUc21wQNmAHzRu2Hyj3QYqmJPiXnlJmFLLAj6nVl7OGJKYw1D79DDsaMiWA
AQjM43lxi6p6zZ5r/IUPEf3VYv2F+fymDnKk/RCCtKyW0FkgTM6Fj5UL4j1ejcAUtoJ2j2QbhVB/
8P/25yvPNRFDhc0iyPW37ZCMijHB3BGRW3wXf0hC5agcSf0tjcOUFu+coyJJR9F+IDWA01wvrJEJ
SkKbrZ+1DDeNo7TewqGMR3NA1kRbwkYucKGlbONndMfYnn+leuEwSF9hl9zL+eV216CDuqXV7Kbk
xWJ7vSf+pP+ezkND0PIQiK5GUgsDlkoAeOFyosM0ZtKaTPAQYQmWUXEA2ABYXG9pJVx6kumc72W6
Uf3Vj0zqrqiU6HQShUG7AvjbJUY/9hYjENYlZEzyh3hkgYV3qkU28w9Gqw/b8koSgvFYojemnXPO
5ZXSbJ8E2GxpbDKvl1N23MltGoNuaTZDOe0OJITDwXaXV4DefJD5RkcSw7UCdE70LaFGamGY+ZbS
iduYNIarnkNKZc3A7wj5AzEpBeuArLPjfDxuVkhdW/oqwFVG7mBmm+oJ7uEJeKYYlZGktYI0IbuJ
RXyKQNPk/PI3IquyA3oV5yEHzhzaBn4RY5dTW1zHF7oY1UZK5KATG403Qp8Nma51oUqUCH78XGiB
s/q18kEPhVcr52pJ8TpAC/jvlgkrFNx8hjBR9srjDrQ2uV7RRJxKPEb07Ci1fEmJU7SewFl//oHi
QQn1EEkDayZuokii0J2mHM8F2TvlBftV42EgkUQWY4O54DmhS+oehxGP1jTJ+xboPV0Z9S3QZ0Gi
lOsPC/gLUglVGJP6Ex/FVIOzWkrDHcEdp2PBKlvzeNwncHSKi4aSWwoeJJNaBbzW9c3z1iFvniHy
EMAxS5o2iUfeVEYTV6G+UPJ9UpPACgyq1xMrBGyU0HFoc/kllOQAk7eewFrYh1a4j2zTwk2gq2sF
OdVQ38WYh/1g8R2v7kDGK4hTpRpHfNu/WLe/e9r87BZjV2eIeFdXKRingJydR9JwD9UubJdKGEmM
3cHfKSC02mpq2lSBYP6VjPbOWEUBWTps7eKYT58FGPw6jRHo9QuHMulunIDJX4/TAERfkVUSDi3z
KrQhrTIoTGG2oFBbx0SOmlv52YUu5JhuAKrrACf+u2pFr84OBX8zPyUEd49Q1G/nNIq9YCMLS3ab
GNe6l8gM8Ifp7YYOVqwBjc6Fp8PP/GvkJHs01e5zqadtdXzODVKqZ87RklVjRGP1pvZ+RXzL2HNb
OSJN6qP08UWZJYptRQWaYBBNBPMmnAiVphOfS8JOjc4I66DITVeea+SW/K9FnXJ5WrQYX0WxLojB
Kkqcey37bks+Un2vZQ6Gdlmak3rXqO7wTBuuQrjaWs1gVkoJakpQdUxQugeiyM96bIWC92ui62A3
gVdnV6vsqGzWXQz+ueheArisVD6bUxyqV6Lp2wi+5mqGK/jW508UtS5yDNhshutDCBCftUJyUUey
VB1dFw2eonW/l9bCxvKbYFWPL1FdSn19oJE5jyKH9tg0rnyyoGYdM2DTQoRw6SX6TTQWt6qyLQ7V
xAvthY/yYFofk21VED45cYPoPiPa34QHQILcJU79w8vZ97h8DFgpGzLmGMAxRcXmLuktjnXnvvxv
dtMZqZePNEOwFiVhDvjEcD0zPC0i0xCnew+x/2+vsUyhHcAmFODSlO1LzTi/4JE5wRZKeeyt49Bk
Qo47Rojhv2lKju6mcn2WipBkZDLtKsmMD/jtiPK2u2DLHKDfU+m0et1Du32XUIfoTaLfGRqitbG6
v+dGZgb6J0XhigBzvmU/EEMYF7JH5C/R0iPzlrX5NUrDNgfoipOX4nm0b8HlRVeniTUhTcw539mR
XTBZzJqQcdmAAkEGM9O15wyp2fP1Y9Zzh7zOREKCeC+bl7Fj7yAuKd3/rSsrBiu2ouACJtiUuvSu
/CdUFrWDznMdjmn/ROPc/7v9yqZLd9l8C5wTjVhji+apHWktXqkwliOX0qXuRZXNopWBLjWrigKl
ZeJOprTUgDFtSJgHJ/jkLaxHQ+GpWPPsDhjR4et89mbeIC+9vvNq4YmArz2otDGO6B28g3Fg7GQj
8qeFhP2z7WZKtCQCfAy7Es7cyJNFPkB2fI+nkqpNNlZfGJDGMWKShY4LTRN8tCLOUa8l77uRgj02
2GZnnGRZaUV0utnwd1cUxA3b+Mf0CgV/SouxIFBHkJrs8Hnq1mBlEPoprVvbTxSZwQVGxzFsLEUL
pYMLRUtPF2BEgYikuN6DKHdFFfNU4ryAeaNtisR5vqyIneuYSuS6i4F1TsxaydayTHlk84T0EKj5
8hd0h4IwWO8Q5VoVCb9AEybWn8aoWe95iDR3Lh/KVaG1zzFmFeziD9fY6OjPb98Q8PeyAxK9O68K
Op8mVI2Bjy/8+tEszy9aeqKrqAVfiYZKuIb8qTab96bISjP0ATSGlo1gMw2nPXpHi2qOVoayhPL2
aIdYXaVoyrsHJ1gc2A6bF3WSVGp931hP7kISEhJYxV7AXPbEP6ApMWZT0MlqmxZP8PJLhtWG80dn
TRrkDFYVUsG+2Gftl7IpySODfACpdTskSfG4FkzISJ217o/AHAJ+KrVL5nfbhPoYuuT82sKPCo9m
sMyuYx/IAvQQKYQSxoSpEwQrCgbe130HSIMlZXG62LwlLivsspBMSpppdmXZG3Bf5vdm2+OYnRHd
vLv38Sz5zsPFa9ep+6glRZtCIUb5/E58zo8/OsH4VGFohhLiQT2wa9vcdS8Y2ShHC1rafJEiME73
QYTf81QlswzAEYW/AVybZ/+H/4h1MKZpDjXjXPi1WVJOM4y/1v8+NGM3MEmK+WEtSLZQgFRSWYMy
LeqkS5+RBjYKI7KzrfY64JmqkF9ATrIvXoKiLK6KhC55Ck/KeKnXI0V4II+v4qWIU5aK98TTC2r7
bU/COrUTySx3+VvU+ENDYGMJCs7CYxpOCTSrBd3cCV8zJLjYxdLIkJEDhBRnzSy5+hO/iif9beQi
+em7cz5EytChVjNSSgiSj/+TGOdSEYMmjoFv4dMQ0rCtPz26Jg8kULAdh42L/IBIMbA2dhKKuAZ1
tCUa6ugVLXrcO8jEvGTlLnmfY4JBsXJvUnMESYjNHBDsWY/5/GxlIc4LrCLylrLqQbGzjJOAZK6Z
DjVaPY00bm+v3O09nj3HyzzpMwjKn9Egir4Ttoj0yLgwN/izzrsJgXJYfu4tWesYMYn1d0KHlgHF
2ULtHo3lM9VZ7D78il4c1Kp6kr3+mO56tvjmskXtk9Qa7yvLR4RnI4sZOy/SyJw+YgIQL7QA7nVr
GdV8jBl4ma7vuu8F61Dumpv20Muye+0w87pjGoZEeiOn51ZzLSZL98DkfoKcPT8J5d6zhREOVZhd
ONkbUzAQy3sN4kY3vo8PVKfIJwqCv6+xnaM6xa2eP2pJz1d/PrGePymTNleEMtfGMzc3EfJlPd0L
GfuZDOUWy04qf0M0ApzfOcmXCZ9G0FareXXwPasYOZcTWlQemhJhWx4JxM9oW0ZSCOzXU1b5YImy
wwrtw4xBa+y2hTd/N+YLDbL93pAwNqyHyA1LFnQSLScmGMd0ajv8Hi1aymVdE48eQ7TDP2ZSOUGJ
eKeTzVD7Z9wHnErzG3zd0qKqrirJHKx4pcU4ikoERw2gviiXclYIePlH9xh+WS3KefTXtNYeTfLM
YK2ZRjBS8mKdIMHuRGo83Ze3pYneg5oIWxsXx31ePlQgdbYsIr54Ujtsjf+VsWpbnQspzbbNzj4o
giezv34IswE4iE4GKX67ySZPhKwkSBSPPEO5pknbS140EvZw0RPS3HoexHppFFL00FOqqxTykWHq
X84PCdgWtWx4SD7ufXtyE1B3HuY0EmbqV8CVeDNYpSyiqad/bUgpY7zAG4L8pMNo+1ZcqxpEyMdU
D9OhrDyfP2tMhsXYmlUyYzBAgHzQA4tjc/KW7KTUgj9IbPiIrRPnYI1CmalAg56IW14bc4nqXQlu
l+ksd5LPeM7WWKxGh/PP4ACChlFwv+YQUdOd5m10efzrWDx9VDO+CYVF++qmX8a1qmq2MKoGrbQ9
prZ8sU6u2VW/557tlvLfJNHvd8s25JaJI39f5LPg26j1dqNEDRgLH4JYYqi9iH7u3PffiL+yfWgC
63BMouJvs5LYFcs0aKFZ2trNH4CoGyIYh+1aYLdCvd1QLkD+cZpBjqtcZQsDFF8WCC+y7zStHya8
Usjimd/3QLvJ4500BUcMhcqfsNTVJO1TSRW6QGA58bcu6H7WjVH7eZcWhIOK8XZ2kkE2Xd3BW6Gj
PivklJXpodCQ7XLrHEwazwP2kt4exARAwCbk3+qK3f/BUl4KJTHVZJgmqlLBhVzhzOhkiQbD3G4E
yFlX4S8R62F1v3VskWj0VZQw1KrIH8oQn/o0vAt9mvKXlkUILii71lLEMxQtaC1lnXV8G580U+Fj
GIEloDJQkU2YSExKRELQM9emNMtttB0fxQYHT63462ue2Fdv4JLepXoONzJ1vRX9YbgJCivLbMkt
YLRvBW3O8H7i6nPWjFfmGyDYNPwVSe6ckC8f8hgYCr2R7mGJX3MsGTWSbN+9yXo33IVruclpm6Dv
W4tkUqgybM5rQGltJgZC3Pr8Wa5BPyK6XWFj0LotaD55/QeLUXUQf+X+6/NgIojfI8mvxyZJ6nU+
yQpyYXqzkdH6cHNwJIaK7VCloxJsKu45QaahSjaCkMZcKE5RH0ofCjTSRrZqM9oLZGmWOroEKnJz
TzkzX14C28kLYMlEcTB0zBnJjJnH7cchqdwYc0ZbclYZTuwjjPGsC1on7PYSw9WxE8VO34F7Ffi9
nCKeufZpKvN3pjC16j041vHELvKjwU7BFSt/UWZeg99hzPwswLbjMu+OcYcVZ/PDv2g5QsVhkrfK
tx+d7SRI+l1m0sq/+KShQWVS6/WytkNeCEW+N/u+iyXwse+RW0IE3NaT/qgs8fysO2nvHxYMR616
CLhNpy8l6owURYy5Whn4jdbbuDZmcs4CONokFkaXYg1mrk1us7ASpY1dgyX0cdpu+Chx/DGx3sy6
ikDF5h1+Kb/FFWwZEQzdFeRek4OWmI9m6vzwuubbXXMYHGu8L3mwauPdekwv6xP0B24jN8HM22Rh
cpTLJhXBvOzR3LTXYxp96IQGFT734WN3uaR7/skAUG+YknT8q8hfNOrP4Mp3LcoxkdyMIn7j+rPl
JbOIyabiQaB3uvZcaYAUgl5Nw58UzlIeA1SqIZ7zDZukZlFtqwGmzqlgVjkygUWQnQTUewrFOD4I
J69AAJjE41FDjQInH1nkV+rSFk2HvjJPwyH7cGSCBpz6xSZiFpQGrN109dPPWNHCWIHWTo/13XFg
jhAZmzH3e31RH4h2PJClCKFnPw3cVScm3Es+cWheSBBNW3wb2EQz4R0FfOcGr81s4ZxECJNbGuyS
lci5FKBvvQyu1v1ihvVDKcc7cP18Dxxy5AWNOvfHdLe4z5C5KcRQVFuR78EJ6VFEwB90ZI1zkYNZ
LT/EsUT/bMFIDxSKeQHO1+eMGdUlEy/cb0Dqxg6hX/Ej+F/MJXqr24nxjMAYU4mI2v7jfIoKJ5Mn
20zWljAFbYVAnKyRMsBZkGSoYxRTkFqHU7SHklp5XEwxLjlBTA55iy+azkPNdkiO32HSpyhXkHjV
ASA+H3uAQGg5Vr7zsaWJo//5E7bE+ZjzpGCW4KJg0u1qxUIXWF47c/JrWmy5b/LuQjBlNHnQmqEb
GBakyhDSmCXYTPcOaKEMEc1CdHykNqLsW+BU4ZLUotdRMUwrFBmI/ISArmlPXHfDFGsLdH9FOPML
kuWc7qq0rakGlxlNHxmhLeW51wkBnbg+0wsg+cwMTNT5jF1GuEpTAynmRcP6ssa7kKk6kUOq52/2
QB2fhUHdKxrgCQEMaJpGVyDSTyGxTZbJSEV6qeDX8SSkf3LJSdKTrUInq6sIOvtiNErQSclZpe+q
MkO52LjOUpMO3zPZZYDvsIjoBFM1jAxScBvZQTSPUmn+daf1FDikdSDD3t2+Qf0urSakkCs/B5Sz
pJuGAByGC+QCOsprxycBNMv1Xc6QUbxc3SQDeDXR9rxVznp43ytE9sOEGn5Aocscs3Aib1HxeXR2
IHhqmSOwTl4SLRaNjIuqdUVlN5DNNJZQ9/yIQOtzvh/yqpO8yk/WTFtjWapN5rQbDOcyLltebg8K
j0p/cKDYSW8Bw25KYCeBdTTS44qurtP53xrxPami4lFzQ04eVQGyGy/wh/t0lwKPUD12Hdxm20F8
5haU/cycQMjdPp2hcltQ1sgWbtIonoTmr3x3nIiNHD5/CEDBbx+rRJ7qvCd/EzgKWTBYraSzkxYh
X+h0Yvog3zdTnCv83wwUwXzJFaGNf4w18Og+shs3AAW+0wMRbhEnfb7w1iPF3wdTHzkEGsKkaCGd
Cc+wBVMgK8AP0dGPzcvM0thJ2Eu4RcF5OggKAVJBL8l4D7QjOfGgUTbycvAuN5I8xVaw+HKmfmfY
gWh2K6sZa0xfZBweLIwOLKeog6mPc2XPBL8OjgXy/Rkw9ecW9IP9kEtG9+62R6IhHcP0Fq5maShI
ndUVSFaxdvLnG+0MQnAbSEesdzxrOu3Xp1bOSoTbb0MNmugaDZBwmYiWUaNoJQMdo4uOKMA4SZbI
5ti13szqhrJYMPSOlaX59QnkA2w0Xda4TuJ/yKp5C+YxFIgqraENwSmGVId4/gfROmlOictQHmyW
JV/vF+jdlatKMH+wB0qVsg9Gft4AATIwEQgtU+rxBvhyJ085Jgo/BBgPaPrZPVhf3O6A/JGeigBo
Dq/7KHaRNlv5ITl0uL1CF1csMtxcrJb9R22Eml38bOV5sSstThXg55qzbQyfNpsGvkUhv0BnhFh/
/PhiAQsoyIrhG+rBxGEXqAwvchxdQBWttB+IEgzOR27AYx9pdEZE4OKmaib/vWIgP0UFjMwplFCc
PSGaTfZVdsJIMH9wIa0SjuhKqFKRFu+Za3Z6GPHrCGM4OWQmbU/reCoMeeinuUHwM2YJnwN683pv
1AARJ9rmKyFAtePAPxc/iKlZV4Ltt3TUtHnAdR4BOK4RpSV3OhBRPO3UNYBeAXuU4KaNUIhJDixs
x2QjeNukJpZOPGofPVdfuHewMpXDrFX937biP6jIMyUU/qpu86tl3aMcUVSTrZx1melzupX5n1UI
iILtpw9R9ALUeyNYb/h5l5YQd5LPuWbF4wWloG80FV3DN4qsulr21R5dq8KDSijmCFxd5fSOvPwi
uAiqfo77Vo66K0J1Z9OJCFhMmEGZcXcQAlVRx7ERBQkMI0EZnszUUtUWEMnyIbe6VIKSphM9PlNq
+bZwj3aM+wnFmDFI8WMkycN8+sK+eApoRYr7/4tOugpqGUBlJxuBCwEdFdDUbAkD6xcs+iJacR3p
qIrI4/yq2Jzyd/Xct+7Nz8hqucnGZAV8LxXnBvPdo72wVCbH0kW1bbKZV5ED60ZUEoiFtPGBu3AR
U05CLSyzz7fQNwwNrkW2mgIO3r7I1j8sclFL9yRThfWs3yHGZE4gv+uHC6JWuDb/UWqto6bKBqUs
0f8cDoasvQ3YLhYDCt6no0ykWwdmsx/O0r1c+1bkqrSoYO49SSBgekD/r3EhJD10WB44JsFUym9P
gU/2/iOLCmbgvktgCuYFVBu6CBAcM2nv22XDI8bhCk+NOwbBziIyZU+v8iv56uvL0PwMNTCoW0iX
mf+W6LrPXWfBGsEnJ8mu4bXHBwhd5r0fEuWsHaCrOFPPWU9/QZos0fNpYKgfCLm9w7EZBypfSiXa
0LqyddBnLjZ2Vjr4+CVsN59XCvy3RIFh2yXiVOUMYZ9hrDsUrpTiL0p/G/s6WPBrfzvW1ReF1Ij4
C0vp9cdSWWLWQd9fhe/eKVVc3fx6hHSnaO7ksDI5Nuop8TgUYcwVtJOg82cmonFol2kxfIpbzm63
YPj932s2GvkkDSLWr2rOMhxIDyzp9VdQt3lDVUmAulb4f901WnBKsKwU6tYYp4kgsDlUeHcEQpoZ
7Uv1gPJ20ajNHlxGycJ4Oxe2mmDmtGaN7G1Iy8KqFdnMkuPq74f7i57CsLG1DvOtw5OR1NkXp5qy
zxZuDMckdr5P7RMigTAsiMS/LWb/3pnUlNQbAOqlCVmiMCPjjTcyRm/zVHPCh4Q987U3wK9rt2Rx
72YvrBetX62yudT5jABXJmmS0uGTEw06HVwCtdfrHdANRHOO1VQSdqjpCQgZj8bFOTs9BVAC74do
+ZT5GO7FrOVmwDWFxTi5KnUh2lZwu6ppmc31v3VkkzwGCRl8nO6RjlQKnnN5ofrT/4NrN/ButPmT
T18j2InyBXvou0odeirMApU+hWaKz91uIBHKBhVg6Gqa39ZXFTRB+Jl8cA64pzTF85YzHwr5lKTc
WcCfD1HkS8wrHnV2kUxNMqVoHO3p3+xa+TKwJVHzfbs1ccdezSU3XgDd/GSJ8oQQqyqvSmnEM2UZ
3+IQCFSoq0GFEqHJxhDVtQImP97Tec2HLXeaoDyIaqKsUpD4K5XnZvVAiU6YIluNTyAW/9Yok/W1
ayDD0c84a8HpX3YSNlzbMD/uTCKmURcYDTG8rKKMu3hdbjGYhPGeQ52QD0Fyoj7FjqI8M/mwYKJV
VhAQDnWKQ1V1db4UVtjzgkVyEkVsumFkftrSGsREvBatp5v8pG/q/zLAtyFGaLokAI+jCu8rjQ0t
sQ3DskQJg0gm6nOj2Mc+VwuLC9wIMgjhCgpPGGaEwAWbejjozhtH//L8OLlwppC7ISsCadqFgkzl
aq1VMCnCeN/U7pytZU76GH/KFXvCzhHAqwWM90vSo1GTdl5mvgG7gQBfMrovHbLMHD/lnI88lc8R
7nUnopt+PYxlYTSNmXBCVnTVlCjWYnMHDAKIu/pVJ6JaLtBuoKm0w9Doap2mN8Jbi3EeXXzPkhhL
KAG14DDqrbTIXR/fU1W1Uz8B0ndzro/cTNkjagWiTwDaJF5khtDvfeGGTLIsARdqPSAs4ynxVU+A
Y+CwG+7pbIGl7JjH9NCV7Y9nFRlikUS7OGvvhc724rML/Cihbl3MLUuUAFty2Rw/GFm3SxdcNAn9
HECEwsTJsl+Qx9RvGIWDxwcKM+R4by/B5M6LpgUel5nPgyZ4C1o+OdVEXWdBk+79bzHmndsu2j22
fImDEY/FKmYmiu4Tp7aQsM16av6QUzj6h+RNYb837u7eCQLEJ6WysdRWTExIcual3lFQIEMlhpbj
7w4QFrbUOfrPlmBSgKPzADkfuWI+kbnGnFbsFBZjLTl5o9nuhOAoq7ZFC0hAR0Hy9UsIMqAxWYG1
+czx3M608k2tVKVomUAu2RgBEZABJ5iUebsKrQMr0xhU1QcuHlIbItJ4LpBzHC5fWmGvZa96JnGL
H8XM0+mmZR7jcH8gLKAMNxA3XK/0Cd30rHeY32NlDBr8B2qpa+883ORvfs1rrtv6dOJ2hYl2RVca
ZGdi/kgpVLz7+Ppr/DX4aFPS/oXXAYMBKtVN+X0GWO03fgDrzqL2AUSqQi9hUpqG17WsTfF84UTl
S44e8RY8EPiDOiDTmde/39ntcabPTYWdQC6EgElI4qu2Z0oxbfu6osDQckAzBpvsYONrM8492N3T
NMw5BTDGpcMgVUqEZOYGM/hAcoaH8NFLtfPLniq+V0oyDnWiaHxZaYhj2iHd2ubEuDsKT8kBY4jw
1ntb/sf5Xg8K6kj03JTNZeCwL7hnjzvlRK+f3MYqEbHKtt3RZQB8+XptD2Gm/XskYBOkD7fUQlqq
+ggz0GeeO5u3nlqV0DTcS8/zw/TC5InoE6DTWdIrAbukFo4apMPmX25Qz9N5zJ7ZKVexNJnRUs3g
L/GxU2Y7rj58OZY3CUqJ0meU1E5SmbW4OLGwLUAOD6D5UVdfq40zrMLMUE7qULXqlZMpq+cif9ow
Kf9CIVpV/0hA2q8l2ikKFe17OaN/wLiVFDH/5jtPO//ZusZAgRVqi0k/n7ZznmzzLjMWH4zpWmoq
e/43fY9vv5MOGSJjsESb6TNXT/b8gIDDJaNbQqY8m++MUGYtTsVKmB3ObO8EBpJJ8OEf4QhZTPpt
jxsCJr8r0XSl57JW2dZROkrdEbsc9Svo8DNoZNcRyKYf52JqWd+1kiFlICohFYG6MhKwVXshzngo
Apxk9/ET+tVEIRSqgDBjXh+xMSuIWg+HWQLM/QZuzzT48z0fSrClvq4TdCxaAwuloadSnQUrg7SI
Jou8PqTMmkJ67WZAPVvVso2eNgMER1HpeqvMwwcf6MjHaXTQClg8KyZnYHb+i4o4Q8A0SEPwfBEf
joZEUc8/0Tp0Jt46ouZp8eH36XiU1ydi/IOZV14jt5bfuSSfbP63gTcEI7L2VjJxg3tt7adUt44C
cuJRk26upEw/hFmIskTAUNjkaPOvr7mOAPXkQ1JYwKGXqYQyDR9/L3p2Mu5+pMrl/VNLeCEB4q31
d5Nd12ArRf3vsKA1qo6bJn5+VV8t4WwBPGGI4+ER/gVUoZOAcZUgXvrj1tVsMll3tYvIyuyU0faq
Ka56BOU07lWurmZVnGv4OOS83d95q8wFTzxT4Sgyi+vDGbHCYwVx84UOES8VO6ABYEs9y9s6UtO9
HRHBKqSfJH5l0AbCQjrGxu+E8zZhOv3HkdW0000q1pD4BbVladOz93PHMRJDlw7FP+at2fsSEHNV
2stnH5p+fnPAeKATOjbIKRuha2BOlh9uq5nypkAoVySjSREX8JHiOhjJGatLiLl/47Fb6XcB3GfE
TIxy5rA7T1TmjZKHfGu1auiIe4ZIp+QwfxkvqRnHHHPo/T3Qao6h90oVjq4uxz+Vc8UM8NjY8nWP
rqayWIv/pHjCcz/dVUjf6nkJvKE7dZE5Yi7mYorhQg3k/Ws3aK6m7w75/fdwQVWh8sT3zgoXvSaE
L5XGo5ROJSwz+/7oK2PImzfaDAtFYZexoynTwAb+8bq5OkvURKzNj5IyGhWqSe//1UfwEaFvOzY2
o7VsgUbL/y4Na4vyQ8EFd5sSptE/WG2M4i6LHhVUc8aGt3OVJ1uChwGIB8Y58XkN7EsUBUGrzjKG
3FqyKN1EWYEWC01YiVRJS/cch+tPrEb7u9XNNMwtEhzC36nIl357zRtTBvAfdVYN9nHTHWcwRRMF
jvyYAwtYR+wKW+Ta6Edm5zVbootKR9275kEEq17iuXP3SCIeck6A/8sCUnliS1a1OQ8DoahEMDBk
fFgFzOhumSYsxOQeA7OZZTGBlyK7joz4N2W67dEvb016AqovILXeePl3mgiUcdpxY2a9hcj3K1hm
u3EHZx0xb+8ACSXYlpZ0o7nLS0/uN01OrYNKau9oKyB5vMmML054Zo1biRPkI9JGYqxn91/APcAs
Y+KnoZ5aAnop59fQMTflk6AbA/rQZ/GL5UOKu/oa0qcR9gH+Wnn29KrvxQJ/3bCaRT5vq9spKB3A
Aa42mNs0yS34xZb6oVMp0b6Rml/Ue5T1xU1GFmSOgnaXnMlZ7VLOTSLEj0TfmbQFGMwJX10soU2R
3tG6CcpeDFYivEiffzGBEuioAlszxkV0SwFaf5D3YrHionG8kxQCpRRwXsaQggsdQ4Wt3caO048I
UZvAHIFNh8118ECxrNYxqV4Q1ugFh0exVgLvLg8RYd7/lNrSYHGaEnvRffwZmu6mgVu7VQwnooBZ
butiILU1EpsajSuBSyJGnH4FRYlM6UOdKDshOIhypsrJEpHAwQWAOygRxiDtPq43Z1YQSPyXwnb+
pNgEG+WND0yDV+0aaHUHt0651CyRH71F4/hqepcRmtGhR1UvPo3BqTeKnYeuFCqatsXR0oUT53oP
qW09cpHU2VBhuviSFIBAVwe4IOlNV7JlQamw0deddu28utB2bQl0EYkXmZvE0xneCBhiboEmOE0c
fjy5zvi46PX2PUBfirO81+MmVTI1pKo5BdsdlcCzUcMzWoEBP3FK+ImKRPOp+Rw6wJAs6w+qK4mE
C7Ag4buMWonypzpUXGbWwmTR/hT3Iupv/CRN05HaN4Gp+mwuty2zPl69EzxYmNUvSAyz6IvksKfj
HoNHx3oZpcSxxLdoZUa6MungZM1Ep9RQPBk9oC4vuYQ8gEM8io7YqJW0dIkmDFLxPf2Um3CcaCeD
TcgpbK1E2kZ4/xSI+AdSlopowBS2KoGj2ryQnuWSeGWg01x38wLxDKIW/Xpq8KNN4NWYQDj9U3z3
BWA1rzmyTEh68FuwvjosuTBmIYdDnmjODI9bUcj75oUnhs+0Ybyr3SN2U1+DHFmj7b1HSnWGvJId
9QhixYqxJceO0yUk9FP/Xklfy4iAaPKUqIb3/U97tOL/EpAvqfoT7OhMy7o/gh6plbgCOxih5VqE
dt92cz+ogo2S62NW+HoRVvQLBDocXt4Bd79rlJEBqJSV0949NA7LHeScgFAljxOIM2Yd+3JYVW7w
qBAaQDUkwDSVNuxcLPhAEpb2DYdMpoWkU9gHNljknefamXQXMjnVtSX6UAVFrE1m9rMeegNu1pmM
X9O8mvWTpGEKHNnuDJnpmrXuhLRwAngjIDBAMOGNkpV0dwKyENxP4BGVUHa5X2BTvdzT5CyEE7OE
RHyL+EIESVgPpOnvnxh0DhH5aXVFO4bMqW3hZ+N/IHf10ulldDnVQ9DV/VFBF9BGfuwqMiTV1dS9
SspQo3PxszvhpnHX9er4C3bscbuNfATLh50qlisc8FZgWUJ41yqPyrR9C438ZYKr9lpGaezPBVMN
yNM1Pk6pUULlNpkqBLAGI6+K5DBzTK/bbqNMQsBdTW89i1ZwetAztt4ekvCkcYFU6HFPFBuOo+xM
RbGZsbcWEweh2UwyEgck9FGfeJtAWkyWs7iDNxkGo8rAIJab5jtQWq9o0uaKVSXJ9g61X8dDETFl
zsgGqvhcwNdEII7i46GsZ9dFsJz328x7YyW3Z4xMnm1CMY6LmMDJEsYi7NwVLdEGgcLa0r6cq8jr
3/CShl3i6Tss61nJA2SN8xbW8h9OyLwTzPjHsx+8RKcP/kDDubwHMF9rytQ1UeAARJat7ryFo1Yg
9LJ24Rc0D5ViCpeb3LeCzIe/UKGKoKjGr+VnLWEr+yvLoxpdZYkxooxGjMX7Aw/O1QvMMr7Yq0R8
TLGsoPJ+ZTWNN642uHLaeSYsDIrVW9WIYpObzfKJxlB2XtpOU5kJUoQFn/Cq38lKWrdL00B8mOcx
g5AOPPisW7yIOtyASSvVyjd/s2g6J9CXyb5PcSXEWwqUMLUtqY2L6Wa2rxDlwwBhF8RP3UC8evT1
zsvCegkQOgKiKwaNeDiRr+zNIzD18cF5e0q7Dgb0iF3kD5TTXczIDxCM9EGVMmUKGc58cY5+fYUl
gEROw4YkBxT5XQkpMZ0FsYx0S6F3JmAWcH6viOle1pKi9mg6ssaR1KUv3OxKcL89YOfJsKVy8C26
sC0JMb1R8jHzDpaD0/inSXZ6YAzxIYRg2TtisQHvtZDnYmnYgOPefzikycqQWKdjOjvM5tlUkSXr
iagGfv9W+c/JsfV4jQIgKyBqq+JKVFbYmFkYHoyDuPIDist0iFRXEdSvbUpzD5gajk7klEIqPOUE
4fHjnxpTq22zq/BFSSwFFkmH1PtBc9stqYP/uzn2wWZfp1xGErwDTmj+4RTRAvsoEmnjsyzDU0AP
kHwpRtk7YbajYJUDOeFUxxX/EkV4saOPrx/oV7lpLNb4B00ZwpswDqE7HYMJcYAbtWGB0Ecer7UC
sbDhb7TPZmOXTANICVwDo7LCRPDRXOVdQ5gIKgBpPk4Xf+QEMz6aC+R07mAJcYa0dmVX3N5RNKQb
Trf+inD/JFx+HInStecG2OhzsyQtZOr+PTI6HSCpG51p87/5EYj3yISTBzgk2YYYVvUeza+4jXdW
DGhJYFSfFQMCL4A8CMO4oQNE6ruq9I3Ir10kPx884PtBiEN1+nrIlGfrHbDBghXsZi2hsVtLaqR8
rsxCngoDmpI5ap4YnVJf4AteRppuVTjvYkc/BusTiI6yQBa5JGA/5u+tOuW8niZIRQVhE7/gMRhV
EkNr2SmkVpqkVsiP3RBRhV+MnABb6+0o0dA3i4frEa/9opm0Ol9ZD2DJD7ENbEfzPmXxD5uOj5of
Sq2Tw3YYKGmSsEWqRvQcFZz51MRfPDf5zWFMeNRwZ8tAhD82ZOT8XUXuBKpBM3DZHO9rUJkqzsN2
owNjV3m/RSDarbW3QUZAoKOhp14ouLEggyzdNOesXBGbjPf93trbDeFcV48jgT+r5dur7Qb3EgJt
64A6kPZYU/Or+or5XZfSZexRdVtJJjGJKs6kRDLtHCEzEQPRCJi7Fz6Y+XhspzBPbPjATjHa6+5S
9WZsMml+d4vA7CrO6I1OrCDLZxnzAJZsSWg90CPouY+PxOZh+B5WCpyh3wMGfZkR1LRyU5irMOCa
WHr7Owl1pLj2KFPO5f6EG/0dShIpRW/+nvZsoc5CHXoyk1SvbDq7jm8ntPEvuhC7I4vBoMkVUXu9
ysxnuHXBSFkss3YyuUIj5Qh1jOEp4WZiE/7k/XptBjW4bgSBtgh3bdy6Y9tMygK6MhxwwN9S3/Pg
BWBJnAG5hH0Erhd1xO7DlI4dmF3UgYV3IGMgwlEmtS+0hbwyzOOaxcckXB58loDzDi6JYG+6G8T0
Pm8u70MGYD7X9kN0d7OYfXmOZ2ve6ByW1tNY15/tDr6l1+ajuCNrMip2bYJqxmdM8Hw+AYdtaeKL
0UKjfzSGwUo/XAfzM18oMnWKHgpbC6iypbhcnJW/K0zfz6aIBbAielBG84NWEMPhF+FxxVesVBvL
q2gM+X9c1/lEWsOefe3YLWsjDbGaTNuIostkSXhpcg/ECDA5XOnfAFDRatpKuSeAoz2QiUE0/nfG
xRN5RyECG4KTxbGZXLP5/hjkj9mI87CahxT2YqalDg3I3J2zi471W5jCeJ4oZyvsD3jPYgtvzMbK
rWyByDWEuB+QqL1I38lnTjzU1JI9UYbJib+lUNSvdChDI6k5Fy2nyVlXS4A+zLhp8OnB/5WeJH8j
ZgGe8JeGXU2Ti2ZzTJMffLoHNjXDN4IF6Xlp2nC8PZQ/YJF7EL1GXRhmBC2/J7UwkWGEHJpf8pzW
bNAqT7IVZzBZDzvjiip9+8nX8sbJGjCv1DRMrXzQuUGCmR/2Hy6n7Li1U1EJdUi36Qy3Okkc/bvv
mvw1bG+b7hWnh3GrZQ7daeNq4Bucj9RE8gKgkOx9duK6MggRx0A/OKPzHejPojPb+M57z6J5pemu
2NZ/0RK5iZEj5vp3pzlE7b1PHqHpZPt744jy8nu3AzhIfgp11lnm6poI1fSm3gShGwg9+JnZTuQx
YEBbgYx2N3s9Vy3SQvotu69N6zFkKhFPkTgBXL2XnMREBB4lbF1skOZftGs+kPqdP8vZ51q80tcY
eS2zF5gLrAM8Gc9Xd5WdlhkB4PGlv1I/NOjdWOhbIcc4sMwxkkp22NqoHt7FYc09Hya7EEJItpMH
VI3NS0Vhm8a8/L0BGoRxGJW8Wn6NhmpoIZvOm1fyQTP1YCr97AgXrE2/p1oKwtWpLsyWT0286jh5
vYxQsrfrxzc1tbjpxLsgVvK9A211cXSG0rvjxyrG6C1fM4AqEVABQeaGjkpsBbl0+tkDjdMh7rGv
MH2PAR4HZInDq0MpvlBP7v0XdNP7ye64HvrVqsO/ngRgkPDhFlSoVw1wSSoX+bvgHIUyGo22wjfa
WO8etAuApLXFF8cd6JEc+MgpmxmrejGnT2M6tLT4r4PLoO4X2svXbi4cqIStU7rkVxtxLr8B2uf5
DnY3RZ1XmVyEWMl7DI6Zg9G6qfhd/veROq2jOcEpCJOPXvvnIsa+fp25oCRxY9tEvtZPPmnJX76i
K9CZAZ/HDbvpRd10Uiel4g11cWDouTUCEGI0JV2/gdJwHmalwMfiBUpvyMUwOay30X4f1oNemw3m
W6vHK8A/MiI33z/OXLKwxCbzp048QoWX/eZwGfJ6lWfcVuELe0GbZbFUSe4bNe6B/0xCnTR0vEeI
RGPzAZOpse5VFIgcb4JtBNeHXLEKZkEeqJrY8IxGh86TPD15DeY1ulqPCoIaZCIrR+uuFWjvzkqA
HCaaR8HMGLlhF07EnNwDXyT6/L5Zo93YHOLKyvvu3cGTpRvDbxMLjwtpPcOVywOPq6oAPoyDaPZM
56q5Nowaxlj2Pdb08+2K38VqrHnv7prDnvqovYvF4eXTjZl8xkVDBL1Hztg6/TzmaGrhdGjuPWF6
DaPU2Q/3hBZrWNvAd6rXekKBa3l+UteFzEf/r6cxOe91lNPrMGb4gDEGSMY0WrsNb5y9CqSXiP3u
buiOaf0ZK8cIJfTosKZR1TNTZ0gQdv17x75OYRdy6G26db5fKzBq3QkUmhlJKmVQyGKsOy3lTLTQ
nht3qxT5nFGt+0NDzKYEl2MCHjxc3gOJ/fTtoBFkHOBZ24FQ1QTvWhRmLZ+DJRxx8HGC9mhFQGPN
tZCOnJ46PvQzUaQAQ2ZLzE8wZiw//8qVNz+BcKLR9xMwlnebJ0aucHW5Ayo7j7063lBukZGBbv68
K/zS4TMHCWBz/Y//TlRunEQA5cpbhv9s6/PGWT7rPZEIb/dhg8QyW83+m5q6ASu1ojoen5+Sip2Q
VaGucG2uXXZrCjjwbpN7Hu72TqznYOBJ+pBpNLxoAHszsbLJkzEvJigu1fKHe23B95HF3884+uso
lTGapBwlQASC0nw3OAQ5Jhz+AgvXmeYeC2wtzdAr4QsEzcYaasAv6GgnuliQAmqXHqwFdG072ijI
ZvWV66jwFyL49TLstx4++FgROsSa5RwC05aZVOHAMR+2b2Qr6WhQ+I+1Ms1HBEvVICxsuin8I+Km
Qu5ThwidBDKBaGmraTscT9KLA1yFbBgibQ81t6Yvlbv5GoaSkXfjdkvn0wiSeaXk86AuS0gnOnHT
+PzV6LqlImZPpb8/CjHpC4tqbMivOgILAoY8xyFJS9IuoVs0nG8YU5TcN42MNwGU864q1U4PcXDx
eLzMXatXb8F47oqncxSGeOjRtpl4af/7n2rIyavZhAbI+mDzYMDaxPFaiJoCcSLiXUBNQKVJOv+j
dwpPnzauVPkeCi33fmwnYoJHpzcb+QOwXO+7+jVfajZ9ts+v4JpcVxBR5bXDoKaIfuEWXYExSEAt
svHzQuaPhXT99hN4pccjXllvKWtsL1aSmUeXyIGKB/iFhFCHm0S4vCsRHYxFCQCf1+3VdB9Sk369
10NB9eoef/MtBfTmAo9wFUUI3oSGw/C0A1PajshUuubo7P8G5DFhSllLS+gj3G4lGrWeuVHwFAoz
CRouDNNjwuAz458P2oAqkhVVun4zNKO9KwWJPkkFvtgBAKJLmk3KM4cdPReWjYXZNIcZRmytMsSQ
31+2EVreSsDmUMnr9L4ff3o8+Ax8V52e6up1p9GFc9fUY8nsaIIudlRAXF4khy4h1Vy/1FjB5tYt
Iy2HZkK3v9LR9+l2qg6F1zzB8PZt1rQtYpJDR1g7gt1RkUp0dKrD6xl42NkCtQFsmXEQlO9YLQzx
LYI5qDq6kIQfmuVud1cWMAUKAu5dVwH1yo5kuI/Wihuz/dEtDyJTcMwI5fXIBd+A6mmgjDhJe7zw
YZbg7+DHlPsGCOcZTVAEcdNZNtjUEvxKprQUY7+z3uSMO4kH55yl6GIpjg1oQIf9uLlnMUp/x39X
VQigDi4bKdJNNIa+Hd60kYycYFt0hinaOD9s8OIDL45+4s1wQ1EyT9CpT6vVKESVaqmolRUirfh+
xnad1+Md8hVH1OFB5Q7kQA5XC1ytLCN39apNZE5+VKAZk2snFxm/B2JCpAux2fN1pHKnhE16sqF9
cpl+EYu3iw9fDSnlWKBCCGchtETKnSA6GktpthHr3e7MFi9vdbmvdv92D8PAi68uXFpx6M0HzNpf
stKpyyLCh6ktBEt4f1cMK0zoXGSNZM2tWf24WY/jivAtVF9Gl+OJLwEbIZFyBXTjKGD+ooNi+CNj
/370ZzzcD/T38DvT9vS10EzXLccAk4xZrfBHDMQQ3ekrkS6kQHHJjD9IjceWOw//brLoy7wxtcQs
6ky7JHUxwo1Ryy413KQl1ggFwzpFE5pVIkV5si/gQmqr3sef9lRkmUgL4Dx1+JxqlHzs9jZ1C55p
Dbg26ODB9Nrw7aO1KeyAOu50Ly71RLvPSsVCPTqS04Ce3oUldi1p6C+MFC1JxxZ2utz3WiF/exsx
4XaGTvbPpgXPtOKFtIuUElAKaLZlTeNZfYfijTu3YXynw8nAIElT8NclT5q2TLYnV/gpOXhOAEFJ
SWIsElmLh6qpti9E4+lGewI0dHrIwmLm6OVOdRht9RuJz5XMvsVV7aWdAomsjHEESXpOYeFsr6h9
2bWbBcNC989pzEMwR/gne9jePbVkfW0ivNUchmfhYSG8woZrGh6Zoqa+BO6eq4EsVI0sI85ccdI5
D1zoH/VNNaxhHb27ePfrg2PJiKZ8yTZVmh6Tb2FBxFP6WyxigPfNC6zHK7DznkPNpEHQthtMiPuJ
zb0Ea1/Z15ygZc1gDGmIX/DIhP9KIuunyHogOG+rM2Nmh9N4+b1nCsTexaO6TPZKV/SPFusRWshf
SSGCDyAW2G/rdKNw8krZdsPh9zzcuaYPCPdlU1bK62UViM2QwRgt0pfZKb3208uXKIHBr6o4ZqiO
3PPFdt8ntkN/2MS0PhhJwb9mRjmyI7CzRtgvx6j3LO2O03a5XscVY4AFZKIl+FJCwthYQMGSfL62
Qa2uKD2pCvfRmQZuyjTpe9fBDnOKCPyS8xswa1cEGvzPXv4u8jRCdnhzGOHFnmz6aQ5BJgaOF0Ic
2r/IzobY2eIC/agpecnXKPS08gZUtsflFBbgWTHGhy3ALMXUQcivqfNTMnggb7B3hNphwjZePqlf
I1kk5XE75hPap1fphkuooTf6qdzjf5Tb4jfsKHu67X9FkYzANKSSaSLVMR8Ew/TC5hR5Zn5V2tfG
Cv1AYqKuQKm0ryw0yOsG1o9BtSlH9i994vvkVmWojIIYvwQ5/xpISYnufBvvFM0+8MVQr4rt2Zgt
aykRg/SNODcYTG9XeAz5d+zz+VEMubSLM9hS4eT4NtCQGmHCw5Vna7fG02Y+VRjRLiLpSwvZJ+5O
azmYRZdy+lyffE5P+oYPLDSbqsFJ1emTTK7LtANiil9XdVOfWHrt9+CDwUtr6Pgywv+SHHLdupBk
Q4phDcZ+i7ekqfDNmnHKOLU5faojrg3txnbQuT9hg2Fl5PMMLLjTBgUX7oIv6LXkN0d1+rh15avK
WZXWdutp9wu3mvsOpghAJYOWYzq/YLHzHoTBKnzEymDmuf48oEG5hEvkk4SDnKUaiCDvYH5vUr8g
KIr1JrpmYygc5tEzlvywTkY8CcVAg3n6EaVmbHyaprdN+QEML72jHd9s9YH0mn6+/bE3JCIdjKS2
o5YpUTKeLkZx2hxLWQkKLPZDlGSR1CzWjaaAvw7w732Eji97X+Cb3ov+9Xt5RFperOa0R3r7jV7q
224ctpSm5oTpgQ/k8VBD1QLj2MpYYQTJsVlxLnrM7ArSNfhRgWfyXN2GqaCrKAV0qj90sInp1SLf
29KyIUJ2J4XTzKZE58D9DxqOsz3mGzVXk0AuYRIZa40Y/GEBD7HCQAJaIjrxS+Wbxo2ZoGPv3rc3
SLBusBD4m3IYH2TRO1j/5lqVWZfL8MlNyps4QVNPaN/pk4XmCfePcqwzmSXbJE/PyICoRLvCdF92
DSyafxovrQOJ1sAC4MLZSR/t4HveCDyYmiRoQEucuboE6gJkrzf7gw+VFQuKvQ36uvRUX6j4WS2b
m2fZ+mYxkpxia2A8/DfJ/Yk+EPXvN2OV8BpTZnG4PyxbcUUoaErqO6nWqu6UA92xlLxjaKOtp+Kx
9fcIeeFyhTnFcSAmzFMVkR/nTVbOgQbx6Xh7xXz6kmZyDLxRvjuv5uK5dLM0QAxgtkm1Xgf4zTm7
TYwq6kcdntFcOpy0zrCw1JLqXYpKiySgULWqzp8HvT7ta92oKkcfyAi+BZyuU1ppYM6owWUys5KR
9auZQy7kttMp9qmIoHWbv42jdXBytUraGjXtzede1b4A4kza8gnXAfsnbOkfXiRDKpsWc2WORH0r
H91eougLvWEtGBad4ZGESxDINKFMekTZKQMtltR4NdhgaAoYnvM/TApRTz6VsYqOgHuLW4R9cZc6
/MU1m9KqIw6XK/m7rf9d8b2XOkPLVjj03fa0dufoaG74FLG+UjYyUr2ylQN4EVjLMpJ5X8K5uDLP
4lUWV/GBcI0lyO6+V8+n+lv/Y3dH8PmJ5TLbvWWTRZQqCM0IUo9Tf3jm9/Po2M/JDKDRbqTvdY47
hjZ+WSgLemvtV24pIJ8E1RucwYGkWC+VEZw+P2yUMwQG1oqQvD3+pRefKW+8MmoUu73JQxIQNuKC
ivLq6s3tKxlIuSsjwIGTkZLEDYdU4j4KEGJeTiUr5DGkPtCNNtPijY26dAavZqYdMhvDXt0L+Sff
TrISdriU+7iAr11bWpiY1/dAd6J1VAvuAlcP4qgY2MLBzetCEtltbtWDqs/patSmvSPEgzgC33mv
k0B8mq6EF5hdr2t9Sb7Q8Xo/cjsVnOsvUJYle68kQR8aut4mYMQbyBp8DGssLKeYPQ1sABmzhrZ/
fEGnc5W6e0UQ9J4JAQE4lBHj+3RRZH1A/w+ZE6Sj0WAFb0v7BnBIVwWBrAaYql3k0cS0yff8DOZh
vxI3ubKbeeUAkUoASiOGLXflXerWh0GKAVpa72OhAsOo5bsRkpGuMrF/j9yW0wWGySQxDo4JdWxy
wUTIHG/AhgtcEKMhMSbnL8QJ/11tzI625E6DPyE+0McgdukQwsPJgwDzT07Qq573yvz36kHt08BZ
A4Mf3mYXDoLhiL+lkrrryIJOUzRD2DzGWTNM7LkbGejcysqf8/IVRy/UTW0puD7dd6M7i1lokj4/
gVybpMvAogyRPsX/lD4Efn+nOh5u2qsecnG0m19SSx5wCFcH7ViYAIFq4g7Ej4/j7cw+BTm0OrWP
WfqMDuhliNjYmHRjWeUDuCbBwu7346QJCFrtfGZPkqPLYigWvMK6J2uw8cc4uIIVcHDRQW351txo
NR/Z44KHRj2vxKurqbUlbX17gxvxg5WO/CjG/fx/PcnfV8h3dyia8MW/C6ewDMSrEMK4ZUGmFQRo
LsD2Hujm+W5mY4FL1ULPE0CizVFZb8ri+6Frz9yfw8TK5VSgn0nOHrQxk7Mr6kS/5PC4SxqSWNCi
CNNeW3Sr1alXdI3sSjNFSPPCFA1w+u7fenGAUvU0Orw+ToeympnPEw0kWuo4KUv1HihPK8PApeYa
gVX2IWsBXs5EDopn4iO0Q5t3kv/yrVV4UgOvBQ5hxkBh+ZdG0t/4WAMlDIszykt7pozGO7x+JI89
/0UacMEyCceCQPH//5n2YYZwnED8IKhumwwSIWUOGdnLnofYtYxNslztVgV0Nb8ZSAovftXjG5wa
NmGtJ/Nh6JVhHO1lpuHBSRMvaB4pLuGkvmh0VJDc9vUnl+sgN1vwQHjOnEil17lammASdg60p3o1
0KrGwvWUugqLkYgFt6CtGnVXAWNJvdapwXuifpPcNp0TSCtnQuDCMxme9ie124Wl2hjSUhlJ+fGs
y4hROxbUqIVDKm+CZhSixConK3lKXEliCHg4YSdmcvBnHOywb/coBAx4R8U8qlxF1vjx/31NCOAI
6mEJYC/S9E34ual9avAzZ7/XqEj4sbX8Q8e9vhvSMBQIQKYfvXbzw4h7mw3Xf1OHaeZcl0CSYv1r
vgBwrdaOkuIR8CzbvObT4teelZSWwgmxw1P9ZtqF3LL5fzrESycqm6AzVm85RhOazFpTc2yGDTkO
Ql+WnnwfumgqJamPVU/L1NTfuLGXSD8Adxa9bDiDCTH3jBerpZCjvkem7H9e/OL/Nrd7sjPd8wv3
VaR8c/jHaUjiMMsi/UBRfXpY/fBEzL+KvrwmZfVYszNyomTUbFQD9Xul5OXG/dPajU0MyZkyTYyN
ZF/6jy4RzrdyTaQTx2gGl3tSQ7G+tpJYFbUIW/W87ZEXnI+/9Vul8zgQf5s3NXrjxzAMEk3v1DU3
9eb5NzaFohkcVEFBEjQbVACXlylG8afbAmOAKsgy2+2lev7KI93LzCm2k9CafdNIn5Ml0Upus9xf
9p+L5a2vcpidapz2DQECrbvyBYGoF9dmg4ZS8YRSvW+JsIvH8YAs5VYQjB8MiC8yY8lcv2hmxJOq
9ebQm4R1VNGpZwriZX2q1QPBa6UcdEg7VpAuc40cpQ8d8/7nwn7as2guR9OWVXoukdxPSWec5wxp
P+T+Hd8TCR7D0geWiv2a2vVNib0m6oTdfRCotz+w+SHmjWYNDNLbpUKm+34gQPfJ4FsBpL/a+h6p
bw9SPL99mXctzo725xryC75xP5ccELLccaDp9VIB3UZ7E0obEzjtGaSDLG4CQY0ecRaba2KQTMFO
VPZTssWbXU0qMrPyJkUm3FJ9JIa7Ljtc2ZnJgXVWNQlRyqolC/AQWwKbNA0oyjcRgu8lHSCINbAU
fUUl9C+BZVtaM/HLuJaR4Fh4yWt5p9Dah9pVqo+qrlwBntSuNBB/+2Uay2hpPRoIJ5Jh+9ufMg5E
7Bqa4YGIuQ2Kg12121TJ1F1CdBflphrPG6CRv9jOVSOcTJ7Q1aWK1vwdX9VoD8RTILQ04sAcWtKF
kKmDQryhX9SyJdjC6oGlc/7sBuAm5oZGZ1vsyfg3gyHiR6QS9U2ZH3ECGGHUZMsX9FsinocOo6YE
vKlZaCk3bCF8ai5Bxsb6dSDxqAOeBB/E6QedM0nqJOZkOC2JJmVKSMuRvDF2keXadYkXa7Rk/5Kp
LdqWAc3Kt+l8Lx/kkX08aBFHCw8gHl3EoW7tkiNetyKsmb1NzHUOaaufSG1z8lSijVHtKxfTGn3B
RwYxz3n4sik8wXyKKEh3lCgb3u4JvrmH3FqSgjjHLL1UuLE8gOobMTtIzvL2SwbBNHMHf2kqhm6n
sQm+qwIsn4sIThqsUOWlC4S7eDmDDOe9e6FDkdRWxLC36oF7zHNnqSS7PTFzv397srHcD6qhLsHl
27Ui+nIKdWxAapJAFiMXkW3YUWKatIWlVqMerbaYlgZl3M8c78Eha+hKorbgiqe+Vs/eA2iZnM2C
wvLDL1ju8Q1+xY3UjKmTEJ72GvpWe0FBTeEDYHQNkryM9PuQZVW9A7VAdWL1w5I7NB27ZP+PpBIT
Kgqfdtp7tMpK4RhzZ+Zvbf1lNtsUGKMwuX5wYOPKWuQhBEFkEAzHy7bXiqnvOyxPZqythgfevU0h
9fNvDOgJN3lcf1beQGa9GIQlhI+f8EvXV3GxE+MzQG8TDuNSAkmCogos/7e6bW9mR7SWuM+bQFnB
s8vSN/OcgXn+DGoA74ES7eqBHftKpWAn+VVQHug0OmycoVX5qnGg3VKp3TZFEalsfMQy4ybr1Gk2
0tIo6xqvHnA+W65WCFjhqXO0WSbhy2zVRdpFWQ07X2gsNlS0VN0n8OYO7xrd82BAfHlb2O32yCYq
AU4oxL/Ne+OSNMA71TNvBaZb2hmjrl6+io5ceMflUM+yhgAezId64yQm2Ys/qxZWZaKQD8eOtmfW
0aYgXhompCllmBnRPgX7BOpMQJIiTw0ULR8vRqY2waRNfFlpnNYrvlSN4cQMr/YKz4rna7sTdi5a
S8KbT+KNBW1Noax5Bg5KaRFY5bgHogwQE49TbOGxF4PFKKqonHgyyGMRPZqWmZB54rcyvLp5Q37p
Sma3BbhkyRVo+s0x1WhNVX3ftMy3y/CInW/RA7Kk2iPneh8AkJYstG7oWUnlpLu1xNwMaQ0b95CP
EXI6uWiw/iDd1CyLDh/1Koj1bADTdIFurYWAnWj2OkPm4Ec31tG56XBWtFFQSCTj3DelkG3hoku3
A6jv/t0ziVlC4+Lk2QiqVvUTAGsDETYd9w1O3KLykIM1I15nuCh+ZbdsFha8Zao5qG1U83ahsOeU
Rn7AZJitPBq9cBWsavlh+/yp8pp1uKlPOIJiE/sAeHdVZ4HpZaMlbxmkmad2iPyLyFf+vSzHfPEM
1Q7S66X07xRkgykpwkrx1jQcgWYTaY4X15MbDfltNoQCM3QiCgygXqXjs8IsLfDuJStLiKlTSDJz
tBfrCUVvMrrWXW/Pkgv4e/ECjZEoIGl7Zu4lgb1HKjhxkofcvAkG7F2WgWqfywUg2HsaVn9ZMAOv
OprzShLXe3qdb2ZGR00/MPzcU49d6b3EqJ+RXYc/r8spm4thGAjRu9nIvsFBZUhUwZdwI0UQslkx
u5QE1lP+eqomQMiDh9h2EMmsXHeAdRH+zhxFLStpWzNLt3tFBEgdnD2eWXzWNB5HsdA6NVBPtuVO
ZZM9yYKRnU3FuETMSG9rUEfeD9imrPogZODKtV1xRBGt657T1XfmummlWdrCccmu2zJzamV129F3
achv2Bokmwu699sBcPRpP8YIBFgh+EHz1ARFua0RBMgdJJMfE7tFw7wOxe0ChQj26jhQ+5jcOHg4
4SPN9qjmCtddKevjfAOi+PeTvYr0k14sw5uHCdJA3pbWxTA9JjYDTydGw+G2cwQe3rWZNaNeDc7x
v/AP54T0Qbr6WpSJY1hLb+Cy5zw4/fGFHALjwMhtnXI+sqxmsjZgR3Bqm1ekubwXPx/xdMljJyTx
fDji1/+97iulJenMDTSSQRswiXX616Wv75r/o9q2iOvpWXXrRVCXVbnuhp//IT6mg30MKvvj7sFn
7RVoq+Uij2uwBF2loE0cs/GMhbdxCAo+66G26Y58D+gtrNbUUrNUd/Mm2RfMTZseh3oMgd7R6fVN
KEJQxWsU2f7wleGyTNlmLMffQ1EVCLepnL9Zxy2CVHxcLm9OItkWMNwazckb2XIw4ZmbY9qea7vu
5Ewjk9U1kYxle5KWKfcz9ch4kcuKjGGuF9rjVUBpx7VgdeX/UJzIrHat4kxB3GfzbXJlejkbD1vc
+ryoGvvMhURVfzFlGXNU0f9vvUReRqN1li5MFyeKslHoauJQDmtzI+kFKn0i8Rzlh8AfUpuRmd3z
BLwoxhFiFMn8PGL331f1SPNY93FIHi9pK1fQjyV1OxiS65LAmAozxyj1TlXd3TGplNBeJUO8xWRI
4mDJc1Uc7BdTKKp6wDMW13HDJRBuCnUErvv8wTAf+uqDpZFsExZbhszjyd1BnuiG8eCaMUiq3FpY
odXpprILqlNq0ato1lSUZW2IuXauel2haP5L1CKSrBF83eeOdsT7kkYig14BoitGW8EPNy8I+OII
0Qe8qqWl14x+kdz64sdM/8+yeQNtO9qTmnDL94TmaqZdv5O8pAwVsUHR6hSjaXc2pSzavgr4Q1df
eGPA4LJ3btYPB6F6fFAlcPAMkLMC4bNnJPdfM2kasJHpMM1RLVvVt7LzkJAyDEs5q9n2j6CecL2E
1khSb5XbPt6jIG9WRDbP1Gia9Q4IaS6e64cCh27hPWdKPTYCo44RWn3gafgoPQkotz95gTkJ8HaT
TewlMOruxv2Kc5TG5cTHbJME+zxcYR3FvJRnnXbfFC+GkeyF2wgbgKqs84SHhZ0Sfb0LGJ/OdVfq
c2dtZ/Ql9PMAFN4xHLfNUqHV81whtO7sWY0LMRRSE3LEaXPtaGaGlMldubjeAkv3IU6Uxvcb3y8Y
DjVJOGTM9QzSLC3pa5uSVFq7Urhx7GkRFoib4bVa16f0v+ZrGhhmSO2DDD4Hj6VKm6w7dxNfn9fn
Qz8S3qkkbHOl2bZM4iqjDIoIo6/Rg6yJUBGEcf+pugAe4wJwXF9AfUMTtJZi3ZtztzvYKLS0VcVq
0VGq/Q3w2mdCepfySXclWYShrLF6e/xMHJUny6P6mXyuhoKSdtYVaoutu7jDlANZQgTcqle5JwYG
6HGzZ4Sjk1QKpg4n/CQAVgH05F+DYxYjLIHEnhWBWKikf7vXgmLSc3OvSZbjdPr1CpbS3btS+jQc
LnEJbqNQ633qI6OIimVpkNJt6ufJhLADfavYbXtx27sClYjbWLS+k02sHCbUbR7RjN/CyRJ4hsFg
HQAuDDi4Uj2fUJ2/bNULMOIxHZXZ6tTad6cLMXJRZz7gkOiOXZVlCaq3ZeTaPVHryelHYCz3twBE
KD5j/ScqKKrr5Tqku8mCuweux8ymewKkpShiJZ+jJdGwF52jtdGe8NjPj0Spuzt++hYfvuJzR8pc
jtxN/rOcx3F26fjCL8FB1Qzt2UKUN+P/mwwTtTIrvtnsddz/GXpDYUB8hKvvQ77PVKJQ/9Tqipsa
Tdt8cahWvPGG4mj981IRTmLMtKpoQ4yquNkqDHf1qJRootqElYYHOmYjOw0W2su/RC4Qh9BNzEEz
pl3VoHHrlAxyrBo5tVbtSsove6ijT+TF784dLD8UV9FYgnsfESjMJUs8ZAC+cE6rKoZdEHQJjBlP
jDKGsGGOJZ8KF33kDhWVEY6Bd3jyC0qTSOvym7tHivSVYJZ1z7KgIicjD2kWmEQfs6Nd6eVKWimB
ttsIo5XohTiWtQkdh8c5ceHvoRmPtm9XjfE/yTA7msyBBXHqnkxcw4L3n9/ElW8hE7rKZKrr5HLy
zT/3hW40Ee6+MGM7l3h/ogopwSM6ENuG0MzR3O5J2LfYNvOIHwbQY7yQkJRfPqUtt7wBlgR9GZYW
3U9ov2erkO2cbLQTNL/0K+bekxaeRhSrNkq/sjhzGs4rlUZXy+ldJKVCkxNrpZr92UCMRaEF7lIM
XK8nCJ0k3wqawxaBJzUz8wh09CUDGGkYgaPA0Dr3zhpfcyjzj5VAuzv7rRBhCutseHBCT9aTVh9y
VUhwD0gxcPbPp/XHACcpiMhjEK4OP7PB04ygFpzicjpUBvCDUU0T1No8yrJZ9IzxNe+lcb3llzE1
OniTlnzXbI/yPcuCIDBtdjw1du3WyeOZNtvyTaMCFTFBGRGse5DGZJoeQgzTEiUb6Rhb/M/AeLe2
AEAiCQgyuk0zUTH9LBGa/EkTgoIMEnHPrYmUPsiPNcN3GH7dYJ83TrbEZ31WrWKP5u4PERBY48Kb
tWAQymAZN9UfoGUQ188uCmMKr+Ze6+RLyF7DkDfJ80uXJ3xumMQNz7AZjxOvLJE42gwOwoqSpeYW
3zhv/VscCYna/dsYmErxpGj4IBOxQKEQtTLAKlCcHnCT8pS7iL/ndA2sbHUZUL2qfdrTVIIAVR3i
q5I8BScoRkNVyXsAYvdW1aPaLR0bgyHfrowNvrWMVwW65l80hni74xkyA/Vosso6z2FGr3oVhZzy
Ulfmu+1JqGPel/zo8N86NKyeZINVhuaQJS5F1hRRK2Oxi8H1aNglBuCp/KLgG3yIqTePd7hmOqly
t9B6S1xfdxsS7+wKGmlv//uWcuhRHTNQExjAY3ZrMo5paT95Za69M0NwheHNh60/ZJdsZ9HfNMbw
g4QD/PTlQv9nl8i+Ho/7rwgieossua6vc3wiSnQUgvUgofnaYkJG2/IJTEYwR8oKLIbfFQGnPl/p
R42AjzSX5+s7uiL6AVGMUu3hCLemmgau6iTqYImHQSLo/iaKLlqxhuRN7h2GNkg+coMHtPPTqrEd
iCOXNQzdk9yMsGMgiplrc032rGTLaA+Wvuo2A+VL5SIqL9b8Sagtv0nATFNZxfJaM8NhFaEI3AZL
vC8wrJfDMNelb6MHIwbRPSfbAapDCvEsJGuI5CGLKc/k9Cei9FBAPZuyUdV/j9WBC+066TBQnJ7q
gxBs2+MK8nyYsNZ6X0kp8Kf4pKGKXnKKPY43YX/tVdY4h1ySFeYTSqNzpuZo0HiBgpA0EEfvVUYw
e4lq+oUIB/LGgkpHm9ES6dF6OYRati4cUbDs8+ZCW2VxaiNFiHtI5ogutPmUwhLkD2NSnYiJ/CHd
PiG5Jh9TYFAuL4u24t7E3jNBTNTy03RE1KYiZ+qJ3LH8PkhzaUijKl5cwqrJbuFu+jdoe2J45X68
sS91gUkzgOY7HJhyy2wx1I81QJNnbK16iBzhYxj+LwrvYQ5mGL/IdGYWjJgV6fDjjMjVLiaFYWFl
+ZuhQdVyhXpyv70Br9uayriO8b22qy3C2bSy7sympfg7G68CJ7LW/mQ5tQboZF8PnthYZuO5GEMK
p5VO1w988AhikuIbv9M0+rDNMyfB9L5jOlHYaWxlLkuqfxBDS2dLw7w158LgmIjV0T+nUdsJX8JJ
N4rMlgZGY0gNs/HJHcM50SP+hnE2VLZeULygtXI3hztb3dA5Vc7WPyDS3z4s6n925xUzpueuWEib
nfJvUVNCMLQxV46VuGJwR1KGOMwqZWgB0bbmiLQZObAzOFqH3Ar0/qijLCelM338EvDWmhj2XZl/
skeDt7o9rw3m+TvysR3EHf6Oh2jgAThMooj9N3ANQwRJs8H7A8WW+2KgATwL35hZlxQqp4A8vZ+W
fvmLkaM0C+nf0mvD32RNp4xF6urW5FJf5Bho/PF7FrjYZUDPKPhsVVfAx+hQAD2hl1JkYYeB/bqx
80C50O9psfj27hADZwcvVgqAwf2/d9j3a1L848/koOYuGBy2v6Z0FHnxnEeC1YDtSDHVhCR586Bp
FlerNyC4Wy4HI3zbTS5ECTKagGlQYeyBDRLFAcJUcd8I7UHED1u34uY1omt47CryUdn9rTInwneF
DxbKLGcvs1OK4Tg0YFBAdICn5tuY0hOxb98GwIJ511BJcPQLoTuFj2SEal7mf9Nf0BDuy/j+YlCn
PNPZU4DeoarCFwDAcoVjX0YG9/2B3aw5XeAv+wdYgLdKbbYjy1ghhKFTFPVd6qwtPcbs7O47+tST
OaF6xRLDGWdD/hA7o5eC8QPLS4jxXOrRxGuun6Nn7RJJEDU4M0Pck3ghzy2lCnPsjwHW5HGuRPoU
AHbfJUR1OTJDSV+v1TNpT8k40GWJJA2T3zPnYzeALNey50g+QJpgHMQ4ZUaCR6N3EqoqLMdoWDw4
vJsCrtLLO1/k/cxJtiInqi6g7/xIH6PA6rXYroDjPC1hmQtHF7EExNsle+Fofz+Y2L8bbC04K9pE
Tz/RceWNnjtSDJ/SnkXq9NgE6kC2ZrTIZuFUyt/Mcbl8yBG1KIAyIE+hr53JiKatMC7qQgZ6hBGf
rf1RqP2rcD1stzZN0LWeN5XrN1Hw1WKy05pcaakutOQ/ivOUKlMaGDS/sO6q8bHdA3Ldmm+T4Kcg
C5PXKPoMlLbLlq0xuBxGZNFxw7MWAwumYmN1rWzf1Ix/GqDEm0lzXg6ssXqy1R9E/UK9HILjuYTR
LxMTIS/jd8NpIH8J1nMyMAqf/ot5c2r6/EyuJOjNHUvwBQUYRMp1PdLQXwoPQgn1Yt188b8qiVZr
LKEVEwhN3yDsOz4Kjut8pRXNgYRTUpJSWP4P8pt/msZ/7RClNTkkh8pKUt49iGn4UNrRVUnfC7cu
wcsVC6HrZLNSvknWd4RVckMniLI3Yp5G5q/2/lcqeYyq6L1pk0RqPN1aTsh+ZnMCGY2t54geXAtz
kSAfkLk/guji0ktRLsSN2IRkusN3irsqDlP12iRQo3O/ldyC8f4KBSfoe6oeHk01+qlF1F58psL0
tFWOlrb9pd+CFIPmvsSItXIBQgMcSlMgPKDsIkZ1Sj7xyDKJ7nAJQOoA49ThbQiaOvQmSbcp9lI2
ul7bY61LAc4YaB5SrhRJIe6QkGz+5aiVKDSEt0jO3C2hUbGIPYCpZ39NDHJj+NDe6jGY/XMVWY2m
qQS+Bw7smTG4xmFh9OdGBXe7UNctnws3zVIQ9ta2Zq817Hxx12H+uclSuiw8pRLeu7cwZg96Cyqe
sMCNDiCkGhb0GWz/lsmS1u2gGkcfi+uCgQ7JqjnOV+9s7HwknV2LOxAm1dABvmNfteZsC20sUBWN
/0Z1mlOujKfQLwYlA+ldGFwr1TMiUaYArLyZxQranVuHtDP3ggr3a+Xlcvz/6Z5egCkc9b/nFGZZ
HiKk18XtUYh1cKppTu9W/DN4ePDm5TN8+waIoQn4j3OoXD867n5cG/3NrMK43HNPSsrJX4HJc9lJ
maD7r+V5VGfTbv9ScQtK4RnthIfNXUIxP46cOaAvyukX8ZIYcXlsR4bOGPX35+54A5rH5oJx9upz
Tn6KueOLeR5k3cvMWQh9cb6fEgS+luJ8gLFHhIvU+e7ChCuFAioVXtSfZ5sGeaW9PL7IzO2O4qPD
SJMpVEgh4e0q/42OSyOOwo0i39Tv/5v3d+W2IcBgAPJkPllrMkVIFbagz4EZiSAgLdYJDBWb9Mw+
W8UXt+YI24nmZs9RnX9Ywnx7pp4g7qnS4TGGbckHLuBHC89XTPPbbkqVMAo+d4haPDT1BRSA1HI+
Xbe7/FCzDsr/Mzq1xiFHAFp2mBnV7bHb6Dzm0DMZCZ7s4efYsEr/SHq6GCAvAo6ota62GxTNJRFk
doOygvI01+c2YZ/Mfi6RvpBAENtjbIGX5Vbwk1+Kq7MpQp5TQhYYo/gEnDPandnc8ildA0P54Ggl
EsAGevEvZgkOsOiqzuksBpzZyy35NIzblsVNfJSi71KyxS/ABL7LqgYCDCn8WivF+vnSb2T5yGLS
qWwggrj12zZ5iscHHYTuEV804rkuVLOS5PWs5gkTB6QtyTRhoV0Sbj4HP1UiQf7CEX39Mtw0n6dD
g3WabkcGWE/97smjBRxuePEhi1YIB1Wh4mApWHIlovpCFkfYF9C02+M4esaKphsNs9feP9aX5c6C
xpRmXL1WD3cZYaumYZnd4f8mkRZDHWVQARV+HXpnOmYXjOWQi3x3gM0lSzdBVfLmJgFzm+m9p3d5
iXhqua9u/VGy74wiO5CPP2rZrPUvQBwuZciYW2IbZsRryzxl5nCoHLstfOW3MxM05HfM0X4h3dhp
v31+LqtpYhD2whi9kLOj2icB0axYnzcpRYEVBkDMYJZgBkqZpUNRarjIgtpqcUety122mRUJ4kvz
WZCOQPkhhBkUZUix+PZZUiuBAqROJ7D05xF4O4kGrZisJcMthq/C9XKkASj1kkU2fYHpP60GFkv6
koA/6+m8PtCafcijm1jIBLVdZpQ+ANuFyq4Pqdu3F8UPrTyw4Ug/J5fUQI+xXpAw5BgK+pkQujAQ
ZzPqbTRHmS2sevVQ6DKtCBnkdUdFfGPNb1btNud/i/wpQBR7/IkCP+SmOewpDgRnND2UuHQOU3qi
j3jJBu6vQJU1XvT34UEfIbymIt/Tvfgf6IolR5fLshLo+VLKexqQnJGmBElc5gafyAvgiBkF8n0W
qnjHGIIurOk7St/9gouw3PXLg9S16fEhEnqWfRbpPLKxVpVhG90RG5eVc3P4bSm5t8s0TuHN4xu8
pRmdioKQfhf7+LAVSZZwqb3mW/qXoM/OZ2uZUg3P1ZZ/lrEHJDDoBkZImdJWwUWs4YN9DlHn4y8B
8zfRwmAPFs1mvKoA+k9nsxkjzyW/nqob6j9H01ygACeMWt5KusvilQUOTjeyf3cG2uM3N5LDcLF4
wXdxVZTPOwPYD7QcJDuaYx+0xOxwih181xLPxpVHJigawqClPMR1uSYbGaVU23YUGNflPH3s7MUD
lEyCkhb9hfkkK37DJns4YYLBMi05F5yR+nLgwBggq8mIA8MWjIjBGDzJw8sAcBxuYOqBUvJVTxyK
kNGtne0yXp5W3Lc0ptn4PzF6R73CW7tM4PGXq3meuVG3o3ewDEuBcyLNY2MVvw8+M5zHgoeb0dcS
cSfny6ZCDJBV2qi/5C9s54qVl3lo2byPJ4XNn7/9KWtWuCXsLkjg9XmniDm7Sjhp5g1jokSgJX+z
gp08q5Kovi/Vfh8GkZyrn16/U5l4ZYZp9r6Hv2b59PW9efOl8/6G97yEcjLua1cHgWESfcsA/jRM
Vv/E6fd8mqEaUfa2qMoGOd+Yi9OhxeIEtdfDn1uM+RVWhZKM8elTos9vImi9Ij/FbrRcuzX09c3r
+Yq0riQleVPyq2rZYkgAzIiAugbKtdUrhMkANJ67B1259r4Dt4HP4r1msY4GyS7zBmjXi7yUJwPX
nMY+HFs9erH9T6ZhDSkLSf2svF3VcXGHJrhC8MP6jvLD/CtVB+9qse2nrc/olDzMLkM/urato6B0
mujSl5o+3enUv0NQWqLTCVWsE0na4AR82DTcxjaRfowVmVNYXGgWerFlJVaKjYbaFZzJwn+ieJSU
dX7BGkOO1BbHHOARxTyTcBChWEtj+54U/aOtu/Ir4qx5x1gYMY4iUnk8C5M8A42rzYR1sb4UhPOM
5hJLDxy4WGeKWT8DumF1EsIQCffX/WILtpibM/Uf2uLtk0yLftcaUm9y/Wctjm6gWJJaXbPDrJhj
nkh2Wt3YT0GCS6lV3OsOWnWBKpqWj5qAv5Xt33zL9h001hHNUXIoVeQxus7clHJGIbojL90BMFeG
3+5X7lc9dAujUwKoEJEZYj/zAFDwBTRmml9Wgk/KXuv2+nYse0bo1UooJtba/0XgSUghJJHyX8ak
Zx24BusnMbifYWTzKX8i8j7Am5K9nfTa/Yyn0r3jxpPT8uYpx7mUS239Vz49Tcehgji8+rIydWVk
YemVva00cq7GXRttZ66uY+zY5cMft36PobJMWQAcSzmFor6n2xJBv/xKFlo76hRyTIdw2X/lJgaY
T+Q7z/ebpD7dWC8amDFoVGHNywTBrLd6NUly52X1shg06s/VvxKhSQMIYeKXIg1OROCRdfTdMZDj
dgcmT9fExh8o9Uhg1KPfB+ypJz8pnh2tTSNJPI1mhGYrpPfI+LZcHNIRKPs6Ouf0cci6CSVwoSRp
lpAIFtupwNrxa51JHLxxx8Q/AYCEjK0VEFhSwg/xbBqARL64w2TkWcbMm4pjxhUC5qABcI0h7vgs
RX2gXr6feyikKsM42CbtwyS7ArqI17nNJiSyITIGTMDoyJqgR2dhtKIfgl98qfO7nseCyZlmznMj
rNUWqYLd58RHGvdu7jTSigrBooEqyD6orWzDba+UFyQwkX85hk2ibZ0WMN48gPRMZ+H2/ygJyaR5
BhPfRA/qpoyvdzUcwnskcLMy47i7JlqXVnfLI7JYQ5MdXK+0UOT6l1gsdWBXJrCJgJO/XslwquGM
9iuJVTIWKw2lKt2AeSqNQhuGe9JcZRYNaFPPzeHFL5p6Cl+P5U2+6NYZS9U8E+1fOV/udd2W0bS4
SBen3C30HyGSFfaow4HihUFWZi9qBlEG0b1LkZQikXi4om1yowk2XfGzfID9A0AK79Ve/AtmE5Eg
Hw5bzRIp8qYUZOlyaDCsMwaHQGt15vc09OP4IFeoWQv8hN0y8Ri2RpqUXIvHR65aM9o9TSpMSGBs
rbZzxEo0KOuj7C90JcUMFQRPuZ99JHBrcZ5fG1tIXfGSamXJ92zWK02xWNhGNJMrtX9vNkaETgYD
eFHA+ewQaSfxSHqwHhWWhuO6cFO9OGXT0XXQtj4hMQTGK9n9kFE6Frf8Q67AUmv1RHYZvA7ZzgMT
OLlvLJ9ls7RvKd+6jGfqeBiNCsjuvurRz2VB/ObZCww2A854U3eYbCag98TjBal1oJ7ZUBoXGf0D
g669ayYiBM5fN73Drl3ooaUuJKgD9XRtOsxm4gqoMDiCxt3cKXibP+zgxsAjuI5xHYXTuQUA6JO+
yo+1hh3Qw46FIPDTw7sQ4QTVsNo6VzTyabv0wNSgf9nZge34Yv8/BzRLJZDuUFmEzcdA7TLfxFT6
FOAzWPUEd62j2SgnxH1Uwf6wH7RE4pa0TDXdaQjH6Uxp0i4lL4nrsNWRskVFRogX7RBie4MgQYEq
3cm+DAM9w1w1y96bv0Ki4VTRPwkYeVYZOz7kNyhfxQbKbGWoziTU3oF80ME8osyBSzJJ83pI8Voa
22QaioPzsWLox4gjKx0nFYDcrxFfEhdkQLICyRp7LfeOII932a1kLQAlpe+luRCpQzUu+GLcuX9R
paOr9sMqNPtxVkDZAI0OxaHHVtpcniY2fvENBfxg68jLHoIOlNacGFJY82x2I/O1BEhhmTUsfXML
N7N3IbZ0ihLAMPIh1kZb9Oo7Bv3LFn6NOx1keXU2RlLdLVqhbQlc96nL7ZgZaeAZV2Wh/XJ+k8hU
ckCUb3y+SzEho/C+dBiqejkDMf+bKZqVSjQ46rrXqVUs32KBvMRpXwl0vl6WzuzgB0E68QmLxl0Q
eaexTPipks5Nrz/k9m/ZyeTjBHwUP8go8Le95IeDIljLlz1SnV7nUhs890ZrUQlZ+w6+uFEa5ry/
1bYEtfHlQIhgNSdtglzJrzBeZDHMshdnZPtvZpudmk3WLV8VfqfKGR3aS3i9nizGo1/GtFaglf6+
idf4CQkGTRUPmAK/tQeUaTP4hm9GF8mFX0GBf/iAk41elE0ggEfiKYsrkuxff7g8pQs2UO548CUT
9+ra+4ieK86LKyBbwyCLPhkzS4Waml3gW9u/d4Bbz9SZvs95UViC5jRHNd9+YTP+tiymgdJLkaSb
RMJnVLre/WhV1c7eAbWX7XQOLE0D1I50JiGwZTOvZWCawS70+zqewwZR3uLK8sgVWyr1H9+Ank7U
+TiupNeyrfvuIdj7jRsInoFrHJ+ZErDGVK7+JRDZCuq0CmTLF/Z5jocU64hQYqe5lTUMrB0RZZ3I
/wEv9tRTJEX6bi0DmzvKKBhhYOvd6H+R6FDcPVB5kgculfgEyZX4J6jwDJi5V9Q5Sp4OYVldbIe1
zX+kACFTbBZ47sYjMA83/8IDcDXGYzYxX/wguzFQuBuRzowhN+Pqn361fhl3INKzbeYdidBfYgB9
k7BnrSW1rcC969hM7lYWVnr6AYCEOiPERdZ/sP1BHfYKnpj7UW7SnGTu+y7AY4A9qcR9NcbfUd1U
SHFk2eYyhi4dh7O7QgZxSC7durRK7DBzeYqSPZ2P+cw5JLM8wrJ+Kud7D6ob1aD0H5inGlXdRm60
p85cz0KjvJ72hHb2GjQiBlH/Rhmfryf1ufHZIrB0/5MOFEVe57c99txXu2NgDAAfUSIAx8roA3uA
K7EP+Sig6H0QLSNHMc1eLmK4PvIS0qSq4uwTlOTitqKCbXZ8cq4Ga6WVmnLGYpPAuL9J/Ec/1U60
gTMVjq1F5DtYT+FfMAJnvieVz7y4M/YczW2od/7wk/yyXfyfA8uxrkOUKDc4B9ZeJDA7sjkEUS7x
EWpGM/ygp6UFuIH02knPnYuIq+y4falF7pWwjiclZ8wOI7+xxL4UFrbuxYAz6OHTySKdkLPWvqOl
debGPAFRa9DrVm4SRbJumQVXqNt69++Vol+uDOmLZ4qKbT9j7s9rYvknXTPaQrbVE/pcghQcqlPG
AsYSOVQ0EiQ++GjZ0Cf3E9iTj2zufylOwd2GX0Ym+gK07W2KdoWcQjuAWax9rfaqiKH/67gI9trF
MJ+5RG2ga7wdW9AvYTYqYlTuA+ZZb94tDqMFzoew5gdnpOYLDFrbCFx9U95jto8N/nUVmr87gWWk
PPM1F8aS1GXyx4xHu+r5E02XEEv/yI4TsecstTaY76uTDkiovItLZ8/EdmxwODDdVWsmR6kE/t3K
ccNW0zWDXZSoQW8zMMG+sZf2s6z652mepDLGkHkvENqO7WkdM+F70Mjdy/ozV5tAy7NlBGfiNefv
cXl7wDBmzccSKrV1w+TC8wanL/oT0d1Bzw8CkGnh7BWGDIHnTjEHBseqOxDafV2LWmG+pHh8De6B
fwTALjh+2nLHKrscate1cvMtj1KaAJ0XAyKSr+Gy64sB/fn7ZduXXqER6/C3yrjWyWfjjVe/7CaK
77q8bjc7U0eFHpcKt+YzjqJGsY9YKWnuQZ8mjem0V6DYkcOm23NTbHEphPMJ3z+OmWTwtivk8MDi
CXEUd9knnQpsEXLe/Df0xDbqAvJrf1CUVbhRQXvBCXeePCzJIbh58gT6NV/rhVtl0kSdiXCm9pVr
8mY4qRZDv9vxhrKFI6CFKT7J2FlHj8qi7ZdBSXk1RB2qVGrokDl4kVrArHypLMOVaZ8ZaXvBs3B5
P74TtNy1B1nTjJ/5PVPi8RCaff9mipIFVIW/4YdzujJEqEsTGPvZzi7xpw+K0KJSBHVRVNyJA1OF
IS6UJoj8uzICtPpCy+7XlCYQPm0W2yv5FGfxaImY6BvwrhbuS4o3J1binxng5jNU1xY5HA0b9VB9
aAG53D1C8S5KntbYzJ0JJ+q7ax+fTq2rV2h5xwPuDIaX6asXzHGfx4c3pnAKaMUQln93AOzOOMTI
1CA7vYsWbqSALCXJEbb6g3IAHFHlJxMe1NRQnpGA/0zVzNxg0FosTyxQWR/FjaWE788saTXweN1j
hBQN2u3O9/IVhKP1503DBviIIPI8VDk6XiPqs7ZTaRaSYr6HM0B4tJbKcYpVWxi5DzrDvH0pTa4j
+yh/A/TNcMqlRMBmARTS1oiBaOl86Lk7e6pWsfsFmIrT/+M2JCjKzhJqTNp6uVJeWng2ziBduYCP
aHkCCAyoiBP710cAWuP+9TU72E8952UI7+eOyRyyW318tTARuCYpyCypuKLVCd5urYK/wR25/URX
uot/VC1Rw7zxpw/nEq7Fvp+ffwS/EAKW7SWqcRg7ywPRKH8wpCTWKs7FQcg5BiRzcYnu430osvdL
+Z7l2fu9Sw2lbAvmxWUttOTyrLnJQkMJoRLliN99aNy28Ua7xOXs3CeZDvGO5maZGs0f3/7+d6ZV
cxx3Dzd+lzShNhxfC+AHONq6bVtw87u2I1R6GYQJtGpapkWPJ7HudrRhLKGO/uUs6Jd7zCxBNFU/
3awj3UNVIHK3lJ/p1pUBf9LMCPvnPDGoVgLAzrQV8HoXIT7zRcVQwu1D9BrczaxKHGpQ4sKSXm85
OxGdCBjiTZ3pu6IQvBQCcW1toAPU/s9t9YRrqPGGBw2pUPCNiwyHanFxLUF1IXsHKgfS/exAw1cY
XJEqTTIR4BuTwsm687VNU4e97OgwaYqEAu3+PpMgTzNUJVVdGNqnRenChRf1l7PoZOTBJ0HsN6aA
LAwL0M5e0Af29G2spTTVHztGnZbx13KTS7rUiwdLD8L5Xq9CbuFyrZqCBF414b8XM8pz82kNfJbN
j3oWt7uktpw8r8TiB0SU9d7XlIAid/VTVJbDqQI28qKJI1BwNZl9xcEga4xgwfCGsbfbTsaEcZGs
KC10GZwyJRsaW63icDUbZl4cvLk1PHuh5p2HuJcUCCOOfRkzt489o++zYzDjXmAIgc20nGLelAaz
/3U3ZSm2+D3V0Bvin6D0QcTzMNJOfCCqh3ncHAe/PNY6CpO0SxUgmDzagflI73x9bRqoWLe2Dnbm
/o9UQSctc69PJFVPzsGla70mRzYNMbxpnHHtZD9HRuXZ635TUuTOu8cACyqVPJQVBGN1MZWYwOa+
VUlSawNxFumOtP83+v24EgSfW1EBeQ/tVs9PRcTleeDkwkKfkFaKAfIqAvSH/lLtYrp7vvd/UAkH
aDViXSBWqaxFE2vppvs2viK/yDu8RVMYDk2jc8dYut/0XK72XyvwvgUGSWgeeFaiONR2EugcYDXk
kkJXSZ5gQLcCdOb+TBIOAA2ZzaxTbU3bw5gephBi6/qbFwG/t7ZXDLZeaGXssHnAFIIphX+G7dg7
Zb2ZUbsThDufjz7sZAv5yYAs/yO+5ROyt3qHa+pSGC6PkGEW9JABDDYQo/hRd5lGCELyuMaLA/jd
aYsNFEkDDSdDSx1WACRPfxjVfhovumeSm7PixsZyO6G35Xx+UdPUu+NmYQZdyUQpc96tQ5UMtyMC
kC9ZB5uQ32+JKd8tlKdbaJytKJ5iRK/BfjjGeExTJ0v6amV4r/QphXy2J3hkxuuPZiHHorLtiiRM
WsKi9Ph9Oqg/Www7M+bGeqC4Lf8roYUeaIXGQXBEqCA+XpD9cOOqgmrHrl0brgGbr8oLrNvKhBWm
w9KQqlCuZRh1upnFwSXx/EepOiQAPCOdLjofsvQ+yPCuQT9YvMwdU0Qpu+uOVFl5/iXmlDoM+1tg
gUkSUXepuI3oFvweupFLoaPi2TZkyaUqy+HNaCw2SnMUOI2FGcJmu5PYzoKHc5vOHs/HGuiHaGIH
ay0wK96GwXAcJL+pxXbZHkDFvdBR9gNT6ddguop/6zzeKI+4prNEtg9VhIygJn29R5bIo1Nxb52o
zvJ968Nv61EAUrt/5IYmv4gqeh6cSQ2zy8hF+OsVVnGsYOFlXwQzGx0qankNAupoSN4YLopjPJ9w
4pxkev7GHjdifFhRqdJ0qgz/kHenYcTySoZIj5yoYqHTZPy3Gp6LeJzslQdl1V4lEMXsmFRMdVeH
EOWB1ugM6lXWDErSqKY5Q8aQ9+0j2bFnJsk9kGvH5/vgoo+LZib1F8lkYyu2TsdZEXYc1hlREBuo
M4P9dpq6azXnF0pC9PHPk3i3SWQjQ8ToQDDQ2GPXOobhlst5wVr86l45oronZpHbg1knlxb004bB
R/acOtiaxYYRNefr1wyojdCoYeS+nIeJnFIxh4AGOqgjJess3q8hS/mbI+pFFpVsQQO1MG3BXno4
oj+PdaKB6d5Jgd1Zc8h2oWRKsR+iMnfwE569gxx2Gr67p/vhnTMi00pN7zVQQiR0nKpChir5ioPe
aR9f0s7CH9I6DOtjeh+fnM1Rzex+QNQwLW754Wybq29JI0rLvvfZUjnmRG18S12JKbtGFav88/Lc
i9K2r3B3Rt016NUE+KrGLojrUjhZEroCpD4NSJZo32aW9/ksmdzZQsPJTtWSgbVB7stjB6irSuLv
nKkIQojIcoNmeYt8/I4sO/EgUhuCGmaEykG1UZ5ouePzrz9eMwrNuk2FhEr7RxqpIPXWoRCNwt8E
KK6AiTa5/lGCEw6eNJ1yFYeNiyBafr0dEFM8QeifN+d0aD5yCeZYs6ZbiTYALB79voEN8veY9vCS
Z4/rt2TlDsYIgorH4mnzK6w+R0i0XTvMkoyiryf8xmEuyDt+g0wO85MJSl++RsV5+TKU0Z6FKyC/
T0IeIKXc+W5M9+/C6u+tCKak7pZgSMl+kKi/FIeCx5P6pUVW0SLm06xz29Egy1JMt6EKbRU0Z/Jy
Y852R6fSUCU3+Bx4Bn8hTfHMQvqBMHNLIr1+4ZGA8fOI8UODaIjTKGiHvYeLx8gM6KJ77UfZAM0R
2+/3gnuDAZDkXV98h7pk2Js5AcS44kwV/32hAbyw9SCIszEQ1iWmQjjlgIyF4nUuKL45LYcayi3k
fP/h/CknQQdCJjPkIsOcgBsaHlQYv2PoPNAajMpiINQYF9V4eej0Wf7woNRhul9ztnpbwmXECa5Q
6VBP70ATYeT+m9Qz6L2xT/kmh2dwLrFJbiP0m0DMPeHHtLfZnXHt4jtK5buQtmijoLnF2JQWLRnD
C/QvJnBF9W5D45UKVhZohd5AU+K9m/4xVofH0LT7nmTZJ1X6T2FyRdpu51w1w2fLPTydRMT61d8G
UMdIiDKSiBtBxxSA/w8+1AmfrdhJsGJyHWmT+dJw4lsrw/Gm65oTt8tUKEDHqp/r115R4oII+ud6
0S+si31bg+8azZXRnj1S4f40Q0xJbABS+AzdUN6GLiUuL1Ys59HHcpXZkwnT7l8Sjimc3U1prGdE
nEqPobBVS6aQr7yUHtR6Paodpa2QIUVtPwjkMTuFURGK5q87ncVPMt7ry6cFYfIWWEPhNadXaUP2
dU1kwqiyrLfZEcl7ZAA/rWWvg3lAP2O+UIGx388UllsKzPdfkwa37w09jEwhTmXFxLYlMHbpkgyw
RhP+IH2i0kzEqz0dBs7+pXSkNurlkqyR0rzX0UxTwVDGaywzv5BfM7IeHPE6HXad7nqbmp3fl6pr
VrZtwrvVr59wvczkd/KBFpNmkgxSEUDpIq9fIB3g8SsQWQClXa30UWf8++X6zkdGSP5KRNfyPorC
eaBJZrN4znHgE1ofNGT3v9t8XH8nTiDL44EPRUjzHSE/aD1B2RwdfSK8Xbr6w2FK17I9BVviem3D
/7VVgQmiLufWVB6E8J2rFYwS19KNsmvrdidmqTXEITA5tzhj74AhcK2JIyIfwqgjA3Pu84qqMCrp
9bz1AxqMujb818+2cDnobVIQnnRCsvx4RnlQ8HI1dFYrpOcvCfI5ruzZSdDsDYkA+b+7vwac24Nz
zLkIHYXp5yyZGbRhQvnr7XGhQ6i+KoUlYUtE8eRyrbaBlIQu1wM4kd4AfI7gnm2SKKaH7In64TKe
C8ZLtDui844j6AZBJCEevUHfx74qxJt7InEU/UtYPendCOTK1Ad2G8p7a8rEd0VuDr39WLBEnTPk
MyfRZzSTkRdMi5lClNnse8SOL1z5rIIZnDM4CqyxBA+cm08zPyEaow8CexgLlpuNYkHbYfdD+TEj
PglQ2cAWMIz2+6eT3gmaz0cWEF0/C6ZPoRVIn5MV9pGVhGaDzcmdelvhg6ELdkmvp9dFbnKRM+0j
PkF1u89Ky8N+r/wGi9DTa+YvbocjMszVzzZKDvrh2BANAP1WvfPRqge4ukb4D8kMYLG7yXv3x9Ud
1rwuq4U4VwRuYyVndfbtH2YoSfkvCD0sTduZtki9us1sT6BeO9MiWINdjmZfKGZTX8YrPF4kRDim
NcSs3FP3c5PR0PMjqbm5hNIujJknZBZoLfJm+SZnK9MB4BLprQX1Aao9jlK0xJZTfKutwyPOX18E
0yStdxZAxOog5yJxrPMkOh3qDEGtwiSFHWZL4kGOX3clwA+hPV3iQgSeB5VYnUv9BEsDVVUHi0mX
qpYfpBmxxxhcC06nXyQGVXVTouZGXhWDnwKhZRd8ATJ25u5Ckqze0ntYs4lT1UnrgfH6LVfm9d8L
RTmAi6rL63yTslwQaD9jSinTRCai85y4IO0AKRDnjIBdwi4sZ+B2s7iPm5BK04L0SCdtyt7S2wsF
3iA52/8tNUn5/Yr1S5SPK6plGloskaVY98nGReUnjndDyOzeWBI1t/AQbb0u1k1dOrVKo6qjaJUS
cQLQtU01ntmCUCOCqK8zOjCXAgdgm5YSqNGyzz6/tg6AaJUn5Q+B2mn+VBLUmWMZlpgUSbyjwDNZ
4RximTTbKs14AepR0NXVSeUvoC3xZxIxEHrT4nLRih6tSilM3IwfAKTg6FCO4PuaroFQ+pPbEsVq
e9DQweeGJxq35IsAWdMEhe3qH4X/9wNZaj2G8nmuU0ThcMWFKD3wFQHOE80Nlndo0qx1hCDwsLmM
pRMvSNcEUTH/vi1AVdBeWnkEbEzLSnE6vTo6+ZqEnJzF098RJZYBTrdtiAnESWeFkYP+oDt0bhbs
ylVPUrA15KelrTjbwFE6j6b784W4U28NCnGD8FMrG1jpijPFE7qMGPbDbGNDsFoSdvo7GpBn0F9Z
zJMRuBPYTqdCTiiPWZMWtKn5BDH8E+SL9Ss9LSrjEA0msRt5xGT6W8SC2jW6jS5SKmIQNYE4+eeT
AGhosd6I3N1FsTve74p45cHhBymemKML1SHCNk1dHLuOm0aeIkTrjId0l+Sl8NK2TrcYLyUSHQSL
qBxBjVGMPCWGxlDchtPfeqqxDhLHI9YduHLS549q9wpcDaRtOTh6aiKi5KM1JprtzVgUg7Lo0+P0
bLcGYQ3L4TPfgjs3KY8594AQRgqPLoxTrMBbbSQ3WlnLsQLzsSWmZ+6ClyjU4J0w3cmA2on+Rc26
cc6glbOqf6AGgEpuiNmBrt52gYwDfeOCXlhzu0z1lkI35XeZP3XAEjMZcGblkTv93HGh55K76rtf
XPX4ivmv07IeJ1yMmm1KSoG/L/cE3PSqXgklkE2FkIUEcsJJFlrtzPsc65NT+ou2+zMWCRj+GzgY
g89vxnv3FT6vpZJq6vlyY00izfupFw3vu/OSZcnlIp0Ty5FRpVfr0adpxOPTnydiW1F6yk2VPN6I
G7BwsvF8jz7V7FZGqNEbfKlbpbFdsrgj9K/+OBPQyKRmkI8aVTJN4v6tBUqCUMwvTBZ7biJ5ftua
h9/jr71aRAfj+v8UpIwcVw41HAa3fY56e28DnASL6WM7l7bXws+SougK0y3iAm7YOReF6sCGp52P
b1HV75kLplK8RQu+j2wUS2z+SiIkryRXlX3hE4Jz5H0vCkIWj2usBVebIj75qABLwG/yaMC8Ad9S
bISFzdTrO54oW048aVEPh+ETY5lD9VkOmYMCnhIRw8m0QQ/+zjsjzG9Egdl21N4wGGESRSayuJOp
DcfkShMZ67Je3Cih5Js+HDjhrjlK9BHzTXNovBX5+8XPlCeuuorvUbC+zg5pii074Ah5U8c3hxk5
g7S5uus6oRgz9OC7phUojANcBKbBc0ctwQYVhgoymRRSwkibNCOdiM7HRoR/dfyObyJN+wXc+JjB
5fkofRhlbW3E1mAiMNRVbWDQb31hMwPDed175FbLYJss6xjsq0RGOX/ht767LCYbkcQ3ivk729fh
EcR+iGXls0SeMA8/kI11fXKHhwSw5Xo3E8c31f56ZmnywEnoJIVBR/V9ULG3vLATgFa7/VC4yDjB
YiUEiDYsra6cnT8yBljIgKVCrC+rCre4gFp5Wdl4spf8kEA/0bJFr2nlOJfame0EASIgD6uXs7wR
Z58PiTfdmqfPLwJp66uKYdI7IJD9IGTtmMJcZhTOxGBWppEnWtCnDfJnPdYbfDLUH4nLJfRyXKlJ
/29HRHnPBnlzoyIu2XM4bhyuhkJ/c9MzswOj9ny4O1poGSuh8b/ASUbtrMOCM6/ZmLywaHDIejx1
td9yl0BLNPZjLiJO/fgpXT2F3tMsiGQ9qOaQa4TAvET8ldosz5LQ0xa9BUBJNtsvRT5lrwiRSgo1
yCVnwdfklte/abVNAx18++CcPn0R8oRBwi25ExoejDY8VIcVHVAzrkXBXQ5h8Jootz7nOauxs2oz
0JC0yvQ+Y7EuzzcOLgb3D+zY9aIZ/LYJ3wBpfqI2l2u9hevj/VukO+RnCoozU4Y74jgj3e7ZsePU
k2kFepia2xQZ0NAPBJsuaME+7N23muaSBbAejIJBFRFnRKGx5N88EbFebXwqrAuFWvy78z0C515r
wlxfGqWRDwF3Fhu+t2MWEXZeZsVh85DdcniSqO2NQkFH5K5Lf+K7GrRDUVRaiL39xDe6s0r9WUDS
oreCoKEONG3ENZpObMXnF6HY/+NLUs/2uhUveCfVEneIxq0N6vZUX0wQXedzflIR2G+m9UCnmFrK
bm4udMuXD9vPvrV4uQbwfHd7SUsRjM0Fsy2HfW1eaRbZssUxdRvKQnwOk0/KxTGpRXI5e2nJwmjw
D9UVnDED8hLmkgRiVAVA0ykS4G1BCVSlOBHiFCYIbHpiLj1nBN7qeN/LqeuIbTysDOXxn4RAkkBK
b1kQHk1a690Xn/R/V1KvwlB/fnoWp9h0UWVv4TSdBdbHkL4LvSF/Y2huIOYdSzURMb2P2FrbZ1Fe
CKV4kteFnzQFyR+vGGzG+tXpQOZMREs66aBYxTwtRNYkb3DqWGYy2ghubFWgfHacrw5IWdvbXCa4
72I04IQUaTWMn2OglPnQ9oV/k2/Bm5LCo43eti1+Gse0uFbxM6kHW3mPJUq92me20TA+kmwFad6j
H43gSW8Y3ESkwCaH2W/HVvrJv0zLLsLeY1+iPStgrqrWx+bfs+rNv31tuHySiRxo7c2QjxCSvnca
lbcxoSoOcG4NT68rtxxfgAAhphdsihat2Bc73D+LA2klaPgsAcRCzZVQK6EExAScC0pXeGHYrawX
CmpLowXT85rh1qKcu0h8Dw77pkQfaZ3omg8nAsQrNaDJN8PREjhMQdveR0cwtj1IMHXQ786OhHtg
G/wFK87HBnR4e7D/QEWbXLnOSQwwR03ZrbOLtvKSbbZrqlsg7TlJYTZOACaoOuD61dfWfSWI/eDf
gNn2J9MNEB+28neln8y3lRzBF8qqsCcaafeIW4Zm+HzDqafLQRok+xXArxBpkrZY1G9RVrRP/7Uw
juygfcYW5qk6IPfjAruEHDBnYxV3VOL3BJgKJ7rsU9OpwUFG5Cp992snjS5Cla0GyA2CGadPFeLr
HGDgNJNa/PdKtHAb0tqJjQGsUwn2pC9tMYhct1MFwjh1nG8aLEq3A8ctzi6r+jlsoE8iEXsVblEw
K5e4CB6KtvoB4vhznlPv1Hb071iDBODbJGu7OEIA0OT6bNcdiVjF0Bq90hQrGffb74sH2fra3GVl
Qb5GVBGs0YIeYQU3hnTKe7abMUs/1DP8ZOtGInqmMuvhW0cGMIB3M/v2FzYk0sAv1VRkHebm1VWO
JVtFcsCf/HwaP/D3To9RqrARzgpiLWd80UBCwMW8ZUNakTR63ZWdtbbpYGfrlKXDdzlYVNLCcx+7
BJvyZJ3f31JgJDBehA2HgKzaOppluUn+DgZT/U7NeyYIzRIqYz3naL/bw/Jux351KjmOdW9/b8BV
+IWMW1nTmRJoA0S/7QzcvFrg5sqFwiDt3m6eS+uMavxfS6p38Gf3TpKfJIxBUaXm2FBVYVO3LSKh
az70zHW+oTXzdAudGTLN/UCdeJPebRIGrmlBdtX6+txARJkcrUplY5qhodns8oT98RvHjpQDSBog
SC8/aqD5HAjbT/w066e3DDJcDa2LiPbiHSu3ITuoP4hpG7wWvpSmxkpQDZyt5jQkJbQmv6BWlN2B
Qr+eJmx2Gm9/zNeh7pCRfhRkGyUxuVQcldL+jvBtyVTiOTCrltk3JV2n5RUI8Q+wpoGHbSBZ9DUN
4CnQxLbOCrOEGcyB2+2A3n5QKiqQzmMJ6Bc7IZw8ukdg64Lfd5mgl6f0e7rciFXTB01M1+JNKZN6
g3egJAyhgsT4PnOPWymOiEw7F152xgjz2AnxeYI5EB3BhvDwPZvW1vIpFqi4nIxPf4ujmveQqibu
HpTlYaCtSq687OaK+mUTnYWIjJfSluv40by5gfsTw270V8vhMjmxKhCo6+H+elkf6z5Jmi9DxW3y
wq9rodNXb09vGbmmNoBWrua/j+SATV/S986MNjTRhnCNwKOB3YOgZQDeHlYFj36tZS2GmvJIBOh5
4fLatPm/19k26q7+rqY2p6iV/G7hwKX3ElG2wuHPyea3khWzI40pBrOdp2uZLCZ0dTFn/c/KVT0N
/4bpPh+14SkkUVHShzmtbjTJUv6VWbmPX5vcG3AHEXvnUUVvnOtV/AnVbPreCqJY7wq6SU3Hqo0T
w3O9WTFR8Flgs4B8OOVkL3L3wxN1dxMAOu2aIs8oKs76CCQouS5W+av5hYARaAkiGp/XtrgSr6st
MCqDAOmpWHrcev9e9a/PlUOzGoy9abXNpzrin7FEcBb0+4k76xLPv072ynx76TV2PooUKZncWSkm
PiGXcBL6ne16dBdaqXGJp6MsGCVY+YefCEBhCp1ZL4PdxzR0HCZipY5+tAdC17hE/eqCkEidBVnq
N6BZ85/xTLjUCezx449iiwq5XKMEmi/ooIpf8H7qq6OfA6VKiRGx6R/bRvQb2UHyEMFa0Uu2Zf2v
HlOkh1DKOtd8P+l3phSBiaMgyrsAl50/l5FO8rr2hrAvwcaaEzXXToHH1e36uwNyOCrYvsnUCeNS
9ZNH7kVpjwH7ZjM7HPgVjBZR8ojJqupfJ+1kQsOF9iU2GD5vuqlcnDmwPVQTUA/YnYD6WJZ9/rCx
toIGw2iCTQz8Z25Jm+sj5JTbQyLj7JGiuJ1bSkH+8etDc1C6Anm6FrCt40rP012k9afsKNOdc/bu
zScwkTMWlkCOCrrNg4503HKMhF9qQtaZxIhdrMPtClG6YxhGGuo4yHRtHbmpLRWkguO8xNtnSvPP
m/ZFbwz6/EsBoguRD9xwqlJtwO5nZyf504G8DshrRdMIA0Nf36ytaflOXHFWs/rkp3kb26ocPlgD
YBJx0htHkkiObg88RgoKiLHhexkJYrGs266YSECuJehfn/2NiQurjuCLT3tQ8JmDnLG5N0kuqErW
4imskOO/2+GU0VM6WCgjojL/U19X2zu1HQRt4HPV19o/hUPxYBIL/eCiksP77x+A9B4h7w2H3+96
MjGNidv9EGGOGX/q6L76OGe29WGkObHq95FsM2LQK0wKEKfEsMrVGSP+ghzVJvXp1GN+DVj2jlR/
IYrihT3nRAUDW5oEgsxTL5IJ/FcokdNlABKye3qMtHTind3awDLfEJvnR0cT14uBZ2oP4fmV8JEv
RTd8KHnFYK9njlFSuWF4yVi6PL8Dzrn6jXVCBL5VOyYLtcQWHQT/mAnpmPqae8VIpIknnlz9c3W4
c+IrAsQgJtCQ90hNT2N4ThKqhGii4/Y/DIHqN7TlxjkFPL0SyRD2cwS+zi5BX+f+/XGCkNUPcUVn
3IlcdpZXEkmqc0pZ6rQob8GlKJOst2//G2SFWGWrUsgl6A4DlkXfmvccHMNDzpXsonE2kheFunOr
vxKWUkgfNLKicYbGd9zTqDOUka0t8K5uypDB30w2esI17cQg495VvbN2cfufFw6xar3hNE7pFftH
L/ZaCMj8+afnm2eajrqFxjjX+wNSrbFT3uL0RT9oO7rDEAxDCUNX8C3QRSe2zWV4cTplZLaG+Dva
S55L+BVh+JewNM4R6epkBOIhIrR0tYAdOLwyysARiVj/WBiS/w15aJlx4S1CYWhO7iOtjCgYezEl
kMqb/9t5fGctg16Rrtm6Qw0VWCIF4Iwmhvc1mGuDpw0aY2OZ/nsYvIfQa2XIGvw5Wc3QOW78URIQ
wH0QVo8KRnERjwYMCgClNabNaIpnRFzw2wM5XUpUZtXkhirT9LpL9c7IgrSdxEuFi1l3JTaWZKNc
6xoOzbaDUq6PmzBBl4/KckDCGoMMMvBdDZhlvB0/iOijlKiINg4ZzDLlZspP64hPm8xqN0C/ulwT
3PcQwb0cF/FbZujEapf88XDFhZLNLWeGMpqspLm+zo133GNgVHN4cSIa7X5eMvBiEa0mUgWNcUN9
jMZmH7Wt0+TAVIVb8P2iH3cE5HzyOq23aQ4iEoOxRULZuaM7Ie4Sm/j4Hr2yKbTztxY9FXSGIZnh
A8EcJlnfbWtZ29q5fbisaUawfdtKoqhkKqwOPiNeGNk2KHnwgTzqmEwVnI77gLCBG52gwqE5QczF
ez/JHIDSOsOPnOJOhzT4JoPWdk2T8TbWE2cr0/bqCjlCxEW4tc09GfXP0tQpAy3f2yThpKDveTie
hSeXHO/+99JLX+rbIGCOuD3pzogcrr9vt93LcdBbmFKzu3g++YXw2UiGe0f5sVG12TpPhSfMbgxu
Hh/ZFW8QkDdU7BVQjWALLVexKlADrTlba3vDajTJ5aJhwnUQ9AJkAtXB0w9Ygl6Qr2eX/taKWQRC
AQAmFbHZVf5HDCxtZQcstG0vjvuBYpZ+brB2xzudesK1iCr/VmVBdBghIgYQqF49UUjmvLvvFXZX
JIAoI4QZW3yCs3SKGz4MJWK6Aje6JeQjjhyuLuSF59WW5i+yQZR2/KtXDmdD+jP9fw0x7q86TeJJ
5MUa50d4QRTuutPNluv9moWUcI7dFA23FKzJY9FUxv4cYEwny1Ad9g/270OeuydyIvVmFp9GzIkr
G3+kWmdJmnmezbz1IoPFf/Zmv5TBdbxo2RQhC4Urra51pm62eXuaIzxuOWSvuXIlWWfZiDqvrrAr
RuXS82DckMQCfKRc6JtQByMwSltNo/GL4ooGt7mBOn30J6FbdoG9//Bd1xBIb4eOm9fo0vwzh6Ys
x4KfeUdCV445vPeziELkbGiQ5D/THHDllSKp91738mJilM60NJWouGkH8jznys/N20lmVLMCWr8F
jSVFicY9MS2WY7OI7ImPoch9Cv17nvoOwthekGofwQNM7YzVTsr4yuVmc5UUGHmeCbtKeA8LVwf8
0v8J+d3tqs7tjArtHzWY+Qzkh6QJvWR/WnoL10fhRMW9x3nkGfWyzwxYmE/jRCCUCnDQDvD0BgQc
iExml6X0FmGKic6ytBKmfC3GGc/OSHIQTssb9fR4yWUitxqJQPIAqGm1jBSFeEteH1LVE8t/upFs
v+oZYPo7PPhfMyArBAmxt69fj9UQzdKcc/bBJSCX5fr+z+yFQ4jfEmwyAGTZIXPEFL1HK2Qv0FCH
OV/0QlWUTZT5te5HdtTvOYkEJUuNxxam4o4qzugl8M43H4elMVIra0Gd1YsSmLVQnFWzOQjcYE8e
ZK8UvSZtHsDd1T51V7LcoKh05ipt/Aqxv17K+BJaOkQ0rTYUJA7eaCSmw+gpUaiUUc8SZe9htp9j
Lqv1pz27LBrUWJhMVz2YGxIVXzdx6f1ms5nIEHe572VGo1uuwhP6dMryjuxDUsx1G9Pp6gKkEi7+
5JqK+Hf4PA1fXzbT+CBn992R4Sw1pN7U3y2CIHc2wU4EG+IMdLvilhbmtQLyiVx3ELrlYTWcX4oE
aqJZZPfkWNpr1Vosns4VrcED1P+qJ/2vuaoHq+dOw2bPMBDheZG4d4TQsEjLsGe15QU4R6r2xa4x
AScG6zdQgP+F/PDIQHyncrGb2EaOBqYAZKHRDS8XM3LlLDG7RviYDU19k1tvb7jRFu2UnBhweLbC
sc3VOlR2SpjVO4gRp2pCvX1/E+BNfqT/pI+i6LUUZy2Vkx+G/UG3lpAOA7EjCklYgdnKscrjcY2O
TsqGCPLCxD2n4dsBpK4S8VEiwALh/njuIcOLR0oMvC0h3Q1b5wt8jiWaceMJd4J7/v/2SwYHmINR
/6DQVP8+NGrRLujM7DHGLW98YPh2snQoGtDDguVqiHgtUYMXYw9ydVAenpEP6KwYux/afu8KZZhv
ga7A+ESSSBG1OSNuMkXMunpSnCpBYJVujRsQC64x2dIqo9InpLyStQI03qrjSQrz2eYTYpUVp8JJ
4C8WnEAGrOjzh/st7xpNc0LD0QPl2wSYs5KX5MQdI+65qR/9mRp1IQSFWZNlna2wHffRdo6+NOGw
jiHcVifKgsVjtBQhRLxu7WBc4JBYhI8W0VP5HFtTtVKiQed3xRCkpYYT7yoMNxLfNal09STv8HqE
KG1J6QWyrH/FysLrECip49sIuHZt4ADW98qEK/fbxZCMahLfOQ2Xn/AxYxTdgBx2YXXVyQgdjZ1H
ZJbDvqIbmSuh6btkcgXuWgwikAyHZGMbLmyxOA5Iy8RKWaZALwmQXJLizbDFOoDS6y4MWUfcO5b9
aM6xMwWjT219jPzxNtLVdZbhUMOzmqzeht44FmXctLUB/HX8nd3eSnAHmCkSSoEVOnWtWJVQNe10
UHCIQlTBAclZde8lCvBgW0Bk0pWKz1ZZwfkMkZ392TfTgyQPLA+4NIEF9MxN7TwbAk9ZU6OUy5ky
2If9m6fXdpN5qFt/sarkvJzm7azDqxRs5Emmcmhz+wGpXAH8jpa1tk33uFQl3nJ/SGF73dP+ikHJ
ZgvIoq3SrDjkUYCWpYkjX3EXajWazBaKlmAu6A14jS7ahehFC+aBWVl7D0OA0z3ss4RD0KRthXfT
UYtUTUH8gvM22gBWNMZslanO6ik90e43w7czQJbiV2Ny7xa6j34lYoLrmVi5FXvyYcVTRH+2Yg4z
JaJ7wpstSY9XvFjKu+1ECDqr36JyuICCPeBN2fEwTBa6oBnEThx6NRBQQV7Zkq+Lc8RqROIgWxgS
60uTLtu5J1XmOJG8In5vtPIYT1X8Bw9tD4zhe49SAK6xYpHi55dLnkV2dor/yDk62xlkOIs/+NR8
mqa/Kv3KrNw+HKqe+nhQnS8sDLUw+RRczbajJnBR/X8KJH4KJ9ISZCTrtR0Bn1OLx6iA/8zKlRUr
TzQzIYbnJV/IuwgV+wlojvK+qLyDXM9U2rhac36eKr5Xn2+4M8iwMeImUPHvJZC9+PBg4xAR9cwn
gL53WjFR/wISFcR4KiABMNL2JOo0rmbCIgqZpPPC/Mz3F3irsq9RJjxtJY4F4ljl3QCT8ie2sRpI
boDTfsA9I5quRlnqc/RwlDEaVLbuQrxCxS3aE5CRh4/3uuJqs37tY9VRJvZBIPgV8NxW+vZ/vjiD
h6Xmvpa6iekkcYLYnRF9t9DjHpnn7enTpV7TFnx+fiR609HgI+IDDoRVTv0XdWIp6aabXXv8BunH
xkvi1LSnktMFsDS/l0Z39cL7cV633ZduEswWUqsPsE/Q7QUbMtA3wTzLcGswmhiF5RFqoke66Zrn
1ZYjAdcgmNdG3ACrlkLM1PoPRwOg5Wys1IJDtTa6zbeGL20DXC72pHHfdlJSDV3XhTAqKpRmQ3W+
oBeBO3fs/ZUk4To/SUBsssLD5l4e25f6TppgcThRvUMeDB46JjmKoQEGgAXPUJo9mqsbH/s6R+Oc
/hddkXX0FisatjqoUfrsAW/OIx7cnXPTKvzh537jznyxzCMFSS4Vwv7YjZmA8YqaGA+aMtj2LIoO
3ZYYORtUc5e/XEQ4/lZtgGAmOUGn4HwOucLOoE4k/86WlPLUlFqEXSZKBUcoaz3vlg5zVuLp5t2F
xUjcHOTaIyOr6FhdRuZaN7JyIZKfmoC4m/zRMvM0G4KS9/c8EBiCGz3ov8RFTTMtbjvkS6dV0lZf
dEi5PX8zh9CnzEOSOqIkIH1TdgQVWgMDsoYSNtt5zZhegTlBfv9ft5YY1BhMatH1W0Lw4Mk1LQzO
LT64njXtINOOEk6q6D88oWruwwzDHFlL7iGaGVB5XYLtLPmGt2yhMV6GY7GB13gI853AADDMSB6n
tp4eOH4XtyiA/IX9dKk/CNj9NzxugkvJujjj+Kl6Yp0f665GjcGz6yOsseK30jzK965payQ0wFN/
bFxVcpkjO2F4E4eeimo/+sKk3WOI8EMSEdBDTT0QkgypxtVoqVizpspXp0we/rUJ92MFh70K+V2/
OXqQ5ukJrWL9EGONiopFWVzCJ1FuOOrJSZO84kUiTUH8vLK4GVl6ihxuayZmtyNzJN80N4MVw49L
7Q87hjbVyKRLHOCblyDBmMtyAmGsuK8/aOxtl4Qe0wNVxC+q2MWtkcRllOfy53oGICIw6WdMX6z5
KDfTkP5isQdy1fDziHwSpYgTCpQSCrFqOmkzp6wh/djSB8n/PCLgQiteJsHYkqvsZ7xrSa2r3fl3
32odoacOVnGMPcDYstln7GD8SZfENb7/ak1VrSgZdElPe4UM/P8vD7tqi+d1QtYZlH/Ej5eoxAGY
q7ySMMFT/b4oaC5vueX/u2DNu6a9e4LaFYdFFsglUdMH6Wi4iMXDuNrn/i7a+ZwGG/Wry7bwupsX
Jz8Wf1qVqfs5019cxCDKXb7+YhKRo2IhuCjYRTg18PI7TD+1Pg9nezSXnA7X+ozY7ankGEL0N1n0
0mBMvVEnO71BQUdX5srLiswSX9kfLQJJMxAXeEB3jODlDNql57uEeH+crrD99F0N7DB4juc8Fbou
Mjh1PHekAyPk5okpv7II4QvVV88UPqjleCuT9c1Q8y5okUhIGvCl2vqiDhhrMfGQyVOp1OjZexOO
UO+B5oMzkL2iW1kSGFQ0B78of0WTnksF3mqxHZ0usRk0aobHeWTwhaV5SlSHurIoD0qv3ceEnOnW
/VXnUluVgleKqTzyZK+mAA2FdJySY9ib+rwzjLyf6vCNxlYZN3qCJloZVqry30ZyXG3NGX0AKC9Q
fqGALf6GUq2iVR/DD8kQIP8tdf2XlIEmW4kfyu+tHNoao94O4kkB7SM+slN5mxhVV6ydwWdXLk5+
Nuy9PCI028YGTVzc0a/rbi6IxTTXQO7QmBZMEu2bqNC/hkfGVPWPQzkWh1+hFVLrrxCKPA2S9Gcv
FVgDNHXcR7IErWuG36mrIjRbOr+XS3oG9UI2m5jqSW1REEc9rBx3KKt+5fC38rQgtvPI3aX0Le++
oJ8n06oUyrqcjZ76GqL68gmNJMeTnL4VD3CsDfoltOUckclEEGn+KYAGi0DOl7dJVf5nFS3nN3sC
Og6DjFPWq5y6V0GAZmy3htdKDlduWeraiixdJ9QeOgsZQYpCkdZSTpQ3unawyQI4zk+jFX94wRIN
7dJw+Hdwyh3OuWDHAK8qb0lZNYVP0jE4e+6Mura1LyBTSlyN6VzqQIs8BxVIp9eA9Z6glIiv8K+m
KefSDM5yuEWMS0CydB5wkvGSI9UH3rcIZoYnKB33hu/uwYEwU44+dbwpzT+6PMJHUMj4PMBaVZvd
yaoiFMbzum3ArnnVXMCGAvePvBB+1V5DJXU+RljSApdngCO8/9RMdjZYUH0xjow5bxgBQ+csh33G
S6jl2YhQcdPKzPQrGDth+fQgngE547CnLkh1EcZWDvwIiVmDekFTC/nFgASkNE7YwgQ7cTyutziy
TRrq8MdxZ7n4oJD9ecVuJJEgQ/5niNTKy2i7ztVpwrc7sZSKzb5ZRlS34yHef9CYiXHdRiX+cr79
kems6+nZTTiv4+M0oiRohynYwpPMvEvFWz7KnwlGocqszXrRvjl9UkRneWnIAkH8ZTb0RVp6AMI+
k6MZ70npSCjVS9l64DBuodrtlvfBcxotSeTy4NzQGfFh7geIPzgT6fJJKccLtVG6kP+ABWCgbCJE
UBt1H27/2YFPyWyR8Auh/vZ0z77yDp/fJ/9YRCL5nWH2ctARfDzea+Xoq9BKnLvEyUvHBznPh6MF
mFiec8bPvvCgWIwn8vbUUT/sf+xZkVX4HdqAd0jg6GfZ05PDRibOxS+9ZlBKXIKVzcTsu8aZYFtI
mlEqizrI+p8iEdE12Ro8N8LWekxf39yOEetUOMqzP3SiRCUd00WeNTtje6mGxP2xl6HgjWfBw8uf
zJxpkM51prHbOfCqeCsuIImJ3a3sHFkWg2GKC7L9WhcoNSGYC1EyzzdoUrrns1xLDXqY1+yS5ldn
N+L1s0I0vPLPiC+c9fqriE6mkffg6TkkZolYbuFE/Y/UsEQ17vAbOzSrGnZhdrog6WP84pzisXZr
xKoXat6TN+7XojTZp8M/AnQf2mbAruiHPs9Xh8kEsZ3YkzzXtQQ5kOd1VdGRYeuClK987xPaHD2I
uvQJL3vWtn0/0nRxQoWPQV4wfFl4BqtU3xXQjUD5zLdQijIdE4uwC97owags5QLldVfcMdlMvKuW
fRuDtHnenB/gRShNLZw+zoXOsZrKt+9wB/x1FSVae2rZyIs+NVpaIKLZ4jvU0iTRhSWOYvd6cJGM
yzPDrej8WmN2so/xEytXz2RXiSww3ZOCY4fDSMPN2CS3qGnq2Y6wsb+Ep0MkALOcQLx0xdiiN6Ij
pTfMOVMhxp6fCSRksVNLXNA7pPb8kJnMobPM6ICIAePZ/q6aqCvAVwFOEaonRoRjngBNtoF9k/qK
GOS40rlZKHp61K4xhhnSz31CSrNAXA/h5JWcBJYkQBs49xGcd89lbpqp08CJlWGquBjym8PZUo1g
+Fd4qYT56QN8E6di0oWKb8JIZOgVscAPSps06TJGKFxnxi9y1kGPkSu/y8xrNXf2x5ciftrlhBP8
9kcC5WADRQpjntL7LAj4X/OjA7ScENTKWXhwQAL0PH3ILmYeH0J1EW1+AjGJaQFXIOeG7J/awUva
NmalVkC+WucGCoh9KbO+teUZP8LgE+N1x09iChefzPdaTR36eZ9vIm4Lq6UKRMrYpLZQw/J+Wd1V
ByBT61WKuPHrAqeq5gGexdK4Nn9l9ugH1UZ7mVJmSO2g/uf5mBmhxrTvKrfoVAxg3mbDZh7EKPFN
9U7p2o58vdNC+LTN49Vo142UqWNq5cEsYw6Z+l+bLyyMQ2LPE7CiFtNPbDTpGuwZMnCelHh4CibQ
CTexvb0mKYKpJmIQeWPRlPhd2jLEcVExG/AzUk/lqbse5drVIpbVUHqym2DhfXkZHp80WoO2ddu+
pkQ0+U16Pefb/YwsAw/hNmjBLZNNY4khv0FAQcsEcn1z1nGZ/zmZr47lVpR/huUDwBNMwm59XNn2
Y7KwQB+a1OzVFHiqtKciEC2s0L4gLIEKdUcAN0GYcVixhBlYIcHvZzw82Q3ugiHg9DLwt0d5sZp6
ix9sLx2z5D8eeUBcMYLVmnAQgrXVW/hWTLcc4rLeYdXZFaW1+s6M5qTYKOSa2zYhm8EHvPDJ5HVV
HTzK/vesY1GgPRI4gXVX5OBGoG8Zqad8eW+cAIY2hEj01tnBIMK+DrmyGJ+nnRAtJpAGV4DJ2nLC
3W9jsj8Ysxd2SgoqntU2lwU/sUakyoGRYzUXR7btWIRt5M82pyE3Pyg5Ww8vqFdecUPXpi78SUEL
PAnbkxt2dH4RxmCUvabrarQKkLhfFKqqtqyYxRLplJQI+Td8Q/6484N0tdNmswq4I+4TAMsBaRON
W4jyX2GxarVJOBtI/JwkKFhVEpNvPphVaczBRnaZe2rWu5m4exLKGi3doPsCf6MXSPui+SWmPip7
XAiMJ4qIdq2mKLR+eKeuJDV2RXoLyG/bYW755Z0EamlqrCwBzCK61VEm9O9cOZspA7N9ewwnLkyZ
HQ7nobZyxuTeCg2p5IJA5iDUPDq6aiyqqDdhTGjCjhjoewrHXLWyASCE1SawlrWwCkssI8R1xk4U
bA+weLN0iXqYiSLx1aTwujlcwAQrPqqMF+tCYUjlj3FCq5ViWQ1fUSWQ0BeiajSgdLloKOYGsvbs
khWyl5+FMc2u00jhqZ02jQnfxIs1Tucnc1t1V7vRugexV3bMSst2hcGBOjqZJ52fxcxydOw6iaBY
Rz4g2t4WvsDZARHom1TifIqWXjCH10diVQoJx1p4q6k9ZqsOsn+n378+vbenAc8znYhpkaJy2nmE
2ntv8qMexkq9O0K4zGr2yfGzoMaFTWQTFGdQSgTZreCV7Bz6IL3Q45WgfhocWS9Z6/YdxUvi/7qW
ynCd6w/6ajYhk7p5w0qbzdoFGMNN0ASL3Oj6mi3m+T/bM31Q1Xqt0gBs9arWFcEz7He8dc9HnZDF
DclalYQfypJwc8RlfMfwiO1MfVVOdLF4aHt8LIA4AwQC3QMwdeDzBFtqAENbBYz6RVPd29xHQ4EB
1U2aqDD9XxR8eevnMRudW+URLoOYjk8yZU/Ij2lbXnjwLPGAsNWXAPHpnCX7L2wH0/2Z9t82HtEL
8UrD260wusTqY/ZyNrNMo9D9mO0sMmAqV5esQBYLrbMQCWl8gtxIfKa4lfVQqlbPSxGkfiOB8ymq
5CTqz+A4MVo+k+dLNoBfaelZAxlG6MdheBaQnNodj7mfDQ585ThpSU45BFQlp9Hs+VfDh20klbdA
DE9N+lROrCG/lrooPR1GIcZ24ZyKs1BqskFkDnpH6+tNhmEqpp7fKA1ywF5vJsiK7RbZ+wJGhho2
9AMxz1h2SeIQ494tUGwP0gfJ21BVyl6vVFz6JOfd/tyr9LyPeoFpSrkQbrBiajh1tm0uvF1dAGqW
gY6PqGmtzfLEWL0gjisLES/brnBA4DpwpPqY2SM074K4rS+pVibOvmcRtzsu5LlcWq/LwFZ1MZ04
nsvvtcG7Aa0uFVBc40OaaTuFOT3rz7Xsxt1A58sgcaa9qQhhUtmJ4l0dF7UAmyAkNI/63vcxnnRR
jKV6xU36XIrbDGJtIoqk4UH7z/c1Y7o/PQlT6hfYExN5oh4Omri3YNR8UPWfTRWjENrfh2C+r2Ls
PA73Qi2FRdybap9CJeTGILtb6NDXIJ4y1mYzuDAH29kfpp9TFikCJM/XnotC48Q+Mjc7caJVTSVR
to9HV+bW0n1rNh7TT1f+atUWt2CoxyNWCHYYpXf6g7TmKB7F0bn7afc+WTAzwuXj4F7i58mSAmy4
94GBJE4bC5z44WPIOYblpYuq6LybVyzy/L3nDpTngnqPDn5P1pcWLveQfKuY61OSC9pTP9bIwfqi
WAPaCOopmsf/0ffF26JpIyNg1LdJX8YQ++wV0FK/Sz+BxxotXmnZmpjqZnwXO30ncwyMdPoRaOUS
Sb1e3cbo22a7HUX4hDnP57LerGQsHH/UIGycrMoFd8w4IhYFNxDXs9WuCUpf+IjKNFgg/Wp7VJUK
lKVVJdLdeMCJDq29akr4Fox/33nZy91JivBMB6GistcdprofwTKxGyrNaderjzcnM5F7enTnnbu0
0g0EEfIlJ5wPBVzb2cQku/ZJnRyHX6KhzWn9RSCGMevJXeVzUy1D/l/culfUAqw/gEQievKsQZxr
ikWUovlYGrqQD65MM+sqdpCQtpDQ2GO1cMgGk0PfgNiksJDHA1d1kEQ1praTga0ko7XX0lB6+S02
HmysNoXVdf5kDOgPQ2R12SqB/wYo5fbDrnmX61EKWCYlOEf7uvp2c1C18YDHZNJG0Xl8bWmkBZDW
jCXlzFb6NC3agFFYSF59ptxy11tjmEeZcRu98lv3sUt6i/XjYs22nrzn1LX2NaNydz6aX7kSm05y
8y9onAowgsajxfZTUdTenS7ZLqeQoiRwpgE+Kvg/fSMfQ6G0CLx8L/GQofU9h8FirRvSos4WdVHl
aZciD0L+hhPYFz/psKOuGZaOzY4TQ1keHru40q7etQtAzIavrCFltNyq407QdVX9c/z/RmkC/8CK
YD2XLjAhtnvVAvJaLtqyC+AHJ50Y0eoeRr5gWI3M7mm1B69CuUFrdPwpkaiewIVPLlaiHxfow1BS
CdBplWr2/cy/FadpwpjH12jTh6JRcfX5f7oJmsXFX05SpIILSo3ZtGSfO6CTe84k7+9eUQ6QtkPc
DpTUrVEAkuZRQNz+qXv3BQ0sWH2bRerPIslRBUZIeeOTUXbgpSBax6PuM1h9vcPeZQBgO9xHOoac
jHv0pXwhKePBG5Wf9rjRAAwGYbZw7O7adr4hKLjq+b6HMGiD2y/i6AobpVml+kKZyHjvefEraWnB
QIrF9oSE30v0EiPw9ilvtD+r5zBNpZLQcnk93zMqnqqUDRiGIkTKt+ks5ZqhT8DKpqQTEeYssTIX
F9aBwub5iu9THOoKhnDleSRViPiJ8usCNO6+tNjlGX97IdzLkBvG0hiUBRBXy1D1iItyruBfOQHI
OAMSCszfDLNBfF7ww2kUWLHGVkrkvlcFG3TZFr4mbJvuuKkBosf0HtSzaLa1ivB0J89zGy6UeiO+
vyHEkKswKNodZf/yhBWXlgSatyDqfgZ1PUHJjfS+WcUp/d/9vevLRMdgUT+4KePX2xF7b9OUrq3T
pxMgu3d0pvOMkKvxkZfsUvjbBINO9dh3fgNXPmbI4h96B7DXZKs/mymAOmU8ZOY+3tsfAu7+c3b+
L83jD5XzZnQ2F5Ofwte0t41XmWIQjqVpzwN+Cwe1liKbm3EeyuaqZVpV7ZFHrGpgCdLc1SyR6qEI
EZH0/0R2fTNXxIiRvG1p5cVUbYw6PpJwFAISh/pKiwjYxovo1UZuaCwRk4r0yRPI788Zi+xzfIoY
mkT0CNJGdIphV/Aw03L5Bo8XKXFl6FAKoWaB2CC3XIQWQus3BkfgfeL1HtdP5mVdJ5pvPheaXD3x
m2AN+NhCECgaPbAngDNmrfrUj66JT+hYRLBLaOrCOZZWBsL+jYJVVyW0AxZ6EC0veZ4fUqtdIhx0
InXUmnm8PLpMrIyGskjRygZFmKgEsYCDUqSEeTjkS9a1KCtIqE5u1uj4sQ0PfWqAlrbhOtiSc7xe
b5bqK+lvBSlj5NyynUyG9AMRNb7SAZhPySuoPVB7/Xohcc0W/sYTNWlpY2ISSkfTFB6rzrI5uk17
25kd5vOa5TVBr3iScIvvkasgZ2RCL4UhVzw3WD/GzN+VJUiDk1vsGvmQmuWcxvUo8SdGltknzsGq
qxgpEFcdG8EwCg5220OD2Ae3qYc4SLei24MvyOLkY6SHY9mOjxaq+Q8omHOS1iq+NcnCkmA7WYxG
ELl+l+YMAkN0pvv/up/G+7C4Z98kj/f4fcZpXqrNVDsREkf74kxLqOQs1Z7jUqO1qxbzw0x7ff9H
r1x7s/bvT4sgEJ6m4YHA0gS9CcH7QcYQP4w7HDpl7hYVRGzmYi/CdhjnOkaB72WfgbB9ZCECgrnL
AZd/ANkZ1HVVG+8zRQXN8y6kZ2e5MTicOYas6wQ/kd3ESafMXMjCc21f3O2R3UdvwMSBP4+VFW0z
HpRDakiuEvNn90Oymtd7ZGuVy64Dn4gTtYJyTqzPA5TZLGDm1jAA/BDmvfZQ6Gvt5qCZKY0+34mw
QQ5Mn1ocpMUFHUQAiYxZFFZGoZMPRqqoUpWZwjrpHiHiMBNxvWbVb+tF9Y6ZSMWHL0CUUM9BCXwt
xajW6NcZKX+5seh+9Fa095MRRJ26BcNIAvGjSXJrjLhHTmuVS9RMDIbTFFiqFSTi3lLb3z1pbouW
qVtrWBLtSrxQx+AchvUMkdcN3GaS572uh11/Xxam5NcJCivjmDCjKo24iII7rqyg5jlLZVLRPI9t
NHEsEAhvUkKFFVwF5wJzZmn/+qk7iv2WlpHAdJm7qF8v4Oi9wGO5q5w7kNHEI+rFb3jeLSdKdoYQ
fD55RWNxMS7+Yr1h3pxvQjUpRHnnIbH0xnHLYDQj5wBRwd9yPPZPQHhBKKPDspkF9vwanhABmLRn
O9Pl7hLpFtRlKphqur19opeyJZDZmQiQiYbg+UqWXmr6HXRahfCXg67LoOPaQRhKKRQS8eo0aDxs
VIKLSOroD513fNzA4pNHa6Dc8zPgYSpuBgQy0XeiGKRXAcGu0q6njWZ/F/J0IYjNoLID81erWWku
l8p73i4jt0+L8JNqsnQQg7RBV5avgXbCUaZFQdMdsklpljIE9zS5G7z5GVcTKuWSbqQBsZ3uzd57
JXuEc4JrlPuFHVPJeIFH296I+kFXyxLC0RqXX89z8YQXjAaE+FIzO/7nsfRWHJGHcfEKysr51zMs
WVIlpevnKJy2SXm3IyRrZHnmY18iI+O1Uqvi0+AfyiYEOWQ1jUKeZhxRNU4+wJuHPxlkZcG9NbxV
SUWs0ZERNQRLk3WD5FXaDQDj7MeBIR/+KnGyCPinFx89FhB9KWUch5fHQuz56OSNnZoEcjbztD8p
UbZ9ZhTXyrqJuAGCXj5WQVwCnD9mG+pm/6N5dbHFiq1j01tcl6w7Y0WGRFzvfZsmMTD7xUQdkfyr
hbSKyEzURISXPGiBorQlMeW8J0nei0/qHlhMJdQlSGr3GqdIeKjFKP0qs1y++YlorP4BZxhqDQxN
89fnICg5fWkLMqHxXiYBxyLr2cPoxVG0B9oIZ6QSZQncAdUjvnbGfkGibzhafaVodt4P5hfJ4uVM
0N5nsb0d7xbkVyTJowcec0KiXKXd6wu5MW2fmfAqLKuKvxiA22ZvsjI8HULahiJNkBpMnXOuMJhC
nVUo4prLxqfxOUlaLuyq8GXxTZaxQqAjySvPGt/dSHnMFhkgxZPIUZjJVR/duCDf/1dwa5FHmTNk
bpGbRHYUXcC/6SkHJmmmgQFDrC/UodD4cY1Bwm7YWnBmMjhAF3KQE/iyPacoQWY5evSkbtPv31Zx
CDfGrSD8lc/4PjWNQdL4t/4veNVRw0KytjJ32dwT2S0hk1lUeZ4DtsNSul2eC2nxxtsgXH9Q1odi
P0FRHsNuz/MDRy3bB/WmQhiEqNJIIOEu0Ol80yWVn4laNiuvi0DG4SKvS2Z9lYGGal0xZVE/AEpL
f43Kcjx6HGkNCSG2hYfRMiLSytDKqW/NqOjvrj6hOZb7jy1cZKH9k5GLqw1Xc45nOcTUZc8rbCnL
J3t8FP4izx5nSu7gIJJVScn9uvvkFri1ABvC3wirueYOlH3+04yoaFAG6NKhoSjmSAfpQNq+9Ozg
7G5eni+koEf2XboBM4v4XKsmVLYBRbjvul02qbCefuF0y0WfdUSSIQOKrskGaXT4imvu/aLC6hYl
m8ZVVZWvPyOpyxwa7uh5rOSqlgfvQFniK9Zjx/P7XpMzdpaq55RhWZu2TXOWkhga9ZzhcOig1tbA
gg6ACJqy/r8gsdYrS3lw3LoOt3nc+RqE2W6FSg5druupnAf9IC528ABDtfy/o5f03NhXtrxTVa5V
CmH5dR0zZDjy9q3yW3XlmvsCwLvTZD+Smvp5qcO2g3WjGlEfSvLEBp8epG02qdzNRFpvpbTjIOPi
ftkK005C2mZh5JWOUOh4Prd+iJDyZ9f/EqqigPsOx+q3oKlC0kmcUjrwqjCtdfkGreMmH1pKplXN
U/n+2e+PYbGpCIduPXls4DxWfiYGPsVcDowE4sivTQ6koldbJoNKEwI4BGAs5yAXI9q/aZfvluzw
pxc8XwC39JXDvRWquUF6E6y3UaVY6HoR0G505Y6Ru7YFOQH9BlWCQxgEs3aFbaBQ0c19Bx07XbtJ
L0Jt+FhExIO5scjUFIbs/yZE8TnfeRFkULy8blQSjxJy3RBONrbzmtPNGFQ7QfYdo6yPZcDmmnqF
fMZmE8/B1oXdZMRAaD3iiLH7VDipufpYkv8NaDB0n8kz5IXxg/LD1ps4FiWvXEWsZBokjcMJL5Ap
V+ic87QhAR94cxuifML3Hm+E8BKuuTAS/MqZkrVbFwf6ED1TNZfUKGoK5jSQIahcVN/JkdrXrXhD
Gk4nz6r56GtY/cvZy9BzgX2CLS9sMcSd9zF4+2de/l92yvcpTHlIM0J8A+CU1HBKtsh5t2qeOMXO
qCq9kNPal5qwrLLn7nMUuGQnR3ViafDARCpE8zjELQvMOfjG/LCcAXDf5oAO2hJ4BZfwmAM3nkky
sNo+ytJ7s0VowGOYhiFe9rntGVC0rlM+c8cZ3ojHxtAfRVAV6g3MPM1YW7gDxrvJe3FA1WxQtPXW
ZQuD8MWxKjZvmWMy7C5gV+3snnKgjmIjOBnkFRu1UfaSTG29WWPZRpBeA5NKDCEmRfOC0yPmrzSq
EnF1/JqjT5CEWcKOt0nXVVFRfr/js9IvGBJH2tR7yFL8Tqkjvf2GOiVthAoHvthVFQdgP/kP9lJn
LqD9kUBx7MCCBcFWfwkJGk42ng9r+R1a9aWX13TPBtKqLmUnIrD2p3Yq8SpbqMT7UUhMO/2oMxTX
YlEyD0lm5URoOSYPCfJdlOM/JuRlbp9VyIoaX+ZZ8lIKfuxSWG3ceg/8NeiYB9DzbZuwLTEr5JG0
MT/Pe/7qbsUkbbFFWCtrlPICxBOoyD4XFtuCqUeQcd3L8uSt60x7CRqfRrKjaAIw+wX2XaPjzP5G
M6o1xD0F3tVF2mXZ/WoL1AvLALaEodqdwLkozdNTjE0xblRSMm2HsG7y66XFyxK2EU61XXmhI33V
ByfEVbPdy1vRGtb06hX0TEm2vp0WcIo9gMQnUeV8hIW0MOVaTBGB2XeyWKBcKbYQuh5irkFHcTvK
bD5Vr0TaBtrnh5tv1Xld621z7ReWWCRCJARa4O4GusJm4Pz7snmylOekA7wFhq012B2Ku6/+0lwm
h4UPJ7F66Jtq5zW5lovoqUEGhJar2Ayj0WUCCRVgNT1ozt8WzfXhO8Ys8oqMSVdcn7Ei0HybbBL9
/v83jhhE+g02FRnGYZGYX9LBUVJVlP+F8VvidsVZf8Wi3YAPN9egLmuBdUtk5q9BYN++X4jaZmhO
tidz0Xq2Jwt7IIsbdHa2O6IlH/ERy+akALTnKMUi6lM7Q414waiiiVItEXNkZnaMOnBYtTBcz1af
986dZ5l36XDFWEfF6XxXwlx3O/QhJ7ljHG5dIgCDDdxNcKDuh9rr1jiFIUQO2ZVOOP2HyVlhesgb
TiF+XpGCRF+VvUGmOavC8eC6lC9ZeUjUv08sc49URjk0Bf5vp8tqbgBKOpYk0laDbqUAhTsTembJ
wTcH0fdm5DrF8XiXyQ9DAQjZzgfUzRDQN22eCAsjBPUrSoykULD73hhLWW9B7Rc9978VgPiWk4lC
EIJiDt6EXclT3XoWeaGWcVQQsQnX/7SBS3RKxdee+RZhyojUIgtJUmgAzcA4g1SMQYjuJZGQ0EKq
hhNw2BPpesZbUChWC3ycoWAG1pNhW95d/yRyv8r9xK5xrCBx+x+ACyjYflYCTBhqfIMAxMTk39YI
RpZxC8skDJP052aldpUihK6epUtZ4OevjiukuA7vFauBW9dV5Lp6lqvLFXWgZuNvpmCsxJNVLQS4
m3T/NyQYJvEGzLuu2ufVhH748ZiRF0hTg4rUbk4RWmS/3TGP1FPNyBbljAW4jaYP2b5/JCaf3y46
pDdWpjx+pHltfWQUlOTSlYeozLYqx7pRLVauVJf/bEmgJt21OvbDiuc4eqJzZNH1/ZRoLovkBJOY
JM7RrEMJkc6NqZ4oDQsoLdIcErfJXb/HoVEtU56g8cl4vrMfcLUwqJqwBxVZMQQAalgxvLdIcFw9
ej17q8b7TdphKZCubd5lfX6uuETxf6ysp5Q666pwUNM4mWG5mcrrHaToe/HOSu0MY/WPJSq6hXFW
IIwnv0xeciM3mvFdXy81W4Ns6s4gqSa8Y9WeUkBMBFbJAKqzP/rmID6EnHg0z6BmFeACfLMDqmGk
esqilTQIXgpzE/2Dx+rfww2ZpGTcsiFmSAhbUkCzqvgEVCUUkxxXNY4v9iUBnKS6w/Y6PkPvCR3A
ZqGMChZOePlLU2nEG64GGhEuqRE7T7AMPfXFu8TP2D0ulj5kiu2RhVuvVGaBwTuJx3+O8cFykCHn
NxfoqmhoX50CQ7KWVht+smwPtZf3zNJEz8shM2A78TPG+mtkvqILqwhYbxEOykysWssOFGzYv67w
uu5sio4FhMESFduYPProRWupa87Rq8RH1hIEhOVIbP7ilF4lPLOxAi8kpgnfxaSvQXn1oB6fQ4X7
m5nvDeoPZ16IV2HQSICmYKT4vHebk03GLHIOZ2vAabN+LBznxi8qKZAQWAFs6H62uYpP0ftCDcDb
c3hFCWfSWdnB0T9ABvhdKQNSiMMrhPGiohMKMPfucQUzaJzsjc3VrSaMvIsrNNNdkE9BlGmcqD55
DX2YQtW6iEvUJrZ1jzS06a6giqb296992O5ejqfE5DVIoYYYQeEvlJPMeHSXutkNuVyLxae165P8
PNnzUfZhpeg/3PjXnL4rrJ8o0G3wc/Ow4vcNQf0VYvFzptVAbk2nUen6ZCzfVF88RMEEy2WQHr4v
pohoqgI1Bfdr7l3DnaVJIFAM2sVrN//FfsGzBQ/0kqhGYEkHL6x1UarwEAZAz8Gw7AG5zW2uM4vM
cOEDVRNsUvJ1bFKpFvikn7MUCuHyxHTnAT4Dm0yyHfVyzo2I2VjfcMVSQIiUDJMwyH2bziBc2mHW
2hExSSUbPZFsrfh/+57ZODJu81cgpq9c6XHYEC5pwfNJa0X9+U7CYlZ23kF+v7Bh0aSWLBoGGj6V
OO8kxC0QL2gCf8hhf2M60p/Qf6k+2FapYv/pOgmKgX5DW5bTIJg2NpfaYKNM5DKOaClzbTazOqsA
B9l+UHr4fdov4viOFxHop9knNO8CauTn98Clqxz4d4urZxS2cnwzYSbHBjwB2MVM/Kz9+vM6e9J5
Ia/mIlfhMZoY5f7rd/WfSxydjV6k/bfpSOrauObJ0ghnGNOy1u/s5vWgytdrQ1ir4++TID2shgk0
mm+6l5uHS+fzQXcQLv5b3r6RL47UVA93UIWuNPRlafcCmDUsn9DU04WOr24qRiW49iGsq4pFZZTC
3/eTq2BoJQ9x4W/j85jFXpykv0yJfMbvE/rF66tb8gXKh7R7FN38u1dWsqF48D09Ep8GZloSHpYa
9UWL3EPGR4oBfmwOd4Xj6fziDj+mdrjM99AqwgQ7PhdMxeDNKlLZG2jOZo9OVJIedTaxUlo5RMvF
9VTLvTNF9LbU0kiuRy3i3+KS+D9ooqYax9kvjSJdLQKisLgJRkaxFZ0q0zVUQgjHkG3kPrBD4ro/
XmitneTH4Z9/Md+bCRzX6f036I/El0VDO1JMzHRY7wbu71nraGpClXlZTJ06z5o0FruI9vy8wuDN
CWTsZQmMK8cS/zWtYI17LQUspEJsJ9e+tVKo4u9xSHqSQPYsclIlRyRkkMXeNjNpVlSzv2FrWCKj
9PNekPWqtGp89xMvW4S42jmnllEyvxKFI+G9JJez0iUeU/LPuJ48/kZ0WqTNR3eMYgR1sjDV2/xJ
o05RGy/uTp1NGQ3RDWuNLscUjCrHk5YDay6PfvZt8plrwMdF0psL8Bmh32926VkgJL+Q8nQeif4Z
UK93T/Lvoc3I6rwocxBo1tBa0+QEaaLWJaaKbkEE5OPKFY7R97ZE1MlXhDa3PIgquQnimvMPs0pi
z0mNCCRz5HtXNAG12uMQ85yXPyg1RFsJ79OjzJMKfzivKyYO9aX5+OJKgXHzc9a+gpAP6WDovdnw
RygyaaDzmx3y1rzr3TJy9/HSx+mBlwXFL5J8NqAAyVDIDjwwFKQWidFn+uOc+rJrd2eLKJyU3Xko
wcz7Ya3ls4c5qjpgFjnuem6Sd6v92ZESqAeJvBrU7yYwajVi+kUMyG6p4hPfFNgNhv5hbJLdQh8a
/7E3Y7dkbYMDmBDZ5sDPPd5ycAfs+VvFaSoAMCdNOA8MAx6MJIuRN8UO3VjP83o2pTm7FcI9Wg7X
aWqbtJF66ZeLyRKKhZsF3rhQ7pSKTMBa25lHLXzFKbXEPHn/mLdNrkDkZrKQOSvt8+hVua198Bdo
cttR7Y79AQXAKNI119hJQTpzWV0R4xPv/1p8JmsOP5g6DVDxMJe6Ew8pYxVESEEnHECnI3unIICC
/JFSFbhMXkE0BBfZWREm2QNUzPZlNddq/a9uMoG7eepWMkYW1/XuPAVmKBudeVSO4e6glv1JlPYg
Z5grMscPNWXfL0/yt77TCV6X7LS9vswn+Gk4XzFx2D4oLLLIBCwvKne2qhdUUkiLEABGvTpHQHka
2pBaJ9aAlfo3PVchrbLBzlsU5r5QSG7tYRYo0/CvYCz1eJnKgsbqgF/pHfHPJm/kL329raF/h4qH
Xuow5EUuO3FwAV6kapaB9wmSYeMlkP8NjXH89cfQyJTguSpG/JYPeWIhKhJRy0zX/aB6yCaqMWbf
7A3Z8OIdgPxOrtIdsOLirk+41Oaby4CQzOHUaaBMJ1J8d3GkdMyq6xktU/C7bwHkBhIWgjiPUmwj
INalwscIo3TFY29EjVzl/K5xvHLBSUmJFDoeWOtIiRs+Euh19B+J5t0f30+g21Pb2DpUJ6RPI8U2
k20WoX+FMQn2EYH1EqM81z/fikwgdb/EXEC6ZDTfVAoKkk13JdoptW9E2UnlCdjqFHdhajhV6yCC
oiYkyplfh+oeoJ4ArRF/PovDEEDuRnnUOIuvjKjzdz0gT/2ESWrexZSayabuBXtl1xGi7uucWZcM
akOHAT2872Xs3FlAs1aWg35S0UZpcGrExtXmUl4/sx14cKWjTzN3GWBQcUpH3MLGOsKXfx0de1e/
j2lq/TcX9L7g5llY4E96cSIj4qvjdZ1L6YaGPpOrnhLhReOwPUVS9e2XPpEcWJoUEZyUX5ZakHJA
Uo09axX+EqJBRrMEMbEKWmMIlGzN9XktcSiQGojuJFFvlP6ZhP3k38nmgQdQoBHERfyijLSbLTP6
LiCiZXi0x2yMCvseQ6OjZGJRR7kv/zaC/kLx0r5s0ReLNMyOHFUPu7H7NrYxlOfhwJCdxBZ3hDkg
KHTebRIk7EpDNGzO0Fn6Cj/bxn2pRzYrCtWcd1TB/9tBfJCxOvbwDptlC3dWgiEafFOymrS6CLbO
TJPZACkSDwPITlJGk4a72zXagIjPdBZfG4fVyqMV09egTeAbE357dWFyAIb8mRROHVYYzzXsoj+x
1b9thJROXeDJOUO/lffkEoELA32lUwyw/+2hzsXwSR17QKwFV2vsyZa7y0zaYPsj6LP4ChMylsoP
PaJJl+F5VYByD57UiI8SsXoi8OWmuIWaa8sS5VQVcagDNDx08lZJ7i//FIacD8vBr48iJuCSllka
KvqZ6WbhnhSLnokUVrc0nK1Fz38eI60uY8vsnkR/1DuSrKPKGA0u+7gvj9CrvLXuhHCzDpbraa0S
8J2srBvVldS7ibT36karO5W4EAKCYf3xHYvp6fKuieRSTf9eJDADvsBwLPdI1OOQueyr4iFEAztS
DcRY0+YG09qKGmkD/MOOa0puRuSmCV8TsQD9p0GTvHQPhL3VHKKRqCklhNaQctAqPtBLRkmJOEdt
xFU+E7zGORsqMKonJlyiT4rf7xyIG9YHmcXV99XkGz4y3V5cCXQLG2dU0e8k0/rknZgs7eSzux9O
1PBWJAMwhqoUuVgt9hYnGfHKbktzn2a6/lgy0zcGNGhDIz6zTr2eiWt+yEwdLPcacmt1Cnt6tY/V
wTf7HRg/N0dzJ3TiIoTvju8ri1/0m/TRVhodgMsWe3KXJMXYwhQ7dMSCNka1JBmwXyEDeuUob82m
fBolD1oB/oEtMcblaxpBYBbfDvyQHTl/P4tcf1O3gq1EOBnaE7ER4rX/5T8i9cJNuohHflQX17DX
tx+IzDowFQZjrumz/5wt7mA/30hk8F0kR5+wWxQ3WXs/RQAWmUSOvh3VHXlVYWdirqN8RJoCuiEM
rv00zd2kAWrMSygq6mM6Tzu84riM0mg6BEirRM9meX8gPN200HtDmvzzd84dGekTukCxq5vIRouj
PGD4kIQ0HNlqGegBtTiwjdVxv+JXh2SxEFY8+shCuPh9EK1kTKVqBL/12XMDoTfdl09+vNsAFULs
ciGwvEC1nkfmDgs8ml3JLJDW8a69noR7aBWzHc4x0gC4g/kuMsn1AEm38QKMcIaiQw5MmRAobTgo
0B1191HdQXuAxDo7zWwMR4dKuQFEsG6rnqSH8wkRhq7ygQeTCRFNxzU6C6WaBfRkjnBvJTp3TJMO
H+wM7IWTMgMpwxGGP+uLLEhwe4L3HaPSgY0P3KN3SqYyeeqMMU9Z/p8Z8Z6m0uFZ41zN22CQOxY4
HeS6l8EkAzPgzqxO30l+kyqDrnR+mibWZeyz2hyC9KP0i3vG+YKRAfE4s5zVYb854eenJlJ9hhw/
0IRVSyQr0O8VuY9P3vttwbloohYOD9XJR2mVXKLTq+cKH+kSJIgcACcv3TPOr9zMr/Oa+dRh1aiN
cePuTdgdXVvUGyeNu7k5WnarFPPE1zc0hIlsOETPTlEV8OMZjFvK4TZLV1blrERUt8pytKAVkhwk
uviCIzaTUox0wWHxdE1ZRVTr2OFSrN1qRWgWBk9BidIAbR1iuqtp49YzzppJcg5aRKX2DXUcJje0
aj+yYagL+q5jWkS2PZyujKcjG8Kj9qeg5yi3c9mby2ULXz9St8lcaPRMItUQzJpRnl3yQ5A+01EU
iboRC0GyCjm/g1876DM3HsRZ0OTOTU9Y4O9+UYRd4jrGN0hN7ssUYWfeKJD3aMsE9DWYMuS7XUOZ
HoZYytR8uq2BQnHp8uRgSIBF4eRvTB6VNszhGpnj2TzPFVvtDyM6K0W79BI8FA//F/csWyBwgbM+
DlUHm8FZBvo4DfS4zPJEZdyKqlSqkozVfTr6Ao1ZwBuFdXq0q++OOViSbJnDIpbQpzmOKf4/h2Y+
L/nGHn1tt1pytoefpkhvbvw7IF9ufzcaOKCzPcVbg94OIZOs191D7yXtvfoQlDOCa3M2BHyxl7oV
w7ce//RNixR8ijx3kVdy9BzSategQa0nUqAbBeejPX5SAGD9sy9dXoC8CoW4N8qRCgd2FhSQZHip
1lGJVer0L6KZVUX0o+2xcWlf1sAsSXYz+1yIxWVeuH1GMk1iRZoQiZ+xmkpx4xdEJS9GrKjLWHx5
ErybowpoURGJAm/LsDFsh1MTnVC1s1G8ysLS6GCo9t+35QgLSW0RlLJa+bdUM/FS2u4CVfrhMaZK
TuUJrFieUWcYIorr1Ee2UgNdlN0rikuYmwlCFF7ywH16k0Z3GUMpfDtdYnnR6DfTO2JHKiqjgv7/
WUR7I06wOjNxEiOkAFi7Z4coTnBinc6NDVCl5orzVWr2b6/vYV3fQAXH/uma7hmxM8k8SfqWoe1S
q5e8op1dFeCv2ImvMOPxasGwXJxGzem4DwtkFAy76qQMFfc2wjaTtbpzTPgsCNNUdszp3AnOod/z
eL7QDExjxW1NcJ6l0Ckyw8P69/a+kOEnfaDBU4VY3qay5D9GoQvYGj6lj5MaIaRIefqAiOXhlT2Q
OAnbRRuKjFMADTdoOZ/d2qTYGmMPGhk8U2CdVYHKbvT4Qb7cM72+Nen2a+YOntbk7D6oJKzXWXaH
mmVAFjN0qHhN3IY7BYGeW2u12+u3X4Xdu3LGQpOWUsQlGcqCdyTKq3d3aB42wlsfRLNw7P7WJpZZ
7gA2VUrkO33BhBfMI5bW1WDmJlBTLXySYdXTHJm5lB2+RX8wbNtHftwVmoczdoMbod9T5n1W0HE6
WwJmiXkKq9wtua28T9JGrT7mUd3pGQahVcxHMARtqoyB9rRwlKxLmC3zhK7yJggkKOL6IQ/rya6l
2hlf1EiUGXtLALrrNVHLwyMT9IZtR+L2UcnOiUToH3ItN9Ia12VTQFDLOtuiuRTl4WhbEktWG0h8
Txvlk0R4OsaQPmKT9A2rJE99LM0qoz3KSHsomN0d6v122dacLfYFh08I+Om17nLeEsTfbUgtVoNX
10cEnspDQnnLLF4M80/TIcK/6BRKwTmlqnamHB9dpoq61EgIXGg3xBK6P+ya473S7Lzq7/ZHdP10
QA8yIUydYd78vvqr/m0Ixx0IncCYAgQf7r7QwzGPHMstucA3p7tz+rUZYhsdOvq1OcDUHstYsgqp
rYJUxCMaRWybMcgB+oRvTR6A9WhlQp1H3o2D/ny3CAkin95U7dvyLKzgQ9JcIdXWy6t4acTCaWgr
jw1GuBX1IJEv99kI36WNKbPvFxmXfN/NA9s9h8YbTgKy23qjhfI/4HDbSnxqGXsobcgYGLXm8G7R
iVEpey4PEC0jUjLOaBIY/ThV0vBO+g1WDd/6VWrty/XbpD2R2UdVI/x0ICloDK6Rl/7ypR0fl1he
o58wGbGjT4FNAOEcw3bQ1AxVChLTcC6ZMcwMhEXmKo9OS30yy76BTebPs51g2UdddYEpzC94DNp4
16pad1wtTSgLlmKdU/HxU0eR1QmfxmJxalGBLakMo9t1svCByK6GrN/Ib/kSVeBPoaYbROR4k3wp
X1zKNb74w/KDJKTQ6akntFbwXGguvuKvUJf4rAxc65F/QhqFloz2B504KnYNvJKKzgrUt9641Dkx
mBV5CuCmH61QaR2830wZf/UvLHK4xOdqyXCdq+kET7Dd+zIQlgVyohvXizq+aeiH1ocPgiyknitj
0pdASPh7miDmDRndbDFaau8piL2zVc8nmb5zVcFuS/hbU1jLjus13asB+CGnm9v5CimPrnutlzRy
h/X2C7gxCmLqnZectqM1+IGPp5F5C0JxPeqW5FcpNztf81EH31gBlNYoOLlHzwWbT0jRLnMvkQim
dbALmQzjrceBsq/0afyKH29/2EUHZMDiJlc/KRkrpov939H7E6LOY0pAZTY8oZbsm5kjop16QyRi
Wmx1Fprf2V5QtsIHIUpCCRJ8E0cxTz74yo3e9pcISmcM7rUrM0QmuevEWBLfaC08CdzyL0W+6hiH
qAUEvXBZJjCOHaYuhyZMhRnLF3GYoLOhlrjXDc20eZ3gRZA1yS10s3FIOILP5Vw0ol1XOTyQSgRN
+qLhTjPvaUC/lwWrm/TXa5L2paOELXBvI06A1lqTzdiJdfGYz/N0sgNMMs4Fvrz/rEJlbRUrAhtV
r+K9DzYZMd1eiuPbmcK4FkrVWkJV+aYYAD8RpZ4dGIjet/DfPSNgxdfMZbrxcCKA7WRtzwuWOdXG
5/5yUyYAgab/V3+3lMB4dh771V/XMo1uEogRw7W/v+h2MWsyNUbeuRKawremDnWATJqNVD8p+ac4
CRnNUQjGMB8FVsPv+jNmhn8vcS8UdWIy45CdPR3FGpYPmADofj68BbnGCppLHU7NGpXAJCMrKU5e
q9y7meKqhIoDcpLZrCwSAJxogQd71sDv0E2kgIbMYV5O6OzymOfskL9U7Fro1lJwmZuBpkiXE7Wr
aY7svo+B4S8LFiPglgVPVwPWfuBlHcvUEdeQfMGhAEUt2FGi1hoPqQG03fxuGKH3ytHfnMQjiJae
c1TuMq8QeMSpsLeC6tRHSOo1yNyC5BzuLTeT2PvTIejKJdB0T3sjVO/Fh91IVbl3Sk3ZYSMAusyt
xSSTNX11iJ1Gah0tG8ZX5RFexo9fttNZx6WdFwcZBA6UG+TvXvH5auuCA6eUFkAcqdsI5ZnAEKIq
+AP7Bn7E5RKHyrqvdncUPwYA9m+f8RLk8BExK2tUEBU2QMkEOdvyc+8DXWXCZZQo4MTIXxuPVAYa
17cefSNSaGhIwGxh6Yj89hqyJwbzj4UHxDWE3M5l5OsFx+2PgZ4CGObqXzrEq0yWRpZXa9vBqDNz
3Dt9O3T87f/GIarMpztCUsP+wsxXFUdLpWRI/4H1cZgFhHhcAx/2koKYBD4rmzP49Yx2zejAoMYr
Z2Li9/Yae1HGq54F+dqjZ1ZJKexKY1HT+3UdeHSva3w6mEakklxsfgvc+HFY0THljNIZtSHEuR1m
7aE/67k5ve2A8sWrTb2wb0tEyMu1llwdloyj1Y6APTzVM6dpB+P7DK0WRzmoGqtAqmcmhH3Leb6/
JfFZ3PIc8RrQC2zShr+K1LiuQRGiJMO8q1xu2sXF6l9WNbOUPxtySvuzNnOjOJ6z6ddolAVy6KBT
tw4J6FvWumm8SsrTtu6B94uTgrsGWVNC3mgHjNswPbLivEMgsg9gW3IMLnkJlrCl2HH0MPwquKRb
sNknjA48cyQhP4eBBsPppJtnEZ9s7W00W1PjYzYa/d0ot8UwJQlDx9jxPFSVYMQEOnAXQ66iGzYo
djR3+5TcEGOOUgRSWPVMyWEXcGNqmLZDLMOSfPrxb42jWd9uZTM/YhlnXqV8GhmOiV7xHYsVHRSl
FpC30pbdV0bFzz8FnUOUdUGQWJ5yr+tsuE5ERLwuKLzVQP7VVfAPJId28Q7eVGkqTQuVjaguyoqd
0Wpw8GxRDjpdoxUDhsEwbv2dD9lxr3n8DK2hXmNkwJ6y3m281xt1pmmLwrnDUs3ksCKx+CS2Kl40
8+4pB5r1pl1Y7SsU4tu/aThK8D2lRLdZm3bsM9qy3LqmlabrJfoyjvWkTHOSRAOHTPUh0UVZWj+C
JayowFygEnPpnt/tnpc5zFaVOFgH4nWADGsASIW6LMYt66otnYKCg14hGDAXkF/yswJSMKJIy02X
4nRiM/ukerCujtI4XeWA6vTofjjHAdu2k9AgzHsCCoBlIHHHaRHKLgmUco2EmQ8qqPMn21lPd9S6
W1dD1a0jFOwiEEOViX3+6iyABMXdu9dE7/iTpUJZv9P0cGBabMWRn7qO5MJ1d1XNklm/USLl1YKc
u4mqNOBdOkkPhvvZlBlq3taf/QquerO+Y9F6YQDZuzlZeExCAvs9n1MpaaPDJAI2WZygD/LpObn6
JVjh+TrSI8GGGhRifKUy5DoGyHyzG7+DydOiEA5AeKrHFMenxUzPOitsEUrJT8FXNTEWSB+GCcpp
2HKPleNRMODbB/mxgeGlsOoBZXrKdflXZYi7b3W+uNnXPygr6RpKUkfURfL3+HvQPOdPK0gBUO+s
jh7B26SgaT7cHEYjc1AGtyTv+F3TzCGTlDO2WnR2rNj0GPh4UCeD8djXzC0C/V5RGhEclsIJY/CX
3pghbDio6RqtzWvrL0lJL4fnQDxggI54mZpZYCas/u8ljFhiNk0FvSNOpxmXzJNTyzSC5DL62YNC
L7nhg8kuDvfhtOzaqR9rr568RRFynAiUn5kS1WnShOVSaQT63+fTR5lrthlShufBPIFT9ySS/7as
6C2h+MXFxgsAco/dodRkmFB1fHFxvXkwPqQQW+BRBfd+1B4hBecveYielDNOMsxibR1K9K4fnv+0
CNzG7nMywyHxUJE/XuDWVhHlObYC/lcFg37GQ2pl+nXDamiRyJUaL4PGqKpK65p+11p5KAabqB3+
CRqJRsYcD0i9W11kMcQ+H0AEY3WW4Z9TEdc7+30b5d32HDKWrJVWY+iXm6rsc2RDHc7gbZHJpWsn
F1swXbySeBvw6D6XcGoHnRxN9PlpG+X3fTOeQoCWqRA9lIMAkTegxZUunkd3gLs0rej0GWl8G3mF
39Zq5xQGahY+QxGrQ+Nt7OR7iLCeflgMQbqqyFDmKYxvAtQWHLZsLfbUwugq/HJFPScMMRVwy/Mb
5DlBZ9cP7h6bcxjf6OvkL8cbB/XChRn2RVEAK+4faiq8Npfaf443OrIQ6Q6rRe8E7WZYVwh2O7V8
xS4DGJukRGdjihxoU+Xm65M0MNNz6KgNO4PnkK4bhvR7LTUSSTZLJnxU7+T3v2+O0ygnt9laTy/9
Frvp1bdOomfNA+UbB0GiiE/FxXAijk8hDLKBBexAM+W6VQJ1PhEU3R4g8OQnZmh94ZzV+XmlWqZc
DLbLQaji6r1oGLrivXnM1f5UZDmtOUQUJkMJL0iy5ECcdk1UE4fpmeQ0tZAuvgemLTtNjxaRY794
5qXtjt0hWXrbJf4yCcCR5eJU6Xds0W0IeDV+1bVc7LRB+C2htwVTkiedGzjFftZUeFPZ80AgzVeK
kY/INLJIgxPb6NpTn85Goi2aEClsQyNPa68vDxONie5dqcGnoWC/j/Y4TCgV6H2GLE9PnnG6jFfC
8OrKfphcr/aJadna9hNvBsRyizwVUtsHE0mqIegHqWlrDkV7L/5iZkAojHlLN9udTMSJoLaN5fsg
FcvFpgkKHzI0KR/dSQJvDA4QmpV5+nY6P6pVUrZmZPQ23h/LJgEB1HWOOxf2UhSz47reOjTeVjzK
xiXy1AEgyRsZia48misuzGfoOw5MtQKaJCExv23kFwOlXC3QE/8/Yk9bhGXdRWtdD4qClYAzkIjw
rGbG9UHK+ohBODe4sM+SZh13ZdSwSsk+VJQmnXSVSc8x7DITkJbII2sW7Ijup2lwglCxL3BxJ8gZ
95ATOvTXoGUrKzJ2t2O/pbcXbOEOpmMqrhn/in6SOGNzsR9fRPSdoE4/d/5qUI12aLef/qf5BllG
Et256z0STfncxk30NDCf0gbEFXX0+RznL4GgWgMevdD1CPZIsQ6DT274UMjOvY6lByDm+1VTExAf
bYsvc/FmjR6CPI4pVAjgWTr+0CAvQDgEVUiqdmrjH8wGBMcoNAB2QMkl8/W98GvDIEqjYhHjDtAx
qP+VFBojAUpYjQ4eark429BKoe4L6Ki5HUY8nvw7LuSDUkGEvTwvrBIbidMUqWVaS5ZDTxvLG6JQ
yn55JZ7qQu6trC+Nrf0b/c3EJ8EcBwjgja2ofeo9zqWQNjM9auk7AXe1Sebwf2uztcHGOzvqtmd7
06ktIzdm5hviBxmYpsHX2fhLOWXC19k0SWGOBz1YLkANiKQhvMUD5AXPnT74HPC4TUhyA4QEE72R
wdV+dbjUDTXgqIBl69VhSxqlrJGoiTno5DUHglXi5iz6iAC0GUr8srTkJLxVolqxTEm5pgfwUyc4
4+HJf8uf6nXAljEvWk+ZF7HRW82wjrJRXh5cDvcf8mjIYvBTK0HUvU2ZN93c0Oi91xOgZcTu91JZ
ngcproe/kfWL2x+pwHgxp7o/0L3M+04U9KPcKdGUnvn6lapmRV9WL+GOxoeJL7qIhahz20nz/KMq
owND+c0K2EKXjWJtnbF4k+w5vBfTH+VnRKA7CFrQypiO8HmI5Xs5FhC8MSKPMBaAdDpF5+FlvFFf
63OHTOcAjSSQ3/H+a+i6UscPYamAdKHKy/poUGzZLJONvK9rhPQGcJcaK5pf/tXDvWBaZ7qTWXGg
dLQwFdP0VX7rLgFecVX1GqrTQO1A9jZJFNfL3sMdfULmPypQZBHsTJVlsMpSxOWdx/AXTtU28Lu4
y6NlfQoYqg1Kp+LhRv5l/u/jP3WUBM7N4HKB/D9jrPSPHZ9adZRex9DzaJ5KSuu+0gOWOlC5wQHp
opDU/K4WuDx97dtBBK4INTS3NUkfkBFGUdT+6SJPfZ2kkOyPV8n3Wk5bsUAQzYEIHEjeNe4ztN58
BeLv+VPI5YgEoyYtc1NyLnn8+8XEBFPM6TBglUJdJgvn6bPD7sVT05vLNDTz8WGClLfr3/VNZVOq
Gvl/qmY/sVdlU13ANdysJW8mjx2BVr3DRe4zysu0ff5CTW/zj5r1u+9tSaZLFP9EJ4zbmofTgDEl
AgR140tTf5AOk1/p+tmnBUkuP8tLEcOeOntCYXiccX5C+4mgfT1PEUSR/LYOW208QiDfbXUc3uS4
a70Wy05j16k573KkFHlvcHIIPnatki4ovwHZljpr4EGDoQxFxNy014tss640yOfbeuaUumPFY3HU
XZwLWvVwlHFrlegJdBmKhsqPHJU8hEgbIFy5JPhUkFNeOZX1ato6iwL+WMbJpqAikIabrozhUlsU
XrKThBiX36D+36/rT1u8DY2kzBHZKKBB6NHRiLUe5fGo+jvhfrlcM5Csq6sS3hDfShw8PrJdzhRo
5y5jlbq9FRVznbkFgT7Ia+Hzp3Xe79UUfBGfl2A+IQsCd0uRjyLvkgbaMcy7VJ81UliLy26g1/M9
88mIxiTa3tx0rRSKPH61Ij14Guy+aET+G4Xsq3pMcpoIl1li5GAhdVSvZ8TzFEdr8Ii33uUY7Ltc
yGH7Pz4wYfrm+BcXSOjTouitApyw1Swhb2xAk4BZTpDhKh1rPoYQYlSVRwvJgA4F34Vka7pmuYUn
gXYmzWnChQ75/IFQ5LU47qd2DMFSoN9/i47J92Hdpwm8046OQ7PL0K6hsj6YuMj+FyLkzZb0Bm0W
SI1zCJK3QzErVGLDsz9eZdM7jacRu+/SYT1eTKiSg44BLbF7fsem77prahfXool5UFrky9ThAWKd
uLRII6FVzniqohz4w2PqW2hGWCc5WtYhZYanzldk/MkhlMB4tkAtPsuxu1SSh4P3bM/Um7FGB3GU
mruvoe0/2Y2X+rJjZNUAGnzS+V+NnB6PzRBtbrZxtfFTnl4aehOLsFA//LMCeQKnHklzC8V2vVKi
aNeqxdMBNlaMyDprvhKdRiw/okaEK+uHA0uME7ZvU9UG2OobKqYXs/TrrtGuUXyu1md+rDVK4DU0
E8az675SWJfvPbkfvVqjQBnlE0tmkFQKiLuDNBLCJaO1PlkHvU8lXi/EndtdQGbT+1ItgXYGejDx
JjiNc/TIB+yUfgkO+omAbb+yyxFfLePrmhwJkHAH10mQjVjZS60caI1dZoSmFCEb6RtHjtWSbnvF
38frR1eCEKOFV4nYJGNpPEdUKQLUNU83/Z1+4qCY8rKIb5KjOHH89D+y83cByWny8et8EIIl1REx
R7mH6TlUO8+i+p2UY9v8CgP0lFAcXBeNayly4TNE33FnC9SK4A2HliKmZItWirvLTOSaKtjz/l8p
knBhjlusu5287MNq9o95u+f855vAkrqK20pdydzRnOdYtHmOTsDxxMvrTsr4JiaOoGBk0iLUMzUu
dSP1KGyr9BmMLcEVVofa0ejB/qSxqeS0mVS8XTKGCuKEaPuOaBeASGdmmybsXdUdphIjOo+9qxS9
HSOB8/1U5thsj1jfhCtMenKuH2citEIXx2BTI2Z2gp8s3jChiweVsvJBI+c3HA0V6oZJtzocRu81
4BHk1LiQisjeDjyf91ACcoLhaBckSBzdQ5kKilbWkExHn+zOIRNSSjHXOvE4n6kN53on8u4MjT8g
mpoH2nltjzZWp0Ao/g5LNoC3/5+EZQ2Yf8fwvkoA6EyEZozCqxdEmZ8gR0lNY8QK8RVK2aH4Ds5w
/RWn8vdAU+h6l9zIr9gC9K/HG6AQgTADKPt7Tf/7CKoVdevxuZI2YXJlWGMWUY0QX9nZg9FRJOTZ
M/ph9Y/8wa5YmRSUGJm22//fXoyx50K2DN6+qm6WQugt57yG7UZBw6rdqOjIcldWOPzl20Uh4vWB
2tJFcc+lX+hRNCB7Dv6HQYCjXeWvnvcocXV7P8Fw2xnf9E9ADa2DXWGgtK65slJ7TUfbEmYpvdiQ
c98SEgb+PbF3HXGm93FHHr8WGnKMU0ELiFN/AX84kyjcBApiGZo7McJhQHXvUoNeInFZRxNB9CE4
pXzeTje6/5NtPPA7KgCDrjySABjvYgBmsSjF3ssP6hcn1O3EjOT/KsB2fDiqULPEQE+LZrysPJGZ
74HgSp7NXCu9q0rtMjxFNnT6xXhwsRlkLfttC2/U1c3LdqQPVAfjXwwx2lIhV9UNPB2Qw2ibPPfE
piGUIoUo9fYK4IPMY6LQgH8YniqL1b1q3MIspmtp64eMhJkJO6aZgFaxg5wNReRRQsqBxH7q1XMD
TUu1Aw29Q7Qt0PQCpVJYi/BQEKrlmvLZ0ixkZB6ljWmN/x5T4aU06ISDLiLbJznU/xwSh5c5R0Bx
qsOfZXwel7tPb3OlHA9nxHT59ZOQUMeLfw/Z5MdfKMhjQKNIiQfiaCSGEBPWfzwLVMZX14J/+cqx
Aaj8vcdkFiCq39c/fk+u3N/DmIw2dX9+jPnUChEigfCqKBp2Fdk2lknHk5ZZVqWSyeU+ghnXOwn1
HViUJ/eOGQFkoo+/7RCmjVAyKRntC/GQ8XCGUzzqsETTp3BS+AqbztyKE3YsJbeoUgEnrP8cKoBx
6pfhSHFumkmFhoKswsXCabJ4TyDCYImjRn68gybmt5aB1+qQmslrm5TJtDEIF0nxI0RIiwLyVkba
fyz5bfdJ1qN69z09a9W7oGtseKY5FMrdEvFpJOTnUQY+8DWjQiit2ADFut/uFLPhZ15PTD6xWYkE
hN6hPkqg/37MI65bkWqUyc8FxaWamv4y2ekLTePaLRLBAl2l1ekHUeG+YSMR9n4K9XPCT+DHh9io
z1z0JE3UY2eRHzDvs/9MP6x/jeIjUlGcMqdAst3c6ItueEghfTophdkYt4A6I34bKW5NaO2XAcuw
++TuZY1PJr8gFTVj8WBYfwss96bsHkclU7mtM9ooTDHPtzyG2hKespcw5mP6PcXmz6BalQeOtXH9
TbsRIUDsvKeOwJMBM05Y6Htbt40tNFteowBYbqYzT1INqucs/wFjUyzgARi1yHfnbgrav/IK2+ee
7k3PhPDgXuWVi2jPV9Y4215MIDQpXf4Owo8Gdf4aD5VQXUZc0JcYT/m4Zm/grl1GdS7P4b5IlGbC
vGTJR99/+7Tvft6w5IWHMFtNk3YUQiDocxDk/nJB/EQZwjWVotp1H7qOwYJPI0wBcSmv8kD27tli
g6fL/nh9IyFuGR9XDtlPBpNBqY7Q5WPIZVIFM2coPN8ju/F/oJWPF6h97vQQc57wqIt520kfkBFm
MgqJIXDsA4IfenUdsE/FeN71BonosyMZ2AcGLECliUIHLvoX1SoMbTohTZ4L8/QYbLX1+pS+U/zP
jIOJUwtj75hig0D844XMAr8Hn/Sjb/HUxW3lhwNxmzXFICYuKdxG4u6WVdhSGq+d7DGBNJb7riE3
E3NhEk9hzGRt8Dy1TWMfK0HBUXu0eVTczC+h39+FlLrD+BsgzQvFCknHYcdSE+rF2SKbonx+vJ+f
eWMesJXG78GramyWN/61iRJQQ/8h5yJg7QPW/2VHfkdbp9/lMGC5UNShnMtbwtq6n68t6ZMxQTb6
Y3mK0T7Xhd6YZccglnh+ZugQuddkc/V+khPVSIaFhDoR27PH2JZ1KYZesoIc4prXeRGIPwDlV8HI
1Qh/DDVr0cYYZq7xkmhBU+s4Ka115YH/MhhQ3S3KxAFjFy5hfHP3XrTxxp/afUQtPRAm+VEHsU3k
cOH8R0L+2YdaNT3+zGZ2OIMDdDogc4vADojxoqohzXo4waHVttDbhdaqFIVIZ/TSGYra7s94NKQN
yszV8jJqd1qVcq/fiW2Keca5gPNre+HsAz9SWbkSOE1s5xVSU+mQ4kf/ZcfwKUXwYUI9W6jqmS0p
SQHKypAnF8DWrlShUHzh9hSxZCRauge05ZWT9GuV8f1W/KFBRHG8BuDPqU8L01WXeLpDBNRIX9Qs
4k5Mf5KK1yZUG484MApyIcsICHjiEkwPtHyyJv+SVrwMFXGFcmMte0Gyr76A9rzNr/9E+3RFBuGj
pYsLRBW+rBlY/uEyNzFQUoHEPerCfN4D43uto/RVENAvJTApm6GzBBWXyM7Ntv0GAep3g8cPnVXi
lzb0uCBPTarPcHzKEHcKA6igos52by3HnRlwKpX90oWSbcdZLZxnJJAUDUayUGV26mWE/HUHOgS0
GsTkrSMMAVPMfYQwn9YaZFDHu6N8Vaf75+fcMdbJJfNspvqaojUznSdGzilxUEN0FJdZUYImceZL
auOlJ3q79zRMY1wJTR/HNGuw9brMOzQvkg6J4ozgXO3d8dpoNMu36Mq6AgrtejDR23uKhg+0QhNP
4YNlbCMkD0MmuqwCViiiIQ+qoznWbUAfs8snLGuTF4l3sOALbQ52BxjnkhbHrpGxxMx/QNxIUTrO
bF+xwTFMCd2LmKtSXicV6vOdcyoWJKsvGo/HXIJop0O+pcCAcp9XK8Eqi4NYFDC1A2GKzfgeug3G
ieza5OWBvNhDwa6wzVu6vpybfM0RH4s3I/2nFCuXq4UU4QchKcNFsJEq/XMfPW34WO5+8+Wx/Lbt
xaZQJMyKr2IwG+5B1hpAsmIqBvXSGCGWABWJ7DtNVfb7I6DZewYt+2QBQ4I+WTvegxurzaBvg4gn
a9a1udFj1ym3u5TttDkiYBJ28HrX5BRl7ZupK8L+qVdb0dJJbSRWkPUowM8axR8iLV/HhTcfp1HV
zaIND8X/AxtLq8Wq2/xiz5ODvENszoxVBZUgFeGf7jRfc0Nac3KwvROkCpBV36Z3EtWJHpcNlIxJ
hdI/TFfvDD1zGTb1weHabRFUVq0Akscz4AWrl4sm02t2bwCG1msqaWACbGLl5evaD3Q2Zl4kJITR
/fYH6lrxnqJX1cx2ljvMdcRoLuOFiQ3VvxYL1Zg2Is7haQRxBuyVqo0D8x1tXI9QBRv8jvsAC2do
aZlhEq4uVEFv6r3CUfJyZXX+WTdW9NYlo++POeIbMtINjleMKQtjnfTeiAWJ6kI8jVQ7nhASbI8/
tT6VH58Zy7KEw+a5RpZ8JHj33m5kmD6kxgV7ZL2wjP78xK537SWPZAFgq47WpZqnXqOEYKmwj9vU
ZUBJlEN3LZtlElL2mw9v1Iw5cJ2JmvdA9sSTdaK5442frIk85d2J4nDA119skDZMGcxQ/78qcnoQ
S+d4w8996JqBKUF/HHkTpcQaoNQONtRONHuF+17pXZsk62OXmMSGVHquocoLoZ1Qww2n30hqzW5c
TV0uhzq+XiahYrMVG2N8ScPKc/HEozSdR03BBIgBg3a/Yqvzjr74bI03a/mKffxPSUz7QNVOQ7Wu
WN2JGwT/ksVFlKbTz5svTJopgcCwNEMFQD9yMH/iO9nRG+qlzPRTO2m5pdZLT2UTQ5WniV1XmIEF
+fwhy7+l0Ssk1i2D47+ZewmKsRgW0U5R43nuXt83EA5uCvB5fezHbtL/9zEkrwxyVoh43wmysGLr
SNsK0v2sCO3+Uaef1uUwOt4oz8ZSNzgYaU5p9Gs5Iqq6hmQdItj3Ci4E2nzVEa0QjV5FBXaug0HT
u5GtP0YqrWVwNCmZ/twJj1XS8byXM/ZYcucWHVEYNOGDlFe+Nq62JI5BNJ7N71gYvuaXIazsufwi
FWHrEjwydIAuYtCfNzP9tsI9V53BFL0h8swhUwtXDHWvCRCmDL2PgwH/z/oZxu0Ec4qmbcwJFJD6
u7WwXMOGOzK9oKTH8puZrOKatMSl2Qiv2oxpS4YGO76mwguiedfDlD+ur1aGu8d3kzD8UNT+q6F6
ADCSMYz26a869T734plYFdW9Ccp4BC0NvtM7wqKMYeogR9HL1aotHmbcB717bubFMtqGhLjgRuMA
mrOPFrCEaX49OVWgre4HaoURgOi5vQBImt7Gd3s6qpCKyavtU4bbgtgqdzFR0smq4SQImR47GPsI
5P1IBGVVpjxLM0+rFubSlW7BYpNs9nKc9jddFCkbQWdmBMaaQPVZB4oZc/x6tS1DDxBhf0k6Ep0Z
gWFS82fgOwgKVn2c9e33nljQ6HZYdil6ZJn3p69pfaKpWs/cKrtR/HSoOfwciWGoaXLcNtLeww2q
QF3G1bfLiU5KW6Sq/ucjZOWBjJXL6mb7ATPtfY3/DocMnakNFb0XJ+mn/U3O81u2CCr1YT+fUbgZ
0dKg3IdRqw55hoct+xZxzbbwb7l9ploIhoRz9SflK+8rEdg9tuZywgdIVivb45+StaPyHh0Q3uvD
FV+CHIaFSEq43L6OumItDjjG3WZQp4BKphM5gMK4tYuzWn41ZZc5Ypuk2podQ7tzQfh2oq3Vnr3T
pKquwLdqRGDGRm2s0ZSoyZF+eaWLmHYYMVVVS0CCHaBn2u33hOgZQ9txz3e98K6YMaL1uwCJCVUC
OfpmKZU2fF59/lTd3r4Y6nigtiTrWtO29Xlopuf9vbZTYBI/Tq3WhfoM5dBtUkQSwJm559xfj+pg
6xoL851M2X2ueX0+mBUBSDrTYmZBgCuxuC0ziojQ6o0NBpGmoKqoY159U9Yv0VsZtuh10SFx137s
DqQWiemzTR2OR4OWXTa6cPTpQoEcNvsrPt1e8J7/rZAZT9/+49cyF9/eLCHYT7OYXBWR9Ty7QmwG
7Vf6EsVmEc0/nePvBq2dzaeM1nvKCU6eeE4S8zIehrMcAVYHgO1syjWU7m3t8yNC5TmZXThAgw/c
E+6rVQkYuaCTzlv2MsFImh7ogDRw/bN8BY1R+eWbNspw9vIPNBDbDUG7GTv7zj2nv6HgOcnVi4ke
2VQMX4oN5MX+9XTzMuy9av5M6pospGDhAxes+9nCfmLld4KF8HuWnW7zFrVrmx4SwBhVNxfVDl7A
fHnR24+KasSxWSKCTEKeNQCxzrL/LB0clPrptxnZzjp7LCFfpaTdEQCXI9mBtBgRaqfO/iWsIdao
wokWRoukjnJ0sd1EUImkexGaPev0W6zssUHyTNCuTioMSwEKAX+1crngIFPf/BbGfKS43ahr83S7
4J/IZYO1GzweDnH03VPKjUWoghDtnVNCWMveIwO5/Q23U0y4YgaIvAqtoKQGXLy2CZJyQZQCS1Lc
Tbo3Sg+0/WDRyS4OyYLV9VnZe8h96yRF62KezzMtKpw9yIoNBp8LjB3nQVjdRj6J9B3+OPqmveQ7
b33dmBTzuH8JnsdejuUZBU36wFzSL5fBo4PO01/ANmmM3MyEWKqOYDfAQ6HWrx4xtElI87avur8G
H+LOrQ/lc4eoCYB0YCGAN/VFvMikXIEfZRUGeM5bC+bh4y75YRWGdoUAhv54X0hfMvdl/ut5etGL
4DgmXBNMClR36KDQeAOt4F0nzroPZBtgJtK9WXZjwByFkw8+NSVlSID7UpptMv6wD2d4OfddudW0
M0TWGeZ5JcH2OLORakpeVFeXJ1q1Cj3dqsij9tudd6EXZfeJN9T0zBK9pMEgJaBe6DGJD4N/4I7e
rhVsW+nBKWv5oDLdLPlfgNiSGZlyt9XXU86nX0Dam6LDuk0ixFkV5gN2RXl0VcLKwgZcnEcegl0Z
gW3EH9yOT/2EUbJ+S8MZ6g1HFeEJg+FxRXyLM+/p+VbFzWMs/SuAcX+trpxJeO/3O3f5wwHpbQdh
A1KRBU34z3mm12UgSrC3yPLW7z2vr2dT4qF0kV2TumxZ9y5O4jI4hRAvzgUF9p7wXWKX8ineVjxk
AiSKEJg4lpvuyQG9BJMtqzV5hsEHMYKDm2tFebUJf15Uh+4j77Xol4kmHrDvcsFteMXN9MBOEdHf
ryM983pZBUwTVDmNyxjEhPKCPeKdGc9UiavF7scgEoYvmSe5KiE593HNC5hIVJUpdi6xnM2He0PJ
P+56SPRMW3w44gksY4/dgOFZmt6ivBkBVJ/WXCB3rFljVrpe5wMQ24TfPxGyyxFEWxwJvdfPUY9f
pAoexScAG9/MOFCIcgj8SrF94s2nczzpOR+15XDr+XSai3l6p/HJAztFyke8ct8EiGJeew9g4OXm
CFxVyhAFu37+LjxGm1XTz26hHhRBzklgvQKmNwz5/Wdf7RVwYh6E65kCwaM0kkGwYzyJ8+0UTHAf
dUGXoBfIjYaBSMOpQP2gCgFlFirt6FcpGy1LUmgr0unSgcVzvj1LmCIo7GLaX0BlHD+NyxTLflYl
CLskPzSchKhdNhietNPQRynDILS/8iULBJeLGWUSL8MrW62eDLzZUIPZFes440WONU3mvj64wevn
uvY8kO/sN9UfILimflFlLFKXZC1rJLDZy2xZpVbBEVHwCSBJPZT77VaTRVQz6a7ItH6ygvm7zlfk
AtWbOymHGXZYxMfQ/iKIVQcV1ugCX5LHZUU7a0BoZKbTk56DP1hkExqk5KiAw7uvU7TbTlW7q0ox
MTxm+aYje7+4Q16tDDT3pOP6/aj8c1ASXgoaQ9bMazc8yhjQ/nRWihT77w893p60qYTnHQOiTUK6
pH8Cohfw1Q59Bl6W/7/IVNnfytnR0YvSaBkawGz8brmN+mjYQXRiZ2Y51v7ea4jBhPjuuCjRxANv
rrboWoyg6rAXIg==

`protect end_protected
