`protect begin_protected
`protect version=1
`protect encrypt_agent="FMSH Encrypt Tool"
`protect encrypt_agent_info="FMSH Encrypt Version 1.0"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2017_05", key_method="rsa"
`protect key_block
BlTcj5uV/pzDt3Ns+2r/sW1Ygr9PKlOrSziXBEbvqCuzEUQdRssAYT6ksLMditwxfhgdVyzf0Scs
niC9GRh7A6ENQVSaqPoWv5nGqZKQla3SjlHZqn7v/zl7hA6S603x1wge8nQzEyHARNd+NPCy9Mgz
DduxT7y0QZXZ1s5NI2qr1kgfmKNSbQCAG2lqP7T8za90wrTtzIWe3ZhcaBYBo4sJEkoMzgExjWWI
HvMKgtKNFFV4c4DDmgoJ+asC5kP7d7Pne5utLtOZgQMjm75yp3ZmRubggLO3XBGuGoxPbImYy16K
B/ZqomXIq7TzNeAuoxWL5WXNkxzXCtRvFRE9UA==

`protect data_method="aes256-cbc"
`protect encoding=(enctype="base64", line_length=76, bytes=967184)
`protect data_block
/nTrR5V86ND7NzrRj0fij0Si29HIXLPEe7KLdB/2v4wtyVyeVyZalkG26668VeUntDm39DJ67tTW
glzGMl4QRCoOGeLfHLuccJ45KBuNiTBvxMCanz+yqOvMrP1LrzeNdGCfRFdeqTdB4opCArUrJMUy
nXp9KPy6+JHNgjZWyAhue21AVbnohE65ciXfXbXcwTDJdcB7Wj5hbv9MamTY658As1CB7NMFgoJE
VYPcKAC1qMsOVH2xaRUDFDD90pDWLpbTD1IWDS0kIiEkgzePp9Rj3H1wgAamla/TfNy6tu8ZdCbZ
fgGqL4HEXOf+62QudT7QIRMldzH0ZzA9aSUemnutcGwVZYbpItxsdnGjsJAWne0uXi9KjLxFG1aM
cMu+FdrdUuF7W6QQr2Qg2KTbjezZjPyj3Kl9fZQ42+tbZHx9FMtr1Z7G3UPZWoDTBJ0LElDwCBM7
z/1eVnNId9VDhaCfvwr5lD5mAE46bWhR6Iepp00d9oFXGSJ6J+oy+81D1vVqF0qO67Dckn3Vjn88
OTZbPawRCqqnJGJxrQsBWcZjmj/xq3+l2QU5tBPmDGWxPCH3W8UKaML376rtWpDyheKCTVA9X8TU
X61N5Ik7XBWDShsOa/g9ePC6Ljeayu/uJ7qClMNyAghSsYWzIZNqD/CbDAZ+GweWBdz9Ym4EgR8i
g9rNoKLW0YbjKdGjBnSDxptQBDggVCN5rUh582xWjSoIB8bDGIDzMM/89jQQ2Q39sxa1LLRrk7A2
SCK/i3/OXusiELfyteq7b0Lq1VM8R784pH6xymnP5TPdQrTyrSMIy2TKnC+6SNqICHTCtjRA/5/h
+vj8TTlZpD7ul/2p1YtT2eYcdTI9oQjpo8kmaIb6m5oYExDuP0VjJYzsVjci+MNWU/DPQErAmqFE
1EOukLwDIsinzbxKvGYtUemG8cxuaDa4HggQ009JqJxP2qsEwBVAutdNr5rdnR072dzuB/pdSlOW
sYzfqNfCbE/T6GizsL30TD78KKSVB+DFOxmiBodrK8S/dTj1VquiN1EV+k+dS3cSN/yeITRJaW2t
8AOFN+lNcodN9oYufg8OoDezqbQM/C5wz+adcDS6Kewg4TgQXU1F8VfpuqL25Y257B/H3a/GqQb5
tPW19oX16IkkKpq7FDM9EtapAxemAQNYg85Q27ZMXGEXZHYNqLfgx/9uJJMbJBU3kBfsHslpswub
DTg4W71dATuucLBBCBaIggDxXWtj6179N2RRmEwP8maBK8SQ7lOsbH3O+3zw0eU/3sjvoqBovuHH
L0A7eveoYcE4m3hcNgadPthst/JuMhzJZES+qvxe7xdyQpUZWyaJIOmj2A+GDXtQ0eLBZODsaNoh
9wUPaIx0Cdf9/aNAt34tSR2pJJR2JtCvtImVbGtzRlnF2SApgAb/mFwvap+HP1mgX6pttS4XDBfg
1KX5+p1fYDi7iOv/xBZuMvbBgKqcCdSLPExIIb/n7MI4xwLwasaHr40119xLgH1/wvTMmLJF8kd8
90DLx/TrAlZwuanoKLvk1yceJKHKTjpfH0RXq3neY/DzFUT2fnMo4dEh3gaihLG3AxrAkq28hfFZ
ErDERAq18loL9pLyvlVdNgbDIQa9BbT4JYcKKaSKmfG2aOWv+ZdJabp/eiGZL555XqtWCdsQse0r
H98iyoO6eCN9umHHz7HbkRFgGlUr83ZafDokkr9HhmPbK7LIDxXmDH/HUCnfeWikgLatZRZ1M0Qf
xWT/ngKG4+FGur2/+CG1lwZeFD7UdHQ670JDYeBdduY8nNP8C42lbZC5u5ddpF+J0sJJyOHOLDAj
todVtYI5l2zoeGRMjPRGt8+oTbhYPQOJsvFJ83Twxe6pGyBJFHDkdpiC+1zxW4bSHtQHwL+G8jy3
QGRWhZ8fC07gb5Qwjca68T/NsTWtwu5o9ZCAvUcwU9QP+0ld6QF62fcqL43hDZuwNeEXElYexjnB
blzwsAYMDrAakjGat0x34zwAY0C64R14J7SZfqZCVAtwhb3KyLilCRFCpB5w4SGuXyqnOF38db3j
LZIaPzHC4qdPhsKwYpf5EvRModbj4C/7+gfaUjiI2cuMR2JS6iiyPMz7SyuAMplNUN69Rlt68Uxa
btLLPke10xKqcCFbm/rLjTXD2kSWiyI7GqRz9aL2zM1F/kUJtaOBr66tIACKpEU3RWDjTxCizrNO
zXEbt2slgcuop0Lq7AwRUETzn3pvi1/SIlhHeVJZH0rHZDRT2RI6ehbk7+4trlG8iTplSpEq1S1v
OGzFX6JLEELxT7fzrNAsFcDmqgEpHoMboN8S7LM4rZ2WuVJaN3q7jMQfFSFO/cJEtQPY/uwxBV9y
mzz9hDQEKpWquyx8bDziXrGVjZCSp5qH8bgqoboZ9/BEj8uhEDc1st0xaRk/GNwnmk5CA2T3EM0F
QYtKG2RSWPj7HQ2ayRSJRXkpCj1CnEp/9f2TeTBjlNqdee03PpADokX6BU5hI3Ookd01FvKMFPMw
LUfDVF2Cbzs6jizSkNiSvQ/0zjEXXYXJKcv1myV5/PEOAnXHiJd+QV7PQfVx8ukG/cGmuwsjxeXN
4ciltOtX9VJxhF6Z9wIWxR4mIu5YyNLs4SChsx5aQ31SX7YkP7AuYbvjeV8UGEMXgzX+kD+Xk7a7
WAMReHr8c/VRSSnxKZZMCmXAVJwTzQL/ZCLNwL6l8jShqj5jcFcc1bu82eKaCEBjuXa9LBzUwC6P
f68sWxkTVtY8TmNxBZ4olSVsj4cj8unh6lyYR+VEMTRiY9QX1HaIqGp0vkv3LrU/lzotZmuDa4MC
MJeunodHqI3tpfVn5k4u5+uog4qpRIm+Ewl+9G0ujKPE9JQaZoCHUpL7AYe68iau3U/LDtF/wTeE
AqU1F1KMrQOH/w7G/XcdF75zJDIB2sNK4TlesO0MlcNtn39HG271OMvaZqG3ZXzINn138UwtnwJ5
wrb/ku6Ir6DwntALClmSh39MTh9fJZIS/2CXiXTzTZOifdFLGwAwhxLV6nICQj0f6i+jleaMAmXX
IztjmRJjju3y7pgUEaMv/TUAhh9Ulb8lKhs9UTgqI16vG56xk1Wry1elk7kSpov7nBKqcd7WmUFh
pgZ1NVsTIx+Uo7lb+gnjtfvQRWf59gxcl6pmRRfyFN6bTMlcc7r2iS7b07JalxwO8gIbStRP3v1r
AkNCSE40Nd+qxbRXEWlRTcOPdKwziEimqD6nBGsU1qHG8wBthbIIPcEhTukEJ6PEgm4ay5Ff3kND
B4MaXL98CgUvLO67V3dP8AVwDYVO0pbZNtOpakuY8lfnS+hFVIocAXsIS1aFEM1Sc3ORtItlcUnt
GT37ILMyLbTeyL2trspXEQVRCSyVwVv4MwvPllkzb7SlMAn9rpgY3lZO9/o2KaShyo1zC5M+pLcd
Py8RLpcGNBuXpP52ed/quAjuJBxDQJfnhPNT6VOKGxQi7YMki7z5XBY44h/ghVDIPKcQRSgkwkew
wi7SvfS8DlxJKW+FWqvriF4dZjBkSk20bdss/NN41sYzjf2G20I5zBGmLlF5saOu7BPjXex03zeT
NOVVI1TrK288mgxAbNaO92uNqCUWqdery2V5U3FHtttr5IjB+hki0iXdEMHWPvQflwLfaTsrk0qh
paCJHiokA6CDmkvAhu4kxSWfDJeeSA6Ze29LiXJToSeugab63TFr0gFuclrjKMnGLpgO+2dYJJpl
nLjiln+rySt0x/wuVNXgjrIzW803ZZDud5PaK8aAlYexsM6etZY6ZslBgWWSgfUwXrFtuiBvVmWC
D1H/H1LJhZMozLN48Cs4slghJCD3aKpRbNZu/7L1cK5ovU+D3uVuXQNPZYdBsN/jwT+bHG1QxS1Q
9jhVXOCKCvQMvIoXDJvvOnYaSlTlRyZ0BBIYX4sqhDe2lkEmfdoveN/W4CDQpXqolKCpv79zTZsG
lru4gfwjY+mVFabhmJdUCrW8PfHGRbHRJqGIchTjo2uV/jtAfRvM2tfeGol1Ry4HNcABdC1xeJ4a
4Q9t4bu/rCg/+ZtZaJdoH55W2NkjxUnopeMHA6aknspMDYJDxBw8ev8vrtN02fZegx/6IpI8TrFs
pSIpTfyMbIYKfkPac5n5w98FlPny/DpgZGBrbMzT7mwpI2VUeALvnpbt2C7wpzFAcSx8JgUdwP0Y
FBlwkHKxr7y2PLuWr7seqJcMND7RVyVttcF3qK6VNx8eLV6nity03IGp0sJPdw0ORVENTP14VZXh
8Irut3+n9nGzqKGqNMAYxdERor/LPKhf0WiBkSf66f7UZKnGqpz4IQ2jIebM4IHGEp5ocp08Aej4
tIiA9I9V/PTltZu2FyelkZ+8UU9Pq06eqiF/8ueRl4XxnmDXpmIyqPRv5HTIlcIjPDfxSzrkval4
dPBPfaYjG5jg/LkylAPPetc+sLcD6ga1l9WEIWwDcQso3CY6LTSzBtXIpP7lE8UM2MZKhT8yK5G5
YixUtjUNd7jlO79eHvkGK4PayVB/0cETMd6LvKvsW+05Ovl4DKUht3PaN33neL0N4U6IBhI2FbqF
h/9p2TxAsFWqQClE67wGJGoNruBnb4UAwfkFPrRjKE3YRyF3EUXeiyd1v32HlaApi26dstzYULJN
Bc+PApxmZ0kbKFRexLyWtTEfpfO3eAUC67OtvmIfbJqSUx4GREOqjcfrEynrSuGiKjp6bvb+J6Xk
RXvIo5qDgnj2ddMFeaVTRanekBMgswTYzeKMDrndGLhVd9xEGgEKtlpsB7d7YYt95xcgvUbERGOB
rwP6UmhwUrLWihxcJEgv1xEFJUnw5oXVvZ8s9JGj6/DRNAk2hn9668UrnvskeGznWqDGZsLZ3DeF
wuPcEjARTbATvNhiYoVuakYTVGcGN7ABnJB/pKgho19iT/tqS4Y6kQjx1SsCu6tYObFgTeXFzooR
xOy630b9YnyN5ofFpXFCTpqGxvDRbqzumn/Q2aCIAx4EoLUFRbSTpBXCzwoAfs1dcwi4007BpJQG
xjjK9W2dWCG1y6P+hOPJf9YODMrvPVNuVU0Jd5ouN08nEmzOfx5/WWV1Xpc2MdMqkwwSxtLoGdIj
93uNJxcC12ZSe2DG8w4zNeWGyMm/x/KbbP84XPna01olVOQOQPkN/YBFYFWun5AYXFddQq/+BEXs
warmRIZenr3JDBwzf0gs7+gPZkjyeWkSAq5dw4QPVM+v34ZEOPkLLods5mVLJHFOABUUkNYVOBiD
HnqPR0GAZmCmLxjdMa0OZQT9CZYyRgCi5oBJObfbX5feN3qrW69RdoceIor85K6Y+J5m64Jt6jNh
5xLAziKq/TMtTV21iyXVn79BYE/icU0kuLsL8hNuBE+++f6NllOe6ZrJYRDcl3xn6COaUSwBqXSV
EtBRI43RUs38Ud0ZDzrLlQkDOgz902QyXuyPauLlmxcZRuOWuGUjXVAMrMbiWDfzBGW5ov0ixqnc
ROcJCUz5V3tLj8EtI63eoVI9L5q45vIA4OVNAOOaMay99TxIH0y1/h452ug2aUOMEs0XL2Agy9C6
NV0y2qZ8xDUKHAu4424P2hsGsRC7OaxGxgZhsFL67y3v06tNsqtmck5odY8aJJVCHBd3R3PO7b+X
AGcsx4VLJ06f84sx2c5Mn8dw1p5zVrIqxSGadKRcaPBZXPvZ9ouk6XRkfFoyoDNnlpSUY5ghzYMr
jrO4MbjcgPhSGhleATWWNZXxtnUGV1oR4dI7aFICH1lvfpAhG7BNaKmmYdJbBzN/Q1OjszSAUT3T
3vKACLVzGsa3UaqsFxB7SzHOTvxXBqd71o0WrMBSWo4KXr8SbN7nJZrt5dK6XQbPqGWoC+PYr5jI
pw+CaeTo/1bN+pxiklQi8VeEZCZezmKS7s0PF6SwxltjfN7wW1D4Wg4Xbc9mn5uqvk9b2ULL/lhP
FGn6ecBHpP1jCeqoJuHbigQuF8DyMP5x4MM7+Uvcfot9fUN4krzAmqoqKlGAzoilw+QfS8kPx0Nx
04jJ5zQgzgLyHoVjB3UBIrtV0Sc2tL4ljWR1YCYYfRntPobWh/0suYRHWu7yUjkS4oVkGELJJQ55
hSi8V2HuX9iA5HZ2bP05K180SQHDv6tiPGq+ZG1BUuGx2aa0dZcmT/nJ6epQ8kiWlCTJz+mRzgCx
Sv9S9n0HYYLfalQ41dk77s0H4E6HBP5XfkwzK94Phxtfp15lHexQGwJTS6YsPkQeO5JQYSOH8kiE
BZawCuTv1MIsZObjtL69FGFGASU1fYuEYtT99hOA3JENCyVLfBXALoR38VieKjodCtCmCOXwybeI
rubRcMYhqb8vH9OpRaQeWAcTWuQ6WitrBdEvtdnFzH1AcLAeNrIyvknYghtJVPHAeuMVShT1h1N/
IB3jRraUDD3daU3htJWKV0SJib+MYRidLL2TsB+rukMF/QqZ9yNipqJrTccYjZYzo0O2/9buMALa
sy7YEBxcLvl8sagrAKno6m/nPHGAXO911oeXo9nJ5/0rEgIJD/ukmFuk26r0E4Q2NSzpDWikroLk
JWrHXWhdw1DB6jJmGQ/cGlocAZOqc0NbRthrTb7gRxWCcWlvNnH/yJ/oPXeY2kMZnBoy8kz0Kg3C
T63aqML5ycnWokQxWPIHpLkRf9s9hHf6oONi6vc0kQQXkAKbmsHF+E3dO+RjbdnGU0ILuTfDVTR3
+3sjPNlrMtwh45jakWfhPAkInwuYPLyHv9WQxtYFpFTNgYoAvU2bZnbi2ctbv1+582QjtltdOR1Y
WdpIAzM1iDStYgmI7jkkbr9TcnxRt/49JMow6nf5T+88+MPPgJIR20Xxyl5+53wsJuZD/wiREi/a
iagyUk45ihBI6RvDkh2kNmwFOW+ALi1kZs6mOgM5RwjoKMDFBPuyrGGqqJlSCZogzPfr4bEDWXMc
KvXXul03vwKrYSeIGEHULHQSh82MQk1r09kkTuLXtBG7GnZeVdD4vBKdyGU16XdSzqUMNVeAG3YT
ke+5r3o26f9fuNGTx6hzbp3YRURg2jW5caUVGykuHMqcQJJATEwf94KrcLNEJz9XwLUquw8cGoMl
5Ip05iOPmo04hvdHc7nUhnQ4TmZalx6YFVmdoMz4mgc2qiJ3MyO/qa7i7eH7eongRzXC6PXJ1vlO
UxNIA+BWPJy4OH8UbiP03x+EsHvDURl40EHb0C6zCFwdDPT/sZrjlkpPpXMtn4nhHBFcrpfOPGaO
JSAQeXqUqtBcbt5SnTEWCySsW0222QEGPnA9VC7phK8B0U+K+Z0kk4O5tyk33HkBiajgZNB4jZGu
l5hGeUL1PSTfKd7pq6Ye35c1U0vrznsfgdaVkvURn0znAU43QSuSfhFJek3VrDESYTwK7qkSfsp6
EgCnFGEX2WdkeWDqC+vENVxKwwcCpsSvxOYg2hpX6sgcVjC3MNHaGY4i3hQbUBftG+mm/5zCWYhm
ARIdb6aOSicSf4+IzpncChu/1CtNOulPyFjYadf3FbfNTyiNEcauYO8D2M3B43sEiG9ROlzmW7dh
BPo+8KNeu/rz+KSB8eyrxgjVU3EtXyGcO9i9cWd96PuevjH9yV7Jr2Lb44X71k3LRaX7lYiOUMz2
GLn8RtcC9saNPRi5j8g55SDd5M4yNF86YLcN7/t/ZqD+JMfF9OZAOkwE+uzyKE6rkxIRKYhA/jN8
oTqgFPzkzMhzAsG1qNM+Y9xuKVgQw9iuT+vVpIm2I2uRT2GGO9C+SN5pJx2q8oQC9YIZj/D0AAwF
cxj7eeT5+6QQyK9kl08M2nAofpXGjUdrKa/L9mfUTKccz6bSPBttO4/sSdujb1CdDmafpY1pfK0i
yWDpC9qOklp2pmBvOGEvsmBFLIi22GoUmPCvjx2JfK4ck9SZL9YIkNTZldcL8TX6H3ag9e43r/cQ
raNvCH1ONb6oWErkeVrTmSzBhoDfSWbP7LQjrpxCZF6A9c+8uSCZal+GEVNiroXy8ThuVzg8wUvR
u5ANUp8kJgOWmRmPdSQvCBG8cHfrTSK7v9vosG6RHvyujTgjAT2M3bOjf154F2p0GKoRPkak/0Rm
hkVLOC/h7bQNd0ZqOgW1AYUW3moAQKu6CPnjzY6wUT8Z7KvmaRAIdj3pknUOpNxg7g9fqgCIXAKK
XvAb0zGeUIqar9gRmhEGF2AF6NCTftNW9caMuud8wtd+liFpjqQibdEl8WK6TTlk6hvflRzpaB0e
DZMIaoWFQw0aTVI+AgCNIwDHR3UFFNQUNppDiRnns+H+gPDk3GJGfi6jGE6McddOxfqd/+WpVHT+
+AA+lQWsY8TsbyHYkh9KjKeAp6ZlznEkUWteWpnreMn+d8gfZ259X9RrBVqSe/xvTLSUlUwVnCMv
xWaBiq3dgnrCcvMrKp23kj/g60Yb0cEIeBhyG7VcHU1TXKZS0tkcrUuP9xR5IvC2/RrC/Gkyixsh
YzlP8/Hbl85h76DSIj46UgYkv76pFG4FQZ/zIhyqNv3JL/kj6EhP00uM7JElNRlAftyHy+wnKnUe
OYtRxNwWveZu4CJgBBspy4XjGJDUIB/Xzk1g/N1FwiURHWpxq7CA50SN/glvDAHr4FiHpEgatVh7
hEpMPAnME8JFS3zUNhUVT+3e071uBTWtdRypaFoAnmNU6Wl4NIyvlOHZL1yy3VM9nO50s8BAP+zW
xul/QxchmKTztY7smJkXkk8WGzLCwt84erYi8YtoGntWPDQbhLL4j1OoinrKo940yLshx6L66TNt
7dF5xFjqafER/o3EIsysX1WLaF/iXKzOME3evTBpBZzyDX+uh/aYOLXS+IcWSHUYdw/1XmRizpfK
iaW66wk1lRIN/Xq7qFPsGOwlbAEX+OvQRFfM5dWpb04W/aRFL4hk+H7MtQCvyW2PwFBdpNQSuouQ
stcTXf/hdRlnii+qo/9O7t4sigO3xxl2pS13CU11aYs0Pwt+4gizuFtY/pvgq4873iiFtA5/pcUK
jv+/4E3LECzAXfMyMtxjmt1Y34ERBo4BJPi5RwODs5LCqpCTRdKchoMdYttSaQ+OGqAnWLM9BIaw
kpfE3iyyI9OK+DQf801fO+cGVy/E4zOJ+TaSBTwttXNNFH62yulJf+cPVT9ZmGJCuw2G8/8YIeRL
QEpiGZ3cVN4DicE/8YN8q75BZR0KO6t8oPwthK2ptK8N3Awy+5o+t8aF+gJHPwLROy9pfHX8qWeA
K60y++9Dx+O/UVH+dNwxmGuhtUHyVCT2I4QEEA2P37t+HULVnrgiK7nZ+u5mP/LaVKt2jTgJKgEq
Hj/hNse4+yD+Cw8MN4wr9/j0g7SSHDY43b2diWMOuBh9v3MTiKjCHB8k6j8i2cm+ocXq+6nyUFgI
YR/HokvnAHQy6D2TmL0jwGx8t09V+VTJZXwcUFZN9lrUhpUE1tirF2K6hL85MwcyLgsoue1tkFni
rlOseh4c2Bne6EJVvbJZKwErhyc9pEXFyV+OoQ5oSr3IxFFZ9s0JqcdZ0lHQZX8Sk2pu9ghzGTxL
kazI9hnZMn4Q/EkNB0/cGoYKyTiSLjQxS7YXgWM4iHiDD/MoXbWKYTRUIXwntoisSNIM0z5yO9D7
C3QzasHgm1+gG1HsrW0EpIysNNa3zi56ovNjzmg49LNA4/iyw6PIg4aYA3tLJ4dkkIQm2Hjy0Cbk
x1xPd+5zemm/v/4AX2Qn6qe2d9uaQY/kq9g9iIG1Cs5Z765sWsRbYiV+DogsnPt6r2Af9b2hQ3zQ
UieQOJ17hcd0bVzjibub63GxOfArTISmGkTE8OUsZ6UprmPZ8NYKu7R2wG4iw60YLIaV2nx7Ucya
Dc27fbjP9Cu35tT+mcIRdTrxC57zGtfq+Gg4Elv6thEqJgRMMyRAP2SrcDyodTqOv3OYboQHbFz5
dLCFASSH+HMgHYuhYRamc7NRuFA5Yt9X+Xv0OTpYxIXChzPtQjNKM4FXwY045M1vTGFTpcvP/o/s
YZfPJpu0v7kY+arJiX+D7wZoJni6uJKUpdt5DuejVet9bxfpwMfTpAA3e5mD2/vc77UnaRZAte73
jAJWVTXqyXsKALyX2PfygjjQ9Mk4cSPdXy0oBZJxyQRl5qNMqCpj7Nk7JslO3bKD42sTgI+7CayS
dEgJ64rWCKWpJarxIxM7BEfcvZL+Zxgw1rj1r+7GOOQsi9NwlbU3wPwrfm3JE2Su31vQ4dzTu2/B
IMv8hV+bfNBzgfwXuBQt09P5I1jD/Zq7eYZUGUYEI2zQ6j8hCGaHp0EWdYfCHzLji6qN4K7+bjzd
D6ejkVrdv2pExjCneyD0+gG5X0t2xbU0aK0n/YWr5NaU56CeogWYQdNIUEzifTuzvkyMTY03e/os
H1FC4lPqTFwZzkU/FvlSrain+zl91fVu5m5T8xx6GAmNGEsqcEqKBlmdU4h7+MpYDztTnOs/9zSr
CAD9vJl6ITe5nHx1jETXoYSxg6CN1YkUufRTSoSGLu514ttNsvDf/q2dQ6EoApmQ5mzqkwND6Rtw
8wb0brIugQ0y6bKN9hblxVegeM39pjt0bXDIxcHx3PkJ18vVThh8kEslyvwAAgJBwHWzRsQChNDg
D57ZtJlct3E2QSZP2DcUFH7dp/I4L/85/lsIH8JTaelDCjojC4WbnNwZF7OD6dSf6eLOdkEPEZGh
Yoev0Rx01ffGWHmKKYEz3vszGRfGqGzjD4SiSEllL/JZ3CZEX01+/DA9K4oTF5JVRGXza2MG1Ou+
1nig7yIM79Z95jy3qdXDDALTFFcstMDnw2CAN58yy8PlRulUlegmPj8N0y2bCv6j9ExHK67agF8u
JfxADjPEUfI1JwTe9r9ccM4hrv1suinwljKMd9JIxNAYwDc5aY7gPZ7QqAGCQgrPvdg7OOC2mUew
Dvdn7RtSKRYkt4S85Wnz1JES0fTuy6aoLjF0v8CGNQsJlHK+MioizjJslicAk4VSOwCe4RolcWDp
f0eZkM0CfRj8S4u4Qwk2I4WYdV+BoOS0f+BGrji/uXzHaWdYgtz3ZKWFlQrrSgSNIVVZUYb2egIZ
6LSePHVTVjZrPgTaMqa99f6Zr/6nyTETnTijafVynDszhRX8NFadBpGW79UIZlFcGeA6agaozHlt
vpLrSjFq9wl9tCA9LWi4tTSPhwU5hEG728LXJZITfoc9e+7HskkqL/MCdvwmIEo9+s0V5nvBMG+h
N4bpg6CTWAKYx5ZnVpfdp7kOHPheR4N/rHK+0eHJVOLfoZSB/VMqAg2uTMF9p9B0ugJWBYVbhCvT
iKl8R1YFWmi52OUvSJNbD/0UYqWAu/dl3jX8S2oXMtuT25bwi6RYct1wpisBODinkFvos9VK0D15
MOCxWMdkSg29xzN5WucbJIWi3cn6MXpBAD3fTW1DfNvuF2idYpKhq6e1Qpd6TctGlHdZNhUezzhm
acXiMNdzr2enjA0jMuR+og8Fr2qETL77YbUmV794zQit1UrmJg49wEfnGFqwZdycUb3+UvAiv0Qu
5svIh854ykwou5t0h4JJqSsMf2KiXUuxEAB2PUAaiiikgtB2MF22/DErJZg82Z5XX1qEVAO/6Muv
6yMlh4AOxtz/A2hbfEGbSvlHBKpw0d2+dvndWa4Do51lhhjrTH38M/5N1MIOFAKP25vhNtNFj2B4
KKEjxC05vMS0Lq1a+gJAYowg9z/1j6rwzL0604TYlF2/xncDiXv466oSEKcD1cLnb8ZLxP6dF987
EULK/nFlZuu4a0LjQ1Oyh4FYjTKqPMU7/0jGHDxJKpdYGqrlve2d2PFsB6uNpE3M6bdqNrP5FDfs
i2C5ikg//Go2eMC8cp1A1kbnJ+Z40YVWJ49d2l+iyqTNCDA+BO7bj/TRtpxYIBA8XFRu7yVrpcSS
mpR/869yIyVCmqUuZsUqg4uYdtqP5ojGbhTl8ICCbp+/vwlMjU2+Jc2mYOSN2tEnZafVaD31y4T2
yxBLMik6HStsF7fNzDpb+zSyMkDumzLi3LFyAfiHnHmy4CY92TUNazlsReoVddfaxlrvh+Uuitrv
jf1LLQMtke4eVneLc9BmI2497JGuW9/ivMXeG/1jCgv7700KCreZwZWKE8Ruu6KHOzeQFkMO3rpb
EPcBA2OITRreApidqihOPss3doZj2/jL1CDA4U5VbnO+88vIUF5mxLBf54CsFrm9zlR00EZvxO7n
e1Gx7OgV0TeCRr3l+yGtHQgWAkLA24lYokzFUQ6BX1DoA94315pXl3I4OCgr/SvhKRgqWmFFJdXX
HxmLfhs/YGg7fC9rqOmbJ0XKc9t5w/i6YPkJqXLq/95V06dBIphi+AIgGACWIuqJPEVvpwvKALvW
HhjgZeXLZWsrC3mTRyAzyCOgqFd0l88OikxG3vblSJMI2zqb2b2mbXyMjvipuySHABvBhHq3JM8m
PQ+C9hzGIIr0Ssd3WWvPTBUcD3l4kK2FKBggVeJ72BgLBf27/u/XdBYiMv79xXJ4ceqd6lAaA27a
KNiLyhgutPWFXDLOUU5vkl19M18SqULlAqtS7hfX6jeyP/o6HtWtS1Ouci8riohXNw5jDv530EU1
b8S6GO/K1gsGmdrFfYb0MqD9wRh0EyRuVJJZIIxg5gx5FpgNc8dLzH8EXUaSlz0JJ1GmCLMtMrTB
RJJW3PpBX3DyMdqcuc6S2k/Z/LjEZKjE6Nwi+BNiGHemY9pOmXIDOjLgPuT5sK1VnAhvlQaJ3Jme
HYZAjk8Lwd2agtEwNQcTT+4srWnmxHZne9RwgGN2BRn1p6lm18+pCM3+bN1dwl6fpvQm9olPdMyU
37t/9R6hjEpG8kNDUYpI/QHpd2uwLG3q48OQQ5SACLCsVLFvuaNDjjiy65ncV5UEPUT507d1QTTp
tOtge4ZKTukXYCUuwsNDZXnrk66NXlEwnpE/uSQ7cyEX68m1M3pNLq2HTGEdgoh0HkulxTU3PrBF
vjSM8Nf5Rb/XwywXKgTVSZ9o0eDaQRpeYN/VE1S0e+9VhsVthAk9hDroqt/N5B8FmpZr6/OPW/hq
ncqxkXatIaKaY6RYqtiiJEDBC9qC3PQ+rXehtgyyyqkzXN8PzpsFoi/pwR6td/gz+Wrnd+NkM85y
69QQaikn1xUsiiwZi+68ZJp/0mvLglLc0I0AQZM9B4SeoAEkGGXIY8BYwH/1aGmJAYJh6Pv5TnX2
5FX4oD0lBPPjKewK26GcPM4gXedEgiusQ5EvKa8ucUPJZfSFHJqMDH5Kz3QT4wvCo+ikoD4GNP2d
vK4I4vcUMf3Qex+wEZoFGLR2BoeZ563tRSXKYUDsd7tIvLEjkNPJCQscvpAGjQvTCZnYFvaY7ocX
UUOiHAWLu8qnJP0wakG8zlFAkw6ShWaWXNIQNvCKbM6Z1QZ50znLj14pDvECVH+rknAjDsEO+Qml
9azv/41FhtmknnH/Su25qzWghKVfg5OOsyzlgrPQd4BzPqnwU1/Ihq9thatVE21Nx2//96Gy4Gw/
mgNJhPrc0xoAR+87jyaOYuQrQd1TS/IC+O1o83YbLfdXlMcQYRhRRUDLKWEbjpy/JccclqFcTDuM
8wGPpKpkgQYQt7lZQ8mAvSvnbfZUZJyLElgrLMzFFDGdarALMS8/tM0eyhtyQhoJHFbjf/PM4zQk
Gum7cy0hfsAtwk+HP1B2riyvFCHhqDVaBaLY6dBMfCGpiODbbfnIqf+orPx3tly7kmMNoTXVvMdu
PvElIa1bvckqYVU1X2Tr/QXwIqkV6ymF5gZuWPfdwFGDRojfrFgEU8MQYp6x13fwGGCr7CY9swB2
PshjsfgWFnhMp6MhTvk3zV7JxUTCuLnPLeiroyznEeSlkRxGKUxzF65lfE3XT3VxBZCsaG18Io1D
NpoIhcgpQNRhvSU6UDGWSvH1JqGA1Hy1gxBw1XYbqT6CkBhMs7LcNhMmRDk4TobUfTaUth1hBuy+
g7j9af8WlLfGaHiJkr28oVjUHRREAMYlPrvirRGFUW6UT7rq8NMLK0wGd3PlD7gOeOGtjDjV9Mrk
3OLqK3+dCz0DDi/VQqvVhghqDJ/JDbLtvhXypIMLWT7p+D6Tp2VV2MhYDRLn+T7UCFA5WIe5uUKI
mQ8mK871tJHwKnCWYLk4vuvyCVY6sZQ2CLsqeX8A98JM7I/Sjrovya9rj9RQqeSlRGqPxTRTEU8Z
csQq5WN9GAssl5629FlNjQYCzmYHTPABgVPgzqMOSMyx8t8ZjZI9RkyhrOnso+C4/peVQGohYP7+
8YfGrVn9lrUPOjOrWkEP4Vdh0jnAFOs9sak3asBnXK0GjxQA6N0msxUflrmTjiLrL1wnBfV1luqJ
mAH1fsaLYFPamSMCjOzCswj1frhp94zt88OYvvHXBUMBv0GLfqUyYznVvDJfdofpUOkCVXNGWI4a
Z4qScVeUWutpzJzXTP/kf6DW7XaAdV27Yx4rh8ApJdKzvX3lqiHdxqGIYaRIGr7vaOI0oDNNSApp
gEjE1zioAi0gpgDG7jvXRiemuUEllDA3QSpgYX+x/GAtaIXQJFZu+7Yi1DeThD2hctvqXzc12UJg
zT1AV+uFcAv6Ikb23/j61nY4UZhp7vqzdLhvamppkbocfPFSGYQdg8A0R62ZQ5BE8zwR08LAkV2m
V1paUgy1L/IsF2z/1pUPh4Ul7XoKkc1EaaJZWTt6I4xOFLm/4mi67tXpohcol+F6w4h3UBe2qj7Z
tmd7muyzDEQE2bMq55UrSqj2ui3VajOjRwN0YeoHdZfx/Z6KQ8WKMGgQ1LlATVgHEWUhgKrJOmVc
zSqR+mvZl33eqRxF7qPTuYiDA+34jOcJtmN2qbC5l8s3Raw522ui8g2x4iEuRtMskBSvdsKjzb8Y
/ggYsYL/7F46+ssRcwMHCYfA23GXO5e9St5OouHAS9r3r5XTZPcv+xe3MtQj9pMTQb6hQ4MMfYAu
EQebxSF/RoM7dcyUGaMjo8eyO8GzuyiuYbNQ+5kY9OC7+ohCVOXGQTYF+IhIpxVmKYc76KihDDt4
V+YsUUKitwP7hek/rcC6300wEYw9O1270f+oZcQA3sCwmRSDgppIgKudX99Q3f6rLTCIN9ybu4Fc
VipxHOlfwhjHx6UUMEw+49Ls6VKmGqm75tiUj8iul3W1QZbFrAhCIyzHdIjyORo3hmueo5rb0AIn
d5xJY0bWKptnTqJKN2kW+xiGHDvPJpJ78hITCFXGOgzaJlGfsn1I675p9npZfbDzIJRrfaW45ECj
P+a18QmwcWzXA2DbLA1GTWx7P05AICCqYBH0WG8tic5Omj1XxFuBETLRuvl6pjHUFzeLsGeA5NEw
MFSH4EcvHJnajDXdLqNTYbSVUp2luPesuGX6roX3gz38ZsCqPjjwR+93qJg+MOTHo6B3gBvAtA1h
Ffz+9eQed6mZZHC9UECr67x3pKR1F2ZIBtoP2j9U2EaZC0Fgy149cyaraiu/oUmJH7PopkUT0Rlg
ey6V+rdvKTTBv2lB6JIq6H+OH8poluEn5Kebun5F0s/r8nsHxYbwOGED2ggzNrkdPuvlCeqpyeX8
nh97fXpuizrLKekbut9VqS+I1RiGGJZtphg2fOgF5iqhl0HMydv5o7CykAO5blUCDMPi9O8HlXtj
vPJgQD0VotWMwm39dQ9F/bf+7JtO1Hf8RIeU+7QCmn8TxNw2XopRmAR/rrtLzc/F95eCDyAJxjuG
Q5vVA5Yg8x4NJ9LbKJu+FOh3J+6dP3E4QX1RTS4M8GMTPqmv85UjMUgG3wqkpGt5d/4SG6kmgByy
jcqgb7Mornv4ChwpkkcuPyOCfzUAlpg3qk9MoBBo4+8fZ9He1olmKddvsKaiPvUmLEt1VYHh/itT
emPCu27yINHHBoUxewONX5+5T4zqLTK6uxPdqcLROjcNPiGLTmv3pmNDkLSxjfLu+NEDJghd9iJz
IPYDrbNH5IcJ6VyTZ1/t4ecC0MzU3WyDMZix5PYxrhE6tlOZhhtglXkencZtaxP5QJr3wSJaLj7v
mXXwRr5XBaIrXch4nRMZajebl+qRPZqIpi9LfTiG2OrLtrETuHwk4uXAuik+o40PiO787BWXWZkJ
Ldm1Z7FdJb4hbsWdRIfYNV7xCW4N/mMlhibCIi51u+YR/yjBPqZ45t0dNyMQcdxs/Cym/IqJ72YB
HNEXVT/ec+hl3QCF3gYt3qTG7eD1yk8g2E1V71hnJiynxo+t/D3q1xpUsN1NMb7t8bKMEpBq9wv/
v0/TbJ+jAFGK3Co6Ih9+Ug/Gpm70/UXQ+m2VZNv4UT1VK6KyWAo8a9N97ky9XygIwn9weaUosdux
2XJfLxYDrwaENzMyXPbdWNa7+V9wAFws4aJZyAyMM9jeAo/DuW8JC2W/R7/iR7ybmXBgR5HJMvpu
tI/RGsJDJJNU9Nopew4zklDCkeEwqGrhcQprjYir7ZYO2/QiDFlphmdVWJhamFzhd5WfCI1oTwnt
HAgI9jeLbR8HVy1gxrarStgLeFV++MFCtWVoPKiFVmTGbzL+lO1325PRptNa4ptZyccFoiRHM5z2
VQJ5DU/FJXLCDiLyg73UnWyjomgKEv/WNjlrszIe1AOjmI+JtcGTtVLrwvm4I/hz57ARpTbq6NR+
2isCRhoVabSQ8zVH4YMI7pU8bvvyqylRUBm91AgA0CVikGdHqraGNWlLnn91X/G7h3cUNhQwAjrn
ZjcgCuu+wiG48/rpgqDMsbSlTd/dZZy03eFFzSayj1IUNbPitea/SXOiiDwJzEkz9e9lBPLSYcQq
UiMUmNb0MVKELKPw545P5E9E1yGqqjC2fIovVjqF8Xm+c8d+ZbTB0Uiwgpvdydl7nPFPUanoGCrB
kANQSnDA6ce5dIE0wa+HHDQtc3mc68pPrvzT6czZ31ZE6Kuio842XsXTsSTCRh2xN6vhHbHzZPzY
19sx4n7Ad/KDBHkkK+zgOUCSD0au+G67fIfShNvJTYQ0yCNs0QRWLKjfEDMKC2jiproYAYKq6b2g
fXRv2f9DTSgbgPIYdnlRtEK3M2K6r5msWtb27Xe2EKo5j4KSoCnUR8QcqZenDNRwQrmRZkQ5EXW1
cOdwz6BZaYC4GvPEI5/jjrreTYVPMjEZOiViQuPcLgYvJlPZ1mthL1Mr1BD1mkLwVS4kyAAM+duv
gGAb73ZabkcrPS6+FYlPL7w3HlBRaGe4aOR2/v+yWrAlCfCg+p7KT6MhNRQARCRituJekerCwyjQ
HPuAPga4QQHPhuT+hoJG7/I9VriiVjbchSxHY6gkaIGjpq2rifr+o11VzqCyBFGxQwbWYYdZewUQ
bwxOYDaegb8k6I+6fMHFHVdiL5EoXK07myLNwGrW3cjojvORV3bXpOLKNMcKR1bTM1DODxnyRaMr
htsoZR8FoHqiHoqeSw6yqgE54XWrohPGLTgIo2WPRzc+D6nX60YMgdxtt8laQFQjB6dB6ccZzEe1
272+yoykzC06jQQtDA390zbbNiRCW139OIWyAPi7g2iuIdHyzMnQy1Rckz0Ozq2DGOUg7RtyNAuW
fZRkBncr/GxMt3y30c6J4h1jqF9vboOAGIpJULQLrE/aelaj6wYM/BVa/EL530J2HhJfWBq9IC0g
IzG3A1XJLRFsEJTdYGdAJBsC0XYqwNDHKtcntqzIujfTEg6KLB1q/8RkbFvFUSyWcqwXhqTMfQBg
FOZTHTmXlun0b31kXK8EKX9jIIa2kRGgh49jLSz22EgRXEOd+Uohw1LWnUZCq1x9efbCGy0/1qnQ
ePalMDqtMLs3K5WXvK0D9TKJqLOIt5jjsB/z+DgmGA/uxolHwiOT18c4vMJ39lSLhzmWKzc7D9s9
yefTIEeEl6H/B5WlwpWMReAgdL0sMSUhKULGbAtxJmkzyygxeS+SEBTxpHhDvcA4mKBCGj53fk5g
4UiKkn3pB82tTH6WtWjdqpauMHcz5wLjBp3G8SFh1dcPyMh/03kZcxmJB/CgZat8NhJdcBbuz4lf
kOF0wtI69+iYIs6fF3rwbFMRF+blidpJaxE9dqD+KtN2Qey1ZtaYeKHp61HeBS67igWEuBmqwDF+
eHPkQifz+0gsl8OJ9YY8MnYtX+ZdaVsUpF3d6KHUbPjTHJShufqGNfBdt98a9R9Slpva9+M++8en
o0pFcECdXLCOScAqlVBdlkdNsxb29395tXdlsdKebAKXRZS28SvztxyLLSTUCONK4F0PtCpyqjVP
sNSMdkbXpB+2xhbmy5oMICoe3ZuzMCcOxkBe4qYVq0dR9+Abhk9zllefi3/q6jFoqHZuKAti71bL
bZTbgwpzw0nenxBZO3kyKzhIV21sjMIiBlSJ/6nNAw3ee/6tUMXEPqCmW/7+SsmAeyDxTAVBv977
awYZ9sM64fbc6JEdFy3jVex6A37ylNSkKg2OsNBhGyCnUnwsBavbQKaOo95GvbkHA64+JUeccNCW
D4SJk0Du55C0Mx0jtyGIrktNXB2UDMG9ysLp31USFNlyhXVbTCVXYaw+VKBBuH714HFx32CDGl/n
lSqZERIcnyp7iLyX3YxPDmhmX6j0lL6bXX89yQGuFSKnJX9bqX/2FUElQCpQeOiIzAmxxSw1PPVo
IT26H74m6mDF0z+9hhCIQbXrkjNL0mqpf6+Ca091I/ce335HQWCLqz/CugUX/sr9CTFLUUbbNWxs
2YazzGqsFVRyx7/JTINvHSmDa/i38SUdqWORCvzgHT/dI4h9uS2UlUGHwzfJDK5oCLr4hJXqYrpZ
i68WPYiUv1svz2yQeqFX0teeKrIBLvfSRTkTQSRW2bj8kJSZZQLs2X2xF/ghdpD0N9TiTmfeR7A4
M+R7MFbuBStz9c94C/kWsPAmO60vVXLRp6e0NzMrMqrkFPSsEWt66LdcjmxtsgjvTvfaEhGmhQik
GLlYoD2Rmnid17wXWSkcTIeup715SB8KVhbOwiXqNU3VBMTvr04zzPyJqyd1XJS2izt00ZCjGvGJ
e+EbCJrk506hWyZYCqwpRWH5cYumLUm2lPN9NDQwlfk1uQUT6ehb1qFADWQJtLWR+BPEhQg4eISg
Iibm8iUbaze6LJN9Nh1j6kyVSjUBnghmuUbXQA2Tru0vD+90UUzYYKy24ZmbV/OMThqGqcryshuf
Vg7uIS4gys7T6obLkFSLWSb4UTuPWW1DxF4qQYONwrodtauPxWj1d5O9I0qzkWC7UPyBdm8QG96i
C86tfmJ49oHA6oB6HuIWEeEtdiBB5YMlLYs8jD4xWyedoTKH4EfSeCssQqIslMLfPZrBqAUNx4Eb
LIjnHvfsYCutzCXryhl9og4tY+JdA2nneDWeaKC5m4HXZOgYx2W4UYNtONc7ChIrxPc2qxTLvWcy
jy+/YqKs/xs8XXypdxjeVP0e96omFvwLHbF87xkB0c0OY182MdafbNtSMvm5dwYUyiipH/AnUxY1
DMvaSzjIloiN9C2Dsi+4nUrcpKbvHo8oQllxadGiMrD7S9sk+oMSHRAixN51fUnXIl2hI9Z+5IEn
kVtvn8IsDxG1PA3k0Hjprpd58/H1E24r9as+OraE8rYcoERyPWL2TMwumrAXBmoHURL/ExaUN2PD
6Qp15jxcwmY91J5PepKF4IzY/3KanHVdCyiR0g9ULa6ELM8nZM0auRD0GNWQk3tEIHZVRopPABRc
JVaJ0SnOvTItlPAsxluXIDFLOuHEDxNrAnNP9KU0YtPurLzBJ4KSacMH8GF7SWoB8WGf3hySm4Du
KmrTGfypcTa4HWWOzg4BJNwuaP7fuN6Qz84qHYKfUg3NYC+qOoTLjRx3tNqf4UZEZB62gKNVWxOu
S7gjtTZBU6DR8ZKShlRGU5loo7mwFCBKcwlLLjhonWGRnfmGR0V7UccNjl7OebnLUhTqJqkybROX
duz/HVscygC3bodkglUr9lVae/0jQT7p0oigEDXcdoU7pDrfuoQSRsrnjM2vIMsHQGBdLkxazyVU
w8eGQJdHgxxHmfwnIt7fkNXZXv6E8DQQxlPPSABdOHz2d7Qx3VmS30TV6WMNwi7t2mvHU2QYlV9x
L8K4WtPpSdrEWBisOmOeKiC6x4kXq8l2ihb5dcmKtgTduMyievNsRZOTntIbT870hjlmtWvLzbAQ
+f2tL+K9bKQsaxZN5PnKqz8GSFiKzJuLM0YObQcY9Tmir4RC8VckYwpXGXyWS6+OUjJdJTgynSkv
Oi3HwLi0uF0KzVUckrQY0lKuHu6nYY/gDMBjncCVEGySZ0q0X8Tg4EiOsc5bdj9+JphBUiOp49xS
CY9v5+1bzKqqxGBwJVgYPId6C8W6V8zuSc2aNIrvbL27sW/uUB95YOXjeeiiQ4OJQlBUGXvg/jCb
dTWTIbpnpQ+sKulotaZqWxLu3mXAnOzyehVliBRhbmZGg4tYYTNPIxpYZgvKLDQ0pnJsjV2eU9Og
2ZFopjnU0D6dQnNxPD25KItDLw5T2JzDMZaw5LP5W5LHGfeZaGGxnCf/xE7lOnln3JZbKSOiJ8bK
lGVN3xKTCo85rAELorlAKsGewurFfjptOg47LafniOltcWcNGEMWgJ0bNeLgAp5prAcjA/DxmRVs
qHlfHsYPEgNhE+5v6kfFuSoI40Chgwpw6QTQnmU/XJ2cAt8/V8LA2NVgVs6jHlSfWQTjp8dYZLxn
XusuCFa5A/8wPWF+8nGUoD4OoQFF/TtlLx1KFjnxoJh13blv12H+Ksktsh/UvEihu+8Xry6Fdoin
4/RSRcjf5SaFlNTG5xFlUa3nB+qKqwG6j2MQB8UD3J/GXW8ziZtJqh3d+SB3v++tlvB64+jvwHWa
VnVKF64MD0UPiBMOIQmUjin0KgokfmRx+pjBHtv4fQSmatL18/YlIIC907jHC/KYtgqZ2d+VNaHj
+5OfbOJSK6nU6aS1EifehD3uIG+F/qOQ3CrNDxgXhafNoJrYvqsoZnHWzf3olPfeG0Py1I0Q3L4F
h3AiNqDerDF60siIQMGLK38uogenLBJrQALFbzvuYFJ3zibTAFMENuTQpWfGUNyvcoO4k0FlZSi2
q2SmkGNBYDi3NyjTXNu0lp0m4FPpVj2Kc29q3rsU8+/Nq7l0VLg4y+BUbbJAcQuX1BBkauVvUHVu
2h5qYhU1vLa+3EmIrErQmb2Lok3QEtc/vJpQ4H/HzNKNaMmIz7hBTHagxSNcgmbrBeEMdUkLsDl8
g3phv8bhRGRMZRGbK3foG2Ga8O91M3RCfyq32JokI1ppKZAuARVpc8vJPAdJMOamt7hc1uFFI1cw
gs8+/sALaB8/GmuNk4f5+RAbNStBHvZGe2lIJ5Jtc6LmpkCtmxprglrmPSv0Yt9XCo34JI4jUNex
xz7KQrhnnrXfnyMl0ZSN1Vytv5xE1d2ACCxHhRdlv/3L/JeHVriVahQdtMGR8Qn4tWSwon2QTWrh
imq82n3YpGIID7RDLxihiYWizTWvKwJFd99YgmCCJhmDvHvSE7csjPlEGnj+Z72KuXzSxND3oEeX
+nI6OuOKxs1JIqjhL3EQu7LJEihqWwNRLZDeV6VWljCc1IzUjssKVQ10UVlZrOxuGtMVKxrpCzBr
oYdXc55b/aI7Jp60zXr02/xBUxygFki932bUkGfFjI6JPFPmpsoUkZUhKct8BQABYWxzD+iFgAht
rbslVIijj+pRDVOIRLDU63ubQG5gplmlPZSJk5yEpTEo03hxRNJthR+RMIP5/YL/DgvWpzCnL9lO
ejBmf7NBhuuQ1yrKpQsCTJdRJan42fPqgEYqA8rvL7whL5XezyD1UsprZAGfhdSQLh1lXfiA7I6t
gFIrHfXoDB/9t6RfUqpFtPeYyBRC5UxTFByJneKBvl/Rzh5MrUfKcB4/7E+v5Ynk0w0jXD8+6k1t
8S1ygFeTC0A4BYLI/s2QWzAf3gmxU9mBup1N6C+mlyfP7MlDITaZTeQ2ufJLA1qTAGMKfp49Pzpo
084AzOYuVD1NyNOs9Aroe7JxDTKjyiUmNeoqsIM+9fMj4rtnXiB14JWzERrqjPZPmmlfc+bVai7L
yxNqDMog5BDFYDLo293c777Uby+jBtyi33K6SmF773IiKhZ5VPas8qu8YvRvNOm1AQA34nBEKoMj
BDsFAnFSsuggWwoKpaUVHcjCwBIxp1aJasYBMpWiuJiMzieaL2vrkh63/MpxJgakKi5y8k3Z3eed
zWytYnliMn6ataV2WLLW4cdTBqlCaqSh7FZDxmP3KP8kRZp76bpA8aKoR9952nU9XqBmBOOBQSBc
7G2erZrO3iNJFyFuiNVjKR9TafL264UPH4re77dtrXn3xKcGDMy2w7cPgIJB/9jvz9pvLrCWRwVb
ZztxtwJ2Vuwvyr5LHjXna/MG074vNn8FuH3kXYOpkUFbZuw5s48jl6SJG3XDWhMzaQqztTCAoFUg
lye9Dvzs5QEXoav79FnSPukhaXBB9zVa+6u7lHSD+av6XRs/+HT357yJ4I+EoFnnDyOlNu2pgl3j
yEwxdaATmHEoVIBwyb7UVnVQB2AqZL2LTXy6JlOZe1u3T+dIRLCx59pMo5A03Cim/elAOs4zdSdH
8Pwhy29ohbWRxbr9RKlC00GnvD8QI6tangv/vTqdk+3jFDbnSZVzZAzAQGI91sbgWIeChmhatYSq
5AI5/rOS9l5Az7ehWl9siWl+Fimg4HVXkCyxd1I1hd4PVJZRrAxrGQgjz3h+IDcihD1EluIDHqIj
7oh1UbRp1a12BaXWZf8j0XeicHjRWbtgrJdKfhtbYJweqlbJ0kIPlrv/ADOoHg/mLurlCLPSvzgi
LZwHuagUXWocdqAJX8pGaGAAUltIupaRewDtJ3a1G/6bkpJyUhSGJ8BlSNQamLA949eD6fM/dK+H
4Ex+oePJnJVHgfcUCypBgFCJrMnqRfD55t+lvJuD4IkrfYA+UzORa/M27AoA4PdxMCeJ8mVVxQCH
fALL0vSyJ/zObwcoQqgRkQy8njqhKc4crHrtUXwvK42f2XjAqFSCJlE2KYnBQvhJdBr88y/xelbJ
4G3hinHYpXze2bFM8ttameRB0xmcyLTFbnc8cZjjMER8t4xKa1modjy67FrFmECvMgr8Ukh1SHec
b4OxzyYUEXaOk50CKq54ILj7LA55tizcuspjjS/ihtWnqZTbK2D6Lu/43OK73eOHRcwTi3YDc8M7
yDwSZQg/z/3V3LW9RHEADUpTrPK/Yrhr6rGIEMFaBJm8madySi67ufOdDyPcwtHq2BvpZIGr0/+a
uV1wpSFpXO1mKNbWgH5qrDviWQBbV8gZvJY3g6x8VBTeabByaxnemeztScTy3NUFsHzHpmR2UY7k
9F7bc9aZE4DNDJRtXu0TvgoiWdqF+w2TtOR+KL3B3FJe1mdNNCnQWUEjBvvv2suwskcAhcoVdeRl
f8buZi4USxx0Y+3K/Fn2HYZA2MYMND8OZuhXVO6nyhm0JnsQEqmjaCq8Sk2TxpAFfQqd36H3iilE
Xg+gb8buoeuvpwau92WpB+ugO7V2OhpnLyh7YyOcHR20JqE8Pk6Q3uIBR+LkZ/TOyxXYjA8mjpvO
l0TPydP/464GKmOgQsXRB6kexzKCTzY1ysWggnYSsAqNGmsAaR22HYJmna9g0qTNxgwc2XZCd2aE
DDS5BdpDB7OVhoZ9dACEYZulvcsm+JpRwDslZQCfDXI5w/9WQh+d8ZrXTpWG9BNlTtIrt0aa49lP
3ghQ0cuKjFGFVO2CLhTCdpeU1CRdeCbBwDq7H8tgWJ7nxk7EI6XoSEnK5oHQ3MlL2fyi0Z5VEo3Y
XOoPLamjHO76Pu0cn6md4I7gPMe1rrxShMlcFDcwmswSACa0EvMiHjYDOGJPsgDrxxb7PY168rC0
ixjrGgATKuFeWAELc+xAkPbP+xNwNkjXUW2lilnLndELY5dwACH7GnBEJoFJOQ/BBlUu8370rGMk
y4O3HtnLDIpYRxkg3LYUR1VKR5Na5t0F32AGf1jBw3pEidF9ejZExNqEj2Rd1CI28FUkXNYaUy1Z
7VhExoryJHhiINETNG0D4yu/nhZl9wtj9qmg36ud6xbFKgWmuQFLmyDq5GokPhg8HzAuLaflA09P
/0owPqTMC6J9qXqYvQzNq1O89UsE09UPxKPH9Sqbnx85x532nzrreOen3QBrCUpZrhY1u9FDlQnC
yxJbWt439R6R0roFKcpz6l0RD3flitJA2HjlKZnWlwA3Q4pYyTUeT7ciiMgxGgxxuz+haq94B7Z+
zZEjMTPiPRyDTFT3JQ6bB3crYsEFuD5pnTf6cm8EsbY2oA32xfZ2hFTmL8ZmQt7TizN7+T0iiSax
ogNHJhWmT2ZR0dKh/igPCl2KeK6S/OKYYiMtFuhwVOSoIkPR3PapZD1qEmogfAVNbDIZ5Do6YcV0
TkCXdhni5aG08Qyq5XQZ/7q+LSNn8lDbbUYJ3jJH5V5iKy07MbWSAuqk5WPYOV53Th+ZhAe/PbLi
bM/2z4Jkft3YlHKyq1JKNBVBGfVkvZ1X+S/6GGfYPKYZBD0eBxBbEYigtLGfVeak2EfZfEOYHIKd
Pv95iPlQurVDV25gWy0gyyB1qCYuRYir6qpXdky1xEmpYcgHMW0ewhqXM/MfZhRgXjiWZwXO3amk
PHxZGR+NqdV4cvNKm5soFJAsrJKtgyQLv2Nk2WRCGRGyKDEm177t2mIBFGrFEce9FaWEXSzazPHs
MblP0wsStykpe4+zq6jFImiGuc2K3QhoGo0WXK3h5cTox+fyiyhsi+I6gjQAcqWCzkvW7h+BBoWJ
/Tp5rARABXUy7rkQtrn7GbTQoX0WudtgBaD+yWE8/JmTXWGT7N/COfpMCk8vNUtOOnGDd4EZ5y/N
1ptUuQeJCzm7NYXKyhx/PTgEHI4abzu1PGLMuZvkTzGKhXyXXiiJcysWEHYVHV1D2JfrPAZ/ILQy
n8+m4FPC4GRpM4kCRgwkvFh3MHydr2IuQpROBsENbZ6La80K+S4oQWxR2u2RXV5gjkR3ritJovEc
lz010Hy0sESVbhnfYrR7N0rCqn3lH5iUaF7nqRiJkfcbrcEY/e3YAC9w/CPmQGAGk8LB8zCMLKrs
JpEj5E2HeY/GwA7VqXEJckqYxfIV8e+JRYU0jNIISQuUl3yMRlXNRY2+472uzid4JDQ9DTBLOHLq
mKgP5ww5IxqXaJAmK3BQLprOgB/ihmgnV2/JCriQaRZBl2kVvQRRpv9zVzEOYUSE4yrZfs62Zs58
/HemrJhxU2yvJ+lCOKh41Jg8UQGklxK/tYPlqIHd1n7gB4OjpIIsDc0r8ekd4bTUyGtPaVck0BqL
rN7/CFVBxoV9xVGfsneX9b4qLCRMq76E28QrG/b1uwBpq3I2wrpaSygN1IkqCR1DYow5jCcz0ctm
PQmR5kJx+jOGpvR8t2eijuu2KGY5jEZ4UHrmlWv51STR6PDLuUMeZQWSnaiWSfzbn5FbTHf/malg
ez+79TEPMzjV3/xl6rl6mCyMMCqSivik4gygNmbIInilyW6bZCs69tQ6RobOj9QTv0e492RMXX5E
PQ78BUFHBqtIKXvTHD510GP5z2CMGpLYp/gOKzHTETHmNdJCz+CHSnC3AhjHeLTQ8+6hPJb0C1vC
D2G6Mod1LOWzOGTRRggKQh9X8f90ZUZaXVxBIjbJM0ZgbrYN3p2Pb7MQAk4K7k0hvav3C9YvM1BN
ilM8ZhXAJsBrDSbD+lqEOB2rwOq+hcNxlVikaGuX5VWMnXscKbMtRdhf+ckYyPvnXl80Jk27szL4
BUItwnUCOcbU0YjX9MjSS8XUsejVE8HPwOO9e3TwsojPS9DYfhggU5jH2w8cx/4hdkvM5x6Du2K1
qU33x5hKHs/IFxFrsNRJUxYxRacXPh/VMdhGIoWbCh8fsfkQnyEDZgIwiPSC3RYNBRup1tQvGpX+
ifD8VfkIwxYdhtgvU0d+3vPO4Hrv1vZAEIlrznvenDwSAyrO9kuP3CS2jA/lEYdy6x/VR+J/Eogl
hZPP64DzKkQsiqd6f5Y6Gk2nVKVmX5gFdR5K2feQ3Tup+oc6NL6QXU1ZVSWdedQ5edG1T0PiTO9c
Bkm6+VjsA+IkIAoDO8GHLdWa6zTuv3X48ApZLA4P2VaxJrDYw1KM7bZOcbI0sdo3i+m6veBIsYN3
+e+xsfwSTtY2acfm+sEDWrVUBFZ8rvKt7T5ei9bYLzxKiefQ2X5504JjcO+LqdJYnTqXKID7QvBh
yyp1rFo+zLOq0jUAcX+VklMxrDTV+S0+WJtHXpvm0S/s26loXHOK7ftEUqsWNPiRY7qyVeVBEsnB
pCYml79fJ8qTThRyBJ2sW9QFyOdWcTqg2Lfp8pxPfpcXPkGD3HnMwzj/Od8s53sKaWawpDtKg6U5
jfaDRASA27v0fzN4515hE1czghIaLvqbX6Izvb5fkQdlHslJ4GSFWf3Y0GOt8dcNuBllTNCgn8+F
hqUIq+pwTiCv/R0CMgYJpQbSxI7S7KEtnS+P7fL7dXonCE5eZjkEZsOC80oEJeLdr8Ha273wW3jP
ejTo/lD0U9nu2fCbAMii5LlzbYx8/M+lAfCVTelc6n3AzNqh6yIe+W0mc5FnrumrW6mcpzOiJSbd
/PvgEVGq2eyCmWCYXl1CSokO2Qn7lwuEmlYkDrxp4vPlrCykmvnK1+DEa5zMgDDr7fldSNqItWwT
0xsOrhqFYtxkxD26IWRW5TkqGjW0Paz+Hc7KQ0fmO4QBmHRE5sUjLiD6lQ2rXAf2jAXcb+pr5zDP
nm+HAnFeBeRgVEqImbJ5VDV1NHLDoOKbdodk12VHzcenCzpH/2IN5fBX891QiInFJAc6UUOyChk2
Ak8HXtxXPcscu3WdK0IlRsYnlr4yCgDd8PnpM2+dQsqVKkYPkdwwoAhZoK11JCMttXceu2mduuE9
sEUMpbLtlYiRThMMs8GvtUwJqguKbLPhdM9PvEpAIScBnbSwUtcO+TezV9ZBVqFLcRysCiSxHIKb
YmeprbZRDHEOjuyf9PZ5/XOEjCPYrXlU2AxY/NL0GTdnXMLuNfwtkSUyW/oJck8Xld2oK3jg5HIk
IwCLT+p5z9QVydMfXfJhgFC3IXnFuTvCjOgvTyP1H25uzhgKr46weE7hTY5z320/P1ughxafeGyd
AV3PmzOSoaXfP9ICie+xRM/6zCQJ3FIM/igVfJgR8T0gaeRM7bvDFEYS7Wpw6BEdH885jae2xbax
QxBr6HYkJ6JD9M6d1Et76H3ZtKIG0cKx394VNYyBu9C/bxj5YBYeoP8IMCtlk8PI1qt4LW5Odj0o
vVrH08UTvW1tRrtlhp8S5O33BGLDRgLQJ8nLpd3a425O9Bow97S5PH4xNFfnwFDife0i3G4ooSM8
UFinBXVwcEWXSzyprbvGqLeOgj7CUh6fPxazddLZxZvxTKNAako4AxwtqqRz6i71+xsdQ6H0BE0k
oEVT9DN5vdBVl0qhhYdCbtK2eYuxDSelbjVUETcJ0UggBUWkN67CZKEvcFq18gjAQJGY8hWSEi2D
tHjNuXGRjDV94UTlWnDrxZ2zkVJnwTu5Nnym+mxtWNK+Xx7XDt+NFK3b9jvRm9vhTlXuAy7wOghn
Yd8iplUT8c88Hob5j3jrbXwRsF7h4I2JGIt8/eCeLxIqTwQk7x14pL/udTXCD/KL3rG1ijgYxkD+
Bq23ghH5Osr6s/BkB8EMNDGrCNLvkJ1LVOnhVxr9dNr7ZlU2ERQyTe/xSfRURKcYaQtI77YuMHOO
m0NeQKrlAtW8QPVWppi8jRq710ACdi2ZVleeA8jJh6Ay2p8Cc+APw6nMKysyoLgeMpHzrvFAfkmU
xTMgPa4R1FRBT4LXT1kT36rPmD70QidRg5n/PtnndttGJc1bb6qn4Nde7+VlPDjuAsz50IvJcIxe
ZNrl3opDDe3SkZZ94BKE9GkzN5OV14PqxRXjP9jNeegvNMXeYKONHDFGLQ3z2vO/xjK+ZxMm7mrm
5OpOFGe2jXZ9IxjWhiLZie+abdnfbbBt6QMEzqdwJzOVSLSUMQtNF4qDY75k3aj5UBHje3KwpU1G
AtGpTjDiXJghD2BOCaIPMjrJ1a5lHPIJ7T63yH2XGomo/hhGKmcMVxmPQ+tY2wXZuLvSK2reCN5X
ONNuuXW0RyKPvCHtCKwBgX1+kqF82s+M6imK1WG8hV3zJ3WkmnE1Y9tiV2sTCoZlmcwHq/bPJ9Gj
vM+rqbvBAL+92rzkhNDi4iZQeLIs6OVD5i8r/iKdGCZFECam8KFcZ7tskP5RIXlKjqv6ni1/QmT7
He6n721RxCaNwo2PMXcYn+GsVSL7lFctiZNSeuNxs+BQ/RmFb/p+VgxctZuvniaNFmag/1ZhhPPn
MyRUUZ9WGjCPZ7E2T7t6NkONywxUtym9jLQ2dRh9qoPLbHqWYJ2wKmJOOAx6SAoKb2QxAdXMYQLx
UpRA4MNTVKimyet8hElaFDVGcbOKoiKhofR6k2mGGpRRDMQE1vLhIa3230TRUX/haaDGDt1TXHMH
//3vE8eLd96Ty/wn3cQKv6+Urk3QVMO0Dje4apLI4tJ9cnLOz4g84CAyDOFI/uD3bI3D0EkLjo30
5mtxtngf1VrRyI5LE9+a+pA4wtiFGMDjLR79Zyb4JLNIXyiCAzEeHCcN6grxX/nwzhc3u+II/3Kq
NuvdEDowhblb//99HYQgBGii2HxZkMr9W8RfEtvJvW0ialkoNUQX/TH61IpwWJhs7+AxXQJ5K5/z
+E6GQt+rJrXzUQL6orMH0bOXF89n2Vo8lpfWvu2TvEvvLojqYSCLiToEv6yN8XNpIMHGtaTZfheq
p7P2gCto9b4jqIwNbtYEXH60BKt293No8zvVpdbC16OrgkOaMrGIJ2+3MjdpBV5ThqweBscLHTYW
yDGiSLDtbzbJOy2cIOXEcSKWCoQuZRYMY8+C1dQBD/2vHys+pwcAOQ4CTPgMxGdT7Tf0QVUOhlo0
yFl1eDa3TO9BRohm2ndjM6rxZTtY9WfLBQRMRSySFdDByHOJRsso+PZODzAIfiS8CDn7LwKOs+d9
ewwk/EDIaTjeJi5c/2WBJ3H7Uhe34knrABXnKjVMFV3J2C9QLS3N/p91WzVqnwwY2i8DZ1wIVcCd
zOSYtz/MUNcCPgLbR7jqfX5aXyjPj+7xBbHiALX/CZBPieySeA8s6nmXCQXSkK706x/VO5PMgtIb
V8ydsHw20zzlIFo7Z3B9ne8CDyJTgwPnrDlJHua3S7cuwnV+1Pg3aiCOTdZDsNwDE/jqTsdzfYzX
ldj8PH+0DziCT8RzJ3Miy6RQcbIugymVEFe7uYlkm8XXZ4kf2NjbpcbhKUVB+1FSeHFyBnvVxFJi
LDCWT59qiBVvmch9QxO643ZlfVrxIJrjGLnFyYil14UNLMvSA6dNPlHjtbMVgetxSmdGmyQIwec5
oYtC3AwZrp/CLVe/hHBsPJPQgRVY2Snt2HHy1fFm4xoDJFl1Q2DEQlsEWbMLADHJVh5A/MPFavUA
mssRlE864kf5hPAq6VwVo3XFtW84jYmtyCA0SuuAQitl0gUeNrpUgj3rC6F01zTWPSTF0K6HX8rE
KL0IraYTe0GNTJ12Hs1BJBSovRORynlO//0h4ff+3dsdKOLqPRJcLygLaULUg9s7QFIAbpsiPLcV
HQg1sMdAAlzONANBqCLNDmiubC2355XLCDP46UPK43t8coStfPBpzO+OFvMGQxaLsTOf2lW1CrKy
dCBAnX6CFEyiYOmYr16S/PAHbSx7w159IyhVRfPQddQwjynRi8DqfB7SADNf8ZOfeLJZM6ucr0v4
Se14l2yof9PkIkGa0wu+wX63jx61Hc2ywUHNX5JzdjY/8iRuLTDFcgHWYUmym1lbB9H2EQ2Tc7LH
xyrcD9JdWVHkOQFGqo+nq6D7T9E3Ru47aSijpxm1eaC19AE06mP7JHYpCoMycM7Bmq5T3PORQt1o
rI8oeaO+Pfc2kB/Zryx6MJZZMBkahrztj80vR9SLWZ/+2Nra1sQ6FajZSf40JkrgnhiBiGrw9StE
B2alKsR5UV2StzM3bPkWM9w0wE9rB6nHmGWJVQGXbP2cVmIV+s/IaoLf6TKmO/aopjT5N4OAdQwA
N656f7k4+Od8lJeIFx8vH69wpLPBERUVK+fR3D9QWVlyM1lRt1p4gegNudGkrwAbDlyuJGkReivY
OAgnBv0AIni3PajLiodVeMyXweSsfWhR4cnEDqjdQAIaNxFQg4gq5MAM4XvNKoLxYWNWIH44hcFO
lImmeFAKO+yc7vnQ0LzOPyoE7tx8VRJU4nmPTdlwmMQ5WZoA90Bkxqjf/R8fq6TVpbxtW8Esw9i8
b0YnM7k3K3ZhdRfm4wW2i/K0EX1+osCPo8EXocWZ+ce8uVmGQZJ/14ZWLWQ6okY4kJaEEnRwjgNU
apRgYJqUNt6iGB9O6aCMHA+slAZqqZAgJIGZNCpGwFO821VCdySMwpRSpFll2TVP5oFDe0X2nLsf
FqZCiAimipPrAkQopYUXKmm+oplEzJLaY7F6ssc5KAyKwwVs210UFbLocUhOOATyclt3SF/d+/wZ
mqkqJBHBM8ceVw9Ni9NmtSJWdQ2R/Fa+pfPRWZX8Eo/Xu/VyMl3ldPw/Gd5y4eOY8UrVK2jStUkK
OP+ie/Qfj8I9gNbSOynaD68oJz3faQoVnGC18o3S5tOSnE+044+Gea/FEsLAu6DRZIfeEtjIOey4
3amUyoMlm5UpDkzj3uoKiMNho4fHISC1DfN5AiLVKIdOsChjofw3zEupoETJjuqTTzxnWNT/PN7C
TVCMWDQt4whCWKBb88njqULFcsjE6Qre8LOGzzgYDjCuf4/drOYEMgAIAGZCsuhPlFDVhxz/HEtO
iV7hui+V4TJqBHFFyLvs8FPbXFle3C5r38P6SCcfQabirhqCtD68/mrxdyxq/Wk9lh4IG0+FCFBq
X6KgeYfJrte5g6IAlzCwiAGJBFZNEclxmSeZ/hBGFuqAUNqF/HGzn9vhFWB+1NCcx6/KcOyXq9ro
ZkDh3OHEnOiAkxiIvtsu397YxwHX1rWSLEBi8vOJKFV2uCRLeZR75QkhQeT9z7xnZJXmS461NejP
0m5BsSGcw3Mgs6AKjpP9EGx2FDRBckRUbY6n3hi6uCmHYSwrx33PKpmwzrsrzAsVOUZA9OP7ql0T
9ztLzlyvZEeJlnuJsYh4MP4itdG89CBtmakLj3dcZUUKmtdrz7WZDCli0mFqkypMzCy/39dSNGnE
TEG9uyTFxdl18/fpOB/hk2jaLBChqsRgbTjHHZYA1AzS2eA8KxTjjYLLHWjY/k4y1y8TBEkwuyn7
04YI9tTgGgwSzRfoD9zo6ZjFaJRIZ5CdbtYGk/jwmKHjY0z07CSyKVk6MBpyD/GSLCQ7Hxkxbai1
WFYoS/NRXaLRDL8CbNMR7qYFAK8WyqnYw157CV5LY6y+A2puWZYNjuvSXhLXI3N4QOnskgNoViaY
GM/oD8feS4Va7hAEYpxzoZW8fdVUilVwqHsEElTC6AjL8UCqrHQ46bJE/cuNlm+2lVThmBBkNjlY
Ja5QfnJPtAUoFuW3TUkQQ142zPFycTziAhfiso26m6WjB2zXCgmDtmtCvbIe1vB23Xtn3gytnP0e
sxtywkEmPoYLrRkxvvFxRIhj7ON11COCF1rqokOg/46ID6Cm7Uh+owiUsZ6cDLKCaqDaT769+Ru7
LEEXoWKiJfBkBs7l6SYaCia7J8N/djV5t2p8EEbzaMiGa3P8OCr/X10EdUm7RxrHFRDV8NJXwblI
/MTRLilK8LQcxoJ1VMhP1DiW8mjagNYfGl3LF3QbM+t8Yo9ll4FfiR4irP+3JyUldHumLuMeSe1J
wBmv/QJ1qbn29brrdYxNBOkoWqCc7UMyV0Yz6b7uPpHuw4H+Ehr0lFLrr5CkqgNaHnzvMIsKLTiW
Vf4BxQXjocXgxgs1wtBVWTx3+ni6/2bKmm8LbhE6U+vc2pV46ExtIMgbigTwU6EvaLKcUaboCvoy
WBgyEBm4IYA7Ecqk8Pso7/8LNLh61Y4FWgA2hBc57XjyjsSesdMUfh9ifcgcv2VDHI60gk65KmTM
PLyidx9jtV/dJCoHKg0RC7fNHQ5SmZSv81NYrAXMVi0k0HNFqum9PUHM2tPq1wzHPa9g/VoRAKq+
AN7daaoIZ5kkyQxcGx2tK00Rtv9GCS7AdkFmiHcZPsa08UGQLkCsBYqst/dHk0Q4/XXLu8y3tYuA
78yX9ONe647CkLzNmypyvZOAsfkK6smUbzheC5GN7K+zfhO/L/PRiCESZawnAR8Sd/Esto7tSku/
afMcm0XrdilEpr3b+GNSH7y+9Akzg8rLh0X3HV55cxtHpY3rq+0kU2p6kfToT2K6sk6S1kP9YSrJ
5n2gOGODaqcgCUKTpMIXBW7tq+URhH/kkuLC7SuktRKeo8xREJxlBD9QFg1EUKwCSdf+OeacbRL0
iZcXKEPxpa3bRujnRtindFOoWLiRuK/VmAzkKHN0Xd3Sjgom71ARhXq7la8gY5NfFADwkP78wzU+
Y6n99x91qdStoFZYhdWj59aNz1yvhz83J3Qf5QvIjWe01uDuGTEu/02qF8MgAyRYeyXp2TT6EW8w
9v+v6IzOu57WLLfW/dmBm5lEEZ+T6ck0nr4tZWoYMs41nIn7K+vgDIx9sleaAu/fACVHdsyifPHR
BV35zbb2fONGj1OskTtWPENsCWo04uwYdaGfikQQd3kIhio9QyhnyXEDz7QDSQVf26UASIgwfcGW
9xlUwncWjG50QESJQBB0cBGQyT+bDtXFBtj1QDkbP+WmHgMkld/0lrPptv2ts36v2LZhhmVE0xNH
W/sU7uuHQmC/yjCLJwzltXm82pEfTauRMkYdgadMdeYixuDky+C4t7kFOX2CjS+jHpEICNVBJfrt
sCiMEbQQpc3KlFhk1umkEDKrImS/ADa8qVy/FpSvLd/8hGVqPMB35YswLyGi2lj2vWuhRpbXYerW
BNL4Nqvy6ThPSdT06nZ7+vOw7KuW7axYKOWQJmdzeygper9sqfFLc/0YxohpJCi41v5xxbV5OR2w
60uORvprYjJHERHSf04CKs4TIa8he8dHWrjjg6jby9Vo20BIhcUDNBGz1KHjqMRsMcU6OCkkkU59
a5eUUePJZ3NJv4gBnna3G1fVLJlcevEwAOAA7ZF/IosJj1ULQZ0JbvTOMpISTjMFdieFevuTbQqx
lwLeVj32H5JGQO9VXw+H8tm0v4ee2MQJfeUNoc0nAYno/8EF5VqWfFFCGNtxM909UAvrZAE1SHKt
AlDRWzbOqswdLkfPLAsbBzv8v7ahHjuqhE5EEJ9Aqs8LmV8T2qzYeKXZ+NHn5UBNKc0ZK94h4xeB
HtA2d6T8ZjrosnWDQ4MJooERCBgNHF5oozAX1xFkPaGYQpwxnANfPDVS6QlcXWzVKmfq/XHKijS3
zegkzSsmAbtUFuwc+i7mewc3aMZBVhQpICvvEj/jwgC1VHmhjcDGb8pe5ZgtR7H5zEzU0g8H99MG
TzSb27tca9N2XvqrlxuoZcJ3JkntVKe+/jMsQtzq4h2Keqp1W/qt0Q3nAcJHxEoZYERtHSQAeMUU
vRFsJfrfKk85szpTzj+t5gQxklsfrH3ooPOm8gS8G/rxnXq2ic9w8Vy/oirQIrhxRRjrbqpOr3V9
v0Oe3PC0BKOnYAW/7AaiaKYHRNsWItrw/sAS49h4WJabtPa48N/9Q3idEqbR5RPYPmGaGWA96L+I
vq2TAVfO+maquzW+neBsPkSz1M0bA5B41/ncLJp0gmxDsUM7Cwv2Rkw0dH4kOgd0a4NWDTkyM+Br
/B+AhcBbR7Sk/SgOEUKDsWxwv1Etyym9m1rxiTrAwqghDH9ZvuPwnDk/R0w7vjciRpnuJAvRa9fk
uYstvBJ5ZgDrbIRppoW6ZuROxGCenpTNjHX3Xl7bHQkxcy2qS1tTW1vZfFviZJXTMaQoR9f3F5Tm
uTk7LP+rdzaS/Dqgrq2Q2O8BB3r0jG8uEsC8YCa98t2JoyRRr4vnCT0CSmNJhG1NbIhSR0fRtqfI
iGzpkP/Cg/sxCPBrvTrtMh7pjdsIKAl5YoYSjHyiiBUbjpG4ae1YKJZsAlwTrO10gCc97yz63v0C
MjkLI7878hF+PHFnoBKaR5eJTvM9lcQ33Ac+xJGzb2YinlhK8QD+/MbST3srx4UJz85oh3QWm12G
8iUQ97wUjy0lvdAztyH9w1LQ+9Y435/pvcRZIaCZT0rFeC9ZKgEFhReQpq1pMwjtxTR4hz1DOtij
lli3P8lMSXw7OBWgdzaywrKBbM01k9NIHZU3abe/oaJUuVUG++kMhJcpks2sjsQeVtI2NjscUIWh
m3ZTketVaDfOTMQCadXB4dddotSygKyZoJ8byk6IDf29ySbj90YV+o/1kgLiQ+pjc3ZV/DEQEv8m
IvIiV0X3F7v87Co1d0G8VXiO3Ra6lqqvxoEcY/YbF/VnVAs4gMXxwS2kWpIS28I23jsIrfJLEvsM
79pBTR/ZbWBHVbR+Hu1J+q8hltyIOhAFZz7khu5Bl3QZgu6vR/ceHJBORZzEiVSHzgaLuQrWMLrf
LbyrT/d2wdUw2gOmlKiIlwfVc2qRQH3MTk7MU9Ej9CcK8z+P+4VAmmZjq90DTDGGvyfYHOCuRC8E
1Rje18/+Z1kwqOZJfT5ARZ6Z+eUk+8uwclP7KVxJ9nLPK2uYbfidSYOTajPNllFTBMN1Kftn0cC+
DK0yOrHJexKT/QOo8cGM9zsasu77O7ukpb4gARQRNiGe2C/c7ds9mcSHOKbfVPiUyDuri29voOQZ
TROpUvciLvxn5o8z5krRK1mxb9HeFLI88kgdQsApt5xCh4HA/QM3anDdFxxVPjVvJ3PPSZwiGjbN
Yq5QyUkGZYrmIscbUii+5+ipDMCqJkRoNSBHnyHdWLQk6+vsuAE70Gr+ammRvRBAahqzutp1grUB
b2sV5ZtfbDbBz5pnjoDQDJrddkrfZTOAnYR4Z+79J2bvVVZHWWWKLDhL8UZY1CG0lTPjndFajNv3
QZMN0krxsd95J8r3uUbwpYnsywdd8XQGjs0keD3OCZOGS89CqH/nne+AQQ99G0k3RzLN4bpu97t4
xqMV7H/HlMlFLiO7HvzO09EPhcPj873rhau5w84PKhUYNvFXv3e2aBLm4zCdGDVzr9pLTCYVq2Ta
8+gNAMnHaXlIcg2v6ecG26Ly51dpJhb4rizlD2Expij6WxGAP3dCPxnHRL824FBkZioxBVVtQ2PY
1omcuqWknP8VyHAYAMDtxxJtpZcCnyr+ggEiE5VmcN0hGf3hRj5JjIP2niQXG89diEp8xDLphdeV
CwlmDhiZA3jzNEnxs2MCsy26gwCy4DjZw18WVBakB8pMxbkaF3mFEzuYG0vJtUUzrmMHmRnIVzm0
CcSfise0gvS5BqqWGkmkYo6k3dOFYYKJ38xyhh7xk7AsjOdKuQC2KwFu9UzMYhOtOBAnbatN3rxZ
gtkyDAmrIdVDbsMQsa0E5VjYFzpE/2QJDD3GmXU4SY6lIaRlNOXBq0twWeKJpRQQKBC0m60A7IKU
v3qXC0Jwk/NlTad+COvU5Fz6ITz5LixhVZf04m3HcTbFTUHALJ+0sQMw7AHyRIqIy3m3242GnKke
wTRGl/hznlzzb/FVDMNS430fNJGeo/GzGsdo1t1Z6xXobvIpFKIqDLEiIHnhWXV0IHeHpsEeeGcA
9/6lFz2ptUN5ddyItxB25hQFWbJrYw9BzZT4r8gmui4VAgcE+doCDp4m9ZlplVh6t+bnKqIqbQlH
sr/OTNArvw78/Pqa6eRoGMXEjIDNXNAq+fQ9zo4AyAOE1zRT9MF7Ji8/96rLsByNtSxx4ZHZ7MK2
6W7tDOemvEVqBYFkEN+JZU9eMeLCqG0oLeorsyksScmV6dylpH1qQIboNCsQZ3/PpPXfbREzLIFI
rwdcdYnbMtngPVqNowSeDcBOl7pxJIe1Vhq/Fx2zDD09jie0CgCC7IMElyXdgWe7kAL+cQMKjIMu
kjiYcWMsyYZ0bEnGVtvoAk/+NhasFQ/fk5zi46XuSmtO5F/Luxh6ugrqZzihZQGXQQdTQ2tmIn1d
YeRSxbj5N+50lzIXIWQRQ3guLxC5nt+iWZXDkv6PdhGEPFQKpa6qEwR/gkuQ6rES0L2cWvxjbT81
mgPaWlp3wkKsylBQ4l5jnwQqMlSDzPJqagLlMy81Ejl+puH5GkCfCzZvT+juV90wkTwODlBtRasc
typerDQsfI3QxO8c8IzAKPs3Tu/kJidFamNz8rfFdweJucDC77dDtCyedmBZT9u2Q2tMrYs/2CFk
xip3KmN7jp8xQrtGKDPwVPuFL/8hNiCZ+qVO9Y2dSFiJn54mqNAoGJ2LEiozxhaXqeaNkmgsJzF7
jUjFfS3+60sTMb/sghQvVBgb4UMKbie0KN9PPBMY5+iV+vxp3CitolYvNd0dROSSUwbyxyOn52+g
J0hxDMRBRlNOw0Iz8HhUR9hEUta0b04WHBXWfNT9zwu6oBhc6Tn/j/dVJk/MctqkdjfJ6dCOXCyO
wrCjvKFnYA5HWQYBMp4iWYJtledHx3miZV/whP1G2SWHLeAspndU0O46igOMFAC9/yNslGgBfLZ/
YPiluQEbMHk/i5amcW3AKvKEZq7Vi0IU5eKqXbmcGoF48SNk2RlSOhTb3YEbzZvovHHVASIkEXpG
4Fe6EprvKiub8aCpHbQ+owjpxJB38DkN7PCZV6zYhTQaaCg+5LFYcMERLJGnyYHoywRKlZx1nft5
NQd2L1pK+VMB81Wfs7udsom4mk3fV4pN3JTwYNvgLrqlIWkDulZVpvXNUAJdRm2A53ujcPa60Cik
gMY70A9ulLAx7N8m2eUONhi0NLjPCWdbeFg5e/Moo238rlBeW825zoHNUfIRuYcqskohSboodfk4
eE+UnJ54FivnG3fJMICdzs8Qav2TEWiGf0gtWz5Hwa6DHab2v8DSfND6RtzKTbf/vG8frVqs3j57
6NsDIxgwiizpyP6OgkjBrkbTjmX22m7nU6uvvbn5MqRBjh2Gmmq6tS4QoXJOhal9W8ioN9Tofgpp
zmNm9uwrmS0fYyU+SB+sFFfKA1n/2XeRoZIxBZhIONVKfHIvDIZZfu3vuRpm/jA1u81XFwxKoewI
Z+jAlP1h+t2RhiopQoV4LLeC0LJlEeuM9ymKaL8nBY4JxB9e6Rob/QolDB0xObOJtRQHYFrZbZEM
nnuRsaYLCSbBBToF9HOHrpBmSgZCLyfzJXaYXGgZvn2criUwippaC9PlKH2cbcsroJ8OSIThq9Um
gFNEezieYcpXYO7eF7FEXvwD4muwWYgAds5WZsS0ei+D0Ucb0gusrooN3K2zeCf89RpOzGA9nSZW
VvVnYa1N/zlljjnLuU9BTxH2BCJuUeQE8E4FdXgBIB7hT77vfKtrS0qXpVaj14/vRXd1MLPLFeEn
tgwaqEObR7nrd72CnI3VBQzMNqUM2Z8B07lqFiXwKslYu1oDM85jtbiqOx/KSX65lJH1tB72CmQl
TjiPrqc1xabO0HSKNLfvqNVKOHiozfXv7zR7dayG++OnjBnmtAKSK4/q4eK0Uv4s/AXY9YgVyFj3
/1qNcDSqpjIf3E7/LhPoYkHjs4k8HPcXvXxQUOsUg+XRrfI3jSFddoNqN5BFBllML8XV+C3ONdCr
yMB4u+kO115Xx40p03TRa7zo5viujzqLrL5zlTl954n7uCxr/QIlhVb0d2CdYBs2iBCPJAgli01N
ivWFcWNr0k+12MDhbVcRfTgFl/A8Rb43+K0LrEsig/eacX1ouYgjn82/Y8rOh3THAdFCH2izia+S
lSRx7ZpxSUWp35phPr5lyw+pbk+STSOq5ppDGwvBBlh5bd1CfkyXGovBJ72weI2h0sHsn58ZtiKl
FZ6BVq+USfCnWHcLL72j039UqgaUU4IH4yU/sgEDfic+0bO5FVaYEmo/Io8M0umo1x9KJax6pGVg
C0hMFQg3ut7oclJvd73SUsq8EFZH1FngQgw/VCQ30TVVArPAlv/tYMe5yc/zd1rO2lk1TVG6i3S9
RIkUHCZq9bagkNB0pqjun0ZoTBrHu7BYtGnFCtJIaM997eb6O4wo5VQaDDuqbf6ZwJyYUJZUUvWo
ynmvm/ecs7YwDx16+2XqjjnMnQCDDZU8lb0kO7KHiSeoH9yRuSzqtWIt2T825ZKPSPg7Uswnv06u
wchiKO+pSPa/GYbDQmP5bU2ATbQyqkJ1pe/0B7kGP6sU4mFbJ3GcjRkoWNSqZHGzQLxnJN4Gg075
Q7ub0LC6gvugEguNBHA3g/I9CBlPAEUZGzzea4BRkJFFryO65CtivBa4hzsYSVDLHsfIJoiZZvls
RjS2Hl2t5cUQfZyHAT7ialHgAnzjI7Lw3nfi8aTnFJJExXIP2Zl7LrXLz2208zBMEp10NbtLNHnf
9ke25Mm9aJOzUqG/z2aBQWjYRyHyy4FUZwbW81HYIfXcpIToI9b/dCag8b9G7Y75y7HY5Oj2xrMT
rWdQQxUz1JpkfuRfoIDoueEVqbX+3nWOCJa4nINveap8p88GXUi0LcBlzpfCVCQp0d9mZphfsE7T
MA/4vv3eaN5SAxtxcBKohhCDnxe61FaAMNWKTcgP7TwDQMwz/GeLh2nBj1zHIsvT9jMDMwveJpIN
QzgQmsDTDl2HplGYn/ytNDcv5xq0/ukrmXGzGdS9DGOBMHwntsz44STEiGJYKuR9k2UcR3ql9SAE
HzhRkItBkr1bXwW1dbFkb0VNd8ekbM0mfn+eYm3lGreh9yKnPtTpWZSEXTbKpPDiBO1RmkUpew0H
TLeWrwVb6iVTx1uZPVqksSC6R1OkIEIEDkgP0aAU9XjWqjuDAvrGuoHln22PFrLW1DLupAnoWG4O
XHiDgEWNbqFmIzN6dFlxHnIXSWb3kDv9+wA8cmyn9lEIOb3lO14GtOl+E2IMjUT0kJNorkSrMAcK
MA8diynmAq0imZ45r5jKePiSXTWhWk7F5Sqq9CID32wSp106qUexpI5B+VIugzGXGP/WRDyp+g5a
Awzk5KoFfZFlA0OOh8kiHxId/pRbsKGv8j8llnEn9uY640UygXFEsxmcObhan9X8C7Z0fKL/+kPD
Z7rxtkZg6qvRtMvzp8dOjDXBRYd/OLwF3GjNae0LOpEZBkEYvAcfNx8o+MkDSnzQoQmL5Ogydhyt
Lk8fBefVbLTRPBu3t0q2MtaruQhQfK2DmK4zI4v2jNYxbcThEBPphA29OBvKQ2YTPE+az5j2LSZ4
dTiOA0OiUfL6tprtVLT0iMKje+KAsWftAc1oxvOc8er0f9KAE4Xqv2EGHK0rd9oHSx5gdPDuqrFZ
8B7rJMvcgFCgl7VXEdayxLuyej71KEirDmrQLFfvOsONbUYm6x0TZKPyd85OpowFHVZhsG+JI48j
pysv3Q2qJZqpAnL1aXWqsrx5KjOr8pbvmueEK4rHu8g8d2IbJlOiJ6FMRpNRAsvwsTygsxKJ1lX9
zwFOBUkRa5qa2Io4mZXGpTQ2UAVhwa3WAuyN+hqKxZx+hp7gwQNDIjEFIZdMFw9f6U1dwpnVksQo
CJl/e7Dv5QDMBVa23bQKcuAbEUQC6XCWzClNqDeT1j1z/7gelragkwTy2h635RoIu23fOZIxAoou
xJuAvJ2PpoJR9Ms5060AdY7rtV0mzCJ7aJo5/pRan05kF5jojT0ynJH1Co9L7Ky7Hwq1mb5wtHVq
L9rMZixry57/nRZ6QejHrnNLi5Ow0WN+1wFyAAptJAdzTjnEv699LM1KJ5/dZNoSVuQldcFVj+FW
iIOkb7CvJL0nRmqBjKLYWTA2zxsFia7nwVBrxOeAoOWblPUxLJf2XY6P8E20rHPBku3l9MV+R9xM
0f5RVdm5Q4S+8PBCO2Mx/CtxI/4Dqc2MRn3royv3/Al3xTFJEGsZtfdZt+0U6yZ8N54MjyVm5mF4
jLuO/ZDEGGxF3+h023gAzwoTAkefiZceDQr7BNAhJDd3T0cQlKDKVy4fCa238i3vurv33mzm1XuL
u06WeGWThIySsP0le3sMAjEsbGUdGS8v9vh+zhHP/DtXHS3fYuH1w5snehYnb2Uxt6Zysq0Sexer
GEhGFuYowjDbHh+fOVyme6V4vj8v1FiB/eEEkhwlYrRLG5hQlQjFk4lN42OzZtpCMKg39o1PjSYs
8rBklbpqDWSEEEHiuyoGmvzpSJlXimBzAZ/GNRlWxdXJLq7hD5DM7KPr6ZN07XYipNQHp+KfGemS
wtm0sBITPiZ6iyY361eb+ZXWmlEMflYRQiebAJ4GYF00+mEBlfzoYAxnu80sP+HRALoaTIA6S2zu
XA7T6nBdAxTSEkMVgNTEoJp1tmzjyDQhJWfZxoFBOd41qB9w4G5YnQI6zLpMyKnYytC25SKWhuig
CKXKz1uinjGjYxkWus3oZ/ut19P57DQOtuA9ozmbB/nM/01CgSxeN8NdAG8D+6Lx1hhduthucSc7
r94o5gV2uyoUyic9gEPPk7vMOXcqFNyCANlnE/dML5xAffzQ6yohuUSp4GYXHHfDBmVkyE1W6VVL
AdE6udmZIQPvhiOsFGsVjZQ5FyJdlrsmLVaK4ggxnea7PlDqJ7QA8JDe6he45TrlYvj1WBG9mg4c
t7FhBCfm67sGJfDWiqMFV2vG6MHcelqwXX8IcNVYym/zoFGMSLauhPza9qV6tOMQMJbz/kP47qUq
jNSIiUnxAhirhNAoASlXVT06yQK8gchyoa+2bspvwRWPCmi9giwm9fYizZEy4cxzuNmT6IxGlT1i
8GoDgyo9SWLW+Qz4ea0N5U/yJq7Je3qqksQAn7a3r7AfhCzKdLM1Ohk3vl35bwy152OmZ5SHIdqu
JBRle2+6kX5JMxIFVvCgbRVhQcDneqlYwPldLoIPBBX0dGeIfy+jhKy60MWPM2onx5N2p1hJUBKN
ACvVU5jPj2YIumMcww60Wal6ouRPXFtYPDuJ1IraaDXI8y4qRZGKHKl3TDjXdR7qtvzwzKhWr35V
w9iD0olnKisSW0btCozo/smO3zN/gKc3O3vbL9R/74fICBQHJB/jaMqQXt9IvKT4WbO6/t5dSrYF
qMQZGY1etO8cii1Ty+2NuUOMH7KAzOYeNr5jVIEoqUqPfyoTei82AVMPYmjHrD8CRfMEhslK4LAq
JigmthTtTXSfnKWTjzNmsGxXVDZK7CbQ/6bAvmXaOQz7Tqq3ZHL6CIzhMsG8EnXnVpiFRjKE7qy8
1bbIQ8V0bpgoe1zInA0MwSbleYsNDn25cJyZENVIYuedadoEjJ/pXl7kxJlpD+axGRR1j1dYRBYv
2lpMYcpeiwxZPVTw9TWkq4JTvOwR5XzzrAEvJF7i7ZBEvmHq9DXt0axoF9jlgFnrl54GKp6xgltq
lfKJOGq6jn8nJaAwnlScN/0oVSEx6GLvBWoS+fE05pTOlylcgLlali1IBaelsC9WQNlmQz7hA7Ht
V8MrA574777Xn+UK94p01y3A3yEc7talkBhF9ikA9rBOUr+wYFtJZJFhkYwOy9mYhTAU+P1ZklkD
BbIyEBIIIxRJqEmcktZliWyOWzoQxacTshYQDnFm+9imokWuTNtMOulowhENl8ED3gdQNSq6IV2J
LJVrxOGxN42b+dfdrIxPwSX1qRoohQYCk4xsu2u8IGlIR1ytgdY8QZCXYl9ADVmvU6HDkRl8YAQC
9LOOmfy5SxvOFzryQ2i5bbUDaOANFdcOCzxTTmL7UMvFc6mf+qF6htYpGyy2vimPYQsUCtVtLucy
0oqLra3dW3KKFa7hiwSbP8ejbNb8BgcL/odIVTNGi8z7VOtUbdV+sKT9C/FFo4m3FATvhXxvDCoc
AJIoWIl1rV/G82cmg1XRcSU1Hdk3QiIwfAl5vu1d5BY2ZI5X1dq7cLtTNtUK9MBjIA1cfatiobv6
kgiLmtJy+oMEqczWK4ybJ7Gw79tkPVNHZZfEHVQfDvO7duZxyvdD1LbkG46gObBlnmnPwMPH3IUI
7z5fVn8l/yC6pcpQAbhLRC6kbG/AAoaIOOtB5pm2M8UTAS1+d9uwrrCX/KogCUcsPOxoLCR5BLMP
r4Ca911SyLa/NA7zvgBeYYETlB6DX2vyzqXA3M/P0npwqT1BoU3zVoSszc1gDLkIaFd9OSDibMD3
SiFpnduGsSwvo/wBwo/vrmcX6RJmEobsFfkkYZ2eL848CHiivRT4vAlFOlpEsrBhojk+DUEr7TD6
Mait+k7JPYxY32dBotv+uPKbVuTTA+2WyPfR1W2LfN0aVaIVR2YYoMRhfOB/lERLANAmTrFhM9aZ
NbvMiWWKyxSmAYZ2Mcd/3ooW9F2vuyAWxzSSgz1S+Gh1027edBhniLQS/j+LgpHKSApn0j3zZiw6
lN1VOWWfpRH6qC5wf2eoHYt3bjPev4Edo7GTVtOpxJFUc9L7xzNolhY+oCQ0/9Sd3PvNloVmffl9
Qax0iRmy0aWuzW9bL3xvS/LhgHMFkv6BQjpcyVH6UiGHvj8nf/VeGbW41HjZmKDdVuUMaxQ4oEwq
bSDyKtl6BDpcasaa2XphdZjS+6wWordG9PjD06E7ucJPl+t/FnPZ9os9IihxI21jyypMyhwtIf6q
cvwx+gFpfB0KvsOf7uu6fcFALCd2OfKAecW8OBy3HWTQ99jv84c/PwTg+P49lb+wuDdcTp5k+Ibw
QJW0MnNU8Msz8WHTuqdpM+7EZ8SkHCA6XbfX4RA8sAQuCHBZOrNJr02FoQ7MVCxzdtHcYsKTiewO
4s4qu6ZpWKE0/8k71XUHJII4B6dwZ/LFeg+BBRpfzlJCUNYH2/rN8T546Xfivfo2ITXugqthVyJz
ZaIBklUzrA45h34JoXADXiwVvr2Kp1tHLwMvo5aQJBcK0zSAgPfJS/VG0KW6Bgv107JtJesKBw+Z
uaVgKfysPUxYN/TRSsGRj0SXOSulDceBpsLvWf4fkNuAjqTNNNJCyXVQNJzhHJBNQHrZG4gHL7W1
qNobxH/2ZuuW9oXaMrxQasqZfVlMJh95n4eUulL5cEyIAEQpTtFY2JYuLZpM90CTDeCg6hCErC+d
92CBx6jP/L+Z2IaqnuiJRt3Qc2ciEww/t1KaN0bKArsXW1sf1LdfMvZo5RpllgMX5sQuQrxlX0lG
bEot8VZ3ooO1+ftMjgGRxNFuPviY1SmyWJC2nPYn/479xrmD+bI9+8fa5W0IWiWkbRxCe79B4YJS
nbxJBKGTDPn8RHqVSri+nyAQnjnBUyKcJUUj156jdRSmfTPLNRpQkrGmSPuUsh1Ios4vF8x29pge
J5zHWBtSNPqs1ILwp5kjLJgQkv3MaQcK/X/Sh9GHoWgcaXsGxGkiN9VJj99T0ed8tdBOVmFfyH4P
W1jUoXBHCG7O9yO9sh+XrVRn/NJGgRU0TMfxGj5PAFDn6u48vsDdbgmqg2T3YJdFxhooZHg5zhjM
iaHRCyFrj/yfZeiAmKE2VoogzpHBR7zY+uROZgbXmK+zjUahqV6p6A+bwbGxj3kdBvYN7Zqq46Z8
HH0uOdZt1yAZass+Oq1AqSOWSVTGEl99wlm3DOO83WX1Kxsk5+Cix5BPo95Zyte+1EU4g4+6FkhO
xKpSlFOmGuaYsKdW91SY2vNUP3xuXFTcTYfE5Nk09GHzIDQZUCDZb6pfqCgN111plTSAU7+PSsyi
edUEIS2LLIdr2vWT+AR9hcb8AE+QQSEumii32LHqcEOY3mvOAenEsJxiu0SxFdPJIAzYlGidaDsV
RFoKSUAs0HNIZf5PEq0MQLp20IjA8gq30qkxIWSRkuVaYraEkyHkegBb+NfumSyQhk5szU8yEXsd
J4GkqIOMwrV4oAbGi8N5bUXs58amVcfbGoQHrInYM1hDFNEzsiJbV3QY0lTb//KDJXoiRA2f1ANm
vZx1H5hb/E6OUN8gkkYcdIMapOORl3bEZjpZ9ABq8SMY4LNY47zJAnDmi8p4NBKH6sZyL7SN9p8x
fwVA+ZJrva/xI3pHa1bhtUZW/dkSwxFXtHIBzFzzWCGRPzpC3oKn2LU2ItrerJ/hmYBJlcG5VMYE
lUoYZIfOLWd5AW+2fwF4ebH2H8+o6zgJa8kiUHhvSy4C50kErCJ04gIGL1k4qAw1ehCACJTHlv3H
DtBUAWe/t+ZR3mRcCiGSu0xqxCtUnQLLYZ6VR51vyrdFEGZRqm5sh04wTSuHbUZTwbehvu89HdEK
n+Jmfo/DlTRBSsPFkQbuGCap3gmm88gV3sXhUVMVa6aY7PycNB4hZLa66Epn2d5BiUmHJoErffq2
eaOz1o6/6f4VDme37YcsFb6YZ4B4HibfbhgnpYdGLvJVoRILYKIY/1akGdqEfXy1WI4bLI4wG446
s56KzVFdjjTXqSCaHdKCor8nVY/hyEpAncIBs4dtBgODNW9lOw1byyMa4Ls9wV09S3LETqWLX4Y5
9JOe3UGJWqnqU0xW/E8lp648g6woy5JCD4+VcdElPKjfVrNk9WuD14uRCF6qWa8G9J59674Z07EZ
eDW81uq3jlk9CYi5CEErtft9hJk49VJudx6PLQraZ1C1Hi9G1LdHqyCpyderUtBQYHH7l/qgRs3O
j+5yxVfaVvR6fCApv1Rq1VMQyV6DwEMJGpZSjKqwkwTiqCTB4IntI9i8W8Cex6CKQSYT7cnkS3hu
IBg2vKVpBI53qZK8S8eGgox1q2pQhUVk4inugpj6vpX97cEpF77ae1FnYM+htziVmlPvlhjzB0ey
tVc5E5EWQWMsrLrnLGK8UsJeUKBnXK4L9EN1xdhzEe85VEZfuStl4etCaB0UKhqQ6BYkbK7RqSas
JW7IIt8qzo75hDrM9U/TLoO2LyUQ9/gLFKcjQ0uqHfzUQWcBOwsGpWbe/WNQ2xSPy0f2bhpBzpaS
ZnRCT755/bytZ0ax16hu2SN5TwQiAluAuoCDmgpUTKw/ab69oVYs20YDHA9tX5s+XLbOdLC+3MAA
d7E2PTrt8rMXlENJZDC9X8tFNJdDtRKf9HV6lq9pHZkBhSYZHW0WoHmisdztFA0qFke7D9X8pzg4
CsSSMFfY/H/MEGn43GOkqO+YxsSJqtObX+h6NqbXkgvFsNiXcSPGAoGSdqU0ZkMhe7MXOa2NCVP3
n9TsCxsrG7tR3wVSzl5V6JVDhqL/aramMm8l6rAt93bnsYDWkXGgUICtwPopf2ib051qWMnXoIwe
cfQvI5c3rLL9TtyPvIGzxo1KRIIRVxM4n9srrIEoLaDJQ5SvsmnI4mgeq1jCOrBgboRi130V84Ne
vJtttrglX27bH+wVzlDxzz03C6kDGDfai1666DE2PtUa+i1ehaWEPpRE3IB9XyqNsCgKnPGYfTFF
LZtnnBOZAQLjXsyN/WQYYc4+TbvwEa9VpXA9mi3bNNfZBuaZG9pyOUZPkbuFP9E/Evl7AnFSise7
G877fZ5edOIG4ncXnLo0nABsjXQ4NMtu6iRnQnk/6JabE3C51gaxIglwycHKlB9uO5YEl9gf4sDS
eMqX4rcdiK2RktEyf0p2yw3uAuTmi1ffDT+m8s25kc9hKnKSDDYCLZOM134jPLUmyaKQMQWBnfr/
Il5gKMcNxQ21wdMJaXNREwLqXgUyetR0CI78hHYoYZu9onrzUCTk1d/ChgbRm5G1pyua1ZA0c6YG
2tP60Ic8S6IYRh1ZVRQkA1ekMcM9kpwDRnqlI2RsKcr1jFwuuMx+Wk5M9nkI1SvDj4ivvwxYvbHy
OuJonXeTJCHcQ6MHoyR0NVBb7ET7OQL7HUxBBirvB35QIK6gc4IwAZSAgbu537Tzp25qHWhvIfgn
Y+Z37Yw9Y+QnFJRrl3BjCGVMOqqorOCkWE93J07fp4PWWIZXubbD8wX5LGcgy+huUxArDY1LH1Ff
E8leGfA+h1t796k7K4lZgL0q1LvDGdIHJO3B0ujqT0UR7UD/pXy1fZdHym1PdRzlqDXYD4WbyqVC
DIbK9djzl0yeRALAdL6Ll8Yw2FjwfJpcfroCGpKOBOPLia0d8PUfHCBULBps5Xo/APBnSFgv1rwy
RON/qCzEQJFg8wjDdpk7RRa+mejrvzM+nMsNrztNsgltbtOQ5CztEramEmdCUxHahB/EyiyjHGwM
XS33FJiWH45zMRPbSzH/m3Rf/A3aMVCngTDKX1xACufMMFC/dr39zESImtguHJRO4qY7ZdHOmCAY
l5/kfdQoBw329d0tL5yBUUsau7rQw5AXOj7Gu/eP3PnVcivaS2m5RLN0R8VDoqfTWQmb4hqid9xX
lvQlBpaA2MdFV2prKn8Ekd9c9db6rc/XXpyuOJL1QZl/Rg9ip1U9j1M2HY+NXUYd9xhPKFF3izeh
7Manjy68psAeJNqjYxX2KCPkSkKZCzSJxjqxvRsMvIoLmjDPHMGU2xZNWrw4BCdQQ+5qHNecNHHQ
DyzFuIgYcf5RKJW+z83nedzeGmXl28hAkYuNQ2tJD9BxCAzXeEItGvRhhibnqG5/alQMpy2jhOEy
MBcQsBq4M8a57KHBZSMT3gFgPGZBxh5icmlDxr/lXVOGof+x2yadnCrfnYi0aTP/lP5c3uxOKRBe
4J3DElZ5VmJQAJEr85xp+ji1dIoWxSBcJIIIuXTEUCRQLuR6p9v2DumAjIUmSEwznpUeqUZwgBw7
ZdovBR9km6ynRUqU+wns8VxVHeFR4HcHYQ3n5kue7dToYrtQvd1UzdpBVUohzofWeXGRyO5sqJzx
4hdzKf3XhEIDD8CvFj2HQGiJOC5pr1E6FRUtJCXfsPBxhauRcq6ut8dTovPd2VHKDRHr2jXgnNEM
kv6n317otrxgfIDgH0Ka83bDazVj9AynF3MGbtAWtd1pV6TR05Bo9xmRKpYm/f27nzvxrWXq0wym
ByTT3j6MTBj5/8pDLKAZfyI84ETiu9QmwDzRqeO2pp7oLtUFBOgnsiGUZsC7UZ4Mn1b5Q3F5AMps
6KFSKxGfFE3AMKYJ0O9Owy47pJ0w0Gk2YIwp1VLRF2C42DlIwPjSaDTzbdAp3UjTTJza9bnfdgQn
yhK7n9LNyLTJf+oAzh206HfbTZMjKADXXKLmgMy9qJYwFT5feBYgeiJWuamQYEDD52PY3V7AlRCz
CuP68MGNWChaZzkBGQ8YbLitMhgXAQhGkncspRMkAbhEsqZH8kyVsrohBtSFFDTLnplrsNkQuJux
mo0wXQxwsJH+ZkuV7ZH9WNvjMd7t09sGUymc8CCzTVa75KYVI6KGCVVdmyb1Xcltd4UHijKE9aKG
XskNs79Wv6sQIrXLlCTNF3cdoquR+KPz6HUPaei3w2fgv5P8oq5UPFr6TNwTNO6CNC4c29aDflcj
3EulGP7MRr2ExIEoPoHIRX1tW8rA9kINcYHyRfuCiU7XWSUhVe2NopidXpsYlCYbLERaWJqszgKO
tSbdYfZ1cwdls60nkvmq2iRLn/eH0lDSZO/0jgOuY3elIhsIu4NDNek1SV+Aevk9s5zco3iRsPbi
I2h78TyfNBjJEtzoGWYAvwcw8sTdjy7g3TZvpvZdr2qOIVKucoA3R1JDBKgp6SiyV2w43j9Di7Jl
JKX9S6PaTRHKIKVXznA38DiE0vM1Z9mg25CK/SsENigG2J+Kefm02zw5RNIzqRrzcFA8nnWtkl6n
vccYUY47w/3vhWADopoAXMhZbGt10AsFcdwdLyr1NUnsuId7cckENBvkebC/bT8B6dkdgLPGUbwR
3zTldZK6Vt9O/P/5dBlL55MaaYJEDzIo+weV5Hxj8GTuiVlIaw5ipldccPM0FjepxYNjaaaJp/qY
kwBr/IRoQbBzJP/GmyqUxmMYIhJGBQJnPE7dGsyqcn0f/8uEdCy2RRh99R//daMfA6SBH33bMRWD
8ALYQVFbpIiiGLTPZHtJ+TVjofUmEQC7Rm0MewcVZY6cfWmXZphYIHK4uEgKxhH7NwNmALVuixJS
/PjlqVm6cojLqz1+q0qU0FOzixNdprCMzbH93BGSjRtnaaOPWRiXYiGHkUhWhlb1aERmRYg9Lj83
EwYOEDy6A/JVNlr2zYbswtvaQV4FA5cnt5AYU3oEhPaGPvy19TFfzvF8AIWbmkz6BPiGehB376Y+
l9ZKYQcwtDlccked9Wz74IiIber41KLI3pw5r0keohPab+ucGgePcOYkLORPnTHDceRP5FP+Phh0
uBWrmRSc8LmakMtvesAeOXOYMTJJHUxZSdvhzG5i477p6NxZq9utHJjPACN4vYjb/7FzJrNoHFKY
xEZhTo4uWlwDGL5FPXg9YnUW7Oz+rMBDC6sMpm6t4lsiHjr52LIY/CKktzrFbOC+b9CDWRFGYC6N
NbrAFLUI7lXoWfpvKNk23ZNkFJwK4TcdWITAilbJN0jd7iWMgxRBEmP4ibyPsMtZ4X0AU/uiprzx
P3Ib6j/mKfsQHj3r/MJcMHc59c0WhGS0bOpHhbj1hi6K2HoMv1VCU8IvJF2F3A1hff2cFx0iibQB
1jXbvY6DTFtazmnzyksl8kwjKrUooFkKVouXTl0XZmFMOTUsvLVUUCnhaCx8o+aJDVp8A8mDwYkm
9+PdY4XHoEO1ghps9xOfG1qONQlA0uYXXlTtNTbCOetho9w8JpgnjULE7siLIbbkqoZF3zmwLBXr
Ras5ja/cavd3qoZT2qZgd7ZrZAAo3QO5voxDtAwBIQBNCfbh+1TPe9JwPuES2aawVY9QyE6sTQVy
j006WIo2f8hrpNpYEx2HWmzjYqBomEuh7o+6B8w6R0RdUmf7J9+YUIsvneF5DwBmDM4HRaaVlgCH
ba84V4qN0uNkVarySHkZ8vtmqFXICEFJS81riKWvGTUe8KHmGWNUxm45ACnXQqMjdoYFCmWDIfbn
hqQulPmlAdlmeVDaMGr/18nJdVAsVXOx2mM3OAIfll6+pA0hXpzTV8nXvwyes6V9Ch+yuQ0BXLZ6
0jlME4ox19jHieLf5sj+HP6KQYjZM3vr7XgkON0m0CZ+uF3bTrAO2bs8UPbaoyViFBMBgZRnyxss
2RzFFbJa2PiMQYXYk4NwrORXIVFsOSSTYyOpgCZxaY15Iyh9ys73+jtPSRpLcWbSepKad46oiJ68
EAe+UUqvr+QLVSGD1pRprQtlBVThns7wT9KdT5me3syb97Q0aYVwCpqeWZg3vWPAmxMlz01livFY
HySftpImJZDbRc0v8vN4tqEOqsnDnPSDYbJUSDPvshg4Bc6wDorKKkK7UWD3l7MIrSAvktW2dUnK
2EJPtjKPDZ0SXwzrTRhyA06/kZ+rQYWcY25X9KhlAHelPscjP4P7m/Lgdj6bKfJdwgzcR6NXor1+
Y4QO33s6O4QMrRCQHqDSchoETrEzSCVWkmR0lvG95QEVbmQ5P6XPCWfaeAj4nEJ85kX2/lG3d2qH
hmp3Y8eBw3yFzvR/fZ1E1oBGzBn1WuO9SdD1vmO3wEioRZjHRulI7Dhok7iaLdzrPqR8+Ne7hK4I
tJzh8yzXNtNwoCHY6IlyMmXuH7B9/UjKwpBiBcJOjMyu2BEZRAz6NQ+4rQaueP+KL6SnMijerrGA
VQAjQRQDqUQ9iDJns5KAgPnbC74YyOb8B5hZvaChxUrp6nWIbeB6YuZl7HWQmMgDg68EHQmTspKE
eWivGeHolsknyG+7c/3JYcf4F6xw7tpKAsoYJUDIHlLRIz3LnqBMbRMV6TGm3uNi1kg4eCnCB5li
iCErPfAUbv5apq8ksa98LDLFUbuKXFnXj9Y+TvbTpIBrsiH9qoQwKZdKy6bxPTSB44WcX7EVh7cL
qtABF4xrwKcQmNrMrP05tCNrWbsaHjRQtQOVhLLzX/6PB8uqXcn9JdedJFmDFonJf/2r62dHodd7
JNEwgTc436T8DqBOON2gaTTColJHuTU+6Dvva8J5Ed28OiLjv9b3UdaXNAImbZrF13GrEND+jQ2q
3pD1dd/sejWJXsXaIjkzMJAE1wDSkLvfxYIrGlcxN2wdvBBhnGkNrJ2uOK/klTOtC737AZ/vM93t
RaeETHo88YSFXJ9jia/LikRXsCOv0P4fQSMMCBk5NJ/EkI1yHD5BNuuko9FL/7e4RrI+oDiref8G
ixt8UHyOFeHG2G7DBmtbK2nF6jjn6w/SlF2I9ABsTY3q1x4Le68Qcng4hw6f4LAY52a2ATFutVqV
4WhMY5VyhHaSdx90Ra0ePmxyMpZ4wllsb6dbVDXq3R/Me0lGdAUSu7Lk3rUvWDRNl8lj1y4Lv3tL
N/LiEx00TxP8PAC0yQwMCGrErZ6AUwI/30yLzZMpCcrqhDlbhPcBImpgykMgWKb0A9ovQ2QtgdKW
Jcw8NC02I3i/uUPzFzvkq7QVF3z/68ZWPZp5rAHi7oNVkGPTQV1fwSJjDYqUnsFu52SGEuRApExJ
5nUC7QZyfU8WYEkZZ3mOnjxqAmSWVBRz9cYiwpaXbtUQybgZbrwJ+20SWPUCkS/kbldSyGn9FKWL
1PM3q2lLxe5cx1YFWusvxbM7lUa/1ncwCBl+h28zkbpDt3w5/C3oBtySBEdLG7AVZtfmdkKxBehS
7DjCLfd9yRLTLdg50i0Ar8HeaXKy6n4947ONMoH7vOg26DXY7VYkpzMoKRp6pyFyQp3BThFpk/p8
NMnfTMTWA7Rgq5MdOMzCEhPCMiG4i/z98+g4uNYbXbDR09B3TNfEySoJLYaMxBaa28fL1pQH1pPq
sXXPJdKz+ZMsQO6pYwhL/gaYvmyj6kY4iFyipTQAt+Yxuctc86vEgXz3zB5eR3BdjnalqyxAFHcO
u9LrUrXAVGIdCNuaLF1UX68h2ytjGdB0/W3adHEDHWGFWq7BsQZ8vCxyvVYVtEftLWckDbbGWQSr
J8VlSrA0LEfGriOHvtzOgWSpBbO4qzRSawCR7qg8Ai207+/Va4ebc6vDxeI7HAU2TABXqzqRYxrJ
Gs72ELsfwv1jwqBv8CUOfCWq5Xv0njxnOJKAEs1qTPtrk9GiZrWo09fEyNP5sI+jgRhVhyvrg7Bv
mh+9n5HiyIAdmYcPbCvBVtdjg4uMJmRmwQjcaaSXmjtmZJj7aOaWZbmKQbOIXsv/O7p+4p4XNZY2
PIzQukXKXez19eh6Clz8BgADlA4a3YIWcrHrqgTD9I1tiJd+q4HaCX5MyFFniTAcCqJbotLMkhBr
T97ROzJxv8j/EqEkZqdpuU19BfMg0ILehA3zitwB+Y3+XYMbE8RIBB1lO622QeZ8T67E/cSs0rCY
MNmeWZk3GyU4ENaDmEnTqGa5BM1z5lKu3FDTh3U+RA7/pe37BlpbZkPCcBPEm3BgRfi964WtCOb/
Bww+VDzzXuex7NyQCNy3/UdbdENCb4m158epzW0Ov/hbAOF2W1BAx67F2kCcpIrPI+mv//1gZMoe
PjRxAOYq0K7nikdnIaKWZU6YeMY25/C2iXOUM5jRLVFh9ODpBT0oD5d0Kft1zQND/H7K2X2boGes
DzqUvXTYOK8/DgAq0bb59cbenPdBpv2R43QMIQXSnero1eUrBBpHPrSpwmKcXW4QB6rtbbbFobCC
kmZwmRaUJNgSPpkFVDdiAxUnVWuexmbqUeJG4FwgPhFbgXL34R4Kqkjnczq5D/47hD30x32SEVhg
cNsG+XMdd308SUT7zMG+f8vcYf+kqTEryu40pKrW1fSJJB7NTi46fVdtBRhiKOVKXtN1rdjx7pbf
4mbpazGpYg3M0+L2u0Q5Oq4jo593WVqKYCwJDrOOehj81+lOII8OQcXZzUz7fsbiE1JKRMzqdHef
THHa2jByhYwcg8IcRHR9leP66ZSSSCYzJ00FePHBHWY5Y5XxFQfcrB0blS07dD0e5JkNaFEqL9J/
OKveQ8/cVcOO0WXb5cZo0blDhv4RqowqH7Jr1Io2iOZeMuZrYTQw33HJBrJmFx2uDJmy7+CF5jCt
HUvIZWxTVbqq+LuTcVjw8qzlPGPoQVWcxqnjhjcICSoILJAIbbaoFAFlz9lVV7KqTwPeMZ+krJgb
bkv3Snu/J6evCxteO/GscfFSmf3hGXgjbO0IP/Th56NKj14YQ25mnoZJ8eo+6/MqOgJCe+lYCHja
/ryr9vBb6JtgtWghrHhxW+fKQn2nN6l/tVxah2F/zExJF6Z+xH8bMB9BlVGmGTgVlpyE3LFPxJa5
/pI0GXmSXF7LI2HXhyvTyFpPenCPO4nT+u+E0iiyNOjz0MfdaUeWntBemowVRfRm/iltg7ku6n/I
WD/AxHJ99YiLoPvE7dbD7Es0vfDhrxQy3N5Vf9YTV6UFRwCzeGqMraoq/g0+UTBgjldRXk0hd/mT
Nh5KrtCQ8AxES5ihojHlZ+NGOXpLaRDIsw4Vo/z9h8Z8qnQoE/2wZ+v3WQcYaTMRuGS3hDEYtuZs
/Zkh+awWFjP5W5ixX8DrLZtWsBdIlfZj5nuo7OOGH4p02O1UG8JT59qyyt3OrAvpdAW1XaJ9Dxwq
4IBkkZwNUIvJo9o547hQEOpU2ODhBR5bNjb1mNbfELf0Blc5w67UX/oZ+KWoF+WuMgc+Iv2kXkJy
cr51jy6b/Iq+g5l/p5+S1HEEHCMHcBWnLW4mSxIOLyRgNVLs0uJ56HZvs1yQ3tL6WlLHSb4vsgjb
8q+nnIDZvbv1U+Mw9KvB6Uj094B7f3Moa+nZZzEa5VU5CA+WVZg2BEJRGkpRJh0BQb7KrBVKHTp5
EuTvPBWxvudXrHbNb0iPBuSLdKNqaM9IF20I6kLm3BGWHKXzbw9hbaDainf3gKTiSDzOftG62Gag
639Z4Dj3mOiKZaUNWpiBljGHVcqMBqmFQIpCZSyarV+MRPthe5hRaHwrYmHT3IHuSe9DZa99OJus
78iFHr+yoyiUTX0tEDsVZQoApjhM2WF4rVe3l8ztjQoY6eXdOnsViUCSzmsY1Nc64TMps3Q/XItX
HSVwdUO4CzcujgECMyI3uHEMe/og+/zsElw4sNBa8fz+TJURBF/smbd5xXmqYlkpboT71oYIYtLR
bCsAYRsKT99whJybdCSsdgJIlRxhmu0aEQnMmqC8idjhuA1k+4itQRtKmjaZGz6pGEQuWCFHLZX3
XaTLvWAAWtFI3vcTZclLs1V9N3Bsof0F2SP3Q99wuxIBOslOG/gft4qqeCkDT8wPHCxMEMpIc6+o
P/jYEGjeNVe1DjYZ2qyRwBhyJlkBFLt94wNWX/X/13TsZalXkgXfTuQeHIZNSO1sf4XSXnYDZd5i
arRObwxMpaKcKo+6Mi/1QS91v3dgG8TE0Rv+Q0ibOgVyXVDsyr6epRbZi87uBqykEQnc82/7Kwmk
kJtMGAPM1UBIu9iX3VUNBJ87gWzdgetOsI4SsMZH7weqWFhW5To+M0PB/YHbrjoBY7eF+aFHTX1M
Cv9hDMGT4YzTHrePtbuiizfilFRrbME389DsDTKMjWgMUjyRlR+U1ne3B6CHc0JHmchQ8HgBenrD
F6s4lWKS8AFP6BVKCkiURWvLRZV5PE5cwK16NRRvVWlTRkaMcvmVk70C2KJpXKM+9mAK7gJH02J1
MBbOh2zgZEjFl4scws2LkX9l0+lr0q4/pOnB8sZppguw/rEGDQb3IdReO08AQfCiEX6dj0AG1IXW
GgmWdRy09CYqwT2/Pa4p6KhDshgFtuWpX+vzf9oTVwuRAEbqgRT6uXtmG/igI8zUCOzZyOqhDh6t
HAwmftH0S0JYgYZHFHS7lv1sbNOx4k/gd13bZ6WovU8MlP7wGBJfJsQIoQ4MBzoZs5DhFrzCUSIB
0yHGX/qt0vPty1Uln0B81KYAGfYeGfG0yFiUsLPPuONFU4Bt/UyCsEPJxzDJqany4SE72kDTFLs7
XdHrOm6F5DdvYmji2GtPy3Qqe8anRotYri/UmKOWzdTWtCXPpdgmCdmZr/SSOOAd8cSR/YVFOIDF
HwBxGbprdQIwQ5/IY/BqwoET9Vz0604wAbj18AsQJshh5QXLY25AnUEAzWPX/0TwogAvEsW7RO3t
fg2ssdPpt8bP53ttRbUfxDRm23AVa5VaK8MUi36fC/Bk3ZlPYbz8dBCjUbI8L27HkYHGwcqJKPC3
WRgq7q3SqMs3WsVxnhgxGSHVdXZ6CJlgrWlnG+adMd2vphqlgD6W1eKC4hITLgqWaINDOAl90ifD
eTFxESZ8uZHbU27DpxgJxkOxv+Pu1C37eLOxnOcv5LpbhpOrNTK/TZ3LNVtdbuD4n4RF0IjsCxJR
EsKctrVTtprSos1d4QGQnR2TQq+4flDkfkfWfbp3N6jJY3yb25bK1kpB1QZOHHodSnFXgVZ0x1Su
bkvSyGupRILahC7/Aes+zq9R+uFmjfpXq7PaRA0xaDCqOETcmCSjcZQX5TVMXPotWlnRV3dQ6CgU
LhWFjtJMVDXMEvpC7zvs3IKX6YUt5LD6i0ZIN68gg8sA6ud9mZfyvhKp3ZyZjYZDTtG09LLBj9ga
gcWqHAI0FWs7j9B/L9rn5pKC/ZIjKm01FaaTUoWW9pFCvfkaUy+ijjnYw+U4oL9bgMZT16DNYHMH
QAD1ceUEcYjOgDA28CTS4OnZ18Kl6h9tUhJizGtOZxJ7hjOu7tW0WSGkIt9Yn8TRa1th6zVaAp1V
zPcw5DSVplzI0YbhYhrREtFuT0VJV/p66BXvy9LEqhP6QzuKaomncgz7XvDzm+0NY33MDTQ5bbZ1
2Frq+qm9xaAOMYCH3jDRtZQEOTv+XmRKfXB0m91/pRD4QwfCXFmOnhbeB13gI8H2PtN7w+ZDEKUd
iZ9MNTVdb3LvarcM6pwJY/9Y9RW+g3SJ7nKM8bVAC0wnrx/nhmMvn06mCHatQbUuqPatBplholjs
8rKgwbzmjCyq6qQenn+27Z8QBQh63g9wiZrc8NwgTwipc7clSrmnoOEwuE7pQbMvWcAUwyl7UMF/
73dU81mzsmbTyzgj7sdN8gzwdK23mMNMQ6hH17GAJjkMjWHsrNBGZSLCIG7B4yT6fS/jzeday0sA
JdczMSlM80bGTzy7CuYVVbeUe3jphH4/nYDVULq1n9AnOjNUHebkTIrLrTAyJ5ZCi7DUfCj6+xB6
VS27GdC8a0yMBIi6OzPZvGVXTXycb9z+kq/HhWJIOL9mlk8OmseMfHF8ioJQGF1blt5rGIwEtupV
LwvW4WQJqNpuxrpYPKJDQeERyWtgUlQqmARRZu7RJUltxOezOWL2GKy72GwqluDn8aOhr4YgQO4o
7c8WJV7WP7AbDBYpJ+AO0PhVo5F73tGONeOVM8kfeJsw0NjAkHYbSspYjCTO9rA/9pqhEJnIRn0P
e3aDawbdc14vqBfrqau3gibj5Pp0fI4gokyLnVV3QeR69tehpfN89a/Wg9BAchHJgOcS7yxs+i9H
lYXOcshgZ/cjVvI3ssVefAjdieLnJp7R8tGKVK8uTxqa8iFhKQRcDuJDb9fElrnk8+FZfBGqsAEP
JyTIpzQT8HIxj4yRV5kZY7mmZbM5qWW/1AXREAIHyNujBwvU+c+/RrvQi2nPS1jkK1Oqingir4ju
uqhnM/5IuFMX1BdmeyVXwnuY60sOf+OteNkuGC0Cpsh52Q63va1TNs0wARcDU6WU83qAehFOfNV1
Qv444Q84M4yPGHkL1BddKjO5x0aoQYtq5EEdy73WeGmvxMYrC1fV6UHP6qWOYB6NEuWOkf2Upsa+
M+fY+0LUv6sMcrayv6NWd+eEMmZ1A07vvAjDBXJH3mg9iusy34pyBbZeh1dFnMs2w9ZvT2cG15OB
giqOSIq1hjNi+uRd0fN8FgUlxcVpfyQwcUs7c0mTz0XFR43rpULm+su6olS/19KHKvKlfabOfPFz
MQsAONUJQyHsf1xisd9HdsuCmJjM4tDxewyKhodOyL+08z4YlP8TaCuJvjC/Ei2ZVoevILMgfSmp
SQhSQaO/HQ6aNAQpKunGR3dbcyqKY4FUe4sCVjZydfdukOTgsmu1Mdjm20VcnUq3GHjxU+lbuE17
PcRHitO1dWNXQAIHh63dtjwaIUBRswulRo4T1O+ZQOOSk3oquOD7MlwkXuVxwWPFlicT6XNb3bMG
K2BLqlLam9oUWtGriLd0RKJ4wd1MHwFsQgLolb2aV4qPhaxuHbdLNpCZSDXfhL/zg6NhW3S9XCOd
dvTNAfMHLpuWy4IrJPHafeeONGYJd1Tc3SSI8sE5P6cOE5mVMS2G4tH5NsgKJ9c0qErskmFNDhlM
dxW0W9qIOaDPVNLiCdzY6rLQHe5q4zj/cRZadHGci/xUcrXp85dMcEsd4k/7Xndlygftp3rNPEdt
/0gIlMxdoRRJFR8YwtTyJEsfL/QorgqEV2jOXn9f+TzOzFjJQ/XQsvHr0UjCjOiNFjYeuKOsi/6m
qgw9pfXwMPJWui7bH2x1Qx9SzUTt6oy+NouQsmxHuaiswcElJ9EJcuOQW2nOAz6482sQvNRB9Ln5
BuepeBsHh2mM/DzqRyw7Dm2et7tYy44aUxqxJxjovCRB/6Cg+pnMakgLzvGN0FHUxp4X5bo1rKx/
SJktP/zFm9eBHTzGmq7JqFqA8e5xZ0e7H8Fp9T1zivUPxlKirW8LyTQEfl9T6HvtEPEIaMY60bdw
3qbHLcIoIKA+/IgnPVjlYKcJL+kiBrRAv92zpvupFlJIEZEKL+qD2aNdnnXdEUdNbi5l1HeCOnqf
DzgaetD9HZDDIhJ7Ps55ynfyzq7Ohbc5PzPxqY4PM7PoVEVM5jIRIJ8O27/E0wA95+aZxupzVPyX
erpjw0OZJWbcfanXBMdk06YPnapz2+u/yBJEU9h2/8KMhJycGweNYcJH9jp2pAuMrusZ4F37gT2e
IJJtjaJC+WRrr8SVinF/F8UbWtKwgDJzmMS7CKtrSEiv7EbNwCd60N+S8UPNviXjPiji9E8RUhAR
EcC1rh1cx2pU0c499U4c1hLAObLWS1n+DmDmAyCnjo3NwOq/gQwdGHbGQsqkRutl0TDB3SjXi1kW
nbwiYqqnhJqpjeTeFLlQUYXpv+sVoStdkmC24V1EX4dWXChJ8HhH74cYSnrsK8zneB+FlhIXjmGJ
x8WRb1mE9i0xVPD3MgfJIXHw7hrv29o6bdNFZITcC8NeiF0t9KqLevBMQ5YXtYL5MQExwvOicKaZ
XCnlXGMBc9xZJ0sq47yu+gEQPZy9RWfB7i5CgSC54KxOovScEA59nzsYYyqnsN5/3W6EgQejotJy
ODKMVDTCfjBUaq/TEuEwrB3CK0MnCRtuPDAJ6NwvPxZQyaDGRJTkbh/mq+McL2xl2Ah/PYvdWb43
zy/DAiGeLQCtb/p+tqPPHIAHI5AbJhVQDaT4odS8zcZ3JyYzkDcr3PmxvcXfMsE15Tm9bpks77IB
iUEGiu/+jvBkk+KJlwggwx1pt8lpQEhKoaqdIn35QcEfBGkm+OyvBXLjG5Abdashkxys791yM+CV
fXBFQKn5Vd4C68iL+EqFXZfKA0jEjJ47toDk8s73OExc7DXr0St4MnQNTjf3CD2CAUOu/I1b67e2
d84IsFekaI9MFUr3kXiTsRrSuRa4HP7XPVlmjFUyVLm0fALsWsi7pLWUsEnBSx7mnIlqRfcvi/qp
2kfEF3GsSDFiX66eucCurBVdrLvSSS0S8a0XOtB8LtgpizTMvyTDsLrxPldCgjPNbxYtVDUPE/0w
QIfwyDvqsP8swD8fZ16HgKxmP94YQky1sQyReDg4nXgBNVcc0Mer60lTEngT+Nm0wz05bntHcVVA
62z9YnHcc6b2n23fXltFhbHIWnt39UdozX7thVddRH6JaHkXbssQjJeIkXEI1S5AEF3dQCJKP2a+
E3FOQuJb5rIEeE96I+m88rYq41NHttfYMGBT2SmajAWTAYe5chJ/jEJx9flEi3HBWAsDSEl2YpAE
Sc4NGYAa+vKslv5UfsZ8zYpEX6V7B/Os7/ivD+NqCgqHmjB8oNAABwibiQSH4JIvWZDAFsk5CjBF
dGnpwYXCbdh1d5Wn/SPyTfP+gWFhwh8EPvBKuRv0UZIl5jVbJI2otuQQNlCwJBP4PTE347LipTNl
WwGlZWiVDL3Azt+fce3YOi6VJ4U57+1PbTnqlkNea726PdogrDy8VQhbBRlznGzo8GE3O16RO4T4
KvfIXdI7zN8a+5BVe5o+0HqlaJtGKOusiZv9T7hkUDDg7DyGi0rnT/RUzFHF8W9a8D4x94znkRCr
4GzXfj2zVuJCLktJcknQjRohg8GsBSCp8c6LpkYDcJx/Kc/wcw/myQ2WAJnt3oLfyhcWkDe7DZRd
fWe5gK+PtForDYqV4ct2JK0jWaPb4Id9Pbx1Wh54SKBYfE4OizH87u1tP4YZgSfkTRj+O4xziDw0
SC4WZxbfXq3pyoFnlSOfQnyC3ira9/dUF2Gp0y9SvGutLS/8zrk6GpeaXBNBpSQB2k2nbpwyywy4
h1gdU9aUiZjRJNZx4ywZL7ldzy6xRNikd0ohMzXJakRoloSiXSjHgqLr+K8NeQQTrEv5QJZsVqEQ
Fq7IzkZKh9FD7yGA47jYDyoosbTedPeCCk79/O05BBec1fSgKyW2EL/MkXQU1JAsNUGGb9qI9LpL
9xvagbVSTFoJjNuG66H+F4THER8DVYV1GQ6DTrjE/6qCxao41VCgMRlbHnlekVpGpvcn00rKOHwi
/pIu0ZZmxNO5qOVOAVVOJ9Jh2TyMNghmLfyLuI9NLGmq+xf8vPRIo2slhV/jHuTC/kKYZiIkPCpL
xWV6HVntZ4zIkhSM+f9/+68l5L1DCwxsYLYbCnR1C6z1lVSrbVe8WrNWSFz7kMOHf6T0hA8Aam8Y
AdxrhtKt4R8jKehEetpR7c3EbJSaq/6RDcPqN+tvjOYHdEK4ZGU1qPdfzblRQD6nShDBAV4/HOyf
k0x1kwy1WaUEM8qMlXtPXo8NBkmVHqSWKcJCO8PTzSstKREj01JrB/T+AjZ1CY0i281sl4syaAHz
YdPF6AQPAC3XtRkq8GAN2Xyxpq8vmTe/3eksxKfNhWN39P7gdLB/eyPpAE1WRVYjZLtUNH3ca7XR
26bLdjBgI+XooPGfrMpBGBRQt0aoAPvhc2NUYFCxd9xpX6rVk22IyBuBlvV+v9X6s6mwuBuWC7wJ
u9YmXQCi6efjknb1IpeShRPmPG0S/mkNFJKb5a2370WOPOSEHty3RtwYTQEkpCMRVg4qkkH3EO8d
rQ6I9RYwFUxoXgPlMrlyVsr2Pg5wtMOdJ/taFhKOPfXqh9QLhfvK1vTayrsPdA6FriRLinsUIVTf
is4dwsILAcEHQ2sqx/bTHx1BD7xLooGEWFrD9nerKRz7E19BVMf7BBUeHhTOUAaGZ+2zXk0jwmOg
LE15pAW3jYWYjbLzjuCw2Cm6EX4q75MDFV/1hyT5fflyjIrdC2N3qJEWNMD88Cy2zuZX6AgonCyF
8Qh0pvuHNPer70lIxgIdiHZ4dqW/0AMToFGL7r5D+goyJFBn7kHQNvSD1pYKrp3F/MXoMRXn7qiU
eFH8aA+rXEPGX5KgNfhjEtlPAF2sqfyuMplQos2XWJAWeJlgLC11vgLPm+QDUngkTER4WsOr3Y59
7zvIN5M7UmBd2X++9+wY+AW6oynJf3NDh/YrzR2vQ4uuhaNztjN+CcQSyrPsOynfyFotdlUylGQp
usjg5lMQ1TQ1+HnTy6k9lez5kK+qJyLoVNpEXe5UmKHdk3sOuSotjPxlzLGtlK3orIpIkJ4IwCR9
kN1cMwRYxYb2x50AdUvHyX+JSFj+f0B1KkQR4dRMMkAP8dqTdQX/oTJN/HCP4Ghp9ryJiDo45xDT
tC3FID1QDpcrBThZKQSADSFrUavHK6W6X59XBJqITAmdj27TM2ibA1LfHvkB/Pcnk4d7RuoKBc/m
JF7+nQ0CytrLg2YVkvSui82H5Yp4frOfJ38MoS72UHin5ZtxUVWWm6DePhSOdHdIdszDwtQ+54Ct
iGNtnO/tl0PuA1JVwZCH2rKPaKjsR239eKaY1P3vKORwpF4A/H8/qXpGjY8WMvYsD94aX7pJZBHT
DJBoSOZ0xCCKBueQu4ZFn9LN46wrhNz2LG+xzy/BABz4MNXKF+7ogDKy1ytwFNEHq+SsPZl1rsni
xmLgdP8PyCAZV4An9VJ83zp7eV4ZJX8yhP5X7TB1CsH56FBWNXDp9FvwTqjrt2CKFqKjM/uaXSfm
3ubjeQ7Ypl20I++ANCW3K/GwgTyVJEYPjhlSNPQovIn9udQGevvsCp/ugKHCorrxVYRE72M6zPJM
w9qTcD5YoeX2r+WpZQVa6Fm2/bhT7Kogx1vmKdvjfE/hpDNsvJUxx7HcGttF4Qd2gcP52G4Vs3SL
9lhoklHK3pMpsGLIboDJUSYxx3yizzCw36916UEooaYO3sz7VKe+Hdw+smHaQfzHFBIdrsbUAclU
fx0ksvJWfY2b0VSu2ThGPONNHVY/W//zpM74gJ8o3u0IyngbhoGrwV3XJ/eHiPB5AZ3UBsKkFOWs
IxWV16XWr1nur0NKP09+lrPmpSpAgcgZXl5/9dKnTo8Io0gfUXMV09woNpGcPV1qS8BKt4Q87DV9
/UNtahB36FG+TYTJJNnFOMvP7/ormzQ4HIOvLbJB9E6Dd3uUnIGKjcntLZC3eJX0DjzC2y9K0gdV
dHhtZ06l6mPGF6a0q4tJaTr/5IKXo4IVwdQuEcc5aDUx6+Gnx2voJUZV7n+HEdI8j/k4IZxGF4PF
x6jeFq/ZJVBq4hBXFvkeEG3EFEaE8w0DjMZBsxO/Hwt0b2n+L9AYUraCrMDWbD6a2u6sQtmM5Gnf
cgRv69+SivNp3Ulkn4w0HKA0q88R/HyKZmoP7Fls9jnQrBfLe+1KqFMnPtztuz/x0DD9GhU9vQKc
lOlHSa2keJaENQ+jETuEYh/SnJppn1IdR75RvjfNcDuJeqeBSZ/rxesHXHXbcd2AU/ebxMPCNh42
KEhNrTl/uPmqU/KbY+r5EASKnEnD77GMEoAKH4JottKfI7xAeDfU3ZetFPfkOH4ebooy1/IdoLqu
bB04hClaxTs1yUBEYuJJUpKtnC44CfBELC5WmYYBwd/6hQa5nkTVl+2NmsgJFnBLkfemg0Q/PqaH
Q8Au12TLf1WOkUTrlMD8cc7XtzdLfu90B2DTBakAYwqPHlmZA93vtL7YfX29cNXhcP9+GWYXQuGh
la5r+cooHoy/TxYJN/GY5tK0fOyjm/qot6jTbsPSPwPjMKsovT0aKN9ALNeA4g/vpjAaYvv1fM86
jZGlm76EHOC/lw7QhcInmiY+xblrJq+Yz4h8k+YkHVEc2NSsjVdDhqRRXQt3N/WabrVsZZYBFj+Q
TriESf07wpUUSN1T8vT7YwV05hYuyWobazChJc0NQMrM+e8GZHUWa+gxESgr+JWrDA9LHQBBER3Z
pGkPqCRxwfmjxcSXcWBL1GW2/Y5VJTTABGLkjrazIL5wpGmlfzFNDomd9Ean5ulTI8VhgGnVWZ3a
QpA19Z7j0M0p2EQk0MtF9O/bMxh/fL07IpCMbjn6kLZ5PF1/b2noJWZBZj4d8hAdng5mwiiik4P5
uMefZND+Y/fO2CVmE16NquiZZvaLRoF1zzGqexNA2aSOvD5zyX/KG5mdY7Mt5N+KxK9IeoF/Uk62
8in0DD6nwFQO/gb79o4pIw8oH2VONG4+1WJ7alaD/2OfQLzn1ZqMoW5OFCVFJz40QNfuO26NXSeM
4NNWOlnpWN3zek4vxyi49iMnzIfsU/yjB8lUBdtiD/l94tgclEwhkp7s2r0gcWY0jImALil5y3Oj
j8Yqko71g2r1rDCy1HgAKSgy2Dic4GVQR1QUgfFwENPC3FSANfcpulktmlTcP3xBexRZd8jrRFHV
kH3Kw5sxa3Gm/Cm8oo/FciNGQ3o5Q5vVHewRjics/CF3L59v+/nlST07Xt7wigfOhH8Q8zw+hLWb
vngWEih8z5Ph9WICxV0YY3UZcSRIO5xVe/QCcrYJCocl3mJruQwfVi5/Pa5wDqG7hBDngRSUCGYi
vo3oAot9+p/eaRmfBv5gfvX3WoJBLemtaWTCPc4cJdiQ1Y/zXElIx6Em9On6USwQA7Rcufk9wOBy
ZLgznFuvHH/V2XX7Qv5+3WUdrJMGSfCpwmP0xYoStDa4u3te2MBYSzjGZA8Bkw1lwiLCbZC9V8TD
T4mhL3UlwEtQ3mm3JLrlBf/z44AMZ1xD6ucXWLfpGuN4JA5A3XlD78BTddAkApK5XJ1g8Le6yApI
iUbFDDVaTaJxUXino6XOfL9Kxh8Gidgj13aPli7BbcMObB5Q46v6zlXBmQ6CJA2xeGleUjllGcdI
H6W5yAg3e2LMTijamS/44DSpypl4SHB4okSl0uJhk3Ns3W21wc8AkUCgETcABOhXYjsXdvwV6L1k
W2WiZoX6arJf8VwfuYRJ1pjcOIcD3/0yhLPzxSVmmcNNfl1hBQRbO6EoRK3lfIt/R7xTSF75/+Uz
P+S51NpQIKTMl8F6T2XBvSbz+DbZawxZq3QoRbNEm/sqg5EUhkYSPTRT7yzczRboAXJJlzdNkSHt
i08muAr3gv7nRJyMmvmJv71/CrsOnVHdCupBhNOgtHQL7jpXKwb0v1syFNEzN8oD7e236KQhFANN
zxpEco+tprscofxV94zLNtuIqPGoQ+EtbcE825C5DZrUJ8l37s/rF/rojrHduQpfdqBo/8LCvQkh
+QHKO+hyoUqNJNV9mMxZuAEiYujM780LlB/YOBvdRWpbGSLVCM5mSQG+kaefr7D3KK/OIsiGGQ7I
3T127P7i/XWxyvEnBnWapzK2tzNMwkrL6z8ZW6l/dfb6lblvfjJqIOnsBBrz0F67Ju2FPXwgqylk
IU6IdbCic1PMyAXV8anHQ/TWxJRkNerAEbyVP2aiQBIVmoxHC4xGblebGA9VnBh1kFBNZmnArtOK
/52RifW/nc/XL6wxndpUqMbGkBnDIhhxvGptrtU2NgS7c2yZyUKTK39DfVVklg7G+/v2LFh33FnV
wg7b03yh7EtJVpGADswrFp2c7RxZd5wD93T9sXRwf3oWxybBIOLwtUiR2Ra9NeZk1lnD0lwOQ5mT
lXX2kLsE8jtfgS4UqzJTTi7Ay7ftnIdpFebQHSiT6mblBx/7IfuLaQEJzxHB6UK5VfQI14KJyD4u
WLK2Btmoo/fwNDp/anANL5n2y//7WVSScmL5vuPZbAtWBwxKarHrt5BfdOgTqk+vVAkRijTlytAI
UEok91igccdkLzCnCUcba5d1h1/+si27hIvNBMnbdS9EHByIvCCqTimhZMetCysJlQ8Onf3GivJg
bZ/TLVINr8H8bTWsYa7JYNmbjo0xtawyzhqIJPCLXUWhumlQ9UJVRtFxOEhnWNqOuUd9uFMSRPOW
M0CgBGB5y2YmK57VBnNic2HqWKTxe4bj02szFmLlQ0Xm0yX2F89zmoorSAS9wczvMV9pineuNIj2
4BEgMQiOW1wfj9uYWgAaCSz7POWyEUcXnMlzs5fNFAVixTZbNw5G353OBpXuFsJyqUHl+aGkX7KT
gGItPVqHuTpXcHLG/Lf28+8N8GK8fokh3+oJSbYf+wWJ2z05Tf1TwvTTUBVEbmaflb0ZTS92FsSr
3gb3zxNLt3woEnfdf9rJRBxC2/7P0sN/c8NsUcLxXq7Pj5I1lfEhyfiA40DwqJcLX2gEsRJ0uzkM
p6bGRTHwGgKbOxuGE34PS1Ib2k9LMt4ulJAcJucbSWBwjiVEI1bvvaaElY0hyiFN7fVclJCMZKNk
H5kvWFxw8wi88UPAXlH8+daYuONxq1ZLO1niqRAmVwMPeq/wSBwfuN641Z5No2icRgwtiemEdCzS
Y/Ay+6Euu+Njvf7H0xALIT9Y8PKlEWyI4xqGUcr6ijN3JzVC6fv+9uOZDRoky85NGFnOXAhcUPrc
IyXLpYldDA+bYluYc6fdgAhHakKg6ZswHe0j2dO++VlOj8YMWi9GHUiPUwJTaM4aPhIdf2J8Oz+e
nVOZDekacgICMwLPqkoo8Fvf0HbEpkwjYxWc4xiAVJaeV0qkWchV3LcbbYePrt+HMQ6J9uU2mdTQ
Tctz8/CbP8F3JeDsaBI33VpM7mDtlOWtJibKaJ9wMmSwrsQPfsweO5XmpWEMtHhyPACFnxBhicDj
wFFdjP2d4iUw43Xt5F4gZjx0Pxxp9uoklP79ryQt8CediZYgAecoYChv8Z3bcsEZ5TL1+c9ih73O
z02fq+cUSAC1y3kXjiv+NCa/EM44rfHD17yWGXgjvdVaW4VTSH6v30gjodE//rBOBL8feveN/slx
myU9gv1jM4Fm+oEl8TMQ2U1XfPLFtpHNrWI/dU5TToweBSFOWp4UMzZYG6cpWlVUSNMoqcRdkuVW
hgdVlhi2cKlPeHvazvw/2fPC3uQp1WcIDcIbNdpMO21z8zbGrvjp54ewkEQfHnlr3kcWrhhMRQCY
6VELpY8nn2LiuIv7i21IdRxD7JH0Vk2fo4aJDPbJQLgAbbBDEFjrZvl+iZfv1lamGppT6RX7TKVl
d/FRqzBMgjCSP8cRsWp1jd9b8Z3bWKP9T3Td1q7vseiyRfZj7d+lm0WTKueiXXu2qcCZJbkbsTIN
6putzmuZaO+AVQS100jyWIQybqCdOJuSYkhlZJRVj5fagB5GlEnYpXG8B7XusHLR9ggVJlHQ10S+
Hri6aXP2YiSo2fYMqCJ6YIuMMyUcxB2qpODfN87mVjcDn1QiSTNUQZ+gWmVY8mIdFgdKFEaO0gWR
X+rbsZkmD7BSfqaX1XcIe5Bhm804D3NZvydq0sC8pKzkDjyDnOwUC2q0dAPHzc/jdzFC4QlUqiab
mMUDR4lYcTNMuUtWbnb/uqu0dpJv9Cd1ClAq9U9aWGHP56srxzpXKkNcgXo+nsfWpaMsMEGUs0Nm
ZByDnfCX9eii8cp7KoIJeZ6J73hVsbxcp6zeeU9oXeWOMXtduED2KFIixo+W4B03kV0zVQuASA5+
Gl5jtGNvj5+xbM823cmLzrc2+/u+K6x1y/Gm18pehPuuAd02wrF0DQ5dYFiSaTj4SiJ8ZsiPILNn
yWxbqh19xa9+Nqk35SyXTPGGNIQdekk4E+9Msjvjt6K5MJYyXybP7St+yK/u4WfwXU8ExUymwUqH
GHBSATIsTLTeMIz7Zf83gRADYYNC3WNQ1vgarYT9ApwavrolcM9Apn2ENxK36vzH+XCpMQR7p3ZF
xjyAEjm8/VUt7afr8PFtUqB7BW5/mE6vSwdV+pBLPZ9y4FFtuf4m6dmrObKy1+ANY/WhNQ0Rypho
Jwr6ezYeU1uwcox+qqxBG/R1lRQ4fsCSQtN3pkpQTcBl7gEK1KlhxCmn8R0ckreV6UpigB+eq+U8
wOvWjsk6FatgFXBIc6xgAkpZ/VxGk8yMXsm4I5lOB2hKdOTE97GEogF6lAaPljcH7JUN2UuXOau2
DySeJcmXNS+53CmBFRmWrlhQuO1kfjtbmcwqVDyftleULJPVJ4n30Z7Pr9llgAjgnH/FOoeiy1Pb
nwKLNj6nORz2/BwJ6f03+ZD6valRjun5VO01yiwckTNnhTdn26zR67QTjrpbX223NkXk3I2uc4E3
vj/LBvbMys8o6N7wi63jez367UIpbXJG2EGq9q40zUEeRf1LF5ii3+pRqO4rEiNsjYZ4mX8PtFpj
x4JYq74VAhZqsI+ZVZBrF0kmrNagRgvKIAXTwgeQgdQgYXOMS1rVcWBipAPK6dlBsv1OttPvEAtW
OaYGInRkSByBhyRL/H52riwSXghaZZeqmkbIBsaGY+82rRowzAJbrwcxrcyPp+KS1UbbZYm46LXw
mDvxTenxnUChaQXet529GnYCypHNrR6wI36YBM/X2jci0ThdMcf2mLjlBfqmZlHhjUkXrD3eDJw8
v2njMMljlA4ElQp3kDqPlmduj5lnZuVzlc+1xdjKQQ3r1k/Sku+JlNWOlyIWdt+a/l/a6Eyls7ve
LTzsZIjOn9KIIfFn0p7piYZu1zxeM0+vr45SZ5kurwCOldkFNfeiCT9A+V4OJ66PTxkmzX9hMdPz
ttQ1rNmZE82dp98s8QTiYkL/3r1TtUbP1w1M3opgDwy61tx3Ur56TydYeGwTxC7AJsBmOYBsg/br
qv9PehDPKXnohsPo2+y3DIJssrTqe21uqJU8Il7KiHrF7yel0IZQDphYVPjWPgworapoC4b2K9sj
JL/dfqqbhLdjI3ktqSJvqNnYwIn8TRs5IRUkd7lwARCB/mMynWHaXTHdXhC++W/blrzUHb9Mdvvv
BYxLG2HIlbwUqFnlKje8nQYIfJucV5Ys7/jOzeZLbnKL0HLkt7qIO76zTe9qszINP8XmRZRKVv7n
SSiSYrJjHjfbnk5GQEOBTYusgkFxHtVpYLuw8AkRsuj6fioopX6IpTUIHV1QCbqV6QuJpDcAN6JA
FiGfeVr8ofg/tFEymYFiileOryndsxV2zfuFfH7jtre22KtIva5lM5Xxchsi/Kywd0qc63Inj74k
mOP1kEju7WwNRr6IAIDn18XIBVdFrkuI2qqdrDuqtBewnBqgSVyWIvUcnR2Fb2pTmpHRNgVfJK3x
TtphYPlBbCh+AGaUdiJ1S5LU4BAh6dCkF2BRfoDGAqSrsAB1WakQsPXBof1f4zfNI7zykzaZ4Uah
Hwx6sTfOP/yaySEk6LLC6jcEy6SLH+cPwzd+78Z1/HVsri8ed+JADD0HCdTjEg/90QJRG5lPWe/9
lgbyWhO+JEPY2I+0C6LdgjIjj90p1bq1eEHVWO6G5NB4gxORNO2drBheGqF2LFSQLFukPP6UbyQI
W7C+VLG3Qbst6Fx4CbgQRV+ldyo6gyoDUY4MKkZxVocb6LV9k3srrbxVyBRwJeuBr+xX+QGWAEIk
DSaJluHzUU6igCQdS1SwwfEl4cg3nZCLT/XP0w4SrV3bPcnuMT4Zuje9/kDnrLn6xU5YPyfZdYGb
StUZOFVAZsWk1JlfRZm+qzRazufXoGOHfXaCYW9aidiZ9W6ji1ej6EiS9i4ajkAOPJgehIHWB2Jf
6CCwHw7BaUUYymqMtvJlaNXWzRganJfVotfOIOMg19ua/tKKNT/hf8zDzUikBdh46KA0/KlusT3k
Xr1Nxd/yJvWACZg9AyQHa8+bTimZ7sMxcAqt0gTZWMhDEQeh5mkB0U0D8sCJR5fqHN2d7ooDVkAj
GS1eqI0x8N+0spgMG/uKBLCUStkbLW2cP16iIX0haNTaUZTZ+oQqRjqgTubcXOa1Byl1y966IwXf
OUkECOTWEH7OVeCaDBaz3cbj/XBS6WTJ2qFTbFiR68B4igT0sxWtqibHPJb/+htUUM8wYNHgC0pL
P9OBv6TA6k/qLPceGswvnP6CJZgE8ERZrXCiC7Ei8h+l3Zd1OE6d/md/54sokQ/XwkDNPr06mDJK
K66bGSlq8iMWlBsm9iqtBataqj/xDRRO/4+ynwQo8Fcg1Ir34dw98hwtZpqr9q/ObWlQDGni8l6L
GEOhE2VGNRqSVNU4C1mpZjwMnBb21pofNlJpxLwm3zVmDV/1g7Lh0v5g+TSB2oLPqqIBUgl1U5oQ
yqgwp2fB37j3ncgb5e/rXD7Nnzi3gKQZMptxMRlTK2A6s80TNX0GZfZZ4zhZ5i+Hk94Y4x9hs6Hb
wfw6M1o52jdbJe0pORrPRYmWFUJ7dPy8vVwWiWi4O9xu/zG1Vg5PYn25WuMTJGWv9WKRFkLuLFyQ
/WY85LxzxdDK6ICp+ydtey4GUpH33rddNCCPncj80zHEZPS8jY77DSPvxbweFmoE9O518F7QjPnu
r6swG7j7CLe3fWs5TALsO7hqz4VhDyzjfC7C2FhK/fVYLJjy3rPQkie8KR5CCNIC0MinK5HkNo8N
WcKx1oTb7u6HJSX1Pfn7wVO0uclawMq/LOsWrhB1drkwC1Ttu3srd9r38E1JXZJCvg2Ikb+Q9S/v
gpH06mcfjaVD8BnIFArZ0dnwFzgQBBF7sew3qD7LQA0qtGItRH8XBXXQa93cBqICRcI5qXY3zsal
unWedtuClXdYzjcIpKadqiIEPRZCRBouVJK1QK4lMV3KIjwY4NdGIgNGPAVucKmRr4X61ZObTxNM
1Ntbe2Mhwk2HJl0VDPhsrthu32zaL+ZgUw+4ufGj4mVmTULeklw9yOjsXa2czGEDDHpN4GgHvu4G
2r0Ko4vrGSWaTQjNVn99B7rHDlhNBvMjavr0GyvQVGjxyZtWKws53TZbGL9fkM78QfbWDC45b1rv
g7420MTAQ7ugy9ayrNbu4nJkKPTnpiE2rbZ2sQ5By+3z3JWO1CGYhePRBQyvuA5CA7WiztOFb40e
II3MtylDM0KCl4Y8WLxt+Ox6dRivEpgYqbv3EAx0r2Bf/1FKopyevnKFr9f7MsYa61z/SUTECM+7
KwWfxNUvP88MfHmSVOsZ6UY1iM5KLP2hbv7FEZ0c/PRsPOG0gYp7EWs87kn+cLsJVKb19+XCgY5U
c2lGZTWnaaAN75ln6cVBqZYC9BYSjAq/5bQ54+ojKhIoJr+tLztcfkpsD4Oz/bNWz4+YWtcuYehJ
MhWJEjW3SD0I9OzXhauOAYy9UDBuMYHXW5K7vH6lE1cHsap63szpx9B4MdpbwJxT892ugeKsKN2A
JkoP5M42GAHjLswkA63nGAHuuRIUVmLngQyo2onkDV4o92SQNqqTmgqNc4W2RsTkWevbsFWK3yR+
s1Gh7memMKTjkjVsC9uRpIa3PLs4he6HYx33kB3dckCDK9CbuObzPNKL0eRgijOj3UsVmi58lKj8
IVPstvIeYmrbiSfs3sE9G1+7ohgY16AMLr85++PPVDQCoPXMNZrrV8xnHqmzFCJs5D09z/qHNX+u
Pn++lWYGyCzvITyOsuFjd8dr4gnswiEkqMuvFxJmxkiFlTi8Km+QvZ3WgpSl5UOuYP6OIXaEecUk
aZnvVsmAlAZCqHrKWsSNPm1npuTPpe3XcFzs68YMnehGxrqPLk1rSppbgcO3nxSOUtuih+dRRsPi
J4aqNoWErMv+BHrfjLjDl1aytfaeSkwyBhTe/mqRNK9wyJ+rE7tynCJDXpqTf3mRR+y6aIAch5re
/sKFTcRVQgnWuoTeiPBfuN/0jOoUP5d9yuQGpKGKbq3Mj0iZQ13SnZ67jOcxvlACYvqtWGU82459
u+TtcZE1Bh7nEnPqj6uhX/seOzo8smu5mAJffQMSkyjBCO2bNpNqV8G/Ppy4fz5Uxv+bYcZteV+R
gTEXg7QdNWTWlWo4wjB3HseWv+c/wi54qLi3l8Rr3q5syQuy7Slt70SdJml9FVVojWEyKMHIEKKt
2FbxEycB7qmUdPZgxV/ytimFQcvXfPpbMsej9xuVDCiPpwyMgEwlNSfIhbcEQ2QU6ALO9J3ZqL0s
WNfzJfsH8X4DIMge/NIkkSvmZfbuED6SqpRTwTXJzwIqK6qkvbsMmWDEOY8IbDXs9/fUMnc1MSqu
4G8hdMqd+foGFWi4/tHT/cSSmEavQof1cRNryOVTUriG+7bnHN0ghW3fNxaiVCW+8cIQgwzidOD/
4M8WhN6A3D7HKhCPKn+se5kaVkx2XBPynQqEj/tVY7jTDTaccV0zN6hvH1qQ6qi9OtZPyXHNn+ay
t+oLuNHDZi5BwzrGE5oir8HBuvF/BW0Bs/8V7WeT/fkHUi0pLqGJ7ALYFJU6Dt0+SkAssJ36ApyB
RArQyUE8Nq9zS9P3N1ufcFhsasRdMRV0cIdXYeKsFZZxNpzxpKQFmsYtXC/z+ePiKowmjz2NugXu
sa5BRFde7nOyuQAmd+pPqYVHp9zVMEm9M4hVIoQjiC04NKXqSkCfvyCnghXVixi5bT2H4ucGcWBF
bvR6CvMqbmxzZ5tYwO1pZARh/LGNLCECVZYU0ynZTdc6lh+7gYREFTLTmHmziiszemgzLcIAk55Q
6dr+CFVOIjjMqRgRsry+iGzA+2eHHF7WVNycxO4j5UGNJ1GUW3BSTNqDfOL+DsRge4RNOaUFPk1u
F2tR6uPwv1HhhSRLJQvORWjXnx75u7OAuG0IfmCDpebyia4EBI4CezVtzChv6ffqxpTUMtg238uo
9swxodJLzbLfIJH6OkLmMtlyY7/gQ7ATQ0TYwGgJ/37gIe1N+gZ7S8qU6PopzGjhHFl/B/cSkhfe
QR5oQc1vMQxZWtdoMyLMBypceikdhrc3Dhv3klwa9XYhZ5YF6QJV5dqftpXIxoJE3S612hRzFues
OStPF7VF2MQ8WWA5YIPH+CuxNyiEITW/Os1fK7ZxVzJyllr69ZLk3TkUNtbhy1rJ9cALAuXzOXjf
xQ2nHrfT+EpP9nD2E+ji4pePSF7GP4a+xxs0Hd8V0Drmh+NrCjRVpB2JI8Aj+s4lTZ4FK/lz4GqP
rIu2r5uhS0UT8wvt1c0pbQHfXSAs/omIP6VOgBbKFAniGC1nLZZhWc5HPrielDwc9vAHe+6UZFDa
3cUZLX88Jm+JnAhDaDQnlfxmX21Q0yGeY2fPzc9X9oQSfkC1yvRG76PZCZ/nw5SGDRkHBx2Z5SAz
f8lP7DCN5XPr+LnFEgMUDsQ2Q7Usg1QIjvcvXqB7HZ/smaO8Y600/314ntALvMp1MsnSsEEgNwEk
9d8+9OIveqnNOKX4OtL12GKKOJaVNC+S0+BxX5rsGhIKejej6znthGVVTZYoccX//wUPkqtub2k7
NotJhJF5NQ5K/D1x2+/ndjWy/N+Henou/Yhr9+cOAYJXu3qNGSdz/GT41eiIPCbjJmx/eLMV+ni0
y7NYFmSSfWIgzGKFET72mUBNI5cB8lUDAEB88gW7aQLEp+p+X8gIRGCQHQLeJIvfGwr2ajDKal96
C4T185Ki+ejzXVDWa3stT9FbZ+rQVbXdHRYDH7sgzt5pKN3aRdQKxQ0Z6wo7h2qwcElS9aVeMO4A
VnDeOybPgAs4USJ8vDR94awRCi7x25trFT7Qx64f7ecG5Pc3326wIzjuDEYvz6UGpi6PyQjX7Os2
la0ZfBPoRpCPAWc4OZ4kWwm4O2Px5T2ERvjwhYzdCOgJCZ8Qx1jukmNiig+Ky1MSL2prh4aFjkku
7m815zbXeKp3bcYWoie3TUar3MbT4p0FkKZ7V3EruF9NEk9uumJNducKGA8vLhlj1XlLEKiKoV7H
ejQDvyefZSPdjxoypVIsYEBGHl1bGNcbUWwNB3DrMFuvyQBZ+VJ5VCSq+47iokNhNRmxOAajPzYn
s2F+vkKMs5/OCbRTiuOBDF6/GR4YQdq2TJjKLNMP1WfZdByTrPcjaLFi7bur6tNbA1mdomwSUuwd
6iMozAsBAuuNPodiT9frcf0RLVG6jAyTxMSiUNs95r6pqqBuFVS8qudHnbHDVT1oo8lb7H4k7p5y
Ikhzo2ofmhs/hFadw/zyGwcG3wObrRoPJOx60Rq/2l+AHfBVPdFbLkxwB7xoibAOUrlnxoKn1f8Q
pMp7/t1ow6JJOUs5Icropb6OAYQizQLiRQCZPt6TsD3a7eLC3ba8TlYwLgjX6LL/qpiyEIj2LuXq
fRIkCZgQ6adO/Jt7Efj4kFO+jvN7OAoa0TRiB+LJIqSWIsPcnxmB07HosBjP7vGIzb1OAabXtwAq
xLHx/YSHUyCBisSJlPqt9kiMq0uRrHn0DMZJ1WRar/bv4dirxfsTwpDo2KOE11p2Ct3IUxUE7Cmf
JTMgZjB/t+8PbvqEAXxMgcKyPM5FjBM0DZe7q6L3p6qSbMmWEqMx5CfZOYGS0R/6Qh5yLgwOjQPd
nV2IbJ1SrV9DntacO6csFN98PJ7oj1sYTyS1n5d01we+qNbBtfwMZLcAfMYfBsYdSB2Kq4ewTyeo
hDGq9KE8lWRlakjLkA///dE8XSG/9LQWhzfECP2jelrarWCgNM9waU4UzosRepl08oAgtmU8/MG9
xGyTU6KFUMaB7FS1pfeZ2GkZmXwGL8/iTm8IY1Ahunzn4ScHfe+ChhmArKL2qyCThmVqjpw3gffp
KSH2klrmMbZrBr/mGC+EB/cGbQkRAtfckIxQXQiqcUWvmbvZoo3HRVOKdAH7V0tB3VZjlXIWcbAc
4L+nTKTsbaV4zeP1jf9yGX9ffABCqsnKsiE/DsRFblC2QF8A30cII18uX01sclAKFHqJz/BHW+XK
i8FRM1bk8WXjiZWUYhpG+DZQ+S7LCnqY7PTB3+z+nZjCJG5Lyl9ivwlnOkG2LN4q4lRVLFIrGfPD
RzJc+/RQGrD2QZXanPt7TstVgmA770CNQ4RZ7+4RpApi8loa5KQ4i858EQOUcyhRqMckfH9Ga59u
bSnmrTI2SCRC9obiq5q0FSO8Kb9e8g//gpbfXEAeWNDgKTKXh533f0Of6x7iQ73n2KpOTbxwP51J
D2u6LjbjweCxCo+EetHG6w64ihsTO7KeNsf7+KxBuHx3EuWNM9m0gqnKGd1SAVHY9SrMQRqwb5d5
4BOPfc4qLWwl4TE7XOnNcqaMpA+Qcjcj8MwjOAs77i5BNb+q5WO4oWLk1/8EH39yadPW1F7e21Lu
89awuge2/VONEW9o9FwVQhAAdYugT+Na37PlXH+zZLPw5BJnFv3WKro7c0/dIXBxQxK5BsoQzLp7
mWaD9MK9ikpaFPxlTHt+2+txqfgkOf+WYdtZ/Q22mLnwQwZgPZ1wtdRN51y9hXVL0weoP8i999QP
sNW4/GOJgkMAMnbDCsroMmjl7ZEKqp11vDo6FBJ0NklpyhppccMoLwE4/iJxBYfS4NehEYxuf5mg
gPJALyOJ3uRJfGcij1os9wohgrA1kxTPlJIRAvq7Y9QUpgusX7SBxn5j8+NjcSfmx1reTqzsA8xI
YNP7wPloiVGLM1/yTcE9PRLo8genV4zTgR5Zej3VsRHXXXQmJra0kY8gXbCRQmgotTxlxoVHItAM
i4ojWATKziWLt1p8zhzeSHD4yHUPEpn7kRlsZr0VOGl/fcOa1iB6awyYOBAFbdY4BdIEA1pPi9LO
ec6S2NQ2sm5qgJLyHZSA+JJ0NEPx5hsxeFYwO82thyAmN8QKmmV7wn/O6BkObEa/GYTSlx3+PcNj
QsjXfKcFdEzXis9Ve0STEuWifnK5HbOpJ18eccb/I16fHBKICZgRt+d+EbK3+hELLnrd+17ExFic
OFfwUA3LE9N5mLW9Bi55nuut0UCq9VNZDVh8VT6cnguD99gc4IfYVx7W6Egmm5CvxmjoLcShnk3l
a6EHQBj4iPmkFpOeUqPz4YF7kGthau5D5mablj9aEZOCcM1jKtYQSvH8m9WtJALiy+Bdgdinxurl
8Sfh8ulYU+HWhB3U/nT6rlz/aUSM0kLwsssNMmp5Yhw9mEOHOju20X9HP1fTuyazrR/KaN8eHlfm
6np294fDiAADjBlblagYOLnnWJax4ywbWiqnYVGH8ivPDN8O7sqqB+Cp0fZzrzeY578Jlm16AgKQ
JEcaKcF1JJb3IBoSuvnI47r4RA3Wl9rEc3eQs3DE4s6sXk2sPybGFQcg/R1r/3qqvEYBjC4tpt3l
T9pAUckgF9UmLw86yERYuKI4wpZtE8QBfzGtMmPoi7rNtwtkR1c2qmme7oJQI9jq2qfSbB+k7drg
F4NXRhd+XCTrFmUvmIJ5mTluaUEuitLe5wEwspUVxI6IxuEHey77nHywYQ4rKnIxz/QeBCsj5ryR
4ZdyLapJu8rbf5sgIVahkp5qlr7Kh7J8FP1Wuheh14zClJdE69BXJ7nVzxODro2b+gU5NVgm5f/N
qwgMTBas/WcOX+iZpp0iD2ZRXBBCjkKuOq/OZ3eQJtYCEK5Ihh9A7YjcXE3XzeSNtVxswmKQPeCy
mBglbA+/wITeNW/+E1c7SJFNF0nW3i2UixXZaRZrtUeL0rmjqyTW/+AOW7l12aGCQQQEOA+p4KPl
HJtFcqnfnFv9Z7e6e2i6TYOrQYsrInJlT4YFZzpfYKJ4aQkO9lgt/fBwSEiTA3ix0toItyZlX1VK
o0rCT51UjbLpWjVWOdwVDU3sOR1pU0Ek6PFS+86H2B6NStW/Zpydt+h9PIL7LMLKo6fJCivwdv2f
BByM+8pSk8s+Gx3ZqWUxi9K4y+eCGJdDknYtGBlyv5LVLQF7HpBqSFl14UhmUK6JHRuxl5ud2zO4
bKEboaL2Ot6eJYp5yI+2oDeKXumJ8jKR0pGIDXi1lGD1iPfwOZ3UVRvi0EhVxXD+zcBwXHI1zRQI
2KbkKHM+cypuGgoYvzQl6Zq3QGYyKIMabG3jakqGDsgRyUiAWUsPZERoKh3MGttC9RS6Dyfn4/Nu
pXxASnfjHYwCYGClBT8iipw0iQCJNVHNhKzqk4uMv5xxOvTEKbBIKCVooiNaSbVI0WrXu39IXA2k
Nl2rcF/Vh3nzDFOu7jKQE3IMczGBzGCDBIqZJcTarZbQCzybqzlTJM+FRYSjE9wJ9w9V8E9ommCn
kKdUXlLHcW21/hWRRRIObozfjYya+D9boGkNcK6Os/L18jvROcO1FXB+qWpoWuttu88hq3iztR1K
ZaF1G/Ou25rabQzGI1W8z7Ixh8gRNQERqvYZ7raQAWYgrrSCZObuLEuhnBQ7cP+fLqJxPoUWVZsA
TPyrbzdDKIVyIpUEfImHDk1cjayyNsgHPG5knJBILZclZO4hrX8L3hV9XUzEXw+cWLgnMpZ2MIDq
iCFAWa1r8ok5F2nZVmor2V07Auge93WiJCowuvZBUPw3gnjYtHCH8+1CEY2PIAxljtCsW5NhL5+c
4neL+i9kaIPYp4f1GKr6b37MeL+swpQKlButw4VftJqgVSlTbRWIsG2WU1I45laxuT1c3N+XWd9u
s3lNK/MVv6dxyIT6ywrRnu4Tto/ReJSXl24to0RxxiucliFSYyEItGE5WdYRZBWXhD0S1NxRzFmT
g1RDpvpBlOK/XWHeHYMeDfxOguDc559b2B3kw8+J/Utaiy+JgYJTCzIEBtU41GZ2oN/vWgU6xLMl
2H9uGNtulzll7LyOikvsfTUrjf9doQnonrjqZiH9N0HR5c2/hvwWi3doct5SqKdowdw9DLdPap4M
XpMWr4bxlMUJf3BgK5g9pMvDnihVPbf04ail2ou3iDOzp7TtxvlzE6+Hv2LBfJYwP7fjolTTy3lS
4a5xI5wj/3a+JZeFB416RhASrswVlbG2HKhgRUBkI9VForLlnTyKDX1UcTYVT4FAYpW1jaBnvFgA
tbCBv8SmjUqGJLoq8IEH7Yle/CSyxbCLRGvgAbcW5jiyAvyo4f5j0ndTamQeNKSr4bKcdUDZlV73
6AwTo9aXHKohlQKyw85MpLC/5jtCK/1QF+xFSW3aKXswQAyni4r9iw4w5l76Igi6OfRnFS2PlqEO
2qD4OfWtBI8u08B9x49bCVUqyGiPUrVwnJinTn7Wb5w1TfS7o+PRaqoicmvNSdlIFWEy42ZcwUee
gU3/ZCvpLDOPrehAp9ilo+He7RU2s1/7Uj09PnyXQqcvcz4h/AEB80WX4U/cYXyv9B4+uu9uZ0sH
SsWxxo+jGXWDA/V0hoAnzQUT5pLCb3xPhHXJ4/KxmnbQQWjPkEEmQfrY2Mm8+73Fx1BSxhH4oieY
wpVK1rUBejglqhF7R17CJ3swRkbqihkZO+3u95o27HVo2L7g2SyPG6BigS8Kxia6hQM5eAemp52U
i7wV63ec+bcFA8t4K/iObGfBKm4IlHaiCNFQ03CVvacwGCvj/yOaJL6EWin5n5Cwghd/fp6yOmVU
+C4X3EHgiI+oOck2qj1J9dkRH4GiCjbuBWcH/Lxvc8zUWAESRZdwXCAKaoto3ixRJAJfQA2H9yau
kEAi5OiY929+xAMBSmXkyznnv+jSZhcNkT59MYI79UdOkEvj0l02xWX0LZx6laajzAqM0qwKvT7g
uZOKu93aWLfOUlUtW5oassCUhI/B1KNiuQBQopbLmm0/cRZmf+V5LmZyIx0s/aPEdf2IMwy5ke/J
3u60udcdHpG2dF13hZN+jCcPZPWpNbBxkemkTa8d5azDmpGW0x3RzqPa+u54uZjedY0M5ZikDR3A
AEilqOrDz7swXsDmoMp7qyrq7YoXkC7OFcab9bU99qcc8B1KuoffUUy3F3YmOE5uNxdia4j45R9f
9KmcT1wGMpokx9Cp/Q9ZMP0C46OG5zJfPEdM5FfvusWun2/ZhVIz+Xxk2o/nniT8NJLzjACZgL2C
L4GVa4MUZmkLWzi+8K479SGQMKPBCGpXJYXBVeYv9o0Qpvhi4m9AkbtmYQJYSDwvR03pMmJQWEmY
F7axW8qe/MqGjfJ1Jc35/fggDCEPEyUzb//0GzDxf9FhcVHXMSzfBWAiRk6f/Ztc9hBLl6Q5Hw+p
6jYXCnJFX8/ENpu3j3t5PJnf82u5D+ugUIae3GvdbzHuLft23/Q0LNqO9gR4TuTAeiuu4lj5LBHw
qOzYa6zYEWuduyyKMtGspUCSlH7elPyTi7ufOTXwSPABeqTeZ4c15N5nGs1A8EFsiZtot/652pdP
zIe9Ho798Kp8kLYKVgQVKl7LXq45HtjRZMuZVSsng6memq0xNmz0DHgzQIJiXTn7pnJsHJHWM/wS
iuYdTdAlzHFShDOA8tCzNEVsPYyIGttIiiWvt3gre2r0XmQEF7ZnvYIlkSu1q/hX0KZ55/Z4jY6s
Rk1fDPfFM+Wic4rSn/m8hU5IVbYGrwMC+vSvNnY9pBuoaYTEKpsfa/9hpL+3/tyNJ0YS2MWNM9fh
z8njV1N4dy3ckHkhGpuXbz02Rw3upPekZQu/+/M2bkuN8CoXRe5X5E8MO+qCAH3uptmUVCVx7+/B
m0k01gyjr7mjGDKaqENH15nl7PLw9zhvAlTsr121d6c9QFHecN5OO8ZdhlFNAxAgS+k8pj9MJAj7
lsc/botWDonyGdKioTcqmVwPJnGtr7xngKzfjxMzLqTOFb4uNM+ptuApWyvfw8uLmrFK2GuusRwq
eihy9Ij0BVGY4t4HJs+rxQMRFpasTfsG5rMiaxhyLCqlS05d3fEwOLzxRR8CZfpu10cpHLjzBeId
rroKyRQ5QBPtw5MRP68RI4y+QnXkZ4gVQDJAFbCkz/+foHQgcJDiWokcrOdm1hP3cW3EtjCF7Nje
HjaHktl5TCfWtMyxmA8S/7grJo58KzYJQ+x+fxoDhv/XQ2durV/25FW8TA1xSjGYrEBKGuF7xSoY
g7qAexKqNwlWih9DLYhvfNKvaO/iKEaS3sHzR7Bt0IHZAtKjPK9zdsK1Kqs/lYpvp3u7U2Wa1kNR
rlYaeg43Q+sEXynq/GVnXgQlU2SGxbdUHw1xMDf7fESChGozLm8G0LbITW0yTbbQP0WdISkaTrs5
bD26unyOEVdePPS9ZnNhP7BMEPe1gksJt/IQIhnHByld/Ik/+yT62uBm/hr1xQXawE4nh6qfohXQ
DL2LUB6OdqxzAqTEXLEfV+n9kt+loXdQI/BiRN9UuCNukPwPXvPJh8geRdq/BqYpnO+J2XOwVqu7
UBsR5pY1NaSP0g9y62PaZU88wY0NK3GLsihg5wM/M6c+wEctPKMl4jbdFn8uGPCAukHFDup/+Sch
t7TaQAfsNAyy9E9J0ezHcI1KMJKTFKJY6hSxcnRuQh3UAsxDLbbGbHEhQL9pC/weMmk/F+FvcVJj
Go+3ftnJiqiVDY8JjVXhUgEaDW8dpYoPK6pfkQ7MR2JWwGWoS3tGivuyUwv1ULPGtKxIzjUk9Yar
V+D+HQ5RZ8TkV/pb6/ZbHrGr1xvBU3NQjWiy5F55sqISazo1gtKZ3T0O4TmEiji3ohKzo2OiC79V
PpbponFQzQ9jda4KP8FnQJKfOVtnCk/U0tycaECqXR8EfVHv4AT9Dh1lWD5so1hB6IyDf/0fgpSB
eHZ2z5cfYr7s3Y3AvcEFRO2pRICix17sG/AtAjd91Z/eWXuftW5BPuPIY+4M+D7J9vAMu0Qr+9Sv
hZof6msdWDQ8RE9M/XrMRn4w1coqmRaRqrWwK21X95qqY4uczxh/NjrRDoiT2EUDCi06NKGrphfh
GWO4oh6TmXdqCy85fvHS2N6hJwafPWl0xfPT0B9aw7JEJzp/qdcJzKMlwF05X6moHo3HVlhj6CAJ
/8ELjuh/nakTHY16hClR/jIxxC3VV3ISxSGeeiSlOEA/KjvfUWCcEpPcAjABFRoglxAJf1Fj/RqQ
IwEuym9MvILhPszBEZ2qXgTF2Ukdqv2T6Cr7gl+Q/6GYRx4dsDieCapskLFh/dC7Ua6heE8RHF8l
IlrS9scODlkbKGYRxTIhFrKd/S0EuS20ToFH75b4CNqBSOqFEfmsKJLwtHYh+47HTynkIEpVsxta
xwBxPZrFFUojci7cW4OLDjeCTgqYhKDgSNGkypAp7G0kn0/M7+qqWcTwnAn+2ydnKkyW/OR6VZ51
rEUHez5bRTjAKydpqhab4s6fpzWcxBx6krnfgoZFz2gppaRFI59ZxU9LYCTn4zWvSqPKshhnIEC9
3eoI62KuItbpG3PdCIcWx5fSLVYSWW7YQZu/KdVEBgrNwKEYko1lsXOPim8Y6FGvLQZqrRQx7AIG
c9AwHVdhgoJXw+1LcvW9v6V+1Md+hdJitV1QRzEoHMMiNFkee0SR7qEmnGyBCBDkTFZY/n9AUIzs
DJS6C9DIHtNeqSZenRZU4mpt41PeRBp5mGVVqjpDGL6UkYUsk8OUh8CgY0ekuVt7cZ8XmGCJdLsq
zoHVmvHvxCd/lJyR1RbCKlAvzNH/RDZV9wRqK/+puVGGDcgnlTGRT+FpMIl6opKU1GnzpUQmM8JP
QZSvEgg4Ob7jIBor7T5I20lfu1P3D7JjJi7DKEUm0uTMj2QqtMUSNVxkwLoqx+A21KzfNWpm9FGR
oFjF+6YEZ10LBAkGwL22L1+vMaWGGiKYxUoB6VizC+kMprqeHWIaC1sKM0B8X6wQYJUbwcvUzcMp
FsmEaGyHNYSFt+FLN4rQZ38apPfQfuNAf5wKbzzKPVGUPRGH6gUadolmnQJjZwBGCKy73AGlnNjt
AYzTp6gUPYBPnza4jW/ktDy3rF/D7qkRfBP6Bwrf5z2ZF7qQIbuF4r1X1YmWFQvxd/B72T70NWww
I5YpLelnHMd/es38118NM+s1txcSh1e5skz17cN2Bo6LCUDcFTYq3i0p8+pwCHhXrXh3jH8FdhFL
ODkKWmbU4Dg7orf30tyiMUkBLW/z8PaMqx3Z9ARVzhkDYqwDowxHWXEy4b0qR8MIqmADcDKh5Q+Q
E2ipm4HEpTVOUIoXApLxoAAXsjzhwKTq1/Gb20Y9HaxGzyAim3OXXac760K/LKwNtG/XLKBDm75W
FycZnSHN9f6qL+zxBVsLKg44a+9G2MmD5OFruKksLoFHlvSWvU2ZRuWK/hbGLNAjsfdU3HiWi/KX
sFCcmld+3SHap9K43kfn4e8Ve2pe+8bsjnMnGjEPK3LDqHzYurQQ33oecEFE3nKTsYWuCuyah+Bj
yFtBILWR2UwgASHRQgDgofayNrpx6CuZu9t9KendepCh3ql79489n1XkU2/BJbnNpZMl5IAMrEyL
LUWQ2s9hmWh1vHF+x2AQl4s55P8keDd2cJJyY123c5THyemHT57N97mvxXSXQ/e4l8wP7ZjiHFE/
OrKhZ5aMtJYPlSiEjOCF+Q8D3orSwJRS2TFZoA4hrHt97p0J8x2/edPbZfJRWTGTrYZrXhkst9c1
rWJS5z3NEUV0hqBOtmq6oWMdVrzBsQix0ilJHGwWpzdgds3tmVsThacM9g7VmpdrA/0yMQp6i8IJ
MKm/WM/EykCZ7gkiZDUM9QYyhRNFNiV902dEopKJu0J4yyGm+P0Z7jgIZp4PwFiu+mUULzTgtPAY
ArJvJZRUJd+7TCHg7QwVbyz0+UoO7htD/tTrAqQES8H+pVBug1u+1xIFgmKIcHlQZ5VgZMOZLXXe
f3JyAVhwHlF/Ix38kPMCu6dtXMewranbB5slcIw08cBG9046g3yesKCsftKFQRu/yYYiGInWROna
CSXES0ElBD60DtkdS3yvsixAjtaAy455AytIpyT2Az8a7ruF+RFpMFx7U7MfwxWAxPflk6UOO3ZM
B9tnuaePgRMnCR46/TUU4P0XroWANhc58Dek3tNAZIaT8HJrN9YmynrONYWb/JmX6T1Z+yZu7yJ6
AX3EYqn6DOQZ0dRg7KO1pCt7Q2v235EhSIkahP7BbcB7aHVW7N8cqNEng8gXxV7QD+NBWNkJTBRG
/E6ssDM8Pg23G+uCxVGp+k8RvG5/NEN2eWtYXikpDapNeefBQiEqL/rqwlWfe9GH2Myj9Ij4otAz
Nc5h/oDAnYeXtwODwO6jq8AbvQ6P2khP7Vzh+xWcjnjViNbgaZwuyDfc6UNgg3bto5asLthKgrAc
6St+Cu0zEm1usJFd2snl/qVC152b/sUEjQUcWWhAnX6TGZ+B4WhZmSQDqbJlwk+xO9RleG3Tt3fX
UgidXdXsLn8MIjU0POnQ++LuJP8UWr3QbU1FQA9LlDuHq1x1TceFrmQeIfhQCb2/v1Qb8i++OOn5
44I/zyYXRzIgpJlxzi6OG+cv2/Qgd843t5DpS1eVLbsj7nSCGgKwXeWdL+dMaMgl/B8C+rEg597W
wAyoAQrVq/TbpmAgosbd8EBishcRynRHwMsoQU1xsIR0vYZuyjxX66C3Ye4BgwkonmlKBTItTbYC
bwjnuerqcMOCY3KiAk1Gp/ZGpvwzba3Fqk4WLMjPn5fkE7/euf0ZEp9zH9apJXj9ZhTUQUG/aOBu
VE7x0Y+MlBNAxQNa2Wz1w0YRzExRt1QJLNJ7hCLo+yt24nYByNdVPPILCPB/iFIV8vsZVROSr1xZ
iue2JzMechuNXARKr+sw9rY0giE7ASdSH4saxTNvEvVlmz+iffVGhYqp45gNVT3B4lX9yFS5tPv7
F3rjGnO/f6qFNpqjHdM7B9honD4ymMO7bua5QyqCTvtGO7xZBCZPydqtr0e+xeXkH1OyDY9MeehS
dxuNl0Qq8UrTmyezwIbCxHmYNZBDxzTTQ0rqXlcypSU4nSNdWya3rSQySiAH8ZYmxQo6xdE73Nc/
bQ+3ESb7nOOd6xUyVzOj3DtGKA9wl8gP65hvYmxa7bwtxDtm+l8cT99EpQhzl4A8xXcNZN3sFfUG
oVFsFlnhyRxvcu7PBaEyFvn+qvxBtIgOzHjrwy92INbi4/UGyXbkTqyI5gy8+mjJGS7yq5x/+bGH
yry5P4J7fNc8kIeOdHtLdEem9hs/eLGcxhIW8IDh0KIOa7xhERNW+X4h9XYi3TBHhmWvCeek5uQh
NXIt5xlUMvPCjCS5VJIa0xLyxD+c17/EeUOTbJfQobSeLFtInDr7gfJYgYOTXTxg8Y6LrF2NTaH4
1zjZk38anp9azDaH+G2+sIx25hy2zz81DUERtE4A9lT4NJTXMnPF+DgT5ltYzmZtB3k47VIJRiQD
Ty/6ufZ3feCiby7OHmuWD+FDA/8NDOzGqyROYqTpqDnkaP8RDifP6v0f+lddKRjMQSyTj/ogF0Tg
IAgGWuZy6XSHT7k4H79g6Ayt6YAWFdMNWR1065ER3kUuCHodENVlNnm/gerZx7pqlYZvCR72Uya5
3wriGMqd2y98nd49sV4Men59OWvpdlR17gC1gQ0SXS4X2NHlNVdsSPFqEXQWYj5/vWgTLy6kYVWb
lMRoEo2+8oC3dCCWsIU/01WLPLgwwDRkLPeYN1w0Ai2PJhiOuHn9Akou7wqSo/0wyVCvOd7s1pzh
/O//6t5SaScnShklzb7KzevOiG7qi9cPFWUgfP3iYBlUNcBSl1Vd0ryJK0AtTL8gT0ytfpTkVwRq
aXycGE4JjI57AVXHHjnBt1YM4YLSPAa6Xy0gWyxHq496M8ei+wE+yB7IF7nm+iAydP0MzSZersoZ
arZyNd8XYoGTIW5FY41e/lQ2SGw3kHQIXCyBvAYo3ZzHrjvimhheRYoQsC42Odvw4o7NLzXHMPFT
QIiuBMrG79juztWfQWWATlgKBtcxriQ4TYOb4covMicsFxzgQlowFJDenOWEcwdL0XKbr0UAxde6
BsPvthlFirM2B6ffSbN+cTElbfqOFOqfbfER7xbAXQb09fRPt6N0KU+uuT/O7KQWM+kzSGI9zwdj
ZivMo9IjM7oRZlgKoW9ynVzFzteRGppe8f4MVtSqLNxhjNfgSGiC3nUSYI7hKJG6jCUsccsqP6Vi
TtF8Id5Bh4qcID7F2sWCQ9h/GLzHCOJSZLKWLGkQAjRcmk28cnii7hg/okzRW22P3WhxWOS09gv+
oS7Ca1QXyIz32yYVehAK7Y4/DxlXxCePNmrINK9XgKG7fnavmYz5nEsgZNpBTSKjHRlLuiNAPUsS
Px2wNTPJ9w4/hnVT1Lb4dCGSgX6H/OHo+mbRsL3Ry3EuBgev3m7/cg1WkW25va9OLt+wwIIGP8kC
9pjZHp09uAr3Albk7m+BwU2rdgfONmhRpmzI7b79vVPI9vnqodvsCEhCA4dBNES/xT54lrnBS4Kt
CVVMRtBCSWQ5BUxARKoS8QhTIkh9WTihVXw1sW2YTgAaAciBf+31E/w7otybCZYa34nrDx/cjEPD
fDn33lp/Rm1nbuMAHhZCABasEcROeAffLADpM+pRW0K3IKrcOxW4w//+Zlzo5VL8W9G1PjjY+b3t
6RKqgGKxst4maz5JFDxj3fZz8XAk8dME4A08jn+ljRfhBKvCIXv7nzREBsYaSb8+taGxzrEpynT+
Fnrs+h1qIWr3F4pvrEwXD94RUixsCkBxN2D/PPpeunyn/1Y7vClxjjGV5IhXdXci6VyWsvMNJk/f
qyU3XwMsfExEwSz+jJE9HDX/O1DNNHgQtJmef1ZC3w7TcqfuYFV/j/eJnwTDsNYfhjAe11AgU4px
KbSCcIM53lSlv1xkq9wycqPQqzk7C6eDlomhNBWqrOrG6t7pbbYfvWO7tH0z9Hc2hOZ27c7l5w0c
TRGvzQSzf4w68Aq65kreG3NFJY/DWbTx/oot/jVfYR0efxbIqAvSs/JJiPKfR6Fb3ORtCW1i1TcH
33z4VOTazQq2yzlKGnVhZjAy9DhTqJgHaCnu5z33X4wt4DKQpVXmnQxbmwc1rwL1gE0OHtH7g9Qm
IhGNvNW2KeAh8R6uAyYEbiWbPFA11W8NDwkC2PaXaiD/xY1Q0wgJLkmEN4vXr8d9TtkDsCtyNr+J
XxlYJ6mEaDHQGUAnynN2loTzvF0KHv4nkHIGERR5hGaXsIIVYSgpK830hUv6fYYZOYY8nD72Oj1i
BEjRytRkluwAm18rM2Lh3ToUWijBaErlWY5g19IzBzLXGSO1aLBBQGie1WNolrPIYx3d3miwEChs
fCNs9jEiiBrKzuJSjOsmOq1ImSFRUGKGHbQmZPNtCbPUqbcR2d28f2M46PJUBGSvXl54snraDjwv
mERyZmMcJBd/Jh//BONWyWc/FQbd4qUZBw0OtJidgJbKTFTJmwRnZ2dAg0fAQythqMP5Gt0L/e3c
QwzRxrUAjgJZLuB7IuMnLiyBqCp/nEvVH3RBj1Qd3NpD4itl9XXOdeqlcnp9+WUocAo21VFGbIJC
YXBDYKhnzKdSPX6eJoNCdnDDuub47hO2r947CLDyEbN0WUN+g9sAqpaG+twSjBqVqQOz2Lg4A86m
smSMD28IzFtKKrTPeOn7E4C7YcpbqehsFsQYD4qSvTrlsRRSkyk4jLWaZvjR/0Y1WofkyW6v620r
jXu29CWZPGwkyjxpI5XIHH4StAk3LgqT81wFDpEf8IreOHeM0cYySPJKe1t0SZt1yz4WFdVamNma
7/hZMRvWv2HLIa8HFoz1h+j0hbwTqYFYDdo9102MLd2UzmSlhJ3FaFVDZKbLXVcIiD6dPWN3qvvO
HsZNeNEWs0lz8VxPUbg74+bf1m1YEBHmi76ItFSkOMGWMoVdbtcxNyD0gIXVa1q0meuTkKs3RHE2
VjjwH8bDZcMWe6N42bIktmsGe4sB9uR0N9TmBfMwOgpr1elOVhtkdIa/8kewDvwhsIz3OPLy6aMm
pbuqAr6u+KKAB5PLt13EV/d/tqMR+xyEvs9FaWqVX1Zizo2huU76cU4Sbp67JVufVSrSJgSe3KsU
fiZwpCefHI0Fc+rFNVQArZEnftV2BlgIu+DC7gLVaCjJZJbV3AgIAGnNorzF5+4+b8IqpYL0K6hB
/+xaZjCINBkVcJ3/CoFZJIZdXlBuudeKJ8uz5BNjrCQHCssnQLx4n4ipJfb/o8RPEFbligMIE1S1
i9qZWmdz3n3JUrdhN9VU6shpnroz1ML+ED9IBWUawRWKOm2EAx1/mYsKpBJhjYQ0yQl/ZEGrHzzt
SvVBLyTHOCKHO1s3I3ngdCSquo4kWO5YBdqcExqSHbd7kyPalyr+wv5X4jpDRq89OY5NN/b7Ifry
dQMlX2QRUiaD/XRGfk1M5oPNBSe4I8eLJ+r3taKlB0zeOKWIcnoOtrSioY0Z5a9rgIBeGYZxh9j/
ap4qadN/d/DUxHdaJvxJBS37+jbfUQ94iiUwHtGLl7v8LIJZVaf2gQHJglPncfGoI9iGITigT55z
d4sADx0zBAanGbfurRvmJAErrJm3bSVlIVioakVqX1WJD+4WJd8VuOZwfWXrkqH8unoRrxnL8XO9
qLdU3uDHTou8YvT+//kPu9E6OSyvAEapHqr+Mir9Pntc3CB9o25e2HuA3zpu7oM8jP95J4ZsUiEW
5Wsgr+PFsXRYt14hgnK0vLMp2FcRiFtRz3QHOz+Rm6+1diEPgBEPXZgeP5CAs2X04vli+tRdmpyR
tQbFPz0pZNz5cJU2Jf9JtIYLM//a8l9p2rykntBzT7PyjFrvDezm5wdqMGQC6aIKlhnbZKye0/dw
9Mt4iUIeC8REI5RXoJSZia+x92sfH5M1EXa6o2FFygSfstt7/cF8Du94sTUlOieRvtWcjLNsXnds
8rnyq7hCCLqFzs1DSk0xj9BOtxTcz0+WyoNRqPHiAhHR+XZmTFJfMLZRotPc9UJH1pnPL5LSFGyE
Dn36XflSvNz0Rwi2ktCLje9vnP6jLBiQf5H/IJAC47COzypK4OMwABGxsm9kfcbip5Sz6dv8GtYi
3kl8yjuAQo5ZXbuzWTIOkjbNignFYJUgmDqDXdUj00L7ErIeMnGaEDsOQyQD+2QytndmgDfh2v4E
uGPZoujAmkyqCeiKqc/4ERyqmc5/bx57R3miOzstrwWca/JBxZ2TRYHEZNNJj/vGcbEeX9n+Bv7R
V1qtXVaZhwyowiHau2iDr0X6Lon27PvyZ0wtYXcymQsjvfhrPbS52nEDST6J8O/jQHt6L19iwPOe
QKp53Q81ZJcMeTAvtstHjPcFhB0RkUulI9W8tlg2Qb9tyvmhtgAT+HkY24zxVwR+ZLiP1AWUS93G
BsC0aiyegqyh7eE6UQZsPHUnk3P0Nxh/BlI/Ic0Kc/c6aAX4EIpBZ8tg8tcwm5aQl+dU/GIUpebH
jciWZIfenGHlYyvQVIg/UcIquW6Rs9RpPHsaK0QZRuCqnDPRBSTFweCTpirmtVG6Lm0kfuXe46Xr
AiybzkQ8v95vHb8RGVT/P0n7e6R++0PeGg6UpujpFMkbetlsF8LXonIYxPeH40mN+KqH+S/YbPbT
m3r8kPeo6ufth/eNwjetHSEsk/IkQdWJlQRQjlI8FrblP3gcrc+2dk8AA8zOCYJyfypEyEsWOfE9
vbWOoOGZJSKVOWTlc0TnUwguZm1XykL3UKdkJDhZFdYUbHIaVjXuFxOC/RCJYLQgGkY9ywlncw5s
cgz7dOXz6nDChbvly/6Bx3GOJTg3A1U80/529PFnpLPTHGqBu2oipVG1oIcl60mBknYIsXbZ6PRf
oHypU/C9vPijKmt8BFXLLIaKfG7WxxVNVmtQTQbJzTe3ZPxEOgIUzRxslc9whtVF10YPD2iK4tc3
LoQLbrLEXeaabfpFyeuNi+I4WFeqhW5WCQu6D20dcYPqVQOKGJcwHNvap+8bRGq+rsgRGYlmUZWd
xPsA+ibeAE1w5zxOXoien/LoYaugiPw6sbx1GzTlzaUdQ7QPyCws5QxPJYpNmd65iWbh/Q7bO2JI
AZBplvfAiohpL59VEb1azAKWH/l5hTytrbDIV5CE2m4dLJQSnw6ArzxoFxuK0wUIfNhVsNQs0yEP
FhLz6nMH12tY2ZJ14ulLEGZ65fW9+u7bTUQs+csvfo/OIjYYqsMT118lWPWNf73ZPNIlIyk1x9WZ
vPz3hrNWfFlD07KJafD7GPgvzm4a+dJKVJqLlTpM38JT8on20FwhEXtkJBagqJlgjpi9oIsDJxoi
NUO3OW3k3LqTDy+OIp3vSrPEg8Ll2am/Htr+RCuLtl5azHB+WGpPhb/vupbdD4F3aGFqjbRwonCs
cjBjzNQBSt/nysybcJ1uIqVQetk0mP0CpIBRlhLl04awOWcH0BYlOqduhsLs7kKlrBwfyrrboziG
iRXXPJLpCfC6bNUlGPRHPoct+tEbhMimPEbUzH8olTQldexVnubKCmLqV8kRiY3Uztb/xLq8t4QD
BDJJkDF7X/NHhZdvs3zQCIylDzWJOd78xLjKn2sE334pgms6Lmtfud2zzqmLrLOU8VmKFsZyaAu9
/JAXKlbTrlb/2znNwcC7TdWrYZ1YmPAC4/lX9rouJ66pieUoM6xnjV5tGLYxVtrsGqis/mdWF6uW
3UNgeYEOwO3kKEhxlIBJ0WuTXF2OIgZqlEByYXuRnzChv3NmTnwlLDVgxvNS6ATG9AMVVR2/fmeg
RtJW5mYwS6os2uWYGiyjcDJCUk8Is74Rr2sxRVmUJVvIzdb2SmgptWL+0/p/98AlnVbAymhl4z3f
lIADqEARgGyqCUGCaku4z8P+ZU0FE+TdZFmgHg8C0BZeWLh+dcSBM7BVCeK167JVxSMD8X79sFYa
tH+4q/5lFWs2SN17xgPGb1qY/PPCZJZ0H71HFrkkyiBb2Vzmi4Yvb3e5wmyMmDWB8f6jf2ZMQxz8
4ff/2Niz+vHdSc2fd5JCo7ctgqK+8C7DSVsJd50LBGWBaARlrLrJNj6okx7idr1HspZwK0L7bHui
VOkYOkrZibW5lkJOaHGgfDpDuHxNvyrm8bNHQoaLBdr4AAaYqveXI/OUC/d71JnSLHXj9CXnVzZy
d3uQ28vo3469GwIZ63qKu68DS3pGQgDd1QWaDw/7aQLrxk+ZuQVhZBle7xVJifGwZtLQ5C82GFIJ
1XkZCMUm/OnVye6r+W1TlXvgZ8ZB9VXiXzbboorV3Q5N75pS0Tx4Jn0lx0v7JpR+QL7CGCAXXoVh
z94J612NxGBBGyq7u9gUuH2Zv6jjfOzF9vPvFuGw9Kc9Yj/Hn0OrzXffccRss/wVYUiAZ2XHJNZ4
PidawMWVPj5LUK3xpiAyLU+66Sld55oyapSo4pJCKB9CRwtAkXSWuEhb3PJD3tTZWlX6TGzldwHd
gg3FFFPQtNnGgF2WDrFf+VWjbhuCdUEglxt4b2+92fn2mS9/4oCTuJ6tVbFQnxEhumZ3au7EpNH5
CnyypjZ6SY1jsLGenjonM/FuEeBjYbjfQsMhmu249jQJRpEDip8bJkgRV9GJTkEc4sIR1B4ysvqS
PVHIbaSHntdpCqqVK/yg4X69K8uthCBjJwKfCL+UNmIL7p8jicNUoHybmNjPIQur59NzMLRS4z5m
WlLIi3t/BzNZ87NsXVK9nW5LOJImhGJ0K8OZf02ADsxBQWB/Fl8qniMhMrYFjgcYiBS3O/5vASq6
QOXI1Xu3O37/JXr89gRbFTXaUQQU0H75v10bnZyjKpLNEL33bqngjbXazcCZJINkk7p3V9wwX2ao
+3905xqnpIvaqKtVojWNE88SKDa74v6mVa2KhFFkwL1OOvcKyjXi5K+3shuiImP5FKGSuH8zIaBW
G2/TIYNA/XapI68IXcR46wKBy434Aol4qt7JYjI2qJFXohsftEmw7o46v+xVotT+j0Yh9RBwKa5j
wATGVxfhkelw4bnwQXAWr0ex7jCI58GnerMJ1jHZQAJ8MFvhiYPNHspIJYRgdfuQ9AqpOjtsVSc3
SoGfIcE+QtYtItv0Wt0EjrzqENY0sDfpUEQQyHPAakalAFoCcQ+3W01iEmqEbHETXn6fGWXPeGpn
4u93Gl5GvSIfZQDP0yYJsl2Qe638ZxtpybvsBWhONUnpQf4CM/owCWcyq9yUQo0IZMI/+j7mM3L9
xm37RqDbWSVfAs3wrl9jGMCXnmpO+ETybDxuGJAjLGfXkgGWrY7JRzqRQsABYBxwCfjlltdM8mhh
GgvxhYBWyu+roEFzLvKyzJSzQ5NjUDS7TuH/1GckNkQXyGG5dvkR3y1idK9NPFvehPALFc/knA/J
4eyz5b83IrsTx+FrEAICxhI/pw8y5x4PCssj9tvxmv5DOJbC5QP3eEC6ycTDGDVQ3x/oHlhWWq7N
IRmZPHAA/Eftknw9pJfvAGB/Xwd5K3dwgSzuL4oMSDGSFhj8aX4qdACO85+4P4ypfK6dvODkq4r/
v7iJVOIRaa8b/BpfHu4IBAqW0RASHaOndLUbxjCQ2GM/wgJyQFbxWT2dg0yyutdtWDCcHoI13E8E
lxhkDDh2EwmPgL0DSbiUfPGYOMuK4NdfvunsTw2AG1jwny1gV5GZxg9UiCgSBq6u1gdwzI25+g61
ZtX2NNmzfFDbY1fBq4ktvsaBPLYxniMQBPTVNbXAxoXjAbTO/Vh9T3nl+6Xh6tmISpHBbn3h0It/
YLIDnWbSjuLGRJpskw7g7u71SjAppPskPELvjiBcnk6etLu8RddVWJT6Df/eXl4///g9qWvbgyEd
cjC04QZ5lNTb2NTCkcly9uhCb+Z1kqkoLHRXts4Nt9yQMrWcB+uYzr69DzGnnx4Z0COX6rk53ver
Of9NfhFYbyBFVQL0apBTH22iFDzeWPCUG1VBODOMza1DzJdmky0qi0j9lTmU14ZmQoba3HFTqRyr
2RooylM1Brw8XvFYODyiG8pEHEp0PbIflaxmgjYUoq/zSoYKX56l1rRZTCdhrO6MlsjVvy5Z3VCo
O12yn5wxmJk/ahr7Y2mMPwUEouARcZcYexGNPWTAWcxkf1HlfiaUxxT/QNfTfMOpguaeVe0IheAG
KpiKgJLB9UTLO8LBdqyEjAOjWX+5dKCodoFJW3djiuVLfttLZ2MD/XLem2vFrSDjGCjHMEBWJL40
6KbmsyrLnQBRgMihpATtgYBG0Ktlzeo1nRoEJMwhm+spFbPP017/6S+laPI/n0TELuyiFB9Qz0iI
qNx8vXVmEEpFx/i8fVXhiL+ECiAyxIMtq37BNhg4q91NXFNUo9BGuQlsgT8ZuqlDkM4JGZ7cVP9l
00U0MItIXhjBClEuVdCAeaGaJxbfBjAn4I4MVCU/KNSUWEjx6QxqkQRA0GKXmWwHM8Ugq9a4IVst
GTjJR3Q9CvDnh2n6bL8UR7il7RWqTYNP5dJsAzoQW398OtR4rJAigxQi6jPNy4KUlwsaN+9ze0T1
g8YDLPhjdxUatIdNJFTC5rzJ6sk5fa5RUI07EVMGW17u/A6w7LaSXmgYGULNvQrJ/rLanOoLlze0
YdNpZ/2uTFz7EzFVTLBxfG4qfWJlBLMRHzCsCB9QbOhfQZEUGTgH4gpSVcNDS9ENlS5WE8cA90YO
IFCDZGFzT86STEPrvfoj9QQfy+jl+oEUCYniUqzsFRJCdJJP4HL+gSCCj7c9n6V42GAzhghsKJxW
K1gDkDUPowb51BAJS2c8TJQfPk83BaL2I6j9DOKMDPWWp106KSlGhyH4zUwM5uqUNvwHECgAA5A4
chKG2TbRhGvgf8oW6jtu9XVB5OdlntXxFREwjRaWNkvLNiBzZgQeAFP5FWGdAkzA7jg3FaZ1o9n1
UcXuiFCuyLOWW4vvDlendLaAsG33sFSuLIcrEZedVeeokGRdDY0NxFnUZ669xaaKxi/hBx5bAaWv
V1pJdVCEp/NuFGBIUp11uCZYaWOvMg8mYZNJNpq3SsqdZwTJutFdZ0kRytKSZLuEDu/4ahgZu2/w
2wdLvh1HEf4xlvB0sKKDcMuHx8M60P6yRWFoMJP4YH/NeY/OttKisc/BR1TiE9a5pKeVvxEF1chC
m8gl5gssEEdT9j0pHM2Q7BxX/BzDgkBZyufAaAVz5QDttuCsPWYvnu28fr23dkIlLG8puLQKYv8B
X4gp+FJbjvNh2LP3SvssqQSXIs+KwYiL9zdkroq9puAXGuYH/Py9E+MlXhFole44ZFA7YL5kMIEa
Cet9nx7JLp6r3jXVUdP/snydqTWXWAygE7uxXrBgnk+fuw917Z1BBO1eQqdTqBNxGEUAiHjTZiqJ
HlHKSLVY4dCWh4KPvfpt4VccNQsLKJjUj05gksCPyWTfO7bU4d5z4HVIOAJjyJsYjxyxlh1Mm5C5
BK1XO8wv9tm1MFCRPFZnpfZKDt/9G0mBt+Biv5DdS6mp7Ob3hpV15dw1I5dJqiJAkfDh588m72r8
aosUFxolyGsFXaJlaad9XEkh3UBcXe4IdKBGREuU8syYQgdp3Pu3dv42i2Dkh7auYAO2XC/xdZ/j
adHY8BOYqdy+DLsC+F3blofyfHJEA8CCvldX+BCVN2nP0IIfmbngd/fSY14fbc/b8wIPZ61Lzfhz
+AmzniaJ7BqrNOiaNgMDhM7jm88+esrTDHfqptAHe89qdk154Ubjx1s9yxhhiVWbReVfbGGX4TF7
kzQVLJ8Wt0bktGMKuYgTBfANMG1jF1/J/AzEYXqxfhhVwOBUTFsYpjrW4bGqXuLQLz7zXFM23B/E
Nukl4v1hIusCZe+jJOqxYN8Tu89Hmj5CiEgr6Jfbr0NwXC7UM3oSgfOuWRi5GhTydayGTD9paT1N
iRncOvZCzQFCT2qQOV/DPCxTHY/Uzrbr1jvfqXxa8b9NxhiJ+2hewtMPY/pRTAZKUBHpI33rJXPn
xGdKYJrQXSjgQvabP/OCSFAKNmwW8rXD6L6hpJDQlhzvcIDkf52hsv82RxyRbW9hei7FRO7Tu58Y
elrcWgHWPXT7pyTAuleqZ8yPs7N02zneHVQHLVzwIi4bZHMWqdBPxNaTUuWY5IH40yvzfc3G0l40
pB8GO16old5EM0YsR/+Wa+gpuaWxBHl9uQe698ndkGbC8BqsJ2W+xvKUhG1WrQH/jDwDV7gcz2jt
u8J06ox8gSmjU9KEtdjNGcHxjpfqKwOVFB707yszz1dL4betwRdT5pPFTJi1z4zXpNJNSVNjhBTR
WRA5mh2vjqHRhQvrlP0iwTmiH69fTPMMwfWjQDcd/l5JQ0W/0Rm7OLE3KH8OZlzC4Wi7z4Odgj1h
VDeFvWqx+7NlB0paU7l1ybPB9hW4H5Dr430AwMJQ4V0dUivasa/H1U05SrTQthKFxx3vUTpLzGG2
VklmNFWrFu21ixAReTeAtCu9uAAjONof9pwGLFpMegZSIcuDyUwh/z/3PkVOpq18GOq+jnZsK3js
OwMtjjUJ83wnMl7uIJJkDFa86E7PCQvmyEd/WGrNS0fbrNTwqmyM++7u9c6xrjYaorzS2OBTKUpK
rCZcJGMjbkkElDxpo2/Ko0n/UpQBImORiDybRrLc2T3HvIFETFxxfT6m5ZDYPL2T9KuJ5sI1+U1T
xHJofw9LeKvSQGhm9BR2VLgxc24xsUC66JWLm3PEdoV7C41zctk9e+YoY4Kbg73lajiu6//jEoR5
HvgzT0AvSgEU6nAjh/FAuDe+szwGsabtZqC8GEVyXqJN0vWoziu+BWEYFCKs3PusiKjw5L5vBbjq
/gDrKIVo7owp10dtoeFdIV0PtPKXhNEhdTL4XHd6hHyWsJYMKgMjQRamI7ddYml/+k9n7NL1DIGT
EFLOmBWzeG6L31ipPejNAuaw5TLrGCXqGi5RFH9pCWbmDp9zsc4e62p+Ds3jlC3GM8LLFIw7dOH/
xTCNzmYaeCZKVjDfckKJYQWhqFZQgvSSdANyjY8ebqTkRWdUzEngBHkChXfM0lVnow+qwXSYQTRK
jei2XpX8KVaxv3wrp6+FudK0tzYCoCb6JAMRnjje2Kox85MgfiYXAarjTfBkpVoZVX4c5PT9rMNO
1q8Dx2Ugq8sXO8RTGVBp7aF7HfohHikKIFL2FQAZ+qulzBSgbvQfhdh62ofBN4tSmyaCBurks8SD
RpGdxs0AyglgiYmCIBMeOALODVQma2atw6cS0rVvF7Jgd2Jdl2tcm4VmYwo1hBtYfc+Ia9Jam/0L
GmzIYWBt3NJKm49ztX3Tw6IehK5gxmEByup0d4YljqiC0D3m8iklgEgdV8JZI4r5Y8GwCp1Q/W3B
5rwk2sz2n8mS4LJomJNK3niv/E62xyf43fPicw5YpPHk0/yAOTiyvq4w761ga5WYJ6UIsj+YT64r
226+0gOWUfAQU9tbBsXrY2rQuKZrSLAn30LK0GKqxLhdRJH42S3BWT81dnT64ubXjKF1BX5HMcns
IxvSfQ/8BtaGghu9hMvi0ZwDezrHnpdKZETozPjW/TVR9zKHlO0LPb1CioO6nXsu/sgR0ilxuJss
7/Ng6a995hAB4TzyVC3fDCWhRs7J7xP3fyS019lpnP4mKtfCt7obJk2rk4tRTqE/PGnZN+3g7SCt
ML64XwV2C6LmwjUQHc7pkMmT+b99vHkfZO82A9+XgKGHuthoInNgZERwi42VKNAJFh9fMYlBbqXo
4mLXyv7DG8CCFhWa8nb+dWNm1PqXoFNY15hdspHMIPGbsGlRN6He+B3lpZhi96G2g7rREA0z3mbT
dqIqfmy1ujHcWc+DM3QQ0Up0NYeoi1HexFcJAfTHD4XFY786BWwUhfsJY7tZU7jg3EzCIkwQJ2Rw
d3iCNyHKFIY5h9Z3gptSu5vhCIBfzkOIfqlbWg/KYJpkuWa82RLn03X98zUHXieK8VeT+LRvwvM4
Sv52kow6VDY0f8tnpu9l2XlA7lORNGoJt/oAUeRwCCpJ/IqOdTr9sgJTKyj0kDYkeNZJ+KFVhpy5
9roOWsPInHD+Nh/cMA8BSZk7JK3vJgnFsy+kLQh7YuyZg8NV+SnZBiz4YxsB+F0rwcIeNrvQKHmo
FXFDmWBi1jMWxgYvj2+b8lrx5pORNhOShb25a+TJwZvwanha/j028TDnuqTUgosHLtQtVmGPcCxe
+Z5hfca4a9uiHMIrH8GBwFi9R9XUABi64b7iPrF+ojSgNxhQCHIwoV07xcFdrIUK4RUc6sL4+P3p
ItHjPjOmhfWPkJPs49zr7r8/ngOWQzB8/z+gtcEDbW/BwPYAEtUYeKxnPt64fIkT395hf8cEhZgR
rgroDMmDPrmzSA7Jnsyqdn8A3zbr34ggtojWIDMM94ADPCJtZXfKYaXgX516O+LRDFIZ/Lg+rh4l
++eHf1bm8vS5A7V1mpIssj9VgADMYvmUfkzByhdYWqHHQSi2pyqR0EFemy+gV5HKlwsLy9KazuRl
CnIBjUkG5m9ammM2X7LhVooIpTQE0CMMhUc0Yf5u3Kxg0BXmtBW3ZM5Jl1MoK05c54E4qIifdYtK
41UfvychGtnY0Sm9f79OhmjXh1APULQSbfCmqrNMO0pUKPEE6E/hBAcErXpvzfwmePAp/soi4euR
vNQ+NmquJIzdliRGEXnOyzntteUoAPlnmuUC0sNKaB0mRd74M4z0GLzsmcFqNEyqMFY7THw/gL40
iKEujYoHFkb4i0LolYvnE+0jjClnOZtogbQWLZv/F9dKjhyYykCRbQ8iIFHTEw3y4xu9SA8JfKzY
w/t7+3HW0zDMZbXqO9+xEwDyks2Ig5aEC+56Jk9n1q+Xe7fJmYljUnRu7BDZanTf/WE3wqU2IbEP
mo17H756hSv7sNN0rYSsUuk3WAG763gDmHtDXZkZhQcAJT7qGz/Zekbc3vUV43b2m2AU2crEgD1r
r2iNM6XGMGYhxoYOSufthKB9MTWmbhoUfDOBIv8anm0bD5lWTJARXQ+cSXpUYhSqOtdVkksgK/3I
YBm6yQ5nCiM6NUREpn+6zUbb2mmAQf+gUpLQ5sp+Zr21uXTGg0a+WCVMNXTmH5fWi0LFtNmdJupM
Ixhmu1QmtnhRWHgekIjj5gWJap7BTZMi85dGc3pyBIMaFkd0ZBrHlU8HAb3miS0PyTZXY1w/NJMz
khc2/MJsSTUOdHqcWNw+nMgXrzRemWafUm/hYKJgTrMB9vvo499F2UAck7lkVGdebbCc1aIMrUE/
UCi9FldQgT4PDUZJaHPoYru4ATSxmJdWVUGx1oRu15NtTckiTFE8XpzFaHGIaO4ccyNLX/3u/gCH
BWkbRi5xbgWaWL8Z1nTxm9VMd94ntZZ96YQRL+U7KvgSYdCsNg/vM3fqz3yFtCKm7Jh6xhK1U/yq
6ZRlemQmsnTp7egQXK+ikPfLSo9+CobKN/IiT66fLZAOGEjeGWvxWPi78iLlpxs7P3PLcvMGB6MG
PI+XomsqygvigNxygj6QKTrLQrh6/v/7i7VgLhbHAEdUI3k3llUtb3ulzAUwXlB99pAQBekZnVKb
jfiyYrsPVQXgYVGw/NbWIK7Z94VETKZzdjyUsJ87NKRak99BKfWq4Yv2uOe9NPeVEH8UDsFk0UhG
sMLhn18ntau05Uoq6g9kCKwhlXtFZTeCVeGbE9fb6Cp9WfJXOJq9k4Bzs+bB8YTXTVftQasKr6A6
dyf+AGiCeTmBf3I68/bwrzc6x8PVwcZvKsdFATMNL3meR227hWKMr/NiZYlURywB7/g5ZNmuI1m8
K2cMc8b9G+P08jRle0wQQd5xq2SGeGb/LTIC6bsOxuaRzH41ftdPzcWte9nxkfC3kXy6FYQ6gp/G
mnfvckVnRU1HWvG/KzH93NnArvUwx7s06jIoyzTmLfa+Rw/4gIHTLvRsfLH3258RINYKblwGCADK
i51rIjpKh2ee85HcvpOA8L13hR7OEOLp8YP0Z+UVLWPNSOVpmZ1D+grl4Cl/jOHf6B17C5Fssh84
XvkNusC/xxrsy7IbasCjNHFnI1TyKrVooyzko0oTBwn8qd+XBer+56MR8tcvL07BF/7AbbStSkDT
VjtUb33M3Z7vGTpux8cgacBdo2ggLfRyvli7vk68zAgZsDQ6kRgDWL4rX/+exA0fC06qsUKA7pWq
EsvW+6s3Zwd2tEMWyq57XmVbOFHpUFLR2OAZnR7YK4py08IDi/oKOk2RhsUzVAqO9PMLcOc4uX/J
dQkjDRi8srlSB35vlLRRfEJ0XzOGQxn6d8Z1upcGd/KBtWhZKnJ6Tkfv0B9x1OBmaDJhtbtPZgEU
bWKHduuEXh4S7l0XIQolDIzb7Qrm/95j7Vvzs1KtfUdmU25DcAY+uOxTKdgGLJoJmSuziQIBNlKg
m0G4sd31vKBacgrLsLDnro+iuOlcJFlSla+E3FXijVE7XTCIpLyixGKw7iCOXO+BmVzbsS4tbaRF
OZralU/P4mE5iJLdW5l0tb89UnEZX8GwoMvYGFAZgQHedcGp4AFR9hTmFwx04yNeQgtSNR7etKrz
2B5s6nbthHY3h5xmMht3CeL3/+b1e0lMwVKa1aZY47xG0cmvl2EIXCDWWWyxcRRkeJpaL+9GCqgV
/0ZCeJgfDmfGJAegvoJTRNyZdXt0qbaSen25v5TaSlyR8OvZx1XpzWyWzJXHu+g0/qWmFSp4WVc+
IamRDwVNP8dH723wuQv90XMX8gE+J0XXJLGVQQV/wHq1vGdUt5hDgqkgGJU4b4NM2LbzhCA2FR6f
jQKjuxLdYruep7gP9TZKMzdPPB6ef/LbDoyMdZhr/pZt6BWQvNeb8yWPWZ8Eo6hDfrEIY1GfQqlL
ej2EteS7LgOLrti43VvGrzdQ9MvS6fMD4SrMH4sCTSjfZbPlYzA3clkHR7+9HDnJPFAGG5CTYexh
A0ilSkNfeS/+X7MonVRFWZVRkFLKk62KkLt3uLX7mUtSbAQP+wv23m0NHXnqr7fjFMWQJPMnhmZE
clfczZezz5dXwkyBZ8Qc2whgmckdA+xndylukAJqcu14PP+577tcJuZ2yJTqbqSMj/wuwyseufZD
8UJ93I2BNwR0JjQ14WDKpMXCMUIGny2tPD1tJl7WcO9CG1CtesQf0Lge0OLc+Y8zBEq+hk/ob+Oh
WAc0Gk7I5Oo9g/yH55kbwC5yiMiU3K9xEL/ux/sAgilR+S0M+6z3X/XRCzDNiFw4MBxA2dxF8foy
4NOConBmcVxQEGylJwbRXXOe5G8ChZO4m/9v+fyXt1x33vXtmyf16IEYpKwvrAwzcmlxHdZYldcZ
0oGEJWjwGapU1buDdQDCAei35LRqiNFv2cf5LGoEwonYbPEvAa1vv9tEQ9OsNbUYD9SWuLG+36CF
n1bCbdqVjVKizDnX2LoWNQp0zdDQBO3X7fmNXLn6DnTuv8FZLkJNJGZijMPv3Bu0CyLllUwN0uKe
MuZx5zZ9u1uf/RO5GO69171Ix2YSHamuh7iqoOUxkwpjOz+D3g8MQ2H7lTb4X4Up2ydL4tLJVTLC
FPXj7ypUzJPshfVNBYg/6zITmsx7U9vC7G/iz0Isxqahv3p4T+iOubd/E9Kx9JgqJqXS0A9gKXT8
B0EplhakG79RqxKnhSuSkhkU5JFSx15ST1Su48+U1HCv0etEmwPRkzhMxdeTwAIg7ZwOgPhUn3pM
BuV4nv5tvNffxnwDYE7jyWHPdcbXTNCOjFJY4OpVfnMnKFRMIwSi4cyGC39Oha+blIe4FG5ARb0g
vrfgPxssqwwvqY8yzq9z+m2z90itS0ohGqYdiovgGEdO6m+/v2HZjsx7lSjDrvpcHMvgNTJJP4Lw
z1KTi9TdeAai94bphvbWUNb8j3l0aM9vxkjff02t0Ts99jYx9YdT+egTBRFrWH8CUCJ+G14Tatpm
JMqsMskiuLr+lKCB+j5UZE09LXYKBWqS6ZMLFk4Vwf8d63+pCGmUGALC9vDaJTMJFKypsD/tyVKJ
n935NBHzN8aPDiSqnxeCKZRbKDZHWlFCrubk/4J95hMiWeJhINdIrz487Z/NLiidr2vjgUk0N6OI
r3WtI/zn42e6Qnl2T1CgCLWw+WdBg7d9V9sRLAFQfnm1dZU88e0PZFAgj0yPFU6mo+gW4BYfsY52
i/kWYYHCGIoHtzPAxy8iXqFCQnPcqowhKTFQWE+tNdW+x4Ewf8Wdf+FLqBNPB/4smDVAMniLdZR6
Mm7GpDAklaM5IJN8vk/TbXCgpoeJBR8+D4oX9ws7krOfmb6wdldDC9gLJXeUZqete5ae1AlieELK
Wr44Qtnw5qObHx2mdRcAWNAJfTJBuvJEVA2Zz9NRu2KOChIw+1QVslHH2Ea9kTLTkQUF16luT+5a
SeeqoEZIqlrOZ7zczFw+uiHVfh+h0EZkYlZv9fP8s+4Pw0lUgzHhJNKS6mZtflpIY21dxDS4RKRD
5eqUCzcS0d+KrUk9lOdYcvTVIzS3szEMTZPCnablwyTlOXSecWuJGqOvKlmqOFz6ZYKvF/uqVOOa
XweGYyOhmRG/t/AjgImcd6IrZdKTQkc1yc6xdA9Tk8PpI6L5Q9CGDy1UkQZWka4IqYpDKIe4lRdL
8UsNRm0Ux5VjQsy6AoXJ9BIRKp8bqjM+xfAxxB/uhuhRsG8mcJ8D1fvdCxxkYg/rzvQWhcCPlpZ5
VVgxlRTm7lsE+SxbMEHXf9+5QTVHFfmmxVgeWEMRuRpd5rX1QQOeTVMfisLWtHkpJrSsXTHmNcyU
sSliZbybmgqryJxW4RI197KRnSDJKGqD/dJEiASg2Zmhu0MXMMqwiL4C18+K51B7jOgNaLYhbxiU
N4Z8AcmFo7zyi1Cy2k6GvehhkPQO5OLrYteN5ZZJb1ja8n3qxX+U0hKRF6uCnkEqa0b+f+T1SbNc
xlgNlhd49XrvOX+DaC+aLfGFTFTHYf6Q5Jn9Kz99IyyKAVysKDNAeNU2V/K8kOwIjtm1ImQoYBi9
v2enB6fQAQo3FVsFTV98medzOUoPBT3EteCPleeJnbcvdbpaaHk0YamfhedpvGDx2lBJ7nOLE98h
p1c0UjIdOLkZMk1rTc2n1vOHDsn3c/tX7J1p7p7nsYL6lYM7WfMI+Mn+M+wDluHqjUyd1XUqsILO
ETneU5iwCo3bTpoOrG7b3H5lbzLp6pwUn4utCR/WNouS+eosVe2LPCFBpvnAN0IPhLyVCHsoQNdI
j74DqFhFOFkMW6uiSzA5u56n4UJWGPNZqsrUMn78fsOFWQdN3rClZyE7PyFicXVKdIGqGkegbaw7
L+heVGg2don2uh07rbeO1C8oHlXso6VP/sUe14yoe93PvOvkUGGTXBfUEyRRSXIWlCEbV7X6nBm2
y1vXC7OsWpXdGW7/DMBCLxIEaxGB9C68Zy4usxRf+zR7pKeVU5bR7Nc7BC57C2HxOQBjmoOVbgJ3
PHKk00JBTxwzwcRPSEsNfsMoAdt0jF+x3FGIQAqxdi81l6IANc4ROvUONVYVfld/0G1X27WABdL3
2cDjVmXaBgT5b+h8gBLg75g1ZzGCwLovzlqfewPfsA2X6JAqPntIySMe41XkypX0pNHuic6v/t8i
rQjE2yQD/PP9hsQytPiIR96ViiBa9TVcbs0gH0WE5gv99IBQI0st+E0ViDndTRYMNPvTcVHgIwht
8nnYOcf12g4jNLddgQEuSIDThJpaLHhso3qcGoOdnKnpeB4PETSr45N/VAb/ok8TDMnaheLF/zd8
J5YBAwBreSRNkZoYYT0PM20MvQ4UtDC9ebvNFXPF0ge22zh3LVg8ULBpfqB3Q+G1Cgw84OUkobCa
m+WQkYCezwILkCTy7OlRl1IFyUSThGAplQ0lYYTGczr3ySvDkwxYGqGfKgTkbXZYGPloIxSXTOq8
fPtBRfODq8U2XOhAxr2XWOxg1JbieCwUyMi/YtLbSJbSEHYaoZh/jrCC+boyUvJ37hJV5/OCKaM0
OfT2H6JJD3k8GLWBFHShchvKFWJGPZpGGC/8Gn+WuVEuztxMYVAoMdlm/uuQ2wM4cTGdxjZkYlY4
F5QxNUGQB3F2Bnx3TKhQ4FVJvHs6Fq0EC3BnGeD6swWLrrjHcdLzFZSEeaExK3q+LZToH72cCq/Q
rawAsmD7R+k75gF4bl0/eoz/o9nT38iGmd01QOZBEITtSPedW08WLOQc1Pev3W1UZKVfEjoxdR4a
xHdKHN6m6yHuXJWG6Q1Sa2F+97eVttyMAvSShTHli4CnxocGP+q/ogZCPBfRbsq/Lw/qGoy11t3U
qkIHnc52EoICrS/vl6WCU06WkDnWD+vQqGhPt6m483fy8u0ch41qHHnr253jiqpc8PpnMLLtoCwP
Ohm8/9iL5MDLZfKC848mOM4JjSbfU7Uc8m8cRHJyr8fQia+jI9e+hM08Ek86l36UseTTRrJrnzOH
zZ+S+r1X8DnMLbHoFczsO5dZShcQGsfaXYYn5rjt6VgmDuzsfSzsAUYF93fcd2mbM08RPgKZPzRk
z739Cbp7s3rMgZMrIgoJEEjUZPeItmoAkBD/v3ygrYmBwSHli/JNEuNFRdQKvNTHQfzMcQZuvZ7i
Gtb3PhtPRDgHMAdon+tdmFv69Fib79hsINuAQHJwK+rRZRGxKkfghpauqnMrMNJNK5poRVkc1b5h
d0UKVfTotI0at39deMwJNqwCE9g0XTHuVU/MdrBm/L80zDMxuSrBT2Jye9ukThZoQs66PFtffhyk
tq+d+cfUshgasF/96j/WM0nq1VPlctgujkuZwTzkJpKne4Y3g88Tz+BxooCcV2v/eTJMiwyswW41
NVZ7Ws/ZwPmWqu++wHatmZHYVfhLOlgzNWH0CukHfv0D07/G8MMugjB5zL9YnshHNSYO8dVXd7D1
qaFsUUScXTJlLjDqPW05WToyjDJH7B0ObXBT1oMcvmDGrDUnK6S6CmztMdYwIAFKDcA0azN63oH1
s5a61d66o/fuEQwQgAu2FPxg9Kjz/jThJ/AtSm7lt798dEdFvq/0g6V+i2at++pB1mLxoqH8+ooQ
f4EEC1fUFOZw3Hck28RopoEkj5DroGbsfwAwuW7GrmUJ/Oi8xZvA8s7MsG87lU6jyse/XK3EDxsS
awYoN+rOupiawpd7g0iHSfgQVg8uHH5CG7UBRF9hMZiDdVKso4TJrUOEtn+cwJfnBhP+aMB0obb7
J+V1Z5EGtrWQS8umy3+Xb/VN2HwxyoNh3AYE6Gpzu2vNU83dtj8QP8Hv3RtW+k5IKV7oxgKh+rPk
/lP+U6HCfuM87yAxqz8sLwKGAOSmUpwTzz3dFNQSCv+X0OacI329qkQJkZk3rRgmPldrHEHXJVOX
5XMFqW8pA6WNbJlk6ooir9yhRxtxofH0Gwnuyy3v65pW7xWZNGSD19eS+EQWCXq1rnHO5HIwQFmr
9HvXIxyOSN9IUStTF9fN1II8xKgPHRZdm3fCVW96DUHJuBdubu5FziXe7jVK1oL9GuBFRDxU3KXd
i2PTXcW3LXWyByRRutt6w+on2cIyHH7isaXPXqBYf45e5ahUx32xZO7hu/7Khcm92vVdrofL2JQs
Ha6U/0kzM8MA453hLCu5Er1WdHqY8aoR5ueUkufdX3cHmhr8Iv8UIcMCrcrwml3tT4xmhhLA1PEg
YKf+tNaUx2yRxcWisutaJay/q/KFVDEWwpD8/8Rfn+Vgvi85TytTmeRFHIn0TIKLBfxvAbuNn7aE
W4ETWYJ+3RLxFXZsW+lpV8o2S+gvZ/dY3sPkl4sDomOhY2PWgvuF9SJAwsQsTwlaQoYZieBZ742e
xw+98Ond6tngLE3GbAqEF6D80A5WDzrXw6foX9y7plqaJiaYjizJkoz4JxkFtp9nrdq4/lk5lutL
jnyumhcXnjpKcJrtbAHY1kEUQbZ28vgxLltYEPlvnbDlKQebusqb32k8kWuFd96lS3trDjWKMO4a
qbp/SxUN2fmTLNSo89IdC2ZAs3z5/aRH9ruYL/YKTLKIIfi74Y+lE4OlLgKGFxJlDlKnomq3lxUj
f8xvRee2pfCJ/WHLzjhH9oL0aKtRI7SVY9ywP6p49SfIIPtJc/lZu/CcvAV+HjDslPQDyhKdSVwC
+TRGsJjlDrBb0IoB2AQQOJ/+1BpmjwjrpIIXdVtJzN7CQgW8//tNWdBvRSARCWk5NfJtwNxawLfq
fX3F94Pu0kuCk+xLGJVlbK/dunTO2/aURfDG85WKODeCnwel8OHoExp+uMH3ae4ZOFPmhB8Krd3l
e8d3AhHZr9Xu2AdprVIOWRl23D7deLd/HFfPgZ+LymY5eWAwjpYNP3GIIAjaJ8YZCetE0tXs1cfR
D8r7m3fN38spTv4CFtCpYf0QS5iNEmcaoAt5x5mSXsdD5UQf+gji2zx85OFoHEVkrDR/5tuplOgl
ti82dCSrsD+8UAIF6qoAPzyZwx0irnAsS5vKj9tsQq52GBlrbkJIrkTFIKQDJ4h+lpWLkDblV9wG
Ro3ZTtGZ6cjsDkNGDYWb6nM5aqhC2Y8e4QD3yj8BMOQo7khjCgMo30clxV4t8hbPsGYgzSgKkW1p
thJVmm8Q4GCfbY3oOH1OneR5cmheDnm6mjI3sTLaVduksIrAmR9YoYSRRJIjn4O3Oo9YYgTzJDNc
VOLRkvDQ3tVAr47LlZwPK36GFgrBXGhgBnQOymrMFFG+R0jv32Dtc5XJWMKLDunHIoqnBCA5jzod
3sWEBLkhDOjuADFkVns41N97eizGG8Sq8SJH+rdkqqK6Fc1v8vz/0vN3hlf/jsh1atnu5iHNf/EA
GeKYVCElcdIDa7wPMYjtntuIjrVJb8wuAyqznP1HG2lZIFrfz8WgK41wcgnIwQVGnFsntNHCWsHx
wtIfps6q5AcUkTX0Y6il7p+7fK/OIg+8Py8JImeF2GTj4M24aVlT0GDcLmkcZo61Q3l2kprrKLea
AtLX+Dha3Hkapl21Rwn9mFdSKyEKpXbBe06Tmek3oNW19QagCI6HNCzllySfbQkp/QZ6QGcae8OH
S/QZUpAxIHNnBzofcpYYfVcMhkCxmgdeivo3TnoKgB8GG0TsrMElsDcs52ckLDy9qseeYGr7jQjS
Jvy8PXvkGbieLinDQtbd5FtQfhTtdT6skZsTelBSA4ZVMHaEN2ec6j37YayfF/3kb97RJKsKJjaq
7tmFVQGQdIseUZH3dPP5eT6JOy6lpS7F1hJ64gsBEYLzkxEdM/+xWhMc/qQF45z5KF+1YTEmxHTB
/ZgQojhQ9HPJUNUs+NJImUil3QeKqcOcxyF6kMTYueeKJrzlnqABJTP2YcJ8gz3yQyykwBziNllH
1HLASaCbL+8bOKXhROdfH7DICnXRcV+OIER5UBFoTYifitQZYJt8eOWmxy9AjT3rE2BU1qMaBt19
++UpirZl7F1T0wCU6HFkCsTenjnu17kg+3ZDTeduF3VkCXwh036FjC0aV0kFrRnQFGFakq0XvBrb
cVm7cEKYDdt5eH93lXGmYTNmENNRDKKbMlM2fz1KFHB9mZ9BqLIl/gSD/tWCN1GnbccV7koeNzwQ
ttr4jId1Hb/ktxmU+4GIrcI7Es2Iu490plsnA0wpD0Xi44NTYJ9iAB65j0P7qKyzM0B0NisPYTY3
uPIbn+sFCblyhdePXRWnHgpQo9lZfJ2V/VIG6yiEuvyy2QbDB/x9QbuiiBGjbX6hAs4ez0mm+7XK
vtgFxWhaVHra+AFzQEm16Ln3y3KNdEyo4btcE0+T8axpk5WThXc2eYWSPrU+zFqGbG4FLEr9a6wx
GiwAYrCKTiXP1SFCycX6FHy7T40TRGz6TvImOEU38nBxT9dyyyjuhhcZlIdZlASs0Mc9dDFEO4pS
nVp/pDW2bFzmDKcizG+qQdeH+n4yV6bX4FPUXOGq8AL2dat5nUNcSWNlJyP+stu3dNWCs3v+5gwz
T+kVnus11ydojzNdv4Sg/WzNeRBM6Age40CqruzdZBzIxVZx4PZv8kmoe6O2FXg07QJq3+jIxLka
1FhVQwB4/kRT+HnauqaSI35K0zXsFzozKx09gSj1EFmErv+k9lOzJKJUuUT13VinQe92k4EvRi6k
fIBW5Os7+IUWDqswbOAI+efNjxhOCA9Hm5HF1ymNkqNOHQpVq//WM1jj7KrYL1o83ZtP8w86A6xX
x1GT6LutNyHB4artQk6omJWfPKi9/x/L08vxVXCizUq7Cjor3W9A64OihftrJlmxaZv8X+czjtnU
x8O/yLOUHVO+BGaeicJCFSWobdTdg/KkyhiOA0Rbwmgmz3XYUpXTGu3Y7n9J5B13aj1pdpgU52zd
sg4rznS/3oW3cFw8z0csZn2kQF+9bsKSjD/ROqxJCIIAsrFwD8sKpV0kGQ66+ojc7Wqo/ZRQbC3o
ga3IMxa+/HYmS9/v9XoI9GAFNJm1vfCRudKzdc3nfkmWjlFSBXe/nam74RgjDgM4K0naMLZJFPD1
mikTza1EWbmDWav/wipsn9Zd6Jv9uM6DITLt3ebNfjUGTZL+RuPzLOEJS/dw+jDFcbnDlUOcV+Bs
10yyfskM8gvyzpNqXVgErkhcZxXO8s12czt+LrDsCHIdAa/+9Ouy1jHLKgvC7AieYG4SabbX8tFd
9eJl0kCvqunmRdWg60kRULQih910gXsMFqlDijxGJ7XUTIBRNlAx9R8gbq1d5sp4N4dPumMQN6UC
fsr12bd3YR0t5irb9cfAHgrtIUtTjIv6nzVQ9oMIvQ93H+OxQQ6fyQlnj6h0xhMQlWJK/Zm1CjKK
7XaPLVJWXCO+McERwLf2zDVAqgeySLCSDvuEQoAWDLmFz3WQf1ZPgOD57Mb2h/RDKvhYcDFQpRmv
CJxDeiAaBrTc8WV5P3fqSCZarrXBY4czL0l4yfJWFfsIM3JQqTrZN5zDvy7WIKO9iD/IewiKvXNP
NaekqRm6seIGbIo2/nx4BcEV+h6TKptkyWaAnLI103fzReny+0NgfikXh9s/T65MzBkHvexW93c2
QEzGHyUKj6D8Fu2jwgCu94u/T84yy1+dLHQVwRV21lZ3UiIQ8nSSQYIqsmzNTFulRo8XwYgnsFmM
1oQQVdfPUdf9NoTBVl+lrgYinlp+zLEUIPOIj954mSOFaWuWLIZBM5enn5j0A9t9+X6/ohKGUCBN
Hkk/Zt3RpnjH6J8pPRBgbVWbbJgVnRvxOSLJbrvSsy8FA+ojFTQgOQMD9cy/9TCD+VwXTdFOGgS/
ueGJeWr0hiBsUICzxcNNDrWEAPpOVwsYBAIJCZ7OfPuaA/JivAkzfq3UaTJp/Rl2rW3loYTgvkzG
ISYAh091PE9vziAEiGdDZQw3b+092YgaTun80RMpfstRNxcHPgmHhVzqhvirdskE4G+0xrOcMPts
qmkTXiBXPF00rZsEssaIcZnzmus/wF0IsDIDfkZBXgBtMTPOV8Nfi58vWpj1Bi7VIBFaqTTvouDQ
0YQ15vuAuSN4YLXiaMs5dcS1lNUT3sU3QqussJV4nThT//7TUYeFs58O2HF/lD1uSJpRDxJoyNW1
an01uTIyifXdRKOHuBH/VzOiBCcsuuc3un/u1HmaqierYpFWg5Q/YVYeb3HGsHVYXDh1iJQ9Mclt
t2prX4ItxZO7TRvp0YCzInlOXmXwkVd4qczK8Lh5KxIax3+Cod3g1JsJpKC2QQnnt8vNYw9E9v+L
GCJ3Qdttl9sd2IXTRBfRDMn6Cc3X/VOIjoPhs8WHy8br306hNEPmM04dEpVT2KodOPEwxpHGIftC
/SA+625LBGkKEfOFLJLpLHZ4m0DChFxCJcEWHyjxLrZ8jQJMm/kSN0qMEzPYbqGVZMifl5cfy/wt
mbtthieFQItEN/MeUD+DyUJARpdFeSnYNwrQneX1c34py/8sBb6uyd73XZFwbdOivRFPDpWPskKw
tith1q4X9f/hRoIqaxQy70KYA57/CJGOEA84fJW2DxTJYnOE/e0M9I7en+p7qrxLvwO9Msg0uprE
0Ms/tOOXE4SE8BAf7s0PeC8+2UeaEpZdb09wKoTkBbBhILjqzNl6FGtidm26FJ+bAJRjChS4r3U/
PF5KCl+2wk2mo4M0/O/n0f3T+8bWBUDGORQCaVk9megtJqzdNBvTKnxYs+3UX2xZc92yogGm1zRY
2yTJ4PXSso06EcFXFxR5faGSRj9HjmI35319K5cjkMuop32B+obMTRXgM1X0Hv2HrGJX4ByGA504
wL7Q+fmgPhBpP6gzeNaPEVEtEAGC//aJ0ZhcU5zyF98llP3UQJdxAyzX1P3LoySh/P7Y431uQuob
lgiQ934pnWRu0ea3rSxNxINNKenGVq/+KvsRaF3HSeAmIM2tuyewZiT/jYNqJ1gaTuQiM0OpDogx
tjb2q+anlU8QnxhMX2RnAI16EXqqNEDKtkT4BVJeUQFC5ToSoQHDZxLjNSKKVSKIaGlaJMl34WLl
QNCKVEdg2Ouf3MJq8/ZqMhqJa8T9cq7lXQEvR7VdeVFICnwOnwmPiImohDYashF3LrBukM6b+LjU
Sap7j+5L3rpxolcZ6kcd3Sx6X5+NwMSevAgI5W7UDVW3ixfzmw3drxZrA247rkv0mOEWieEM27q/
wQsIoQYsmKSJMyax6wFURX1imvcSOn6VhWMwbbv4Z5qg3H3DiLHB9QB/oLLwAbnYizmZCKYjx+FV
cJntYCIEI/w06FfU7q5qQWWum+ZN+g+O+PxcxpQMLn9FFAnX8w6PqLX5aqIfUQKOKVh6ZbgflNbf
7WroZGngFqeAB2FMPKA78gQmhBemZ48bVclujX/ICVebKX2JUoOTQNnnxVF+2osKrsbhcTRruYe4
tvKy/dGulG0qiKqfeyBtuyOyYgFUvohV4jzvH8Adsv1W/nxf2DGQVqGR4qxeXXdWoBLoKGqUTTLt
/GiC3GsRK58DN1rkjaHaM8QgrXNZLSLrzg2XmmiDPG3fnvNwju6mORZ31BlgHUCF7HboDJvmxDN4
6yYrK1T7xGn3TRJR6YZzmNKUt4WWdNGlQecYdcPaQUPw+9IZkezbRGB6qTg5acXRrzE57vz320MW
5f6EOxx1SMXqbEJqxIbamWw8dDJrNJ3MieYLTkGk8E4BUX5636ttSn4xqPyeLxsvKZXtuEtb/o9M
j77/6IAQXCeth0ejhVCnQZZBp8r5kNUQ/JxYTSzaOCqvB7CqB7zSQhUe6vxk/PyD+C09WjPIq5iO
P3q1X+tN9NDww9TYJBFYopiaO0Mn+RlQjUJAXRQw8oJuKeUXVxIZ0M1wT9J4UBmGzWjmsQW4Oh5l
kDMRKnY9/41wrfONAycqJXHcWx2CIFvC65fgNC+tHGtvuIIhLee6LcUVLDGBJQ8uxnsPxor1aI0a
aI0zWgB5t3K17njboe9Tw2uIHizrH046WhqMpoeB2l4eca1tUL7YfaekbKCjBIuMvlXf8WX/a0Jb
sls6ky9HGP3RG7EQFZRtj+o0Z1lUcEeoJNV3zTRvOdT2aOm7rE6Htc1+f713Mv1frlYvv8R/1nec
s+Q5DM/8wltdEYY5nJqb7FF0/NwzelmQTUoeWjd30quv60jM+MJwYrvHOwBxX1zARuifmAVi36t7
sbRX86FsVIKcNuitM8sSdpz0D+CKxo7Tb6gvelqD8m5Io3yt39zf2iJDsB8flh8NiTn5ui//9q+7
oBg5MuPivINHiFM8LWZBleMlkWs2NtZ5GvB0rZqOWyl1c3PvHzriCM7/QR5/OPImjTjvWm4aOEPh
2aiwavGptmtvNJp8CmHmNx8v0CbOY/cJadVQwEcmAnFku+798IMj6y1O4OkvBttV7Cn2ZOoXeAs2
lpkJWZ8RFZzp3p0t+ayznnvPEGvgDgl+QVeB1abr/8LAwpz2dzx6cdRshlSt9YI2I4a2fECeyeOC
0ZTaRAsmgtK6VtvKYXu6xsjBZbaMlV7i4i0BdmF/fQo8gUgcuh96HIF8gP4bXd9fb2sr+M+RuAYX
3yJtMdEUAO5b4vBizTaiv3SwGcrkzAtBH2NeCBIdYhez8fbsK7/dKYU6QcMw3Kdhdo9Eldor8iM4
pj2EUi7CewktRHLDck9f9C6u5wdrkTD0Y3kImXFrcrLykG9IiLWSxqE3irKEnv8uAIyNJuX1fMJJ
uvZUjH/ZZlzcUHu99RkBpaTMpnGGh5JoL4Eg2d4x6RlgBxzIx/e6hg2F365sDau7lE5zVG9mNSCQ
p5+RC9It7f9QnQUSwltWcuJ2HHj4juvfLtDnMcjvG/TTknASwjtf00sAKteqIFNm54PFhi3AbRGy
31mn2EtrJEXsYJhe2zao37a1n5wO+X7v+vPQ2kZEqRY5t6BnnhiZO+AeYZyrg+E/nEGDbb3mm76y
EK7EeEAh8Jsb3ajbb918XJBQi6yOCJ9SJTik6IOLcIRSI1CRRyb6QWezwpYqG/1QyvV5d8B7pkWx
pGo4tHFqcEESLJiILdolIb+1nuUacTRc7cLSIMJylyS1GMf69mNhL2vXlWvpCslbAO1CMO8p7jAs
fom6eZoTXFQgwu/dYil2P+jJd38WTU0YJQCkCWwhpMQx9AhYCfsoKylca/P45ybkA1QWFZMRTatf
9liluotbM/7xYvHGRtRONbTulTRX91FZWp8+I5PeLP9Dz2jltSN9olUa3My0iZ43sE6Se0Nz8DgK
gLwuXpXWZDPZF5KSh1TdOjjemgwrA4W+VFocwDA3om6ObliNOVyDTJByxRj2yEKhevISKQ1mim28
rraW3aIdVgVprlYyyexYsxd1maJZyvlsm7mzkHz1Fgwcwg2DlK/FcmURtzXjAjojEbKix28FPF1h
o3u8N1cmaCigj1fyw0JSttAd0vnS1RNQxWSZJB8cpam3ITjAyG2LwiH4Z4KOPyCktyV3pGYMcQbn
lvjKwo3JzJpTNlaSGO/3noUxIlAdXntEaMxQHtXEfzLQim+x5baUXdUqQSydFDsnS4vvwRPSOrPK
w4f+lDMprJlWsfzM4cG+MdapervTaJkM4p5vUljfTVyymMSnJjjFSL+I4C9ILRbxYUlqVd1/YTVv
nQM1K/v+CS+Q8t3Qkbl2PmbS370LC3GkNC2M6Nj9fHA9jztRBnqkiW7nX4YZaVBn8g5HaHjB7Zis
6LcriXjRRPQSkeUjq+/ly/QAOv582G96c6jh5B3IVjcZ6Zl6rQ1hKAdniX+BCgKhVKtSSZLAuhWB
DNHTRZJN7fnqy3ApAhS/dNcStX/3WMLa0h49GN0jPd8GPJv4t8v6JcwnZAAWy2RvhyqRtPQJqh96
Gllkqoe7vCggKs8AHJYxxx22abpYvqCrEVoij74v4frFtLsn8/G1QFryru5bLUGWml8zOO8YgksX
gi739EzD9Rlfc/3iIzM7SKlPhrqzoa1qz6nm8WgRU4f8yVM5rThEJVrwdyAmD5P8EpYGe2JQwAxQ
3TbygLavWRpcFdd85QWkDW3VEEXj1kIUu2Z5kHq49mY15QnGsc6rUErHsyG51OOOuFERL2p43Epd
fV1LWGyQHy5St/5pB84IwVSK7tZN7VuZOZ3KW/zgEx0pmsC/munzTsbnojSX0XCzrCTgNfZfpEcJ
AgV1fCqccB258BHoqjvF94akdeNpriK2x7uGg88xzts7MWmLkS4src+5PppYB9XCAKPOuFqFFl0R
LrI/NBJo0J6Hc7Q3m0QM6b+H+eKwEhogwGKDA8NyTvJJ0UU8PaYZ7+N7J09Jzq9mfDAeeYFE//lV
ho+roF7V7JDTuXAyb1NT4AK+jVNjn8kmRl16P8gngNhSaMMZaJFOLluD6lGd8MJ64h3o35JTgovK
/FS6KXKbgVS1k3jY22yGk6to6SjAU8ZQ5uQ9XD8Bnz6PtjTd6CEs5mj3aebqVjvvFbWe0ARXcVR4
06ETgBGstv8D30XcyWCKCTkM+Dvea7NWbLBJhhm0gEorWqQORcjzugH99KVkW8lIr85qkxQ15p1r
mBE9D241zF7xswc4iH27bHqOGbQF3qnpGBN2gs9OmBm6ZMgFdMrbCvkE/HeWtYH1R/o1Q83PtQM+
liH8wFQz0Xpnc2xMiwicI1FllOOE+mfsKxmV0EAROxfMhU9nm9JJYO/C7UxsUkHmr6lBLOhIK+7i
cKQWaLwKajTCr3Prkd6FgKHdUnb+534WMLyxm87fg/qwHzNK9qtk2HBtCZH28Gfb7B9Abq7AOcxp
jBmGLpSbZrZJfa0nZ0kr4K6I/JFUTrqR4CeOqSnRvNVsTWMkej8+qDS7F/5t3yU+GcawJtHanVY7
5MdMOzdyE4ECgjUPMSqBV9PxgAq7cHvH5ly03Ovabkd81/brzIGUxuICNdR50+Mk8JNcmaIgm8eP
to81IP3kWqEKZS13Lf9gf38G5gK9wyniC3/rnIDV+qcLEkvXaVn23ix/dvYEW/WdSkQCncfAFB7S
AsLt0Ck1BrEvtlpRDsH1Pj+MCBnumof1N1CA4CLpCV/pjQwH9EfdcQZRCuyLzcuUydELTPQA81Lj
Lwgp0phptDoXaFxkgWc2+uycS0iXw9OTKWttWJqu6riXrUWf7DcqKkhlBGCWVESDE6Y/VZQDdZ8m
pNP+2PdfABuUisOifsT2TQYr+bzzUyvEO4oT87vTTwie8RRRZ4qYHD434wt3aAu3NDu9AmtXHjO7
GWnyuuPCj/fWrc6aNtljjmJOS1sDVjs0b2m0StiG0P63hTh/DAnxQ/M9ryRMxlD1VkIu+Sb4o4PO
hwmAuflkZN9Mdgazf64V+ZsjxkXY/BYlomrkiH8wAJtoRzYC9BAixobGswGAQKvJpMhND4gJ2Iwi
/cqulHpikotAU6W/zmH35Ag8fPyOUmBFPQDI38Gd/g5ekb6GlIhqeQ1sInrQQ6cz2GCk3tsphKoY
hQFGi5E+wdH8JK31ZagJgNiZI3rkSX8l5F2PovP+CJBl5JCp/IjG+e2UanWjKZbSt9BXsT9qYW40
ILkCGIxR44k7z2KNSytJd+WKF0rmVjTjwEcd4B43SAnkhZMRjv39mq88cxEqwBZExGTMHEzV3EA4
VPLTf1kftWcFIMWdaGzeWGnVMC/CzablPf6NmTltdSqUyQw1P7grKZOZRDY9EEI2IFx9jFQLfKMr
U8kUJ20XcJctoaGFH64sPRM+Tuyw8ktzn7OpNpIIyyn5ItrG/KZwYuwvaH5F5aCoEqzAfiiMT4hW
DlF+gE0CancTmZRDWNqY4mxjtTZvjdIvHb6T+jvAKXrtlU5sCcZ/T6RHxYIK4PIHo87J8WKZtsW8
cVGj02yTB7yEEIEynyDfS7m4cu7YQoNcbyPTWTuAf1DGrRDMZx4kWhUkDiLQBVMwuCd1+mwN67lP
rYBwSqEXMiukSTopQHSg1H+cWi/Bv2k2zrCnIwM5UZcuH0TPt+wR4vmeB/JNtw1/PSPrurL6eUgG
pW1oM3F8UW9shUeSuPIDabRrwNixcyG6wm5/RkGA5oCQfGls3iTkKuXzop9TYApmYSjX/jORgsuC
pEka+HCWxZccW0soa7lTq79QPuun/PYSllna6MOTDh+26i8zXaT+vdBxJklx/+p+VeFkM2kAItPs
aaviIw1XdCzV95EFUV8OksunQKMA7ZqkySgMf3mEut1+Kgq0MHY3a3x8hO9V9CW38qWCR1wgQM8k
idXJsnvjKX/tzQHjVYnLLer+euQFDmNMYlmoak37vok+I/Dgnll/yjL9q+96Jh7Br72i+TNv+DUr
/IQqpa/lSihEADfQQyUABLifJHUqU4cqXMOhVC7yDNnxgUTkvbw0V8FF6skS04REVfJKbaeyTxgS
iiiL3WRVHx3P94mrH4cedUTzy+vOQXCc7y6//FtSLP8EXDD++UUNr3IWveXADK77KDzwUA2AMWsp
759TMZ3c1gIoMLX2W88GXB6aK3QGpchlFwC6FwW1NxmyF7jF6ixP8aMdRhhkXc+608f9mBeyC+UY
1Ro8pSpDo6VGGAgY47oOd49uzpald0ortNUreAKk5efNnmr05nYqjAMJxEsQgmVkiRoDFfh7b0TK
buqxioa1/vPNRwVTONPq8b3LlP/bg3Hnv5rBKlxDLgb1dIq1XyvhNRvjmi96V/0VHq2lG3gKnjBf
8khq3wYim1vlsOZEb+o6KhyLnFi+Rw06g2ZOhQ3+ifNEuEGw9haJvLdpN0vXtb70fYJhychBLry1
lM/GhU4ggV5rZv3smWbtkB5TZiNCdhVsi9gh3Uyk8BahNKLr8dK/b+CuD2M3VCxZzIc5VFiALngA
ZG0e8DZmFDLQvaJpQfbsxstCZ9DYNMg55AvyxH2X7NG2XmC79wr693zf8N4jP2KXcM/hMF+NrjEo
l86it6mP8RRJqFFQ4QtycYPSaQkDW3Vsp7TR9vKMOmfTF1vZ7L/xcjdC1nC0MR29aasNubrWKMwr
xulAdiNmOFIumUTIbM1AkfnejdtfmtjB90j/b9aJBftvB1a/yCmlXyYkvdAgI/Rk2sxfLu4vBszW
3XyXh0MEQjleq7Hs/U0Vj5mXPJrHcra2VvWEkJ2NqdlCWHJzNWwS6EkHLiHAOHb12/dMN2zNkzbx
YFfWE75Alg+KU/BLedKy1CXXt4ZadGfis/KEvztrfHZYkorIWYL6fsHu3X0gwqtHkcaeNUK59EgC
eWKE/MmmXh0l8Hqm7RH4NcGPud7KWy4hiXMVDccaq501TQDxn2qHe1n112Tx+0nNYVscCjxcOb6e
mc2nBGd8srKjsgswEQTSPccWXEuambpOBvn0XR04FIv6bjBiYzWk9Q+0XX5p4jONei+V5XaNsPFZ
jQuts4B94gBQg4RUW2XDpGBqg1atil113S1UHinvud9cutYblF7DsfvPzqoYMCmejd2KqSSg+Dak
7QQRYtZqpJS2KYYjkPZSX0x6/wl6hkHadIL1madl18k3N6JP7IrK/TbEDRVeyJQBvkoFEpoC91iX
wIa8F+siqakOfF/lsPlUDNvelocyhghNZTmZqDXGJi9Qch/x2n+udygk3982MxkJHyF7K9jpYyb+
HKnJsbUnNNU35ihwR+li6wyu+Q58F5hf4DyNzuSc8yUn1pCQh0LDCScHydD0etAwOvumVkeadVVg
zNhQVJXMszQiMBkbKsCjKIeKciZqI7FoFVi1VNvBF9Bx7L7Y2/Jsxzlg6QO+9eEL6hmhMFXVBGaV
tVGgwpWvLWn32KcjpQ2P92EtBQyvexAntQNtiQZ3RRbwcrl4GqUk9KKuAJSY3zLqcV+SuE+w5u2w
wbYBV6Q5TRvaN6zfF0/x6T5uQv1SuG09UeWlRkojXNZos5MKC/kF1+Rb97wgbfr7+CwXWDTSvvlb
yc/gqb59pPweBsTMyNqzim7MnGVjxQyKv45Ja278SnRjc1+6oJzZGzfVHwmFWATvZIDpLq89q/4A
mF4WjHTj5jnObqqLzMy3cHo2xjbqS64AabKGvIWhUVCeLl/NFhK/UFnRIu6/Unps5CWwovrtIj2r
6DAIXHUH1SAAWiyPyt8Tca41+M8ivbplENRAb0sXAFQZk8oaLD1aZbirXowGCNucRWi+dlCqYHSI
OGFgAgR5M+6kwcr7hD9Qy+kL38vI6lIXj8yVLe+wg/gldbyuo+dWVgXHHoBB/vI7j5pocEc4RLDr
sflsHjNLyVcP6ErsAVxFzJIsefGUxvTqoXZESqtnZ6NVpUXcK7rNqwGT1UAkiGWFiUpVHcJAs8vq
O5+zf7IUJUBekrOGWkuGhJzlwj0/h0/GMQml95zF/KXQ1lNdGZFtkVTasOdnui8EgYm0BSNQxXqh
fZynQ/Y+2eNAVq63CtG87exHiB5dRDvmGsRYQpjtVcHjp2HaZG4enN7rYO34RM79WICVIB2MYXzM
4+hmjESULX/U+Mi1b5/EekhAQqc21MYncGDvccyUroUUo7h1ViE+IgJ/M67/YQ2kLd1gGbuk1kM0
Uu+LpFvbG+QnhhrMLV3JcN0ScGHZzuYpgH4n86avgECy1QqYoodtiD+NuHBhDtiV6AXs3P5weE1A
dngUpLqrysKygYhQxpkCfFBsa4sr3ZNeHHDVdRjdAJbNS8se4dcJOWlqyt8PfLryfstOijMF/HE0
zd+3jGM8jJEU/TKbQfatFEA0Ue3We+bYsEyz8fJZIGnf6Vt9xiwuhk4m3xVP31617eLNmjP/ZRa/
w7/7JxMC+avpqFIM/AjIyc4o4AbNK1xQdhVrgDDj4NlLT2qWmvxNzd+sw2YkzoSVljPVIks+55Y0
Jyn9onP5RS52kPXbYpU1MtdXGX0f2cT9cV1Qffc4DCBwNhR4ndoMr3kDJCqxpuY4bV8H442yxRRR
/Sc6LnK+1V62WyvSSuNTTnTideB1x/c/3Z9IZCZcPDA9yDIYBv2Zx7ToTXj1LPcMyEEq3PbG+oMf
UMCWeSZt49WvjoaJHTEU0RGtC06QvgyvoFEA3++R7YZgl7xs6nugqKrPDYNHAAPMfESxMyZdNAiN
SnXk3TaQRHL/yl9XcXgBQH5GKRB+9LIgyemctKL1mgUxoxlWvvn2L58ECP87avuW63j6R38pr1da
QCVa8Qt5+PpCq/rmJWJO3OX6sUwtvrso5E3HYpZtnIAwQMEnK2R7asx6Q/3Ie8/wx2nXrE3CHX1P
zsAFEGsiIRLHre5V03ugeghR5jMPDQckB6Zws4PkxAFEkJPCQK8Ek+M+42F/AGp/JCZdZGPfUoPp
sKEkYF8tJ4HUoF/TEMzIY2gLU4vLiab00PjaEDIjmJmpxJ9Ga6fLISdpQHl6DVErO/iZypxHDS2/
hi86+iLCroNNtmbC6wCG2/xY3pcaqn4c4SMXBpAA8MZHIjlzxa9p6gxoObDdPP4Zb7RAnM7uEcPd
fcOjOn/DohGI0KF8hsDFgL0aqCJN9RbaI4J4fOH86glYOzXiT6Z+9sp5eQhjXsyfhjZvsoZaCR3P
wyOmS05b05YLzuEi7dVn1PlZ52gkeDlqASMDgqj6C3pVQR+eVCHc4xmyA5DMbYbUqsPIaY5OZWOg
JchBrUcam0udLeqg2haEC6OqDk+dzyCw8XC5OMM1CcW3j4FDNEu6J5f/wTaHv/JBG0UUkPgo8bee
4vSpYliRrYUVDhIBOt8MhyYJ7OzoMxLHFPrKFvx0/7J6BCAyvbWrC9LLI11DXbEXz3WEuixmFMtv
4/qJsqKKlgseXZ4AFFW3XooZc/ZxzRjoo8MJmc2Jq6ol+wep0N7y0mr3ED3lc7j0a2fs3mO1STyS
wGVGU5pDsCBzdm0ciZF0IZZ+hdLXhy6DryJJq/RyCnNvN0tg5rgGguTgSeK1UE+23TXiNksH80Xa
57tCFUkCYK8t+NrQwK9tmM1dX/VcSudhmGj97Th3sL1olITP1mF7X/VDPSBwx+CoPNNufiHG4re9
ZS7tlyYMawwQt2MYb56wQUo9vdRlKCf2NFndBWWvd3SPozfaBqz9QkdFJCm7hqoiHZNyxrxi9o1p
fYMtklO2a4UqVXL28HizyQKdyNKlMvWkNg7wnfe2zmFpTOfQ8+DpOwierEUqqnZZTb22uAbf1jA0
pSvKZwqXKqeKACqH6YjEyiR9hMIqBrroyE5HdmAmb5T0vvf58Kdot2+wIAS9jOnVnbV9cXWxh+Bj
qOF0o77aqyL6i+Z2FxM+ij4Plfd/wsGUoDW17YDSoDDEn2KaWSErP0vQQyPWfkFmnLLagrqG3vBc
pWaR0x5P8ZFArhPiqgDeryjaXBxakwptxDwIJ3CuOT5IdJrrXYH6PQgBP9jPH097qHrL8YXp9QQw
7GMLMv9eP7MT8w5wJ4wBL9NJ8xjvKc4VWMJBzqp2BK5ZZN/B2vU0o+2rCwC8b1E+r3vkylnJ0UfP
G2wpWQ9tLLHAUQFfddzOPkHpmprHVk9dK9QGvpIWHQVdKHQNn3MjABVxSru6+h8mZ8CraPT41NGR
xLNGT1ndXEWEK+C739ItM7nT05bNuhnQO8+XsWPHcctOz3RPAp/qoi3+KPkN88VUey1Yag2+t6gn
pXm8P03Bxz/20iF+jtzeUJDaDTxQNWTTgCc1F8D05JpXlgZ4jPSMJlXe4qJwcCvvlkdzaWa93BZv
5UjsdOv5TgnQdMKFscJBcFc1byszpacHWuDsUqbeBtCAqArV4NphYKWa8moM1SMXO+H5EgUz7vMy
HBRb96lTCg8iN0do59wmoUYri3Eg+gFsEDVxNR/Ivtmv0roud6sqaS749yU/Kl9zmMGOKEiGbUGG
oNll18/lQLdQYpND/M8YMwOw4f9Qb6u+Ecg4Q3jsbaIoaeH726aepup6LouHOhoPCgH9gnVUuXoH
rNTQHnSInG6NbVTADdOmtTHq9MYMlyP1Ngjg+E0xnHFDtejL9kgBCyURQEVGZdOhVZAp2P3z7ZKF
1a2n7SqR3jNzbCYZ9YrZjru2SNudwmlk3H4S0nkjIdtFP0EqGcs4VML2CI0IEFKYiH3QxfBIe7MV
aGome6kBgd/gJ5yKZE8yc5C9vgdeS14p5XQ9u5DN8z5zaqNtw6sRpE7zuCjuk6usATuMbm4I46Pd
RN9WziK4aDiuRD4+Vptdoca0xQKJR2NZEZb8dQmW5N2co2JTiY4Yi+owaCKfUEx45QxjHxeRUiA7
GxcRA3ezFDGcEOm/P75y+/9ScTKoeHGQTnobGqdDPY4dJvuA6NNoy5xiYvEtcnBvxhGjA8+74uqF
CC+bLO0vbuF2Ec+M8HMF3/XSiXxsC9tDc8M5oVDlMFD5MH4Kd0CS5Mq67LPtuVhamqCrhWfVDFEf
Q6tCkgxk9IN8jcIQHFkJjrof0WClDJRBx9P05RWbk3WS3I+yFX+MqZ5MqbeNZ/b2FEXFsIfFvU7f
ECJP/WsgmKEv+5L4TyuSSZdRpWfg0KN3oBlcsGxHMo4xiv3FbpDNLJVq9/6RR6ikyy8ruDf0rvNy
VThhbqGtXhszCzEFDLaABmSYnYYD+aMwT1J8F1txbhQFBX2Zqv0j3YscT1gu664JdDwKKKiuNPRh
iP3rQw2Nhm6a1LfZ5mGwX5F3fArI99BBtRdDRb/EM1kRL16f+0dTGDob/d8fMHNqqCeoD9obNPcc
grRcKrKafs9Svf6fQp0ZlXUBkqEIlN+xhkA7j5HZGKu1uH6/IKrfz26vR2BbQydwUGUBJDoUA/U2
P135BdlSYhQipqMf++PpvncK0eA/07A4Dto3wO9FeteB+s+FvP7u1H/nnmOdp0+bllva+lKjbwqo
cxQPCk+jUzrdjdZ1ErpzQW/+4vsUFOMKg7uaSZiAkRxU2tiI+gPoUq7AhbaJHLmZspizlclxe/Mb
D7vBBTWR/kG1mrK3AhMs++DrEySqiDbn1KDGMNPBepNi877wugAXSYZl1EM92D0K+lhzZ2fIQGmG
6oL55cQWfcvIZXHHmMpkAebAKU8eJK1fx4aBz8YmQlSUwBs1bTvNBJrkZUfpzWAIm3GzA8FGzhn1
273cZHngT7QpaZpp9Ja/okvoSrbq96sKR2ya9Tje70aeMJDVOzO97a+6wL3P7+VOgFaU8qM8tIe1
+ioxCBxmZvQJ0NyJ3Q/DHlHbWRwJPTrRbhenVFGg6W/FglG408WVipSTtG2IeBFkKEajf1qRsmCm
6GpsSt2f8Ub2FCk32hEQox1uEimUwc+fmhOAkiSKOEa/cQaQUGizZI6BvfzDmt827yvZjNDK2kkk
1ncyxUU7nVeimvQgyFh3IfEn4fMsHo+a9EJrRELVP5j7HMQ4JUhLLvjSYkUWEUXxEmXEq65pqVGX
jl+E5dQfa8+4G33NbWQZngwpsbwW+LvQ1eW5kdyLp2nbT69w5NpjiSoVFmVDuyOkFYIMLgIv9axf
4LDUZO++pyfOCahmlOojM0Y0Ji8JTcyCnlU/4vwvCoJeQn6alovTVQZgRnhD60p3W3oqyniUiwNB
9YLxtVdjY+OyBjajMFCbcnLvt3UWjsTTBwlRTVRoNeQ1uHHMbiJGRKQK+wm/ZmAUtncvpVfZuvrM
ZjLezA87xdjEllcrQT8zJJ5mbQmvGCUFY2YUqTUKoWY8LGEnFu1XoPE6MrlfrOEb1j752Olwtwsi
YyO+IItq/zzoxX2qrkG2YDP7lH1fHTvTpebaKkGZOc6tvr4+Td1rOrwBd2MhqgEQ6tvm3D88lzfq
QN/aIH3ssrBOV17kKcJxh4gRdBdrmL2a+7lgsDMUa7kUctTJAW3bEVGu+/MI5bYMi5+jnB6O/Uhb
0JXnxLa3ET6dzQLMQOYxfTYNxXptecoKsXGwZKDapDfbcgEww26qMFGZGzq0DPrqAy4fd7BIy4u+
NgaDbqA7cFwwC2b0wPE2zGjxlrexvRDfL0P1+a6FTZ7HBIaKT0jMKNBK4y+C7eEo8Ug20AH/7OJk
WAi1rFOq6IwB9BsWOvZUoxVfzsNA6CWeS5UQ2z3m3Bc5zAj7Axr7xN7sMD3eHapSQfo/LRXjIc0v
cdHisbMhDC8WB3hi+WbNBZJxRbFusIkzV+qlITEf/YUrGOxOEYtWBDmALzNtzl5gyRK/ajk+5aX5
PqXz+Oag1MqU08x5MMDBiGSEDR6AniuqjhItrJ5qMzh/xWX1Hv4VVFeuvf+mL3uKkdeIyf/I168n
BqOCkJqCSyxd4UMRi/sgd3FDbFVq+wYjblfkoJwx4FMt/1XnAJWaGEsc8tKKe+1VBpi8XFKY5+3+
VBjxgI64dqB5TjNHTsXWMLuaTeNSMle+abWYcTHobR0UPhINkI5Nsme90NMBhqSm1JDBgCg5HQGQ
ov4RHL7iOyL06IEq1niTT4+dx+t6CRck8053iQ7xuLavFdFgkJUGEtiLedj8/9lh3GlerfqGlJwD
4h9UYwn0s8bC3+c009iszzNfNpiFN07GqYKJPM9h+nqc/wdT37dQ4hSDtsCmEWv/BE2czuazTkp+
122VUUcE08JycfDwKGSPGe4ehDJTnjn5cP2+1/9c8sUY6p8YvZ4Z6caDTJvz9OjnJ+rsHxK42qAN
FveIUePgPUkXFgO1dNuCJQnNu2naBhDk4G9WwUtslfcL76H8bO/kLsjXANhlpqX8SuNxNITbHCqG
IJnyo1R4yA8rF2pRqvsMuU067Q4XtCvc2dRB105ECwpcHn6C3QhixdciwdXL7dJpmGanR2jQvPRY
QFmwTjSi4mMUCLyhlYn6A5zNLNHjN2+alpPQt9AHULfwlKjTxIiucuwVwd+wdGhcu0n9UMQf8MaN
YnqmcFQceqhlImYuyG7mLq4CAaG9UJ9hl3DgP3vVgu6Sh/vbTI8YDPuBXE/MZz+cuh0abiBPBsJ9
wlfSdI+HQm7VF2gsIqJhIqQIMn7oMDYac0ngIuJYSFbdW4OCcat9za/JvWdFxpYY+a9da1k/Il+u
PCrBMarNAF6FLzr/ubTu6ItnzK21kO85owBsSnLtuO1mg6iNp594YDtP2mV0q4mFBOKuaFrMYDL0
hjSc+o2Jj3pwSREwrIEINSNLaym4aq3WzBw9X23qP8f82wkIIVhWNU/tB7ElC8jqCCTEzMviNq2M
qSCJ8Jn+OnHEKt1d9pgE52OvGPR691ODAOpdblVhrViDtS7LWU4C/ZUp8CwM3yW4WQkKqQ4SDmS+
/o0lFFR+0TMk0NI60WKl5oZyyEc7o/W+/d1sqxadlR9iaGPTUXt6/iVhP4N9+ESwKxB8vYuV3mXk
0o3zBk0ugrbcKq2DP9aU6ZtXKU3xPN3qQzlA8v295wQjdvmDHzCk5+9vGwETPB1hcFssJPx8623F
B/tq2/Ky6z9dQO0VRebkJD3jfLOZDMP2tj6eyaDXfTuMPAku6KDL7P3x3IIuwdRbw4Y5eBT3M35y
V1edlELNShJ9/RDxI4NGr3EbaSIkh2j9k2lY0CT9h5xIdCa1+cfUnoou/DNbUQaUGTjIBd+vRSx0
spFrq7nlxKkvhBZgxhRmp/DURd2Okle2FA7StVXn47LjH+E9f4GLfow7O6iXx3hWjkGtfsN8ESo4
zQCIfDNQ0N/YUQA/ODb4Sm1F1D7E8JTyoqOBgRcFuRYSvpw44bwRTrAYdZiaqWvcgeMsLl3HA9vs
FEImNmYOamDhftPtuvjBVFadqiLdeaCE8GT9kbO6WhWFdGxhlQNfFkfW/5IcOIrdH5PLMIllSq+5
u5HYR8B1D1ApySLlocjnDMYDRL8Nxrnh4RtbYoMGkx3kt40KW9+YGnqiduXaX4oLDPPrPoV47Eb4
FmvWzHRjIDSn1hKJjhnXTskh1AcFXaO0j/LNjJyTYCskKZSeVNF1zktDUWb/Gwf052Lw7Fr33JX2
8PA1jEzkY3wY4W3Ek0mP5Qn5XMhKMcDqU4kDSrlov9oBtqc4/J7l1phInTZJc9sDLK0Om3roHpEP
4z8LI6rXGtgr2yMaiMFvEEEgy/z5N3diTKyKJI7GB0l2gFtYWsPlxyGfzzCc167sRcPa/Zgg3/5a
H2Ui+pyVqwk8KYhON0hI+2jrBHK9FYozTbHar9VYbawHjtXFwvLYerxQDxAo7w9O6T0dOK7OgG//
CkfYMoweJRASoavPB3zmRtsqc+ekkOoF4Vrec5AGg86Rmh4paOLxbMfh+34GJxfeNr+It3cg7OZU
WOb3md3XJVN4/y28rWbczuwd1GEKITCGmcRhRoIbbGZhv2ndp+758qxkau6SJuzvw7ojnEObeGpo
9D42SZSkswwjNnKvG8XPvO62z+XEpPhPOBJ/8yBJ1XQkdGJUnFcYsBKjgpdOMWyDLMRxlHMfEI/+
OLYg8kxpNLvDCPIw80qNcsrP0MHNRNYvn87wusZb+wp7yV8tKdQEhPoHOH8cuJVzePyGy5IkGYU8
yvuu+ez1f3FSWUbHB9+3divKMUavHMoaS3o2w4dAhubll4mN6I5U+T5kBi/LT3FgYSUZ4y+/vkRi
P35JzWBdtSo9Kf5AlWx0NaPfHbaj6C/4XPg9mR5hL2nXIxPiiGr1T9uoaDuYKGH/KrfDykkPlw/q
Egp0op8IdB+YZ6JkzuXm05WVYHbB2ptrIYaNTezvAcw3zrIiuV4eCBSNYafNCEUo2kJp39pWnoSQ
bPAgHNezjbabO7sbkjiiN/ZyPN+lriQOHRX+JHPDfaSI6/oUqC25iCUQxapp6/6lncsMhhrWAj1r
/ioosN0F1Mi/rlbcsDd+BaTh7f8mpiFXdqAYIe1524OlyzzAwTpeWA6tR+FIAgvvgJMLxVTj3rgd
LEJBtS1WhKjBArnUXX5FQHZpoWx4jkhSxG9+ZO8UPWAjj6tvU0kLAgfuZd4zw9iKBr59oIIBEvDQ
yt1XwDpGwMqyUfniMOYJD79FBE4WEIwtCjKmtDOGdDI+bfTuWACSoyAlhEMNhs2qxh62HFORH9hR
VyNfPmjUmvVLQoEkrdep89xivyGBm+E9i7DZd/6SHHcArrxxpuYfRe2YrtZ/1ZB6tYmis0+FXZYN
eIkOn/rKzTe4aUICbUaaxAIqPzSoojPLH3O/oBb7xyGzUcbwGS19AQDkK6QAHm7Gahi9d4WyBjqO
xbnXb7ehU8LSSUg9VpRYogpYLGSFpjgm8EHF2h1MpmVUV4aWQ4LSeOsNoIzKiXETUbsoLWfulzwg
uYr9fszIAd2ULHD94+YQXawHCmaC7G/fy6u8+ew/5mcRV9eW+bAr5DAFNiShuz3KXPuzpEZz8P7q
Uj/EwLYZe7y1A4FxOMM8KyGKjwARaplk9BHhtZf8xZo6DGXY8JHYE1riLftuYVsUf6q7+n8gJk9w
a2PPqjPA8TwtTPXyZG2AhOkZp8sLK0eVAMC1zVFfKy/lkTVYd0KaszmrUSl6dFv+ORXoNtfFRzRR
3hMBIQw8J9bEqangmec2+K7K/nsqNkEiSqTCq0Kx7qKVn/zZrD9FVTrSkmYeG4LkrDIOzUu6eonz
3zsnrygMxnBXCYPqOBBOAHPEDEjtxMLaK0kd6xx/3koLlokyXZowfPhEA0ypBe+ktBJO32mFceoX
AIOiSfy/2GJ6JVmFYa+OT46KmZvnlvuxmkTCrVElR/+g7WVkiCtV1vF9u1ihmEzrcgTLdgmBhc8g
1HvA8FsUx9Lees9f4ins203/S9TSSd8qdf+1JvdIVzF21CDfZ/PigLcXzI7hRrpBFUntuwsXKVG4
Obt1l1EddW741JuKY/YEMrK7Ojng7BsZsKN0t8qbfQ18BLrKzMDkFk2l6sYPZqNJWM9F/HUVSUxV
fcOdRY09KH5QalcpIrHBycZ7Sl4HUsbVlWg69hUXYyx0RcTvjhFgc4FR4N721Jb05TGrwVwZXq4k
gJyrwMSoHKEQqwrEA0JMwv3baetkzGu1GSGgvGFQ08D+juhqK3hehopka602jY0G5eOiG24nKtlR
Wql+9YbqRudEqzSpTOmf/beEMv3xwbbTwcWZplUbMVEuKUJ62LEgW8WjE+MJr7c7WqF7LeMQjy/7
d4V6fpW0SpMY5tbIXzNsL5AOvn7Rr5aXvRBHSSlSBnvnu3ylclAbqARX9Oi3K6ThTmr0N92FrLlI
8CJdYmdNup0ZxVQsPj5zEuLdQ6Y1Kwfw8kiHlvaG8wpSFyjP3sxt0Ifh+c3pEDi3Qthtfv97gbto
fnenR+cM3+kV3q3sxez/gDSqnuBOFGDAPYvzSKR4PEFlMhBtaF6P2BOPY5iXRd4ZxTACk5lvW3rp
W6AlmNgbptgo8YMmcdFg/l6Bd3aRFO4rZyC15JWvjhe85TEWdaQUl2wTtdVjNV5i0ZUZ/aIz49Jn
vi+1Mr/cPfkVgK+fBLxG+fXsB0T8dY8DIYOfwBeLvraYLKmQTYW83XGh6zjps49v01B/3gME1pv6
E+LRIrAA/wCbLuWEe6OP8ZNCVUfmOG5lCvdjP+SbDVoJVMM1XUhr647tDOo9v8tepxTIZpiDpM0A
vRubRkKSM9DVp7VqRVboFTIe+810fv5WYJYPBLnu9P/PlYqH9Fp4JTggAz61cXhGS2Qx3DK8gT4r
FVE3M44lg1fQbyaYtpQGe58xXjK2V/UxQxeY3qQe3lO80bNpIHzvWTBoZw5SSLpg/TwZxIN6Oa1v
x/d+EZr2OVfnDY8CEsUFgf0zI6TYrKaAbaLrNBNkhAmy7rdaT63VvZSO4eGFt+qXoM2uaVkEgtxJ
RT3opb2X0+dQJgfn8DZwHRRH+7lQgv+qZOCwEYsXEcGHhPsMIiaPggBlO2HXh5sOn/NvCpp8HcFc
wJ3NLkhrjzQxHyA81mALl6vrd/QAxndf+o41ArHChh+6OAhjuESQMvuN3f6//9SlzOK01LHh+3G1
uNHMWve3ZriE+o8012V2/iuc6Rfxy9XFZCqtkP9vmKet5Hfrn+7AuBL6+Hk8w3oZhpEYBYB3NdjG
8e6m5d1MfgfuU7MBj6LvXYgeMBzfbruOS+vxiKD4JJ4BH/WjMiz4gpyItZe3a8ybSkIw0Os4qgGZ
mAbwdHmNyegDhty1D7qjEOdpoII3CtSEFYBVOg2IIbz9iEE0MVDi51UaPsOcomXqgrIc7vSNN3CP
h/zz4Wy0obC6Uwjh0ZGi43kiam09bElbuHa//MjkxO7FmorwK4FAkD6hYwSlbWt28COgmpt+ixfA
Y1OnFD3c7tuDmQcAFQ+luIrGADjiTXzsAnfzLXFLAUDfCXILJTCSIdlGmsKaJxrF+odcGohqaJOC
8gnoQNWopfyPCiUdCxkgHi0fXe2x/+rP9f771OGWQXuQo/r0h5CgRQ/egL4Umt7/dVrxLlyZpnTU
vID6jzPD4JaSqgTm1EnYxbHp0wwDe1+a7Wh3ocffOmV3AN+tnbcmVpVp265ag1HNcbqBTrcgRPc/
LnlEMl375EM9exO2YL+I+rEOQiR3sUVl5EZJ3MLGL+WEwgvF/8BBjF6oNslJXRsxbpgHQsTnaF6u
dyBCNVpG5lmBBexOI7DjcAhTYfw/ow+PF1JKj9fh0cBoxKHva4SbLfTIwGB09twNc++noTOoalZB
MzofGzGnosPuza41qOunediT9rQ7J0CWByLI3iwPgd6psiaQUvt3biq3JWlfpJ0y3QbUWeN/2gf/
HO6oeYLQoXL1vHk5L7p9HrOgOs34V6u1zyS38wEyRdddqQoHOTr05YUfVdS/pRZCwqM5RcLmgdee
TqnZ5m585+KFMewN866Pf4OwNShwd9mU5AtVdln4PzWEUMPwgw3vIo24EBi9xd3sCvGyIca7dAOJ
2h2SFIJKMQE8wNXWN6spngldvPhdaNvcMQBg1HxNHP4u3s4Ogin4ZvRJ02fgIiG/mEJBKS+aMmFx
l8AqGM6y9Fg6nsTS5kLVwGqz9bsa8T7lBiOiE9Fhkq0nY+rJAJQ22p9PufCDLIplixmxAPd/yIeq
35aYGXDadcE1jb5HfA9xwioswpeVXol7BL7Buy20UgXi7I4f9x76d3aUif2s8LlHBBCwFZlBQ3MH
pq7/9MQaH3tllyRr7lNwCV5RhoQOTj8u8xZx/guOJg3pOWURx1Cr6VjX7Jd79E7sisjppCNV44p9
nLWYVLZ0HrLF/bkWR4HclOxhK7wYD9nv0vxUGYYzyj/m+dK/GizaxtJV/s0LhnbQpnnlpuKMZkNm
UlBSmPAEYWBNcgPwCEDEXFIwXrTvgGw93Qrr6FWQaqygLArr93g5ej7H10y6nhZKYoC/VScQ31UC
j6/M9rNhj5cG9VKf4pDq6uoivijLKkAIYr1BNzlfIjyMjzLsBdDLOpzP2EghMpRh3FpbMf2LfzXg
JnGOgY6NQy+kBw1IvqsxQn/jJ4Q5sTIVt1/yRq8CM11r8vSeAvn0P6lD615skqEmnZsaSXI/1NLm
24DRL24JIuZFXjpnkdy861hbBdYcrTyLL1jMfeZLXQhYL+kQUdwawVkPxsIL0eA/OcxB0oafwvkY
pHY/FmKGPIOgVSErxY8nYpoufStCM4lREVbWW2P8EvCaYeX6j1bukK8c+Tjs2iNAFM6Xfx3d71dE
eDDyXT3X+BOWKIJamyJUWwcrJzOpvB89eGqTvQHRcHc8JV+aNW+9mYgW+f8eIxLAD5D0jQgpX9Cx
6vp6rXFb1YyNyUGQrOdVa3KYmmLIoZB7MBQD9pP8HkXN2xl+iDCoRZ4GU5ONMEVJ+tiOkXDiwMV7
XUb2kfwCEa3da6CFwrf9miPQVPJApuBUMFKtuFqeCUYSBVDyA0+DOl93HqhAot/0gdJuW5jbz5Xn
tq2nxbVSJiYQnJM9LislGsmt0GENb/eDhp6R/OL6jCh0Pu8jOByjNxbAiZXpd1Jn0qEWhYyDiDc8
uPiCq8Xxhc83XbIeIrP+YrVsrdWJXt9ptrrgznppbY8UQsKvKRq2ZtElDkVeWJgDKPfbGUJ3k2nc
HtuKzLN1zwqhlCnSEL35TV65avpmTlHJbYqFr5Kg7Dtj61TIo2gVQOL5dbrN2OAYIbPn/fKdLtv7
wgWUkte15A3DQKKT+vIR3uPaMBTgyqZJRWXtiuKcOBt8Xi5u3c816sMte2JpjxwoEKCaAj1/ronh
yusrCCTqilGTUYm14La4KkLdg32Piz3jwiyPO3MYeJBnggT6GgwqL/3MNPPsZyzRKFcF28d1YB56
Z6VoQGZjGs/qHJVm+ASR4DyAaw+LZIUZpDL2CHq0PdH/tpYHdOreEJOFrXBZROrBHdCeFtIQXRs4
3fs+auyRUaxPZfau6bbDJ+6E5W5UZ1phUhipnFqlLs+XDDc6FlbfRIbBqVIXCYewrcAacpVS2f0c
620vJ1+oGa+zMpILQ/00Y4nciqqvfpEXiSrHIx1XmHUvIR8mdIKCPRdG/9/eoqgLJCX3RaJgqLhb
p3Ract1QP/xa+MwTlhTuio6tmqFokb0i1tQ5ldbPWHFIXSRWnHyHPaCwsLWjQjHWKC4XG7QuIh47
kGLtrXj8wMsc5fXvEpwR18nLjgv2ImhCqWeBg47mnbEGXoJsRWDr2sbvxGDlWizEu1xdyFkmAprs
7giyTkmax10Y1mZWtX6OdpUf8gMrSvvfJTP4iD9JVXILbMguXJT5mIT/0sLQphePicaYoG2hPUKb
4FudAr8k0d9fP50cwP4lhVph9XS7rG1IQgQBDiPyD1ZCvHf11itXwzzdV/Rc4/WBJXNrlOWkhbLz
5g6W0cVhO4ILNiFG4bm+MFn6JVc5PSjSGX+RXqfScO+y4NjntlJ4dfbwC7n4qbQgQhDami+ZHa8X
puEQiBgGFF0CDVUyK8xKgZvWp3wD6H4rIVbSc4kgSN/0Gz9iXaiAMgGXDQ66YtoLbqMO6ydVb5pn
juvfTRhkp69XjJf5tc0xPFFmBUWSkrDbBHWlfLOg1lTpyApg6PxvrIHyzsnL9LSzhh3AuDn02l4x
oGNKg+QpDEw+uMQQNC8X/QKcA4F0v3nVxfpfuAra9jfH7UlXActKCbNt54dk+C3cAB2lVruYZI1q
ZORmF7Bng/UPrrVExXO/fK7NVON2PfWV2WmSy1iWjqlZ2a95QQvhV+1R9L66AYxzN7ReU5sz+4uL
2qKE9fdJ0Wku8VlmUpuGi9zMC/ZfAsHGGmh4rcbytvoojBpg0m1oF3BPUItWwRr9KLy2Fopycv7B
oYwrPjbjDGSF/FL9JbWzq5HZ+muKTWBHiN06/4wY9yCjDnpjH09B3jQ9qWcAdz6BDu7YZfNcGzPd
sQ9dk9v8nOm83EHij7aHUHD+zOtbL3p41aIuJMakbaLDwYHRxw5aQzrzF5ugqUU3GogAT9eKvNmJ
AmvsB2z04xR25srYiQUutZ9x9IxA1JMJLdT0O2/y//SYhgrXvd0219aoB0BhymIh5XgiGIvWCnOd
04agTO5LLsp1j1gJb0w0Pz95V1Q7QZwrGS2RnHZwM/2ZMV/cDpx66mZmrdvyPlxIaQKY80v18+UG
WaImTBFlpJUhFhZC/xUpIvvkVLiwi2ZhMFtNH76UFgqtISUkEHtyFIYirWcgHavk1cDfnKXmycmG
+wQXF/WbxOedOAV7T7sFOoPvOHnNnP+wS65XER/vB7W9MjfkKHrolN6/ZSn3Yk9kv7b34vjCW2GJ
SIqmhF5PKUoErLidh4f4oDfRJS9X+gj6Nr3nn1c6B7zYEg37/j8kMiXpYS0ze5HPn5cuyozbJL1C
7o5R1GoKBwJYOfMIv0FHG7ndj/pIH3ASrQI/53tM+THDVMOlBr7ZAJe4iaGm4wGajpv1kkogPlVB
l53YcLwpjS8yuz8TiCrqQV7LKuXCPHYOwbAPz0fBs5/6nk99t2xomvf4y2xggHizmmNtbUc7nO6B
MwAo+AdVCzL8FuYApPH5oZ9Czs9AsrCdmqqzdqFLLDUAfr8+QbXicsJFJWJlb+n/rlzMrPNR2DqU
s1kp0CmIsw5KLk3fqe3ER2P/1VtMdoOUa6R8FlHXct1ObrH5A+7fHRR/JzUjz3sVWc7BPhCx8d12
doCv2junTqVqhYM/9DlvRGIDuMIu8Y6Wwxhm6n5UqgFugMnxbABCx/TajZT+YoDhrqvACzNKnVGf
5sSK/I08EPiSFm0/0M9n6KGcYrOOtz9DYXVSv09WNCGnE+r9Is0TNaVc4x1DHmo1R0ozYjTh1Atk
bXVdU3raBQGEV7OvQbZb6PV0nn0DFW51zhcejtXUN7tbAR6qybyRudkOP1X29EyqMrVbvZEGxf0J
HXQoGQIm7gPMnMsnvc6S9KTxf5tx0hWHTW3++O0sEhvnT963HMLozMM/lT5aMHqsiTZQYa168Ha4
cwYyXpuUpFvEYBne3MR56h59ktjkJ1UvilQNtlVayvt63eGq+ZIx8jg251KZhFKzPwdKv4+wYkOT
BPN3OA4Uj1kCUhTncgUwUN01HcU+jIi2pGAIVBJfK5m4FgPVMTqTYftYgylsUVenPPPriBAQaknm
2EamqP0Ibv1UDOSb5ONnhHwIYS5rDU3BtXcmbvcz1vMVcZxxyXVvCF1QfMuv5+vb+1jR05heXn71
WV2553+n18PDbAGherWMrCl8AT4GFijMOMhwmAKd3tYtiNFtk8GHRG4iI/Mjinf6ulN370Gzcg4z
z9+Xat9gAyMcID6dKnA6dPD91a6MnGGZE1wKD6N3xq7XI910m0JxwW6ehgDv+LJVNRNCMEirB26/
YPQpIH9340SMxKXlB2eAB25mVQcQ6OH8daDI9h/RIJWx5Q9WC5LdaNWBxaDfwKyFVK6jvEcEPpOD
BL1YNoeKH6xEUv0FBeMV8qBpAGG/rb/VWzQKljBjpMUZpP9f+d5dD2r5arP2zJrNCXMSflMortXl
L3YkFE1JD1pXhM0EmSijGpqRJA4j6aqlsm1HQiYYu4GJTDgQ9Bm8g+rU6UkITUuDHnu1NuYDctbS
7GmETPdDeJnDS6uGKqQ4jK/A8jpivdPEEvDG7JL9i8sEUZpNr00fIK1ZZXVpwjTwTVpArJwzcH3g
oZFABYjFkeKDQvX5bvuIPQ9xNemGUQ09aoAnwMf3naSumq7NVcY/JKyUDa19/M1/fZ1w/C2jkmAY
MRS64xSGIQPPZsJvgV0GdNnQgnfo+wLmoEK7bIiQ+bhYsjh9DKavbqgGBQ+CbDyRYh7YtVpiG8UX
JRW22lWaB1+LiLred/kuFzbnrHfLQgshQvrVM6dnvgBn28I3kqHDs9P34axJNE4/liE4o0VZPevL
DYAUH1A5b8kvGN4pURWJjFsnzcTNYhwH/E3FpXb113wNkvUmThuZR2GUnv2gq8SKRYQvodXmM/d2
v++HQGj2e4B58bPcT90tyyQcb0mdhXabeIXjWPG4npE6izcpb0yuQHut+tVgcKbyaYrkfYjnDOuC
oerpER+W2Z6r4bAXugGqXn7IsMVSLVK78Wmxe54gQD+iNRi7XE16GdbiGfBbaWzFsIZ6PJ8HRn5C
3dS2L4+2efVYw0oWhE1Jx4cEimBCnrxjBkzvO/YmXexCCv7Ouizk2jMxOsmVZkxjndBlho09zQkG
P5GofwOaEy/nAJmdDXycASIy6aibAstZWNqFzJnMdDC+aqqTjVrj2xrqYJWpz3IbB1WTK3yahVKq
8QjFG50SULra3zi9XrfHtYnDA3OAlERX4rf71NAwf+AcAhYhQTk+6+g4QL9Q5Kzz6I8qtR2Mr25z
7/MqrZU+I2FYYyx5/gXPksD1byUt8C7AlBJ0uMkqYRmuZuSrivfAoE8XwExGtnE1vB7fkQcKFFmD
+y9W1PduBN5inPQ5mzTOu/4dea1EoCYDyhW02bPTMlWKLr37NWAucaLjM2WOZC3iXOlOtAH5bnC7
Ve4l8MJu5lWcDcPU5avX62ItOPJws/amj/9ggmFAQiLBvKt/s6k6+8opBxFOpzKF7r7Hz0QdTOli
GIZZQplaujtDhanQJCHvrrnV4SDtUkJJ24PwLiZDhLQYDlTnOnpyF08kYYwjafY0/TuBBYU/gIwU
Y14UzjNwoA59r9dNn/3z+6i43Yj6Fxe6dY6YtfkXv1QaDbDyTKNAvxcM7B2lBtCd9oNNOTxV8zNr
d5i1aO3BmDc2sZnOpFvj7dywGOK2NaZNNTE1x1/n9id4jsQ1gDp94wlt9FEnbO+e+YcencoLVVM6
B44bCfgffq7nyMFPZpTcswGpPpGMb/6tS9LqBXDporL/4nFUVRkgSB/eWdbPwIwDpsRBB0HV+BX/
yWA+nDC2Gxfw3v/fOuuz4CDAnLS7VRKGZUtviUzru1J0iATcoQmn+Sr2WNLwPUL/xgPZetG/XjgF
ACVpL2s3QIxRMVMmeHeCGJtptr0FZVS/YhRuNlV4rdw/zyABk73mUmxQrK4eDa6RgmrxQziK1b7j
5T6/HTBwO/LfWHQhxkRhbm2X4wbpctQWmVnSy5xjgCx2R/OPyaK38czE+DjmX7j+yjfZghU8+eCH
QUptwmmcdkCYp0VD/jQzmLPfwFwKhFHCgwhwIU9Ekn6ZFHR4bnaSssaHfg2EOFT6le8dkf+disHn
yesojyaiaP++q2F3axFf8xmP4QMlyjsfg/FgiMmkpc+Jq5y+YSc0OlhCSVMW/rGK+Eep5qGqFRwe
lpZQ+KSYnpjOt7SPOnFaIMmoxoP+za05mSUtM3oq0bm220yY4HrNAjn9AaZf7IHBoAh4WmXYWHBi
0NShBSisAhC22Dx1dn3e99sPD4PWCOWi01Hsq4QWa0foNhXrnTjcmeFdEm0vwC4GZqWUeLzePzMN
lycUPkeV4Tsz0I0kEdJAy0pCJx4kxRWtHcnL2uWL+O0y1jv588mjOepnQsMyfIYGAjILk3T+lo4B
4p0Us6KAJn/quJhnujGIhsgu2htkCcJoSooJXt3Klw/owoQsf+IGJD39aq1V08/5C/5z/IpORZ8t
iUVMBwvzZwS7iF3ShXOHIhpZozxW4fd5TA1TmwQGe0SzJwBJD6yncfFT/kgC1mBS9vT2l5pa5/0g
SAYUmusI0m+Xyoh6LDqia/NbgDxvtTLV1HFD6mS1byh+iO5ioW4k+XRxkLy8TSjrI3RRLQLoiAir
Lh9y0e2p5YN6Ccg5IDjbwv1SywozBvedi9DWOI7QheV3UrFGwalXGSlcApH+mjOetrv4SXuXBgLi
iJ7SnP39fDKUG3forPq9UDSDDKzP6SWBV5KiK0QxVXEQQoeWk3oVocjBpGV2WQfql7gps11U9zN8
upfMCzvF2jL8XY6nAynE3BcalKXeZkYrzI0QAq8V5QKX649gWAkznh+/gtVXFkFneqhAj49SFLyr
sebSgQprmTWv/sSK7V5A3azGTVi4C4F6TgbBMr3ANvjH5WkVuSyYcAswSFI48Cv/SNXhI6CQyCtP
9IpC9xZWwhdvVP3IpFanXr/CyzAzXGdDIxeP2PR1lNWayRi573PKjOLutStnq3Cn8PRPyx565CUw
cnAvCC2Qa6iS1j19IVZLrWTh+EoNAIOg6XUd1FvcXAmgLTXrlOc/vQ8RxbO5/yQ/p78jfky0BbJS
VEtu51z2aO003QjGgp3tqcIiQ5N9g8RBMSRMFN3wWh12jsU3MNUMpNyRLBny0OhCLMPYMlsr04GQ
0dY+Z+XrHkqpXVl91hur1DGDPM/rGdDHQXjVnKc7HBSVobrzmfw5CaXHgK/bh7kbpiKWMHgYeEEd
DAMg3lBHjRY/sUroCJ+ffpQDS3yBeHtlGSY767Pu977qyIcgvpxQU73iyjnizjsD5NXMjEysBlKb
K8MRe54km3+UHB18s1m2NYKQhaCc6sPYeYIw8advxnEKQi0EGbuE/SpXfbdo8s/IDCq56gl7bes+
Y3jK0jTGSBJXYdRSH0i+tA9E0b5KRtl+mwoaHFzJQk4VbBhaouVlLg0gFvgApgzySBVA8CrjLNaG
k7hF0QhwFn8C0v+5fAFezlQeZvsGBxUvw8YgsGLiNWn1+gyO/3+Fgn+GomOe5Fucm9aDYc3fwrXt
xnhp2/jycctirCX5amMB5Ofz9nIc3lLRCnxTVKP6x0/VIAxri/TIg9pYFNXIxuf+lTLWY92IZ0dK
a7nogwcHaqzpGDmgjKYIZbQXVMwphQJTXHeYERBLLMrmI45t55Nb7XNwvnRUtAeQyZ5N2UKPvgmp
+oKMo/U1+DEY/S3VUojivnsgiB6klHVzmD8nfoz01WqSo/RIgJ4TCbZKGY3A71towcSQEmR5v+m9
OGaW2NhWzm06Jc0oEXm3VkPw3eeGuIvsNXiLkZwj5+XlT6h8kdW70KUcb5uZ6ClyowSe2am5biCu
4xZoc7SQqIGfaRBNpQRElGoixqtfhR6IeLsBEWRd/vRyWLggU+cD+8d2H0QIrVRJpywoJZme7zyF
NvtY3JqL79FV3FeTo2YeJZPGpQzkMby8fvGpdcVBfy7YdMv63WsQsNu99CZ9XlwymELa52z26GIm
kfAEjH3dWSaaQiH7MX53iEdtqmblvkgRFVYiIhWJg2iXQjmvU3sgIZ354GIXMg2p8TXjlxYwX/om
zjSn/hO8BdcOtGCap/jibnz9MvOCboW9w38OxRc9LXdUqiHlB0WsgaTo4r/1QmMJE5RYeicxODRJ
eP0de9dDKqq4Ez51Za2qwvG+FM/JfbPYzh3pVfocUGiZ6S2lOop2UeZW0+Z8XJx+OPLLfqCV0Wti
jrij9HqAfswNCGpevewr3DMQwS8aRV1HLF41zWz2Vjn1MfDbMha7MasbDBunK78+epAAF8WhuCJu
XJjbEeobY68uECJmIN2otKGw0vBG+6y947FZXPWIF6gvyTr23rOkcY6xnIf49eSnVf/uKcutLAA5
mu0bzHT9Rg13o6XbFpFm3012VC5hNPfDeLdnm7RqEjpY9SdhF3+AY9A4LAalg+6ksC4OAJPbWD0K
vyHGKKwp4lCQ5rwAMKEl60a86zeaQLc/fCUR8oTH4B1W6ww39e+bTqfCn8AfOwbC1xHgBBcrdk5g
/w4EggBqxieqnzM29FR9IE6+nab7Vp7jveqCiPkpsArQxFdVhNOg4/FDCMtktqVyMVORBu7gOgFW
OlRrDiP7wZEGLWvMjNU6Q6QJwNXC0YKSYoDJzKXHBRHn69NS1a8gi3xxXdOyjs3yP/VmqhnIjwmP
8urxBlCb+Yh9Dkea2ZB3/ArMmCVSPKv5FrfdGzioxxcGdU1HRpvlfsE8nxwhSNuwCeoPR0XAdJ73
+PuRGokfCG8IlMlOFB894TCL/7LxsmcPM35mRZ/eS7TE1MmnTUQRlc0p2eIP6gC/M3vIsuVy7XxH
nd1kagKAr5TtfS3Z9eYoCS7io98LHUvJP3xY5LSx9zAfiUa4W0b1FHW21igWp9Glvob04uYHV7Mz
CdoczuPNyqTDoa4ArmqoelEAopQEBtbI7N8+JWDqm/t9YB6TvlOZ32lX0/NDyVM8eKMW8ubIi3/T
4mXowlD2bXVnHUcXFR9Q/8g8ZvHX4IpQ6ZiW3jleVkdonpc365f8Ir9D6tz8tfHjB9wN97Yc3P7g
vnu+kmT9m6vXLegLFK5Vd512lLR8ZWV8hX0U6GkJR1ernut1hwwI5A6Uf8cgGh6o4uVBnYcdxpNU
pdsualD1nFBNq2o4vZ87SK3WH5HqsvVBeu2qpaxjVbrQm5tTVbDWURgqLfHAyL3HFNEKXL4eS9wX
9pyDoYakV+WJAMiNbA+q+RhT9ImvxmhF9+FkNf6Z/iNHcO6/fve8PGtrhqC1zICX5IWdQ+L8yY44
ThkB3KZRHhqpaCgjNhDr6kv7mbo8V8kWp459QrHVRm2y3U1U7qswCsFHfU37r3TVkezo/AlY6oPP
5x/fX1LgIucanAc1zZ2b25CYsKTIGQZ+DbxFRAAUQjSvrkn1e+VKyJMhdEAiK2LGEpE2//Y3LY90
6jzW0Q7BrTZXoQz68h/iV+d9V7Tqj0QODYIRfKXZYeVgwmbhi2KUAbhr6aN56Xo50ul1j2j48wn3
ly95IKf2z6Cj9P3OewXxTdf09M/rnyL3uoYTUlHvJMLwpgO5hRsL1q9NHvyYJ2jkUi0v5N6e+miO
5CgZxxFRR8+dv9U4Bx+BuK83LaKiZ9D011Huq/wMupKdQWWSASQHjBgTsGsjb5v2czcE7CQ7zhlW
8b3QbT7ZAe12I2hypfNP8p7o56VKtpBfkWaJrpgHt4cwnuDzJCZLZJbOPJ4RV9w2NyiIHeynQm92
smH8PufOS6+lGP0tS2Xu+bC5SFpKOMOcWNO9mJogxlz4cuanpJMMoAgwuwLmWlm/EYRp+MR/gOU2
mGD4SVkgutcagG9NWJHU6CKQs3p8es2tDbOhfjAjE8e41zUeM/Kg4IP+RlNsMEwsTrb+C1hv40ME
Ae1xmgu+wTO+KmUCamMA0SiJ1dRMa/yQNHd8SFq6FZPQxeiU7wu7H+04oSrwd9k6Xwx+XXcLzCoM
bdqQKip1IbKmBveRK5z03UenS1EvLsMHBBDZtL0ynNDhX/vd+ZGzi6yOxuogSgKwVMfUCFVFM0H4
dN0PZhcCsBvNSuwv++bOPwKkKGjGPH1AUwvTA2c73GB1vrc/KJXskFBvZwIbDEOrC6pz8/HIpioW
RofLjy3NeflmWuodH3ihZAk0VwfJuredAC+2O8I++Sdv5uiAShr+zCExYyoiR6OeUt685NqURHIq
cwSpwbHEjPLTiNO4rFXFG/rDRoTe4J2ZmmlzkToVyeBGd0fy6rr+7f5jJB+4ak2vttb8QpR7pHTv
Held1Cj5aMuKiDQNC3Pi/H7EXyNKyh76MdTVXos/4GQx4Y/2n1CmgwBURdoi+YvtBjCcOqeYKt5M
PnPdc98avBbz9LZOdfg+ddGxs1Ri3L5KyCPDarrRXmPazHbVYRS8k+pnslGpV+p3UT39EtEK/zuU
bYsszj1JoFwRBnyHnV3seD/9BgUfQ/YfVYpjfD4qBnaESxzKybDSSxKkn+/HP+wsq9ub3LZK3dOO
5I05s9YEI8LYa7K3jUenqxEHpWG63j5h7R/U4SkCmt47O2kbO1kYNVFZeO3SzB8Hj4mG5Rk1Wec1
r4kOKzZnEJEjPPQS4FAKdu/3tVjNwihBKdkyU2ljYQukf6+TRgfjF82kkG0KZKelq5En4BrAaRn2
d+s/eDFy3RG8XRb5UUhPGLboqTpo/aq2LlFvS07IWWCsWquRzXnJoZ4w8FBct0ijj2pyWGpTASEw
CTy9dJYqaC32HOUW/tV32bBpbZuEy0d5srRhOXNL5vSzNMHs2NZW/eld+jUda+zufznJHG1JkER7
uBA88Ma4nW4IrM97UUmleULlsT9GnY55xd4nHYluWCcFeqEkBCH/gaeDacyvoq99Vc9wlpUGEMbf
WIn9Fv1oPyoA6MSRFsFmYIPEtSdsVQ5RGRoERDo62v4rXqqXZW5pvhaiS3chTalQxySBpAzH4u4+
GnSkj9H5eCm5VeZtIBJd8QgjFZCg3wsVtgqSJebOVi7UDG2GGteg/Mfq3wCTm8UbmLSq19Y1ijpT
TEo1QzNIlpo+GUdyXDSVjg4DO1rbc8Aj3tDQsY8/xeplnIqzDaBCpjFjZFIcYES8F8+Uw8wb+/RH
JqpG93lFMU0iehIFZ3HrsLWJKx9Jr+XeDwDQMH3r4VED+bhGSy+gtPMfixIUt36earYrr1igc0sk
TKHUMzvHTArAkF+Bm5EStd4TpFx7UFEbYIM21lCT5kPkGlldQ9dsM4BCBWXiCwkgPiigDCFZ6EK7
uOIye94PquyGnI5i5ZUpLK5gw7iBUT8o6xwKAvhPqwkvdX6+FGf8k4Dq7dqEzg8lM2hhTqUN7o9p
P4MJa1ybWFiCi/FEqm0QTTuLgxNcH/CcpN70I9IUcccsPrr/SEonsy9jv5hGoiIhHAedDEjV/w1A
ihjaKtsLNOOd7nVO4CwxI7x1weLlrDdilK31K2pqLYxebsa67o/Ge3i+FEav85S+XNr9bcZuvE2b
BovdtxchRvjtZdvzRS3px9YxHSOSwLlFJgUy26jKSWxKAHFqf+qWoLGEhPnU+z63s4WT75oM05zJ
Wkt8O7U32Xw8oNERNPaRYeTKKSBe9l20pHa27e97yK36uHo3IJMH4/NxeK2KZCiBueH8ETBgTKts
dBtusjhh4P80blr+Fhu5JBgLVNQVpGBxFWj0cBpij1pjCtNpsYUaeeqUx3MIHuNAfGPtnan1w5CM
hqYDrYvwnkBMTLITgly1J/iluU4MfMbwLHa34cC6UpYfSTtZpraGnM2MYC8wFRwRPJDcllDqw5cv
w28TJUBkYzaeh13hLaoszpTXcV2XARSNfZjbddSfI6b7N2f9Q9LKzGaRgBylx3hhwCKDWQWZQC0F
ki7xY8+Y8FPpIQHhyZ81WcFW25huJuALJfvaxWx9GEbh+iKz2TZE9xL6VQRM4+80eSNU7eBdRY5/
VuudA7Q1iOA/ZrAKrahRkpNqq22r8C0QHZU+qDKcg8Ivua4UbV56sel+g8id027oDB32u91imPFF
VqtAPt3hcj5Pqrb8/EkIVOHwqoiDiI2+LCb+UmAAUlD5tF3ZsIhIHEVRVIYlwk3jCJVqrJLcdIl1
Mw8Yi/wYZF6fOGHIjXOaZGcTPFyx7bmB3q1mvIwgy2p5DfyRLtIKaDfKMPKV3TNvu5vWj6G7D6U1
UsUFehuTBkhUWIeiBbCnqtUXzQbNUgTKJksbWXJ5f2tCoS0fw5XeyO9Z5eo/F+KU6DKoq89Id8ly
cJRspBp2lJfd8y7Kh+MrIdyRr0MdvD5wrvVrwzWuQFo57Qx4CCNcK8uO6wXw0DSGqesdqmyFNWBA
HGs8cx26JyWoepja6JZuF0ISlwKJP0/4/x97riuq/As6gJ1fuq+I8xYVFy8cNYhSxecQEAEaiLZM
qJfNGUHeatn8dx6QAODrTt02i42eLJCi4J4XK9GD8XeYPsNRKE6+g8bm1fgCvK6a1v61+xh8ZEIA
EVUWWIxGGBZbFclwhfJkC+VwEAvluM/eHAnBsBBZYz+0e7qpcLPz9sVvA/IaWq0D7OCRwHvS+ZDK
aFNucqioU4jr4GemqUjuD8qtxAk5GtgVoxEkcfkD++GT3Oy1Y7P7f2HtcBHN2Tvad55xJzShagtQ
bYM7BkPjXIjHpDJbS9DRxQfKJdJZI/06jrIoEJgtGuljV2oeEeXMW3Abj/nUm4WAE3DlOaS3xe9V
2YL2cb8+ndwu1Xv6v8R0DEHkRJbLo+LuF6WfuYlXqIZDmP8c0s5LjNz8IR7ncBYr1izvNr7ZGztY
dA2J7LvIWvyJ9/OgV2HRqqTd3WFlByjv9pAIy/c3unihP1lEkRJP6kw6QiMaQ9ne4vp3frCMRKYW
0FIvwhdiY93tY3J8sLh1pRmu0ZmERaXJ9RtN7vM8qDED5JAr8gfrrJ5skO+JyhV+Fn0h9IK1QQTS
znGxxk5JygFYjp8M2Mrk+DnvggL6C347YuLQWhqgMqPNQEidWi1VPIXugGfNnfgh0Xugy3De+M0B
gIMl088NDr3GPUXWg7tU9/w16OslfCZ9mXcc2Y3fZjwV693mPb2dhPsKJjMa+dAsVyH7BvxxPP6H
sSX6cMTzZEUI4o9Hh1I2IDKF9CuFdS5K4suPAqa4MNE17p/AOvuYFJNADQL78rHEOA+HSeJvrKgV
TCGxRibY5w5sW8rrYIXHFtpN2bkoV+mNGH2UTTSvv11X0M4sfWsKjkEHkVoNZ8eTuI7B98XJbIQt
c1riir9pam7hSbrWUnZ+j7JuC4Igxk7178YJrO3LjZgyHnHsgAug39JauCOTHnHbT+g8PklZPMpp
IjuxDAUP5XipFpJmFx6TenNdia7qXxoJcB6lLJ3RG24iEdQs30/yzphbIvgXvQTlwBosRWN/6hz7
WstOczxg+zpojmcooK3sd0OcyGI2kSFIfPihxmh9sWT4t0MtbuMdK0Z1AQ8vPNzqabcKG/ysI4XY
GTe9stEUFgp2V4Gn4WwameNMGFl04Yb00ERAN27hA1yORlMJ0dBdL3ub0KxGgxP5o/5vZ35dDbfS
gYuOXZUg+aF2/bvL8yqc95qcL2cLbatScrPvi9gY7e/jHzZwB0LKPZofGYI3UnuP8RSofBJVVDel
KeYA3wyIaV3bto7Q648bHdVWuc8PQhDRgsUlfBhP07JNGxQWBiR/iIIyDi96oLb9yh9/OIcm7sLP
/OOtRZrbnyLzET52Yys7SToNUcVf9nm00YJdxeQ/R5KxPrYpm4m8T6UaC64Hf39Nuo8DOyp1IzZH
eGEmaRy7HiF+FQKid6+zZ6nfua4cVWmmn0PZl1CR04F4JZr8hOPSt0qegJ3ulPrLNn4ErhPCvAqf
OJPf5Kp6PzE4SVMqyTS0bHH6oOriKozdznc/71l//tiV7A7XDN1nePgmBgMTcFRQecfhFbDxEnhv
gIoePHk0VUxJzDF5cxd1nINlfCOrPhPNvvVRr81plWHklaKIblFJ1FhmtJFr11TWjZ5clnxeG8Xb
w9wgOGUGiYdqM5GuCZe9N2/fQC2hFrESIAO02RRMkpyWzzBhB1XDetABavOqj1CcO6FraaUUv2lY
xmYWty9rU5wLCIvNkMCwoDoRdok0TlO+irD4Vo2SD9TMQvW1q6nA6fSfimSU2g9jJUfQ91RH67+E
Zq5CTRfixIhP1+esXK/4JPxtExhYAYoJF7pVR5drGxibwPSTzbH+sYhhTplWM/o7TPXjDchVB8le
7Ig0vpFN7Tk0VeBL78wzFefIpSWu9T1M8J5Tkpp7WQnpy0cLi0dliNWa3brxFcChZ4ZaekwxfaGY
vlGe0+pCeR/F7QT7l4vTRNrteL5FAT2N32NQXWxOtYKjXJ0YhtAULzJ7crVDZP9gjPWmijmj25Km
e27cc4GtolJwOB+IAi1WT7bDW+O/ouHBnFTc6ysn9YqbLM3t5l/wA+3ZKJHyX37KM9mB/5ml0ycG
Cbe8InfJ03s2rO2qFLJtJf9Sc/1vAdqE7iIVLiSciFvBrAKpVQf3kC0smQ68PIuWmjm0OGvLH8JM
4DNWXFZRnuVTv3+OM7+KgMjRUQH3K8DVxV75lI0tUOdWmgm44QF+prqZTkGu7VJ6awDVGpmJRhKn
mm6HG/hRApbMr0ozft2xNovcmDHm2wr0fq9XsxB/yMn5lqCFBrm3bfFzSRmGcODf68fUquryPdkA
6W7J8GdSBoxcQOE3AVmUazRH2Mn++/kzULQ21kYyqUnznQqCb98v3pTEMRpQQDNoOU+MzlQ69NOl
SbZtNUx+9VTf5QI9osUzkYo8Ls+gvVpns5BVeJIsLcUuXhfcASbPAq0pc1Pu2oMLaUqNbZuDGBup
Zoq2gYxTWSQMnU8BO6/nvoPX6dj+iMy1Vlzbdv69jYrJf+Cf2FmeJmp0cyt/ZKGS7Utayea+1b0k
1PrPmz1/sj8yVuMXoaPtN96eawPm2O9e22LISbf7Cpd83pbD/zxIo6i5NNJjFQheTvTs7EfavRwb
eFpoiqEPnWgDF9OaI7jqiYgKiRPB9F/StCnG/it1okTr3NyRcLovy69Ba7eSCEHYSJZRnFUirAZl
vZmEpiqTLnM6LdHIQTLDKq55cCx2COD8CmI4oai1kTuXKjJs+Pn8bomR+sNyDInTsqBAA3UG1bnh
uc74lGTd0fGPS00JJilc8Ag6yGIeNf1xVWtp3dch7/lK6ojMyf8QS0TZ7CaMMrliatJ0JGBqMfEA
5q7g6l8I6BbdkKZOobVzDMit/X8Lq9XrDQZY0Z2dLoGwnP9iYp03Xd7RE6FaO0MbKkik8tx8VKkE
KvZcVrK8JLi4q3e61Fekty0UngSm0AtDCVxH0px8nuVP1EDssnYuADEjA9/qM+4o+p/lnKE2bonT
oocc+dCsxi68h+Cd3oCoz1tZOVCxdq6Pdgzh1azjczqGc7gk7tv0oUP2h7+9kNHkcJAW50y4gQJO
X3NisdKCnib7ZHyeGc3sd/9Elb9cDjAXwyQP6LgVaxdkTHasr5koSFDH8jZ5jxEzRVFtjEjCNPDH
QxnYxfhbWlis3KyZ99jl/ZlvvhpkVxKUQ/jHprzDLksayS0nFAMYHs84ZLVWIv2k481HysShQdp3
V/1VIbQXu6EnIpzVIBaGxO5OI3oUVd/3R8SToeMigMNV+4GKTv5P1e3Fi3LKw2bPOq5gA9LYy8f5
k4apqfROZmIt6EnU0BSowQQtYkCfE9tpTr13DZOa6r2TeE5qZ1+ckvLFEehQRVzFc8FtO2pjx7Tl
CVRzHASza8nIj/Z4fx/QB2M/d82N3EEU0cYkvCeEFHLc0MWyqwwTNpg1S84/3uCfwlcOE6gzBMz1
TXLuUUrTurf7JwfwDd6t4LR6Z0od/Vg8jV6A1fK90jbAQchkV9FlqufPpI61Q2lMiyy530TXYSPo
aUA9Aa5jV4vohS8O6TC2cSUFZsZuw1PcYHbHHBnZeS9G6qs4AlYEILV43QodJCZshm9BCOiALOwo
EIQyWVtXh9a4xX9Fnsej18UuXteNaGUGj7Vdnv7LCdwbDkGoMOS7Pg5AASGGYdLeNJMLTWf///Wz
JJC9D7fzpif9wx2+NPOEVbXL97oJegf9aF9KCwCrVO4W10nueOfPrNr9pqTiMgvbGG+dkJXZBzy2
fhAPs7Wfn1wKSIRFyU1oKkLmGkLFFumttELNDI9z6sEoeU64Sf1FCfqaEcvRBnq5yqm9R6PDKMOO
RKFV5C+Z/t93acwzOoU2IdkJPJWas4JyRecpmumjh7k3alsX5tze3MlK3gC8qh6z05rt/vk8psqr
XYr+48CJWS4XQxaRRTe3wUOv09THeGcUxTQeCBc9bA2DoCpxl1vRs4mAn8UgazL5X89zkcR2177w
9l888cr/5742gBiYemOs0C2WYXeSPdoI+dwbpegYHngxkhtn1/5i1zNvsEZIWH5bdrvriXxrety9
W2EJ4dwNs9RDzsYd6AU85p6tFQlM4Ie+b58/j2zf2Xo9XirxL4R66RklUQaGf4dA5LLRJraJHPxY
ppWfBMnY2cWi1Bnh9Crw2x4A8whspyEiToUwtIFu51jZNM5avaWm612c4VuSbN23Z8xF7wkSGQ0y
UMRu40uMhl/vBURrmIviWlhl4PSUpj4YqC5nxIYoMW+QTyDIGaEikwwZJ90vB8plOdJIlLLcRtUc
+IHPezRXWFMSFMSnoEtvjbitlSPIbqSF8TfVlroHHXQbATbhdi3Rr+DZ8pc5fu643eDIV2f5Gzme
FN8ERAzfAfzenTv49UTGyUP3FG8V7Z5l8GPQduR7xerVlZny7jT9DkLKqHv7R+gVxktM6AlAclmB
kfrkQo+db4rloj8VyksNoU05gzec2q9cNrpoa905IQhlpCtxC0kmxArSfZCDVX9YwE5ZAOaumBNh
W//hlAF/X+B0PrWurQcuNqPDA3VSh8138vf0jl/+AFgByDuX9UMeIfwCfPJOjoWKxgFG851tamp4
9wK+SikDubCQUj/wmieh+MIiei20bA+wOHRsA3K6hCZmuFZboQ5sEKx2H2wuqAzj9VeBajr2DLc4
oB3a6UjDARVsETq6o1juSbLz05WWdAIvZtoFc0SQKoi2NgHjP9C3TduGArVZmATWDC8HhVqQ18r0
yOGcdIONMqRL23Qff0gY13VYkwP2gERg+LI5IKPihS3sYHWa8PH3iEcGVStWFA3RV8K8TM/NroKu
MQuXFcXKHdPqmL5bYwk2U2/+AnJl+OrWZHF52NYeIpU9y8smsfvE/NbZiwQhc1zAYZleg3dUb65e
PaedsDhUu4XPUTDlyqndUSdC4RkbSMJH44w12gFFr8IiSBolx8mKJYOAAw6WnZNHqCXL8JOcEzyB
53SDxmD6pWwOEVgZgV6y3MxdkWsCUREFNO0xFHLfWNMz41bPgFFD2rjk7lG+IDUm/AzErZbEFIlf
yZWWA94pWcov1WWkiVzQmRylJunFQ0W473WUn38X2gfXTfJIlatXTrir92n+W456++paSOylFdyw
GRYOTdqqjbFOFV978ffv7rEF/2IXmDwCTE+OE/OEneJxc3Rzx3wqgIbaUyzywbkJAXIqo0z2iD3K
zV8TyoI8nVi+lGRM1Jx9mty1GRKwFQ4rTyPR3R00KuC1DegbYvMK5D023tkm9V5bqeUugU25OhWj
asLpdKMGsJCTz1tNSjPK6tpdKI+su69o3P2sdYY3hip1AV0kW4GoRDJZ/I0XaxrFLJ3sUYy5odet
xrymtCXeI4EGeUeuhLEIju4VQQOEWSE+ykaUElYYId1t3KjC/r2eYXV3CXnktKXY0qesSJm5oAIg
HIClqA40Zp/dpiut5IjTvNJMqF4tpnZQr0+pH416RiETdgTM/rP3ebkFyLqSUvKwB3YQhnA1dCkE
OKn/DfsXFsggCVQYqwvIFNXhI9z//gbI/cepuw6wNrnUkbakRZZsRG+eh+klLSCJjpf0+6Ab+8oG
C9SqET/AXVkn88WX77kcEYVJ52a+GwnrfG/tiWYhXgKaAzxJl1gPspjnRoONzAmRujn3F2m6+kYo
zza3oSvEhzEI0stGjP3tQOhLF/qNBAzYRRtZs8tDxtiA9ELxyAgBTnLUHJ9SvPDL99+gJP3UySQT
9dmvzS30rKI2q8ohq1edGDS4wMowMntwjbUwBVbnghrPUYi3XGBHaeMGS3CKvB6LLD19n6XvbdlD
5RmUko7PvoTrjc0yAyygvg56WByJNohcjRB54GpxQvqI9O153+lS18DIuXK/Q5cqqd0KLLdM72Xj
l8s0QgAdaOal2roLelmvNa3uUxHoUkwpLvrUExV/xCJ0PdoFrzmfE5b+xvwYbe23LfPXteDnqLdh
MCSNTlq0TJlyj3/VSymSNBU+t8V7r73pKmrnVy/3tFcjkNRe6aYidRvQl4qG+50XfJiLn3Csv2jr
rdifKGjF4ywTLSVkFX/iQLrlF+q+2BTgjR2TwYx8L+sLUo3rr0BsRqkRY8C3N1T+gmBdB3e5cnq2
3RpBHPumNXsSkFjE6chW9z+p4eFX5zAgw/8S+2oD0fnG1eglXi1LvJQI10WkqyFIFHExck/8r+Wa
vDJQF2qtHr4/Y3xevQN5+8n+qx41eQjclwqTTbaw4m/CsK5y1n/M8ytAdWHS0Y4tTXprycs42aNx
ZY6HjLaXlBfwUJ1db85Vf7/SvQX2BYtlhZBbYbB/0c9inHLxH/OlNuFRWhRjf/ZvISNFlyrBU7Of
gLop7+Rh1JUu81jkPIN+b80iY5WhF6QzTZbCME3pfgzU+dCEek9J3z3UwEYTerYhwXI74tsBTFgS
zOhWEU734qkpSTnqDqSdfbQ/E4wE+r46Q8IyhJlubJx/tJM02XbhyPazLTsFfaj1p4lPQUFnEavp
qV5LAvfglvkDueQpKqOWT95q0zMpLEl2FmcAP/UEOD1p+hZYL9gMrn6y12QMOyfhCLjLKXxa0AKU
1Bbq6ur1gYkwWE4vyHOW2XUGO8Rpxfr9IURirjXMJ703JxuyUqR10hl1w0EeH/rKWMmw+CVI89NP
jU4hZ8nYtHJxU8Zz83weYTs4hOMrG4DZ0Nh2l2tHFniT/pKScT1Kr05BsW0XwFv8Ep1vv/u3Q/rI
RN7mPpmkBTF7/MFGsRCpP6S9JtsPWcyMHIsuzmUQhkgwjeGCn6RTW0tbdINqyMU0f+cRrvAFfQzo
EocFq+F9w5Pc7R7wUM92FD9wEacxjpMCJec7b8WZR28djiyRkRZmIBQP8QKGQDlIOS8QOINmtule
w6gfd1dztEjfOwCRXODxys+vJCUoKcG1vQSCeT84GurZ5QQYEGsF1ez9mqpEZCNUSkkCZhjVJM0T
rqWmzuL1d2F4zf6pp5QqLY771t2bPd+pMH9ordoZNrE9yRFyAXaInsHH6LcnNly+wYSIZ3RTpWiv
DXASfJ+056+VbeSLpSpeTEQ5YHe8QwMhmYO7bPLSU+jauiYmX1xUYqm7t7IfVuGnEc/21agnBzQu
7LS2iiIuEqrDy8yl5ZlIDiPl6TUdWSuWgUdJYSAi/nWKYdo+ilw87QYWhT2s019PUse+gn0/zRGe
SORaRGE3ShYgxa1SAOdYB8zPIyULojqmTcxPijYs81cY1URCIerJ0i3komsz8Vlw1rdVPXsWKIq5
CCEejFuiDU++N5F4maBE5aGfD4exaSB4tdHWN2A4u0ivkGfGIHIOoTZz6cfNRKowdngi+UNkXxK+
vTcHUc0L+5Q97OUM0SJnz8U7nIxSzA6Y8SE/n6mWKZ3p55qwi/kQU7iCk6k/jcmh3FdQLa7DRJWz
p8Z6qCDbbvSj1/Lsq0ZIfzkcrpoHEOKc9hAFZaO24GG51FmddJYNrVhTP/yLz/lBRbfaY/XQCn0G
M3Fc+nSKyg8U6qNqPFlHrvGmuO+KbCa9ykS5LL8uuW7eWdLsPwuCbJMwzFr0x782QsqKzdbvTF3/
P5QYN+YXjic4Xu7u78GCpr4Pe/7xHd6fWCLRRcB2GKFYpCKMIYQ40bItIjBbVv74xifhtz19DbEH
tqsAEFfl6nCGWxD0SVCGrBwvwLIQvOjEU2hvDzcw5bL7syeeHZyXSwBW1ZdZI+XzIie9ixP8p9eG
bPwvaALCNVkazaxcIEbsQ/0osU7b+W4/R83fisQKGxv35o48N+j6vFYrF0cH7Fh5P8aRPnnxiaI8
utc86XjXA1Qde+eYQpm7raP+zIjFrC7MaTa/zgK9tUbe/eKF5S8aeqi4g1Aaf/tmp+vzdagQW1bM
9+Y6We0u917FAv55fLKORazOXxbSvrOvArbv/OCDqFLH3sBaYaeUJFFo1SKyo9Uj6QCwzKfTo+8J
VvZ2AYJWstQcU6uzgczP27rm7yM6P81nbCuBcU/FqLpfR6ocIkbvyTQWx1pzb5ILZ5Oekfx2hyqw
rcNFy2BDcbTA4QyxOXcaduN+QT1ovzTW7paryLNhT6PXuZbrVcSPPtIIt1AfSmbW3Hq9J7QzAGGg
8VpUP4T3KEeuUNoUxHl68A8bvuOk3gywz4SVQqtICq4G1V7dILSEHLO4Ky1bxABVWgIPtIlaovzU
smcs1dxGxS7z8/Wdyo+xouylCd4rxNwQ9uwhwt2elu7FRdIUjyWKWrnVxGCKstWb71oO/fXMicgV
IHYQ5VwSqTOEmVQFeQLGYHWK8bz50GkL4Tanz6blzZBcOixy+lfAMqZj7SvKUs2gqYRlqVYhvl7U
DSf6OUTNRM6PjasjRDmun6xjWcaSKhJ3qiURgbUrN4Ao9/13nxSmb6Nm9gjFV0aTr6R6m8/uEt0s
w9q3kp+cr6pgygciLpyN7NUZKcRK+1LsIpyBatFR5P7bZ9/W6DoTj/AWMqONoiPXV8eouN7qNKv7
MBbxK3c4oiOg+8zydRhnnWT5FjwuK21bE9XKfKEs5MomuXl8IwEHuG0F66Je3Z0pdofalpEbR9/p
JKaAOjx5Z2lrBEt5WpBEMtQR39iCY4dXBuHBX4te57TtwWXm5pENnptYyagcyPuOTFX0xFDjEt3y
YBen70Y1TIZe92fqcH/A2wzJYTWRttqvFyOLOsqPgowUhVkt1J7ySAn1UIa4VPHXgjirFwdobSWL
iRVWanKpHJNGsioHZK2RO93/d9MYVpYntR217gUiifu55uMJdw1HcLdxf2bzS+oeQ0FGtEOEgDSe
1bbVR7yAnKqOQRrFdZBB2jcyGNwTIrr2e/z23ib+L7EgScoXATKQ9T9iOw8CtDztpR2ZmhDVUtn0
EKOO/jHg6D/P8pRYkyItAouc7IpwdoCjjMTPinXwcepXapynmk5RlHxvxkuug90f7ROfpAt5nkvc
BXUddIvKv42ApzxHG38fb2MrNdxc93/+bxL/VRIJ5V/nHPDnGf52vBPzX0c9WYdtPRx+io6Ueiuo
UFOO9hbCEYoT7GtYKJaV2AKT5dFe/HurGXP1W/rCicvfL5TqtFT71/6dstMdYkP1+gPVWJem/1Lx
ATZBbWIv13SmMgBs2c2bAMIxAf3tuTWuvktuyRkmJyCr647hrVeeOmiUoQAfR5j2is7FNrEpVvz7
TOgFdybWWuxen3k/z904KbBvAAnEzr9EQdB434WP/cGdSZ24CaB5UXL7PpiUeSvJ2qWK7m4VjQ+U
pjaleVBaQCc0S0JnqDdSM/pYmZ0dRI+izkP+PlkZaX3XocGOq/PWy6h+cmW3iAyjuoeR+SduQ/Lh
V3LROSLUD0fqQVm7UGkHidbkxlZDcKZNQbCOh7zHYH94/piPK3yPGG4k40bmHpxy2QWV+Xuss+lV
lBFTP5WOJgC+i2ohZxhnKifj9etSZH03JKhZokVGg0eaTFK4WHgexCAin8csgyNIEJRMZKcNJRBs
Gmy4je4qOu/KaTddhEU+xjUMXpLSP8Ks+09U/sFCO85lN9t0SNhfNWjVnNcwDqu/m8IcnrhQ93rT
hjg1wibtoOEJxyBrBbiYVccHgpWJOEVFwk2Yot1F2jv/MNgDEo52KvblbZU2y0DeGn7IHSNRUz4Z
RDKxLh4lAaXzK5GsEHxNY6Pr35Wjocxfgc5zxxKg4RRrJJSA6Gv0q461VOwwVibr+frvEIjboCu1
qiGU7M2lmo1IHtwo9eRAIlJSeSZQnTu8sR3UbrO2vrggIolUJMxfSCZ4RwBOx9Q1a1I1Qzjv8F3v
Nxn+O3xyq2UJ21wmb7h5AXIJnXOOzhmi3wsnUXx+ZCIE6qiYRJ61Avbop3T0OyUeJ8peFNeTuuUu
s2OOYLkPzmRgmOGg2moXf7HsTVZ0V1GTAvjdbTYFSsJWM5HQLFMsTrwwpOqcJTiS7nV8kidqtqiN
B//xjkOofhT2QtuHfNcJzg/dw8CXnXzNnEcyr1x/OMihgvggeGnEgdSOGMaYCfHwoujqLRSwFzxD
WF1XrpNHzzEQTROjPNCjZ5OHMbfP9P3HzK/ivzIYKV+oq0HKyru0RtD63Sb6r98QvxUVXIz448nk
GenJViwMFU8YO1iKn1jcnfpAIV/tFU19Xu1qrryL/9w+WwU+7jqehXzD12GNgqrYM42YmTkF+Erp
w/KL5n6NZcil8mLmg+yGJTaUo5WMdK9/t7gnfEaHOf++EIRYyFNsmZN/FFNYi2AGOx51vnNtxKcS
CFgzyY1OIIRrFMxZq3FI24csR2TXQ0hzqxznXh+e56wbcxCPVxpEPg+LUsccwOJLYVjX8wq9iOJv
3zxEZZncgyY7iUtwfzKT0IC+hy7iUHIp9ho/n7h4HmEaqW7RguhzL+ArqnHgLCej6OimutOvJBr6
BFtftHYBHqzkywXvGzZcKs/aJL4dGC7LO0BIa1UFCKvdjwgb8lFahOzz4uk5iUBjEfhwpYzL08iB
C56e7qPg1877WT8ja61XqtAZiIKNKwtF67SrSaXZgIlB2vWQ4OVFU5grp6MZuSvi0I9YT3F2G5cv
8lJ0zYXBrMbQyAhba3iC0ht25kbxWWog/mFsjBr/9eo9a9WW8zl6m6y4nEnJ0IzM9HNkDzsEQkBu
RwsNnvwUODBdbQiXZ8OKeH8vhVp/x4PNBoCFAQqYnVIThUaQdQjLCLuBKspitjXGTuExMnj8J1uX
xxtlSSLvYE4YPAUDHAb373Z4Ed2Ow2E50PSG2wBFKfl5bN7FjG7Grq0jXRUJebQtDYXBT3I09f5k
Wf8L/jbkvP+gXBjj1jCW6dnbzhQmazhGALiE430H7tRMaovPF7POsBM8XKXgn5IKYCsrR7eVGrQr
2YKhXDIBdRQigTKluM/MYwsTnmyRP07kflhgzLa/TTkPtAz/5fqNwBf7nlCNXyhQ1li3AQJIFMG4
+BG8h0vwsPv7WIHTTlTHppjzAKmauHCnOC+WmF2tDlehY6crmoCJpCIV3yppsRaEwcui8y3+ZVZN
4txxG551u+4Q+ZaywKgk6AgnotQr7VMBG/TUvp95k0CLp9i+ieHPcdjv9vFhTqHx1ti5lqalO+/a
hia//tRxX41v0qor12xu2E1g12EUETJONeSC2Kv4Vu3gmtlOn5HTbANEQL1TvL9W5XOf4KKU/+8E
nuXg2G1lVJNlLtS9guWarJoGUVmfVhiDktAIXkiiDhS3ZV19oVRLY5K5Pq/Y9xmWnZdmC67JVKGF
a7LF0RkrhN0opFoMgPY1J8dnq2P3graGPQsuQwRZ7AV0VzmCwDNTep5kNIM6Xaisg1Hsw852/IWC
VH1gpKZpT2rKHm5XGquXzK8fRoDI5yBmpf1elfDUm5YlpEZ8fFFVkX2S7rGcwD55lODUPdzM4gsx
xPKS1arCfzMp7qRLOBaZVYbbXMbyWrhPJtCmhmtGhOoU6G6kLSCRdrc4uE0ztro8PqpPiziRGf0p
lwGKfg2+u8egb+X1CjS2ES1zA/m5yQ6Anbll//WV6SheTQvw6TB337nMjknaBQUWkMRN+QY1gEZG
5+j1V00J06m8TA1em0W5ar5pDOz1GHwTyJ85HmZ1kGXBtI4INkoaFkabvnWnd70pfKL4+vfDXeWp
xfhXu0w/FFAhPn+PzMUHkbuBGjJa+2aGVNUYZAbLrpeSdXe+8obq7O3Mj6yvZEVoWNbgf3f8CBUy
ZQsNvFaDf2pXwIdke4wZgchZJoGNpjW8cB+ghJrADzz5lo/0w4ot4efK/J2RzLN8vLnUzRvmh9rs
kGblofdiAB4suF5EfUGrqX1XG7NlI8HpcyYRzxjV4N2D9Oa6A8fZ+s82UEcMVpq1ipEfFQ4EUY95
AOvtZVoPDpAuQAQdbAbUULNzfEmpzGzD/ptzN/fHAioevG9zb5ickmtPvmWoSHYYQdp7TaQomYBr
pKUJJMjF2eXu5ZkwED4zyNzYCU8xCl391EwQmwuzPQgrsirvDaMrvAxfmmHesrSQywG5SCHkqpur
0ubgC2DwqD5rosiV5Zfsrbc7wtaYrRH/rNfKFy4KuxGmG2W2bdI12jKXIntipxNX4VAxswbtmtnp
/wCHHtphOwaMJqgQZfgfOzxAiYuTwdFEnqD4vW9rkxY8yujpx9WgH4ENEQr2DzRiTSmcMjpvrgx2
wWc5MSM51bieTWDx/ChfEP7/WaPN4hpxiMW2N7h+u4lI6pMuxcObvVcAjJDcn7YE+i31D391Sjg5
b8Tw62UjrvYm1lbce8jlfkAcyhJzuanu3lJEHlU38szVU378injqxYo4+WP3cDq1/M222VGIlK/I
B8dO5HV0ct0mdKgZ3tag5O+ula+ARCnMdVGkhwy3AC9NxgjlASSdx9nD3JM+ISl3zK9FDyNOaij2
ER91NjgnaAD4R0BVQBvOs3UfF8lAFATOlNeSm5+OC5DiSUvB9Lx2ZRBEuwzLzlHlK/p/TOaAjZQy
7p7ISX0Ef/XcmYt5XcvcQsOZ481F+I41czW+9bG0bJr4VBX1OJs6ufg+2AEkba7/TbkSDQEOV6FT
KGmepj9ADo00zIcuBgUGEpD+4GiQ6hpkQU9SbBZsUdA8mpOWH5y2Z3nm5wOweutWXOVf9H0JHazf
LLKrjitqDNmwAuiFfABn52uj8xER6iD1pqLQ6FrlV3t0ZcDOlaodwEfQx2F3JpL1csMZSfruAkdK
VPH2bLiWZVR6K7MeGo4boSWt/IS6hQxTi+l+zSFkOiJh1xnMKyFiEJatLHZX7EdC7YSZ0LIJltqi
gor4h4lzoQeXYYA60s21QtePiRFoJNrW7d2YLqmcdDX4xjYP8Rplt+G/c3Ip7ud27Sm6xjlXSAMp
SB6jYWtIiZ/vFO0zm8anxTLdjQ5yhO4W1pahhonGJdTBiyKCWNVxHy2hLzRRXxkJky9yh8XGsYCO
GkJ98B8F16DR62vvmgaq66FcCEwWvk/SobX2qz54fHpuKBH54EkuJzFL+vcN63cf0USR1qxMbJVv
t+aG6+qivKXNmywkoyV6tsgLvtOfvN56GwMs+4QIBm3sLYA/hx6QrjosAF3QHjPyVAciIPR4fhBs
D5g7a3Paq3k2VP5NS+U8MMXSxTJrEBbnfZvAF2mXNeTBZvwWzR1AkFN1tYXlXorM+kl0J78K+cAF
dEAUy5UVHfyV7ClcGl6fuPcvmB1Sq/7kLueEhMsQJ7rh4FaXmHFKXySQPOxkLRZ0vbcH6RDq7LJQ
hXnN/DWI7p9jlEBLIoDQe4G1nc4+T5jWJj2lwcJjAKjn0iOWMjjHXciz6S0oY1Y0stf5mv4VoVsd
8+RHxIAigSEepxSCASI2AkXWm6aPIRkLv8ZyDKaz5wIh2cO1D7GVkX8ymwZlROMSY3ClLyXqPOY3
XVDUgkT5CmYeopVcIL6sJgNXJE8f7m+HcmJIoUWfCozq1MzQ+tlCAhDTzn06qAe4e3gPD1Oe1sPS
y1yC62+AuogDbobinlclKsWrmPX/nSy1Mm6jTGXr2zCFSweskrmUr6m/yHH9G8x6mPospfzJTbX2
OQ10P78zJgUd1qMv/PValD3VlQ8GnBWyTKh+bB8xue51KpkSdY8RmVUANSfC/f9d5huBaLCoKOa2
tNBFsA6pgczICaKEjug9w5swJCyTpcyBmuN7iAJ6rcJICiMJ2edxAr4KZj7HileeCkCW2xetg6QN
OvbtoD7s5WQUQVgDyhxVqeX2J02oDa0FiDMWeYqsdXvkq1WkmLGyqhwnekyvtHOd/5BefBm9lbbH
qk/8HEd0yKlNss3mmRksyZVm+C6HuWxN1n7VspzaC7umtNVWD0nBS1C3MsYyYiTzeOIeLxBN35nG
Frf36tZx7wKkwR2O6GneH0oAh0sfnWBlJmX3rmaVHYQoif0MI8HwaRlpLUBpPCv7FsFZke2HQiUu
PJojAH1ltYx2zmyVXvNgELx3n/tKRQDg/4cIj+XZ2jx4KcvCu4EZi00kZFAmUZhjLwrEyzrXsQWb
a5HcQ5BtgO7J7MmuAzsY9upYwMmukQYGVQVWwXskaRlGNAN3nxK1FQzgnr/6tQc3GSJgozvCIFTZ
UFgCVwf4E26F/B/OQeACR2QqtUdcGqYqWPPU44qxTZ/ayFS/Y1wv1fGbQaPHwRqhsdIsZ2hKDxPV
B4nrE/2+sy3iygUQWXzkMKiQx6eXlDqADdSUSTdn3vhmpIj5yS8VeBPdAFBbyN/fRTivjLw7ubtg
fZBrOKZDzSkBogK5XwXOuR5WMBidrwc6dEmoYoYj/HReyBKYH25wujuzdaDXcMzr8yZd/AcHj/5F
hJy92CE1OILiG3Liz2IKogF3OGyXd9J3wmdukFE72tIvImLURKV8TJvu7+kXOLPQt/t130ydFnvT
o6PpqsyHSdU8TsDbQ8lh8Vc6o6nUtcKnHcfg5p/w0MAPqu0d+ovRbqgvv5cbYJUa07Eo9jn53tCa
3tTJNDTPGP9eomjL2dyp84Segb31MM7/v3LyOdRA0BPwoB/3wilxjlEMI0jA7ERwSa+946LxrTw1
KCmUdZtZ4sDJQV96IT6pba91fjrbEbYeWnpmTZIzerkJU8sVDqFrsblKZVuum4n3iNdSWBei4eZt
If/0DGh+fd+eW9bpm1TZHkAbpSbE5oJbFLkaJ7fUj8OoLbj549L2W3bAu0Zh7qvOAOCzRn5EL++q
2iqw9hpgGUJnATJsBuh04vSg00p/nwGQxGMd6I0/9z3NUf/mfWBy+5e2KfSzjNzMbHQpXZw+JnwZ
DLDKRCbIhxt1GtwOgLgkyB3CsH2bqxH1dMjrrPaw9pN5ga9c8A8w82fnMZf3WciwgHs8bP38N+no
6QKCQyEidMo5ImpZTtwhGf70/pHNRH4yLMDCOh/HjNFuyC5EbQor/FLl8+Z2cXRDFlkD6Woy1jCj
QF6Qpt/PwIhuMDQgOLYDEZ+UwrA3fLX2DXzJrhSHvuHlwy0hIoJAjVf2KzLF6HXEbpd+xm7Gp7HY
jcBO5bI84Dq1o+Rs+wwNZgNvGVp/toGu29sMmvTdEWoVgcMzuktsRoF00sZugwwS996QFiwuRBbr
U/hAcm1POC0APitkAO3mh4UjFFw2AcqJ05Q/cazUJdvCCOQUFkoxMAc2gX/Cyk9WwLjE8/tLbgum
q9FAwtilfcfpC4UoiUNOiqo+IC2bHfOg7BQI6Cs8cMQtOCJ20Jmgn5ahGX2pRjk7gnqPcsbSBevh
ifiIJ1Bw5GR+XBHqFYgVVeiclwGMLHWG4p2P5liVPhN0v8h347fHFVf3xCVtRoh1S5X0aza523AB
K9lvIfofIcik6fnyo5j5I7VdhLwzeXfV+4V6Yza5vBlyEkuu6BguDnaBvZTXhSSXaOlf6wqChTxF
or/ZQ6NLgx2D7o4uY2P2znEfrA8nA5d3bRqvbLJgAX8Yd7kKlSRiNqbWcvzRsYT6xHaGerJ5bds7
X5Mn8CocwKy90GvTHxxFRuunGwg2M/ewaDZLtx1smuUaH+ycf5v+fQZw/CUeY+hnCiF/2qbpf4rt
SKQX1olxshzr0vvfkGsyr/5SUTGPnMkkj2aTMQOJuzEtLmCXdwIuYOsxNH5zN/uCmAbsR9G75BWU
06RuqnA7QH2Algec2Z5GNSH59H23+hmiCOT0jqNrI+4Ao/hfIJKyaGfTYFKt/Hh7orBb3Ob2npi+
Pvl9CLgyKSpwWdS21fP4gXBQA4jjGWAMgXIB4+ChsdOr5faDVCb/TSOKPpPfia5826YHx6XZh2jQ
leocucG75MTZnUKuK0ssJHpGv97KMsRtBH2vf7lB6FKmLP5MCKoBvmivgbC9xP8E5eYqyW02hCBi
G3sTNn6WOyOvPMCkiutAs/BB22C9DsKSQnVmEh7EFP03uQib7CL3QmL7xU6rFJBoT4kVE3FtJN0E
FCxTQCwFx5rlM9YB+CiMNC9m+ntEs+oT7SriPJ5Lxah2SIxwJ1ohidZYpYhVVE2plCGX0+ixpgYR
YIz5U7H/c43htr4ayT0pvgskuNDb76k4A2T5ZOSiAdMTBj1U4CLllmzd9yNCLj0ALsR6b2Ep4WjW
72nZKjYn5our8HTKcD8lCcr/e0efhp0S5WEoVHEu4LlKqyJ6A+UOkGPV0m0so3K5s/1nhDJ2OnUS
Uwvho+jl9NDyA7dBLGebFHWeiAChYWQtb3+u69RjuEO6tYp3XN7bb84P6D17/avokMJJMlkSd/NX
M536mezwG/wlTHgyr15JLz+Qc+tfF91CpSM9KrKhWmyIw67APNADKqTAFzBMMyoe+K8M9hZodRGs
NxHTLefnxIghEJETugIsc54qVkR9YL1pCEkqtDSCCbjuy5G9bjwpCsWLPtkdaffyl3CXaT0SdNUD
ewK0J61xT9j5aHCZuyA55mlLCxXciYYb0ZLTeU9tFju7z/koNd4tk9XaeLzNLd6zIpJdR8DQC1jq
Z7FY+zaNu//LPYpBWgEcwQNRzBXYIgpU5o4eaNTpEaIWBn4KCi7nsuc5V9+ihP0KqIEue6zSuONg
psD+5HwIAqCeCfGF2YOqGyvmvyA6Q9u5e/trkGCMx3grQR8wNBm5qlKfDbbDxirsOibGH1psT0Ny
S6DiyIYrXl+ls8TBf5AnHX6b8AIItuKPclL+zq33Ib4LG01ANtf+H8QYyMnkvt5ceLsexmo0l33K
hII4L8wMtBHJ70Gt5az79I9oLCxBJ1pOM2VEEYr9ox7hqXi9mdr1PE8eOMOqpLrSkaCv12NJa9N3
vCTkXPinXBWdTFBWDVl5xt6wQjPNgpQERkbZx9gfKfTQBjfk/PEZHBM3j6OwSzT8KYOELoYo85TU
6r2C8xIsfpEeCqeamL4wKGvVA+Pv8oWZKCfn6WPQkEDA5NaA08VB0gSID1zPt8rQVyujv0tHbrvC
1r1ZjeW40zY4gmcEqzx+1Y1y9WeSbtDkEg5A9BYWBub8SQalit7ETJq0wbxb8tT1VsAp2rIwSpuk
Y5qVZ8SzTd3WaFNh6quqndAkozDGvVFg+m8Y/rlrh6NOASDDzNTsOEg0qFolXwbsm40N5U7+QHZO
Qqe8CV6bkXzDwelnQrZmCEQixQ8V1ScNbhzt1xk4Fe6ke57BMIJoFRvGG2zetMfCMGSom4cdTN2C
Dw2oJer6X0Iw8JmsxGdz/Bh4hZM/8zoxQ0F50pymqhHt6tSV4fYmRR+CQGzJ1Q4CKPBWoJRglCPz
/jGF7/TUMgmmZ7ohBLhrRLIAdwo4u1efQiAH8s7TiPw6XzkVttFZs4AjjMeJF66eXjuBT71fOkeS
I4DGqvIPbRtS/czwNzbSQfG40jRKAZcimybOfKdtVEIc3q7u3ejbtisapPK+jlT+9bkpJQf5K/PB
FlwF1YW5uzpDjxqk4UXuK8ZnemBDf+JO1FhM7y44hA25iRsDDNqsucIc2zWEp2bL45QozeNR9AsZ
1hBgD1ely4pxri4hSgHtpmupxYtF9X+e924D4brvCKkn6uixzy6wwf0mSpqDQwXPqiDxpDa3xpW0
HNYyOoZ/fuPhjMsulWSiADEvrye2Ahbb612k7KkmgiwjOg9oN3XIYhEvw40CdVGs6tRhXiFRnRU+
Fs8NdXOcb4ZW/3kSkD+B+zl08XdZqoeY6A0cbU4uL8e6RauEJksVX4rrCORP1sTEQmEmQJNRbjSs
K8dJbHIs8iny4I0yU5PbYxtDB/k5sAnPHVzh+P/inWisVHbXcJJPHiZmn4G0w8spiFrC+UZUvTPs
wZZBHBCQe5jxYk4v+Ro9OClhj/elHpPc9a/x8Ng0G8U8sr4iSCdzGCsRI+UDYSMdDxadtGj1jToy
YpmezK6WKjjmajFPk1j19yv8zBLXZ3+mNDfYqiGQePui1GEL5U2bFJzff/mYyh/3BitG4jaclL2Z
9D3jSf+p0Km8lPgYMBwkd4ZvIHh+OnMWsNHDT5D+5hE7exlVsOGF4q2O+QbytpxlF9F83wPKa6NM
AWsMGIlmn5Qvc9SkClDM79jx/TSwHSGbTZYpk1mrOiz0H6hHjjpH43KDP6pi9wS34iRqaiunQ4cx
TuD2mENRViTKXDSjK7vdRuFXld8cYZy72ogDBxJLAMfcDF9t7PMfwFpHzel8rCG4jhvuG3OhTiAv
ogWw+XMBlfoZVxio0kS7ugogzB0XwZ+spoPzBtMoyWaFlYdFrYmFuYrWAWUHwL4cN/7WctDN6ayk
BXnjJaxN6SJ1X4XvUkDRtgF9MF5WWu9e0txEcNovBHWPPaj4KRQyPvNGJe43qfhMEPJ01IIHEkLl
x9ZoLZODb1AJLtm+zzm45j6FNZUPcy7W3bbqJb3Kv8h27ET5FRgrPQ+wCWY7qp1m2bB1AyuCcsJI
XyRx14itPljbnY983hGkGP/zsi0Y9SwapWsCAAN8u930IsVksCn39foTuubeK+lWZ4vRyWrFeEhD
T4XuhcRjtuDQQXiQT4i14d34Cd6RnZ5HgCAK6evppeaF/bN3P5UIxaYkBm2mLslemr0pCYIG00ZH
vNTZ7CREUhlR1unhvkKKBE6Hz08K6gwcsRN6kC6ZMs5KuIZ4/E+xlxz9FU8SPjpGwqdIlNzgd/LI
pMT3zzjtuhOyxhvZAVQGf5L7OC7yieGp/3YC9w8ZysNGJlygry3PxRzPCSa3jSiSvBok3ne0DTXK
APfpmeRkyYhiYTUJVr3G/UJwWls62ErXj9j0c/oMXU767y6OfXiGC8+0C3HRRwa2IeZTjGCPo32T
LC4o06BbGbFe0BltQxCIK5UQMzinnyqDbj64NDCXdFwwXh5GrdFVKvZG5ZG8I6OVhhb5H8nIAU8s
1r7tKRM8n+Yxv8CJwRKeZabS9Ei+AEpytd4AlI2QBHp4FyM+xHvmIP7cAfUmetTMV77HY4ttuPEC
bglsSXNoR8WMsDnhFaJdA14UQQkdwA4Veydv9FNsJglbWNUsk+BmtzR4pacwq/wkyExxsagavBr5
LN7M+FwrPav2QjaQwvHr5h5hKr6Uk68db6r54Ym/lMEGbo8e/ee9LtlU3m1OYgp+xrVObSehME1v
AOqdS4ZX2N8P9D9zKZmkw3CRRXtlJ6jLxWa0d983uTBGlyY+///pSkbkRTD0vxplwW63xhP6VMU4
cbKYQjK2v3da1JHpnh9y8nUWmS3h9DARMsa/w/FTs67kI/NrDgb0zpuEmaHuZYUHJx+XTWmGA/12
vhpFgkdcIr0um7oHRlRSkz2euBMICBrrP8pEYS/nyBPGuaApkfSobP9cXBvo4LEdkmpFbc+1amdm
tzk9fkSHGy7ogxFh9DVjOFPYIKbtCVprE7FMRko48AtutsImt68r0SpKQiyqrWnKtGRYWsW/ptTM
IjW20ZQK0ly0MDDuI6RAFtLsv3KC9/sBY9G8k6i7y3a3hTBPSNOKp6JrByKr66woB6jAyqBil5qF
i5LpbwjuQ4TvdGodCeS8B+f4I3jgv9tstecyjSk0/9O+ORvviJXhQMC9LsHgiHUUrsW0/4U+yaiI
w7rgb3VyS6WpYrqiEXK89D264FqVhUeY+/V3CyzdTGbHVHHfTbM31lcnTWOlOVImusUMbHVJxaf7
/62RS7mOuTzapBy2PwjIyYseMm+a8gSK51xbfKg7HJsLyZv4gEpd9coKuieW6GNx22lF8n2ObWti
oxsig+LBgJojjWzyQEc2DjEUn7bfkarJyXqPunq+R7cUWqsoEsl/QI/TMpVTKVhJNSKApYJSZJ66
XdE+qxjkLWBCBRiYyF6YQjXi2P60Uy4Xk92YnWk6sbs1npflJ7oxHH2kqigbTayCG7m6DedRGxQu
nh3PYKw6W1oq9JiIT/DdsKHAy2Dgji9NPV34cPXvmRs5ddahEtd/yCULQblKp89YAgDus75W5/QS
VdvW1VYbSFUO8uFgwLX1iPbTrF09q85DifkcbSNzK+Q7FTVMfiw+Z7xtjoqcHLp7WeIgBy1yFeza
9t5SOVGgMtdSkdVVpDfLzVLzRoggXYt2+mQ3B3gLAje9lSYVXVLWAD5d1gmU1ZSxU1f2unr8SFai
8Lh4d9PFvzHT3qbkT14nyrRD2llB+7L8psxBTLryc9Buze7SCcNMQZ9vgTsc0DlCa93sSEWwXUc/
LdhPue6A5DanyjE+surv6Dr/MxXn+qSr63pU0D8N5nrtghWcm/kZlEIxmhKQgcESXw/66s1R8DeW
b1i/tua4aGnsqw1bqgH+4sY4qtlMtMh4SAqIvUwtnvVO0dDoIC7XmLXWU1pGQ74WSG0fooKfbPpl
vn0DOHi66AxAIEqawPCxMVJb62cjoIAw5aq4dU6+fxoxV1OuE66gUMKwS27V+8YewMVY7bImg+4o
tZtBDoh9X9vIwWxVdUm8kRflSvzdS5Zja21+Vx/NrfPQZhzKU88UXFolamzoLBi5xOb9cV5pz+91
An9ANMlQqOGaJ9wMc6oFLhutfvuoqtKPsDl/Ef8czraMZVTeNj7/OZTXtM7G6EM940xb9FxQSXEP
QLZFx6MwiGlPiHLXjJRIpJ+n4EO7g6kuNtQj8fIELlZy2JsnIP7G+tlQevgTe/Vt0UUfj8L7OjgP
xqIo2+BVmLqsLEDjgyqAGUcEqSPo3fvg2Ks6ZdTflo3EzKM+kVIm/OXg0I3Ve+CbKXQ9Fug4yJgF
/7vSyLbquCofrV1nfj0nXX40aZyqQukkgrTnPrb4iVCMZ8web3UxIqY5VVaqSiZ3Tzgdsi/PPb9d
xtKuuNNpE3fs58MLhCaKNuP1zIklJmr5PgSUOJQvlIRtEceI/cNM2CkM3TMr/YIfBaT4O0q1Cryn
8iYCaTq9eU1XlYophl4wj9lg3mINc6nvDoo5eYY7BqfIOFEiVaigWFOGHYGozrE+k7X5LZqvNoIY
K5hUx42TUR53cOgy3+tJ8vCa33YEI6fDs9KC6THc38eG2n1V+b6pZUYZ6P/N97I0OUeLIBBOkbbI
qmPE+cZo6iFPoC/PkRwm8jboHGKjS26pjlsJDRiCqp45VAXtGEEVlf0EbAldGYUEV2khIknIF5SZ
mxEyNX78Rd5YGeydsllEpcClDo8XCVIZGoffEI9viq6MxLr7nxyVJ+Q3nkBPXO62q929ttghyceX
5ko9SCxCd6gJdZwzWYYKcdkvcV0AEP2UtFa3B7hJ2MRjB6W8phSqyjQ/xjlUoU9u62fF4n6QNZeR
ZpG+cSjbS56xDNp63gCh0PBwtSYfXIPtSrM+k5G6D3ebYFK1+aHGvnyndKEIMtbvUtZeYrgobF63
fODi3l6qIsWXFOQJ5fOQ8LXigpzE2z5RlkIRdoaoJPUtFyXvWV+rs4TFGU33lJmY/ZLvjnmzCnDP
C4MTvIG/TjZFy8sUTtfq3WoqyYPz4JtdJl/zWmXt9dK9BHXei9YImNszpkEyzx2wI84h76FOPeJ4
lLrcatl+tspo/QAAJi3hnAh+pf+9Mjbn0Mr5eHDqTIKgn1uf86e+yBisEKTrOgPf1l7ufSDsRajf
/adtvN1LfLzriPvoReaNI+ALOigkGzgvzm6Z1tXDyCfYRnzvrlG3QYjPoB3Os5Pii6GZvGirT7Ot
nGQaxpFgPcuTYJc+Nti1qSub37nr5qMd3jQdSlvUhsSQkY3IulFjALCfvzwifU0AJOmij32tiaKk
sSh3jDxP+E9SVXdy4QcuKD2gor1w65FUnPpxneefQomp4TdpjoG28OJ/B0jx0wclxXdzzKPIPEHR
1PBnJ+6OndFuXss8NzrySZ64ZYc00WqVA5zl8IE7cXru5RqyxQGMv+A70TjU5SmgXHWo2d5UXqkH
QK22iFonafGUL7vxLW26DOYnqqYCyN3Qkb3/eCOp3hfwusnmBW91UtI6IPhM6dd1ZyqsHlTtfiUw
FSycgH+5ql1p12zlmC02oaGt/FV2E/fwomnsPOLz4prpuR2gGxQkKGgEf9opFWssXfvdQrIGDPQV
18GYJE2GoUgAELU/gcKszQwi910vmiXJTElMHJuuM7igXMgXMHbuazRW3QZjMk+LaAmASVh8VBLs
aJL0ni/etnweBZ0fotOPG0U1H16uHbfF5xminrCF/+yHDinCH5QX9gpUBfqajrDQk5mYWDXeXSpH
PjRlfrhPneDb5On7ipXL64NrRmG6Zl1aydXfkbcBzCw2aKnlUMBGjbYDk47VjT5m50DvkjreusFE
8mF6bWIToU50UokqHZgNe0l2lGH2P48ilMaWAgiQlkWhmRqnLY58SAZ/p/2PK1m727TgeMGXEqam
+oMEcAso8sa4TcoCUUhBje8pWVsQnuJI67KCehnHw3jvRqZc4PyPfUqTWjYaxFxI5q3kxxgjMY3y
hMAMfrWU/touPJY16YWV8G/H+CIEJ5vpT19+5lOTO8FbNkZVKMPimVCNyjCKPwikP87P2Dl6LHk7
dJ9b0AGWm2gaIfGEPdg2B9YTnzmMg4wXQ946Zln2LCwtPAlONRlPR+m2T/NQ66k5fLLve7yp18za
tfMRzSHL+WTSTduT7kNj0T84cKh1tcSzVwGHMDZZONYNM1eJ93rVc65J1uXP4w4m7eN/b95iHs4Z
jsvxwuMUUQvjaVFOfFb/zNCv79MyAEnP+aQIz5DR/MSJfMrCVBlNVmKylhG/Z/9tROhYfOMVcWAc
zhgtF6OVd26xjM9AFjwxyYM0tZsBEFEO4UUBboB/fuOQsWr2+4sI+wZvCQlpozDH/aa49cX2iBJ+
I/TUbCEOGJ8SVEsXS4eA2DVeEVaIBI7AtHtseTVW9lgzsodJvHvCkOvCe6OXOx/2QjWzcwrHPKvK
SjmpL7LgMA2AkkZ2rfm57zR6uMSTSE5IHxnEF3A+uZdv8XuCTqJR/Ib4aMTIwH3QcGHv0/x9g1at
O6AEQfANgRx/9h9lybqigRb5e3oi4xjQVenX5vu+6OEW6gmnLxW0jl/w99W/zRDBXzUEq7qpw1JI
9F6AWfOsWn7uhQAR3L7Xqro7YDJKom8yC3Wumh9TjlC4HYVyI6KUZKDv0LwaS2UG2jbH7CAi3ZNB
FZdSj1EIvsFYHRqPYEHTsNVYJyKs9eHb42MlNmFBNR64YGxMRRvtYTUnLxEyMhhGyEF2dvDGtIFr
Q9Opu25KsdugYwTIaZB/uEdOj2wEYnojKNTUZ88MyGO4ijN+QcGY6LTRzTcsfJddUQhIRZupprBx
WL2LL28QtYzcsQk7096MkFXrmsaVRgVr56N7OzmSZsnOizgLtZyEAW/Wbg0JDnzGzeO8AmE+l8Xf
yn6k4B1GSjTk+gA+BsKuY5PaUuTyPDkaC29EdKUkrYhMJ90nwjDPZbC0xZdxBeO2/SOD028LLjU7
2H4fHKE90H/GaRUfceuCwpFEL/A743eBAWgYuEmP4Uno6lQkhCnGgeOC5EEvNeS1lgQg1oBrYe46
r4F6ImBrpsa7w5Z1tq+KRmIT3wL+jjEjN8k/HBAqqUXVSOigbZONywZ2y3a22xCntzENbwBTH+WW
6db5xy9LQT5chAFGAGL/kbbtsTulfjku4Re96c/52Y++opEFcINU/x1NXxSQBSEzqCmsTIlIwKRe
WUX+HJ0q37QAzI+AFTRyjTpNntsywk0Ak5pc8bkebSngqps3ZkHSUHbhstrt/0SsKk5yuLt22R7S
jtDN5nHZvX5q1hJWG40RaUCXP9FqA7AR0Si1m1/GD4VCz6HYdyvckBhBm6mTHHKAuFKHBndPLpnA
smOjy6YP4OcsmHVYBujgjydiIkvCdZFCZHVp14rdLN7GWzrFVX11C2Vmifqhr1QUqCYdqquOQpoj
pmwcRSF5YGpL5HIO+kWjLZLMak72mEQF8+hiJ1IZrvulVoxHfBw8v9BL3BeHPoLzZRzIe4lPERtW
VtwT7DiUGMwB+C3PXln72hZeepA3Ko5zpnrk+FXDUNkloOYQvKk3gBa1FkVxt+06YhDcAGoAz2dg
OEOZb5a8Z9FrBh3MASLGWqAUXcL2rjoWsp0x4+2z0Lw/9pbxOYKWn5/teaSwKvEXRQHAwJ42Eyar
lwzLalNtnN/XkFaeVNjSqVSVYXfuPFhXqiLHdox0kcT9X57280ARRHfXJkosLj0nyl//fwet8gyW
RgTi7ow85s5g0bzjwgXXkwQTdcjYtY3B1mKy5AAr1Do4Y2laLolexYiACj0sqLUQ+/osTCrBUhTt
d7OD+QYEafJTZdkOfSAVvgEWOspC2zlpK7FFy7OsmRkDsCF9HYc6iMV/cJWrKLamugrTJitMQSZu
H+pQgY+RkZBZW8i91A6fWIqdaC9vC5kQcJP2TAnudw2i0jRbbMLFESR5A1IP5Bp7Yt1WMRAkvl5c
VzdJGqh3DB/rybLvnYM02woqp6ty5HWdX0WBi3pJcLLaHP6wxq6yuMwXFSSgUzT0R/NG+6XSPbcC
URNDfla42eUE85+icobs7fVa9NMyhOs1d1PrrAfePoOCkjoR0r7kHwgbH0CBTXrSCy3gvx9zdDe+
7Fx+rSVd+8Nz+1GjVBx9xMIO2CsJXsurFGnaddxwv7UCe56vKoVTlCKwz4qbNXYPhNx1y1cQxKeW
XTTN+lUlSXkBWjdQ0j9RFDBd/JVsf5iwf767Gs1TZ/ZW8pmj7Jc2bmTgbDZalDAHtao1WLINv44t
p+DyuVo6b/sRAGjuz4nJTxPCqW1r4PqDCPNO8B/NK6ZvhtmmExu2dxQGUzJ5VH731QL1f1Uv+Kvk
dfWVqrlqVPqnVADb2pMpx/Pgrn+WVDsJ4p7m0QY/UfuL6DLqQI27SXM2KnjeDsHElmbmZ9w3/rn0
WUHkF0dd8EZN9rtm4VnV+joe+X1p0xLvMtEP2c+VTJQmEbfa+onUJq7BMfPwK1/pjV8aOJ+LIM7U
fleyTMlqEIIuFUY8ZZm7estzn+l5xS4pX0QAsZnhOzmSqYeEUF/NSvLjhtCqXNSzxUcYQfLzeIT1
m/HNeYdvq8j6nKkofhnmylouQ5XXJgIXC5qDAAO2BxUcl8lFD2EzUZ+Sf8jYQTbnLUkLRVjPQMIk
GW0Y2hgfcTUfBQs5ZJ5soIZbj1ewNG9UgDugP1mtWAgu5CxnbTgWMwaDoWBXJ9pvJiZg9fgbwL91
hdHWxETeLFMwlp7rgPAcLrm3VKD5jw/qlig2tAIMKHaHOJg8VvA/hrF+8O+8KPbu6q4fjPWK37SM
Bfa9amTRA25+Wd+KxNnbMJQzhKg/2Xj5jfx/odMJdY7XppCfYWMcuz/DSXPo8TaOj0uaZvq5gnSE
6xwhioTKNVYQjZWOIoXw35IGMH3YmMlnrcBIQdo/WViwAoh5wTui3KHSuUKGZzXP8f2X778iIQVf
RsIhQI84/0d8B3x6di2vRBjqyU0UHZUKQ2AIVRMnN3/EjwJJMrth0vb4qcpqbB7jCEHr/VX822qk
Te9+TixX8CcxpGybw9fB6MT1HttWKMgF4bao92/0CxTKJvS2b80zsPYbSR7erCAKygfLvhCck5qQ
ZXKPEFOFJltl8k6nBBP8midTf5tRiOpdlkWx2q4N0wMx878vf2zkArtfYbkAXEnZwaJ3mMksh6Tg
PksDQtc8+wydeu5VpW6HZlGbojE4sMnScLd5I05VACbfvlJHsWAvJQW8FBnP/hKLssSYoj1sxrcK
ey/RsosUdaVPrlifHM73SPEDRSDhA0MawxV24d9a2gySwflNCIvZJNrsQ5I9MRGZyb1XeCqfK6AD
eke5kY54f7r8n8WpUIVDo29FhWNV3IrcXw+wz5YV94xdCS2CYOryux8caYy81a0YwwmztFe83C+T
lzRMWQqSG8ZmizI2j55P3ap7uXOmuODO76UwBU3oEq4sPwACjs427Gd2MZW12Dz/jx5yjiaSFr8A
HAfsSRztXcNSXCEjMApXo+MfT0Bc7YC0xESmeBtZij7Z5fxuUNXxXxzaT8mc5X1QUbt8gTuYe9iJ
vM3486DYgfSrHSan2BzBi5qIZ0HOBTYG0cfu5qlWN7RvP+5pMuyhlqQaK/wiaR+FEvjOXdwWC+XL
AL4rf3TgTIYQrMFQA9TsrAMbpmJZtIhGavyF1RUTMrpM+Hyr7wzfVIV5IU29D2JbrWW+RDgjcLSM
Nwl7zc95kdNXsrUZNFqjOExO7FGCqeEx0BiJBDX0IvvfXb+7T8GoGh6gxgyzBIufezfJzdtmTxQl
nbAI4g7F/4pWVsJ6p/ZXxlPuzR4TMxyP71nFJRcWUzcDDdmTxQAodJM+sCcvKsq7uWhzby8Jy3rP
rYU21W0EbzemtSRUDb6jvVlz8qa70fi0KmAV34SYyZ0yMvflLAfqTL7l71/S4b2QfOUCO3PqpKb7
nbTl1P5qDqeLDRcIusAiKrtPCcHakG+n/XL+YlwMFTbNL7+NrPVpofADWurK67McvVtXUSsu6zd9
yWXeAR+uI/QfN05J8AKgB4PfJrpvGJvl9kGUb7B+mFyPw4Xpuj5eFJhhk8M8BkPpqb5FokhQL1jf
OPcHP+X96MmxQyssq2ckMc3jnyjd2Tw2KNih3gYVZchszqoXkiEoin1Pk1wHkuiV0622Xcd4Fw20
PitQ0f2tboiiuYos3s15L7aAqzeCWalgvKxoXa2pl0n9KCWbq+tOLBd28gfxoT7P2RkN4eNgLfRe
c6w/6h3bTCYaji8zqoGsrsvlPQz++Tjiz8F5Gf9aRo3ppwYzAl+dRLvYPCUB31K/DKiDr+1hkB8t
E1Fp742eeXtMaEgEUWsWsB1VWcHguXw1U0XI3D3FKBigJT3wNCGh4+TtjwAC2tM+Tcjcatqozd3R
MviBIqAgqvk6ujHyiydatL2Vjuh2XPZgzlivfvXq4VrhBL177wMUVKdqiqmnSdNLZlfry/zD4UrY
Jdr2e3kSb/bmNkFDmxNiu930vtxiVC/CKhwBCHCC/V+OcPo/XoyGbCSL64IHuJQOKzwwX4HCFKN5
AfW6jq7RinpCV1XcryXWXafQKjpqj2OtXRnO4O+z19E4Q261crZP3Re8VNkN7PD/NNHJZdOo7Psc
H653y1Tx0Vv8Trnpn7A541fjMWiAmniC9J6ZVGqS1Vojq7TZQllhyGj4K5/OH1pquje2HDUd81mu
Hyu7Mm0rdfjV97lpGjOP7OolBPhKEXm12ruCJ0ihyK6BTJxMp4aZnqrmjFPETRYHX9rTajVQHq2P
6GOXrE0j+ZmtO8ccFSrh8FTATEvxU3SqgCNyBV+OAYyrRB6+Y17drNDHQrwOu7JBKCjfoSgEq7PU
dasQ6E1QAnkYlACqqp4JkS1TLCdZ7DUqucWjSUOREH9Pq0miwV9+GrdxwWquubez1i5QbxrgyhVr
IvtLCGePq39jdLXOsDUiClpKMiUDw6G8iS6BCkg2FPJitV5GIIJ++si3Y21DPdkLg+oIhKoEE8nA
trdRIjHOLawcAtDFMMwv8jkbGTovyu5Eomv5OnD1TpxXds/51nurvIMcdI4wX3flSFrJkh7HfVvk
F7wXJhWRh3NrVLN97u8GVfL0cS5dNQVaoH0vdW5S1/2mp4iZZfnUPnVoPURQKtsGViVIvY+Y7Xsl
I9aiV4f21RBJDaK7hbIpG7fs86XZkH9YiYijSjDXwCG9733FDwlp8rRDYt7uGA88dUkv1G++Ebx4
DYuqh4/wG/q4Nydscf3D1tNDqsMeyaI/xhQGmHjOGGzpSzippn0xt+I8L3kUO9+HNWKexrpdG8KZ
oV03gPHk0+t8S53WTTRW88AXyuSY0QIHdczHIVSacBCmJs/n8EuoH9jaaIlbhdAhymbE71GwGXa/
E4qOPP62uo/KIKVEN2IKE5TQtl4vGFbPcITs7uZNDQ3JBKFEZnBNsA39IjjOhfQxr+PYVUFMyFQR
Tjs92I/zFPUZapKfmeTEHlAFp3zdLESDd2XieX0Q6/vM2B1QrgTf5sS9ajmsIRX7re3PU9Xh7zRp
rBmZLgxkWBUxyP9RhdtEomy4zLx7klHNCCbUYvY5Z59LT1a6n2M/DP3jnCdau1fWlN4NQOf/yhcA
031alxuK8H7Tz8fFWQq8PWWxJfmOmJQGoBIKZDilacOp+FxV1vEUMvjJEFwwZG4kG5CnWPlmSiP1
+ltDRizkbKQ+PDdnrEdnjg94ZVDndqcTcRmbZH5lPiYNwlXnmCWKZaJ/VQ/ymnW+F8WzHpNX1VnO
lanbxUN/5yGxwG31oPli9hIP0nt0dZO8ioU/QhuIwq8e4NpUIFS1ZfJeDbmh0YYF/EHtSakls3Pk
ARGRxU+ZVS8Q+8ejROn4R7kYmkK7KPjBIn2FASb+Py8gAO2hp63KYTYtWdYTUkcqLkdjzpfkogG6
oLQmwyzRHAkU682PyO49lAsUIzjgyshev1mb4rEQ85kSgXSZMUrZpWbGTzdWndwQwRxhTddE9H26
I6Qpk9TAlMs66TQUJhgJ23wFXoMY20IBbziCw8rzS6xoOJDveakwfSd++fwY7hTyW+5oWCOlnP+D
f9Fv8q8qMBe4hrmcj90Q/srM72iPTqcnaZTb0M2m6d9Y1kUiq+Wh8Ki85K1WsQrUGAskZWsF54PI
Px/9EX/u+kJh5j/RpU/O6pNNjub30HS4fXspOeWMo/5OQwg509qM18m9YQxt3Vkbt6nCFelM0hSy
nvwyrwiavPwtPvSWax0El9FR99Cljxgxsboc4iqmnSBp93seExDQ4Vs/aaSpWiphmVA0OpCGZjEH
cUa3fD/n9/+5WUS+NomdaaHFnqVCok547SyZmCZ+6yJ62umIF7MoDlbnFwIqHlTByD+Jt0TmdCb7
zjUlKlGH7eqY5usw1BOxhKILPdfq4Sh3uBqlkt0tyuDy+mdvuyEQJZk9Kkc7BLCzou3rx+xMN0ye
FkToOSCtGvxy7F0XD/FhI9+/w1nx1HTOnBBMW7P750zUOs7InDa2XpHB3UWO25XzWACgFtjJOs3T
Dlm8Dtbxc9AVS4evzbQIis/S6x0X5+UaX9WoBBrnoZqTakUl4f8cvNfSYn0BNUm3Kl9lRz3VARfa
z8qBsUPkAHYn4j3L2wNOz3Kcr78EU/H0SMez6BPeJ3CBfLA04Obppmx/PmJcXwuuFYhV9jOLewVt
Wa7q2agu1H2CDNc4d12L/UfJDWua8Lz8wpIY/87prIAL/Es9SHqC8Se4ay0eqy5qvvSMaOmexMx2
UdznEtx5h/lnEc5CwiXQbH8dr3xQvMUygz/WfZaRM2FzvnEp2hTe6+K1NYVOKj19sTgL4fjK96Dz
KcwqvvO0KOf5aSySg/2MIS077I1RtFOfuTrUpakd0sSEPiPidqbBeQwSahR5q9N4T/LSksjJmC7g
fi/7XIyA0frV5GCPLOrWaa/C3Gn64PwfPbWokMjT5ragtLDhVAnQ7u+aYALN2CKYIzK2Mzxh9Vdt
E27sSoQER49uAgd7GRC2lMsr9EpWJnPGHCNwDdRas41ky/vpOok8wCRD5B3QeNZ7B8cJS2byQEIL
qDLri23SfTheg2uugxUzd+s3P/Mj6uvAik9dS8TkOVFjoL6THwnHLi1ZahXJS1/z2gsHeUxd/0yb
wgYCoJpCm1i8/Z1ZgviZqWEXNo8gUsJPEfk3semZEweHfQ6S9y604AO0qIzCuZbB+bOlRoFv+yNd
5Zrq8POvOY7JRCYG9JDjwccVBC/k+XEfbpkU1CzJC6Muqk8fnnyxakwwVY+TjcZ0JpAu12Lss9R+
fz8v/B6fbuuoevu7ietdPVq/QXhdw0LJJv+PYCERlv4UzO32TFuI5gZ9I2AxqCrxtHO61nvGC36z
9ItjJPHGmjit382CM3OJjAvdUU7mBkWdpLuMhrshUByU2GNV0ixwc8HIj8mLNfIGTjcYDkBjetRY
yE2BZKLJ5UZ0s3GHQzoXukNnQIt1W3AQDufsJpocPVjPFocR9dVAocVgsawVxZVdgNGIO2ZpDoEi
Wlf5+1sL/QLzUw55zzd7G9ODfKoccrAwYW+gbNKU/9I2gbgE/WSL6EbcE1mvBSNpbP7LUGcSsObY
Mi1p573wyVZi8S29AE3TPAaK+IeHsJD9iTbA8l3c+DBr6TXWIiptUBogp6eRNFJDfk8GE9isxe74
DWhYyf/pQyuYURlsMozNtVb4Z6WDPVWjT2rXhOKxsh373eMetBCoOYzKDAgdQx6FYbcy8S7ZQ7El
JJgIDnhy3o1kj6SjDE7WHO2t6DTvCZJbdEstfwKM8dka3JzDxIeIZVcbT+f7xxsrsK/Za/YbTygt
5LR7e0EOsOT54vO7lWw62mhkATm7K6mI82x8rfPLS38gsxgejYZallGTmnHA1njU17b0riW6XF1z
aooFH54IdThrRDVVkvsGrV5CDUOM/qjZ9RHRF+6j9L8KNTX87BfLaVKFY/3VwNM2NBXBnyyVL4Nl
4o6EdoEYYcvTeR17L8XwKJ5gzukoQdmYZ2p56871GI90X8QqTzLNwRk/iFuaKvtXSV7pHlgTr/M1
0RvI06Xn5KjF8GuzSJjY6oWKmYQQ13cGQ+VIeFP3eJQZluk+j2jw9ST/szGMMtaUsqCGotpOogAP
tql7g2QDF0JujVCchtZKoVpURn4mFX5XcUfcn1gnFCyP/uBYBgDcH+lTfydq+kYKo5UUEyB3an/L
Ab4ZMZQKZDo/38A559pMw0nYyr/DdXAAOD2l8uw2vyFkxWW5O+Ghtp29L6IXkWkkaldrQukfLQtb
t+jYC9psL5Z5vryskvtWZijsgUYI+Dzde6ytztNYxCkiRgx9KGfy5Yz/k9oRi34lubC5l2/pDmDW
rWF7VgyDxSaFK6GZS3AuGzT8PP+ox1dKYNLyAZelacIJYR6u6JalrfldOb/xIENYkr4G9fI5TOfj
uvmZeaReiBxV9shQojNHmwZIsr5djxv1+5M4I3UmkRqFKyRZaz25jqRRA8V5/nVA+Bg/OoCDUHYP
yRRJNgB1/uwbj/BIkjg017FI5jGoIAtSF3OqbA20+pGj3LHvlKRwLp8/VyR+GZeKuZQ4s7fvjMez
PG4xmXV9EuOpd+WQGjoKdtwBy3kq2B8e1uHBINFv3fRlGJjO9ZaLdHZdETooSHij29qo5le5ihvY
eOkV8vCAzVoI1Ipv8FZQI2BKtb21bw4WItUsjY1EZ6PBv8Pz/sdmIeqjw0V2+DHKOAWOFB6szTsU
YML7SvFLgl1WNRjKGFJO/oziTVBqm3KnRNGtuBHjxggvkFo1OKduXFO0K1gDBGyqcRsLmlmoGPgn
sB04CjgUo45KGrpyu4sm6jDZ0B1Lc9tg/V37w2tjbT5LAfaItzRrPNulxrz3snbbbMIVV9z26MDG
1qVePP0qK5JGHS7PHqPQwa/8rKX5oI2fX2LO40yBDs9/Y38+xN2d3csQ4zzClLi0SQUSa/8GpCal
yKHSMWEKZF4Lbsa3zALJchTtKDKeBggeKeDKyWrqIhb56OisI0R74rebJgkUBfjA1cWND2nHtpWO
fAL7Bu9U55Ud+/8cT/rO+xPrIdPTZ2y9WdclmahmIRV66TiXvb7ssYoGWEkYhwt4uMFztJR9gyb8
cMb7zFupy6EwKyBKvSdcdlfKPVy6AXZO5poQDjpA6XuaGMQcpbwyEUa0HU7i/UXypaB1NBB2t5oJ
byXKEOk0jQwMWjDCGAO1fAsADJ8wtj89g7GY041oST8Rz0kQmM/yu/Oo2xQCkhiz+EOnweMcesrl
CztvDsJjGOvPtqvgQvGSUCEBIglTkv28XGmsXr+S/1Vuf4a/rHocnLBHLCY0Wnq3d5ea7TsUF5tC
LO+YKmTks50jKstnBLzI+639/v6wMNKOFDB9JoI8A0Eb56SOfjysLNG9u46kPblyp3JvSHw2vZ+Q
JycFjDKCpMld7GAl+CSvRGE6p1ZJhVy2L8bEynC6Rwm3P6EW8Hw76QE0pBUnvfpooK+lA7wo56ZR
T1twX0/vzWJbhAAwdjFmVEbgcJmVX6iNpbGci8I2tbWWN0yIBuc+Utj0iPAhGw0Jb+wH3oM+rHnJ
VQjBzoZkRmvgpHONWuWSHDT5rawU4c+kcemKclIibpD+pr+KfSUlTXGRSWYYSljEw5fT2J6ZGHbE
QkUPOr8DxERui5M9F2UeZQkKmLFtHj9UzrXESjFYCA397kvqcV6Kqb9+CRHScaYm69Q2qasM10LN
iC/SoV00r4AYsqoorZXUQ3gzKtvYv5S++TExKCZEYb0hHeGCQFSgcajqY0LfLolu399cC3qki+++
17ufjVaAr6xxbwvHOdilp4SNt+QTWbX6IZFCYucPpo+cLpreHa/a5AwyJoFV+Yr8C0J5UjjGk5Tl
SLiNOAWmOv2iPFn6A+dgZJhuh8Wag8gptzrgYN3EAVUdHg8IRs5D6YS6c+bJdRBF5gx+FRPFqBYs
2pPajG5amyriTI/fxmF8nAik8GRcBjhkWHmg35xy9OgRIrSPej7Wbh7ZTi+Ic40p4lRSogcY2fcb
h8Fhd88P71LvHH01LGxJQEHNUwa7GwVvwIe2J8TEmaQ6hyf8SaT78VS/RbZvd/D9MyG0+wB3gpmy
e7Byf95ws1k/aI3yu2N8++00LM7ggdOd8uV/YbIldDv9MML7R8fRlZBEnMwH/ItoRNJcub4Po/Tg
gsWmPVqSFFEQ4TDHGjsqv90wToA8grhKL5f0bEI3SoPCfpR9M9TmbmFsN5n7xn+OqCfKJaqiDCQA
NyuxW3um96zvndhy/7Q/JsXwQuw7OkGIDOacY6zl6TRYl4MMSkDQUKe4EMxi6YIWvZYm8zXZH7FX
nDH79uX5OQsy4nwEcSgE4Lrlf8H9MYcrEQl+VbpbJS3F54Z/JR0giHLm79JTHFLZJmePfz64/lb6
dtc96hJRNTu/RaB2H6O3kRt7+hQk6JzaleYziwV9KJAeUucpuwSuCDe+PNXrtm6uorUAp4Q4gAEL
VfstjAqcxwCl0aiMNbaCEOwiLKzhrKWNVfn0geaMHN58aCp8O9xA6+xjArW/MCbh2qC2QFRaZm9F
K/IeqzbBdqN515cMhwFRVC5VLYPTkqZGwssO84zCwqLsFIEZnpgs6sFnEUGXExduTSE9N6xt/Ral
FHAmNmOvLbu6cCEN/1fKuoPke7Bd4NkHSQ9RlWzX4xLShXpg12khUo9Mc34LAO1du0PWQVa0aKdI
7LtnOCO55ua3Q7qku1plgkkRbKPvPh3MHBY/OLBqO8TJnuOlt7gWFaYZUu0nuqMKK8YOSCJ9j09G
/0hk6yN6sJMytaf0TXJK0DJ8VlidzBK7tAtypSj4DIL4OSIr/G9r1BkCYyhBjrGpZ94vpzDOalSX
jtbj62NMVcDRE7qs7z6m/8fvFKBGC36slfEsX6hPe6mbiWUG0lZayaAZ97kKZ+c6vvKYfVpo+99m
QjWdg4jI2JYMZw0YH2CiB7X2B4i4M/3LNC3aeEdXra7+VqA9PFr8c2HevVZ0Iaq8ssdl+8vAy04e
/h3wLImdyr4XfhQ8jRAOLq6LRUPlhEwmatKU/2LREtoxspq7KDVpSpiNaVmKdBi6+c1/3PP8NA6z
UU7R+LOLLhqjd/kMNQ4+3AGhD0GsBHlIQaXoCQaZK0Q82dS9AGRiWUvR4fvIcHvg++KNFMyxGxOQ
2+fo0mMDvtCHSPNn81P7AlbPnhWbXnFHMAtudGnlA7FtC0reGNuoiXlvHIy+jmG5PoQi/dKKLMjF
3eKBmS9AG08CT4d6EbV3yVTcGowhxF4uYcU1s5vMKqh4qjePv5UMJkLBmkyo46Bl6eSXRDfs7+cY
yJHLNW1iLixVxYIF+jbnu8MC92hQtRYll0KGaX4+TeoN7iIghhe/9Wb8D6unAUE18kTxSeuGnEI0
p99/BC70mFTaxIn1P5t8ZdlENvwfum50BEVe88PEfRB4qKrUtiCT1Xv99b3t/7zk59aVNCBbcI0Z
6g66hz81UEe4rA1hUKCy5S+aHV1xN/Qh6Og5bRQo01Kj6EadWhw5gUERUFU36kfVuV2vjo6j+LlD
AdqewJDDEPkxnpZ2t7UFLnuIxih7aSGdvC1hiUEmsQKYE4co94wOwRzsoQhwW0+Mq0wEAx/Sbbhr
A+wyzU8Fv8kkLvhYv9/UGFYCBAbZXiQ0msaTepF78U/PBAmVPBoRlb7pAFaS3atbJ3ZK/b5K8ueJ
M1n1+5c0T+DfHLUEmaVep0gAe8KHFDmnqFRjEpxSM27z5XD8o/hu0tr6zvqYY5roYlQ2p3tIyASj
DdBYYt0TqOJ6lmScn6Kl4IZaoCzkto4fX452i33A+JxqZBCw1m2YiS/fCLp890WR88kzjaYwVcQJ
lRwZr3X2Wu8h4TxPDEQoX4ISxQ1GnCZsw5SkpE1uY5dHY7wKgU6U5b2ynE/DpcjNA9gUFYfluWiA
IhHOmRB55LWMLchD5iPJBVhAZb1a296zDV6GRI4Dx/1+JGiOQCZPqow2Lc4GmzZBFTnqH0geNHb8
DNtxCjjKMC4lyQzFZYbtA4Ps8uq1NG1cBtTaRSgYjEQpsFkcAYD+La4340iUqLvg5HKAOt8MQK0B
gTnUkxPw8qoE83K6s/hhQKZkDUmtzUvKpc6KwCEOxdCw07ze2RHacKaujgYKmGhZ85xwv+GgjMkJ
70WQiHAu4qO/zsr5aP9/+HD1Vjw4E6vTD3fXxRkT2Kpp16jHLBLe/n9vVxjE2qEXRUnIHIqxeJmN
UecPnkalVZil7VUXOF0gi5jPPPZaK9r4XyiRV65sRi+QY83Azbtks56yKubxLiMWy9qpZJA6ZcBB
E4IWQ0jerEivfdSxo23Jt6+hfER+o74h7NOXNlrIBKGpaOZYrTWNbowdU0ytEeNwdPlkLt9ejclf
yR1JShC5VbDlCyoUsJdqJu1kjzyEIQeBUMYn6ZjqKI9WJn9y4BPHV2tOS0NC0uJDYd30o9bHDfbQ
S3sm0qYkz/lVliX1aZdxYBiTnspsR8Mk9g32AbOydqeE6NO85AxjNAMtMr9qTOqNTbaN8GefPv9r
hdseh5VgRQbYJzhrdeGirEB5fQH7E//GatZ2d3o8BOYCAxI/1rHoN3HACki5i/zF4mHmWwGr2hBI
WinN8yqiY+w78th7zq5Gp/oOa2K7je+XCn1ImWi6Dg2/VGRZYOj7PQR8xUWbmpSeDP4xIjPYZiBf
7e7WsUX0BIRtFS7FVW9FOFZ0GTEDCNrv1rG6tBrBY18QShnY8ApIE3/dmiBb41dQiXAhbWXOb9Dv
KlmKkFc6cl0suhKsxThAzMAdTc46XpKV5bFdVqQgeoqxmO94jWDX0HlmjSht3zouW5pZ+s5YIGav
McsSRifcpjJCjOgWfNQUwLjoTHW8pNZQaiCcBnEzbpyBjkTFcLlVNp5AZwJ7dBrp4ia8ibqsnnG3
DQkYrXwn+YVCPf+rTVrXQ2GVyp94u95zFoLFErgXedfRN6f3Uih+0RuQgqHC4G6UZ4Le0l4NjYh2
OSGFzAaZhH9V4GhSfkVuB87Gb+/aiVwXOLmnWtOn6qpkFCmRFsM216vVjS1/kqDQHW3QhqYA8L9F
XSLSetGj7VfRS7jfz6aZ90YjgeQ/Sxxvy5MZZ0+R8zArLcraWLspqv4A32pRCJGXcHE2Yao/d2Ik
eMoSK080Uyv9kop8DqTnlqQQ4Rh21kSu/GNqaId2fACpMLugAQ6UgwufJ8m/fEFpoAoley+ZzfI5
f7x+AJmh5DoSd8l+WW3rW6sBOgOcjusagDqLMcEii48dn/5648zH9MgtdmS+2i/iw6IiLA6i0BF+
PGtyS/25mNE1XcnzcqR+BpuihCmAq7LlUA3HH6cCwBTPl0gM4GzFNhdHNjWE7rWOQiPKqe6RlIGj
7l1JncXYmf24lZBjICefwCOi/+QBIK7kIydb/9D0tnTGPm7Zr2+7yS4R/+vCsq968ajGu8K3DUOg
5PBGtGOnvfgFWwikSQL1bTrFM/uFAAaj81rGOZMx3VbpDXBECYrzPfUp7hWnMCViOWM3mhQI1T8y
4bY7spX4nMs4q/g4RRBAHeWjbvcYh3gdqIZ1LobKyGxqjNuZsijVbg1xvTFZgGtVUclf2rwvCTcs
OqH//ecDgEXNpPY/tY3ol3UTzXAF+3gWS8LPqP/sTD4ddcqSjud1n9rmceQlp8APFDm4ZLRWyk6j
goHEI1cNdSUzVyNydRdJdTvLdzrLle+eL1Od0APulUxApWn5zuSotVE5B63HjrL7sok/XSo7eLQf
x57d+n9MV25S+5pA9LwSW82J4Jq9FrV1qrb8wA/YkcLSqXR722nFs1KUH7UzIFYWN7zYz9jtO2TD
z5llpCYFreGKvSswLm1Qu/AMz5h//KdZO9T4beKdkcnU3X1+vYmUGVsitwUCm4AoFm4oh5+4kbWJ
wxbyX8/XoK3bMU9NODn6+33rSE04QmuQZbjQWaBtPiPcPaJya4PpON14hILut/w3oes8NIaOIOyk
PuyrZ2ERb/K7lI/fafr2zGQkQaQ9tqVbc2ZzG14f53ALy2K1PE5q7sy6kJxB3CAYyb2TgW8MbRM4
l2uJWB/Y4dAi6JJYkF71ODonJu/LCXYViOLx+klqdiIE64UGGtdk31pB6PGH/dUdv1iU5uKXdQY2
pJaeWZZeREDMVAYUCqdUu72Cz0zvYeW775bnu9PX4w1dA0yosGfpcOdjKwOY2Uw/4JZMM2N80mFq
E2QGSggKvQt0c1v/kwDQtFAE8d2UeH2BTBwmXJWL7UrbhU6RaNfy4YHVhPAIrfOCP/iw02RFKxkq
gVir5qVEPOsofm/obDwJPf1zpLdhp5Lr3wQdir+7yMfuQSFe7mfql5RFLI3VsRnaFI+Qr6/1m2Bf
6u3qAIQGE1eTf2glp3KMWhKz4iZDVZbvg1XLDnJHNmPm7krSl0e4Bt9HCIYyf1ZRj/DmCesctYgb
cadvI7DwOWP8DLMffHol/4Nt1F0bKGMyIV0tsS7adSJ4T68Y4Lt5icXVz0SKRunTxs3KIGhvSDt/
Lz4mOjZ04RWqJ/ENmUuwzgIKCjZqoRZF2wMejXw8/mwmJ7xCEGNKmfevIhFVz5On6ulewIG034CS
g4Nuv9MfqT8aZ0mXnZP8/ELnjmHn3Uf1/TXrGKqSbQOkrffaLW8RRIGDUlGJFVIx5C/Lo3pyY/Pd
DBDoadxFXFVYsV3sXzI7lR81r094OjnGNF1M7sBzkQej8KIagsSIXg+yoIU7okQ78AUVe/peWR9W
vPsZ0XTyw1tAVTYrgNTXBBn6LVkZCdL7wgSEbnJaSHLZepuqmdztj/sbbpJVamBxXi6K/Cf5VzuJ
thuQ/p+cAbCuV1W/euV7QLHr/PxlBk5dpPBKt9Iwg9Qh4A9zquKOp86L/gxlk9H39uuxX5jxt/6x
vn9FlOmhQFsQNCkVOaCxc06f+bRFkGS2CyDvvaF45gqjG5Lb1pk5v5EzomKQhR9ans18se7bE+eW
mITDQEhd3DNTUR/6B9Bi5oFExPXXzkOAZEQDvubSTBfiPKZ+EOKyaeD/Y3KygzFeM2zjdUnte36g
CzTmGbOVDCsu6zkgf0Jbz9njuwI0zCCaorp4irP5G0O4xvA12I8qAiri7lbtpm97MD7VKkg7GasJ
s9E/Mf5k0I9c3U9IOskxkCVSyCv/pL3maXefuTG3hrXOhcD0abBWY5owKhyEuY/+yzvd3CodCywe
HUZzwiAGcH2N11BNLmSBEdDehcZxsLwSRdAo2FtqpT2L2Png7+E2pnCXOfvEHdH8mADmer5ebwK+
lBjWqvyNyDoWuopV88QOTm4AooX3YLGnL8Njk05wKFdx5BEwAgbRALEzivgBFe0+NncdXJjRNjkl
Wu8pG6yWGoOZxlqnADfWhvwo7waKYbkVRJhD3m4PqOYitF08EfN1g/QmIPX58IosxP4vx9XIvA7N
cvCp7BozP00GYnUvPkdklyTpH0isDtDS2jfopliGjA8mKoV2Ioe6iQYvDIYkIJcdxg7vyMseqRkt
afPgB5Cj6IENycjaeeFNT69yYyNUrhcESvHm3QBFRu1/mxbdDsAWoNUj0kn06AMc1oRw0WTOicrh
cWvqn0US+8aJS+3HMHO/MHr2ooINqnvbQXrQJGKdmR7ybViWRkwkOnUT78uHZQ1sgLEQK514URdC
os8uMtiMD2F/1CIBcbr+6bxtsjM9GwgD2MjOaaM4tWsCmc0nbm3sxAA19OAkCdj6QLFJgILlouGC
RXidRWS1hZp8sADnFuWb/8ki0qnRiIgz/gUVuKKFMt7oFfR22QzG5ZSoKRBG23+Ii63dYDrdOw0O
y4BkQ1kTg6qLRPj0UBhVt0XdZ2+gE/aTSZC98pm9Hx1Ub2N4tbCDTUpb1136b1MYfjY5cmxMr9ep
QkrYYw7tcj0MiIM9AlhGFWz7oxJkDF7Zg0w412fBowakLeD1JblJZ9B7U89aNdXPSZR6qh5n8FpX
o086ZRYPu7XY0VA+rMvLyyqU3nSbOaMbsMS/olYb5jNGg/5BUFgOsmFJJ9oTBOhR2lo1hBDFqusY
ezxip4earqSiw9cbjNZFuVxpgOAoF421k5zRY2YvtAyw/9HAg7lWfV62mJW8go1ihsiXaQHLIn79
HVtmS8kVntSpJyBL4LHGClbvJK1o6aT4SJeCmYJLf9CLzLzQYrD+ZnxtEMuTV7ko+LKVAARc1BcE
526M8zxeAgKjMcnZNDNq1onWnIxlc1L1EPmGjWineiavObd0USxsF4f7j8VUkkG2jAoEbgOHuMDH
0dUHovrYIc2kMM+wvAPr3Ac10h2T10YzGIWRJLceUt0g0VlhXtHF6xbevQVdVAE7f/ipaxiBpHAx
74fL2rBtxFH10P94IMcsnEJi+ZbRdRpnmjgI+Tdpfa50gqHhRBi7/N4ArQU8lfIKHeZm4RD1oYH4
jPGjeF2mPoBfNSSQqJIIwDhKN79ANL8H0ly67EL7893bQbv+x/m4GZ130+vGr3Efa+PLs134RON7
oMGCFKuElft7WwlvIq3QQeC2XebUyGJlN+HHP2LDaIgO3HdiTsS1iazjuyUWLFUZ2bzQUT5Dngqi
s9FLa8/TQexTM4PWjg7jW9gMgYTJI4Muyk6kK6VUmxZs2uXPGyLfk+UV+VmzQoQVwy6Szn0oK1hI
D7X2doUpf62fhlVTbw5ii5iU+/I03y7xSyS9PFNDBQqzL1IiLpSH8frmTw3RP3+ya06zH76zxJcY
u+rMzOaheZgfCU3XxwOpBYnKNBu/U7m78PHsNqjlUSC+RIpV1oEqn6R70YruEXweygOxdbtMy3Km
AdbXNcYmQbTuFr8HozAT/Cc1t5Emmfp31uNGIYIsj+XIlHHEGzIemG956KT14lUPfwr4lqL8f1x0
8uMQ2w0cFKNFTlGw2DkXytKpMKBuAPuX8s5/forZC7xS8lzVBmcnkHJYhoAav3H3VuVsvbU6P4/X
8EVeJ3PwSUTp2Foa/JRhS/MhXLsY/qksygjhUmn1e6uqI7+vzdDtS7HMfe89wFsoeD/tuPcfA4Z+
mVEAl00JBv8nyFA5jH9GX3cj9oX6qSOdnRcaOKEsBGuVwm8kRErv8ptwfkLQv6WaGz09alQ91Lyu
sxa9fZTaS5N+fniRpTMSKu0T5tDYF4tmA5YQAIo1GslT3abRETGGX86kmFaJarupXJJxdCWRL8qd
Danyh68ElRGtHVy/WUpTM7T/0JZ1oyUocK1kYITtxVsAwMGSWAhqcKfK9exr6YwsR+HejbUMjDyX
dfD80xfQHYJdD1Q6NGA6hpIQnJ0q8uu789S58RjuQj/XrPdgm3Ugp7PTjpQu4UzaKCM97HEzL4dN
ao1/l1B/tpjVZPdtZ1f2ZVrfTeQBRut7ye8kRF8PYrBUoUfB/u1/wf4GF9O1DAtyy0k7De6BIoo+
neGXEuK7ZnjedXcTmFypSrlPvy0LXakx+zs08eoOZGeJRg+mONx2h7xgrVpw9DWiqy5mnZyEnJzT
YytfXtpOtuhGfvM8AVMIZBJJi5oaBKJLFxwAguGDCSic2oTsGi27QskDs91CXRQt1ACu2EDokCSN
Lfnl+SIJzuXwlYt9aeKlv38IU2+x8q8yBWqud5iLzKO0Vk/GA9A2AtFj0ZY89WROEIRQvFgI/alN
ids5Inykr3IuyXDt55RhrRNG5SaedO1rmDZf5RfdU5kY/ZE7k+b+lLqLvGnF81qIHLOaRelUZ5xf
cZhmqaNfhXMjOwKaa32+Y6egPc26HmGzJWfno6KXcbfyU5S1Qc7+6N9SUBca4yFqJAT6u/EmgwGE
Pjv4kIDD4QXN2nItwGAhw2dxDgM0pcDm7WZXXEOTr/7FirmKd12A8EKkighjHmITEGlfDqZoub4z
n4KDiBHkOiVKTh955NQ8TU+N8KMMSFqDYLm8FHzJQpLoU/xcB5MmgUItnUaidyQPYPdKBV6Ioygn
mBm2AutYIquFq0PlpyMQaw8M+ql2S897AQoX3ETDOF+p/WjtpvTDAOOhL0AA1sGxhBTppWCaGL6I
smjF/GeoUgTq4QASwHCaR5+w5kG/ab8lDz6cyvA45o+IK3sbniKx4mq/78zO7kcOrRF6dRojMFhs
prslLEUFHii7vFGjGw1yyUmYM6GI3fuj0CfNBefycAESbDOnZ/exfNx8kk6pZt+8cWMM2gElfEcG
06nY+SDu2WIpP63peSIFufhqfX6pVQR92bJlpgJ3BS5KRmeJS40GrVrCemvyoqLjntSTm0E5AXhq
t156oAviPrrY2/a7Ltab4WjmXvSxemgitIQ137XcIsfha5nX5g7TOGGiCw0MFHWp5JETN9yyVRcj
TQGNRA2/xY+R40Ie1Bd8oYmkOvsGC9uzhdP80PZ6bbaukSLoUweOZAcH8/xTDcsckGyg9Bi14IIF
Ym3ESgwIWWGoQHNxa+Jq3hn2r9pBj78J7Q5fAZz9gtlTbiDwnghoS7onNvQGXYENXTp0I9oJguWE
/4N8ljNMNcjCI9jN2/yqb7X0dx+B1rbfNa7l2E5PFBchuTyDuX5gvaS2UEC3V+0/Fz/CpaCXoEyg
Sb8r9UzddKMriXTDltlHSBzCYGp/7iVZwniHQzRIhDbyHsYWB+uD1GqlkSuOysHcP/LSIbfgYKFA
5MplbSTZBtTx0lnAns3IOcbtJyxQUJpDObWX6EONUDJQct0dqHxVG0Ay6LLtbif7HMMnDNbqZNTW
y3YsasOAiHlRDJsz2BBwPjKaF60lhZh2vuSHuMQhYMsOAASLE6KqBia0Lw5wgfMwRDLc8mPG5BLY
5m++oEe6uObDv7WTCzzHx/tIBCW3V8Yyh34qgPuoiUR1npiWxuSpCtpL4OVrUPRH4/XS6T0eJiie
KBFyzAPo65qWNk+3Zdun5gn5jS6Mn0GlzrLTYmD4v9gk57xmsZ6GcLVMgguo8pBL7bB5Vq0rpURL
nGf1hwUFUKEJWzB0BTokXQ3zMzWez362k+k1LWw3AdEqA4E3kBq23JkaOJN3VAfE596fC2lRufTV
I75aNpNmDsSUMjmjhqjSYgRmDPQvZHslYa2fM3nqw0dZhccEEz8u/Dl8MurgsDN979wyDS5vwVlG
GRHMmGwN5ajakMERXZeJ/cYigYVCVzSN1DTqSm0z2oJbshLmKlD1ReQ+FjR/s3LDP3K0LrdjmFvv
vZoEltFEPxFyn8AVsZxJP6px07nXcDEa8yGYQvRCWf2PRHWmtQoPunYbmb8ugHVHCnPtvgIm1hWC
NWTwoEyXknqJa4CsVQRwp9wYrMG5O0e4T5XFZlMp1V7stQMxwleoIW66A0LP07gvztMc2YD+N3Ac
3M7CTzbHFeOuA/KZx32GwKM3uJUSORv6vxadrZp6X5jGJfxBMnQiynAhp+v1BRJ53q27r3N4CQ5i
s09Ov+6piI0OPD4Jw0zgbBaieaMrvoRt6XfY4uwPRR9CLkhcUGYFbzOsUa6djOlkalpYFsk5mVAl
5n92hN5lPu2w2ZcP27MLov1vK/doxABTuUAIlLgh+PsNx3rHtknSEtNtSYk/z2Nfj+LioWXhFKdL
ZFJlYvbCBgTlPY5DZdYdg0Zf8Nvjyu9RubGTsJ9N3KgwSIb8t82AdabE+mleyDDfqggpsJwamVYE
mWBi9X40NnWofLP0g2ayGbxgAvyyRy6v3H9z0VNL8qo8vDmq+fJ0RlfYM7En95OfxC+QIwMQiGOd
Q1Gg5nCg66PlHfsPp0xe/I8cKab6YcwxlL8J+DAJAdyYprIh3sxcrgkvTx+tYxnIzGKZ8UXqHkkw
TPWOgPJrjmLBkBmmW/f7F9tSTUkrM3qcWx02I8ovVyUuog6XneXIu4FA5dxm+Y2Mro3Q3XCNf1z6
b/vnIVAoeJd4p4sxa9mDjOxq3fre2s53t7JUu3vFvmPb4nIWc0aa23m/JI+YeRiPiIvUutYQuHrt
hY6SYGPDfmEjyIelcwDAAfdutzPjlYvuMFS6tEGzsCUP5tQ6jLnLz7gt05xjyj9/uCoM6mdd0IjR
r4ULjAqSsep08LlD9WHRi4aH/vv7GMMVt1F5/q2Mj88BLQrCTiuBU63BR3Sv3t29TPyX1HuvwuMZ
kl3vX+Z6rEW+EnpNxrMeu92iGxWaZWZ+ZS2HK23pEeTCZCfn9Axb0TE81m55Fuvrhc7LRKiYnUF8
558a6UfTeUwy4G8QtJzikEhf8SXZE0pajk9PZtMXzQBmC2uFwgqHEnNNQKbwu6SgJH+OI/gJ7UF6
4vcYVWovutZGtU47HtKR/UqYBbhU3WMxcF/UR/Nv/Nh0XttaEzVWqucGBY1Gp5PnhMoZrVou5Ol1
6EbybQZbk7fzKk4N3+Qk2ey6vwdSmzj0JVvd5XPidPbCQJVeJDeQbEieX8LrHUnjHgW6hLcVBtAe
Rr+o7HDfKKnbdIdsHh4MNfQyiZzrDSSEZmS/q04leyu0VcTnLfGxPeAICdbyoPQDmq7tEPsqLzq3
6HRGf1z5wU9UZdNUICh2g2hPMprJ7Gu/0rXrx/XOPE6ZH3A1OGl3jkXtI6UXPDmdTfJYFgd5xWQ1
IeypfrS8DEn4rZRFyKnx4ndtmP0SYW939puwdR7RnDmBeuosuzKpguXESCeu4zVL8Cw0UE/hWHLI
V7xvoQxDQzx6Uxsdl1wKlNy0jBCKP8LNZZm/IjTmLS10RlyyGSihHP/sLl7Feo8Ci/qYmOICEA+P
TkY+LK97n4ABgC4s3mD4nNP4SLdA3YiqFiAv2s3YgIgNCOSQtIs4xFuM1Ed56Lbjesr3diC63ZC/
WJes6Qnh5akbSp7ZB84fQyscJq3qBlxAy8f4tlWZ/q8aqfwzMP/snR3nojnbGQ7Vgfcl+Bn+ZoEp
t3S0V/B5rT8R6yHq2CXiBNTvaIIhnk1TxTpRLk5psgtzhJigJIJfGkORZTdI8euxYoIB1dEmQTr2
cgmJCldTsefkUQectz8bUAhTWLp602hDlkT7mkN/j3s4Io71iNXeF9PAslc6NP9j54cowyB0YR7x
fvBakd3OQTNddGoUEAaxelOUn8rCfoW23XbZfdhSGXa8EfSoDn8O5u8nZNDQrzMkqpdTC4biRMM1
c7tp/BNPmkkdYtH+/A3dAZwjUSraDGXf+KiooWi/NUQ5105WHfEmHqCGf1keszkAiAdqU2PpEN4d
LZD48emH/r2YbbwNDQ6AOBmpcDsFQKU59KBJ6/UcxQ2U9wATjA/UEDYwubmSs4lI5ACOO2HtYmrT
xZGS+ARc6J290lSOPE2lw/2N1WGUuaEiTM+NR7/SYbmvYDrr47qI3p/+3i+h66AeeLbsrDFIj5Hl
1DKzpLRPrLRXNEz5O//P69AlP2wI0df8bGfaqSeN0qh8CmRvTyzh+fzq1qq5ARi0gSIyZMQrJSwq
xQaGFyM1wQCQwm8ZS7MC60HiLEbqDdZTlnStANK6iAxyZawPwS1X3GFSbRcvp9XVFBLRshUSZbyg
lSpfJlbcaIDKpipYVhROKdPdOZZS0lz/BOLP2s4N5aLhB7OnaDdOV2BoLVzR184qiU3+ohfQy/5/
csl+sGlL5eKmfoBTQBgKMvqqn3RL0URPae6HXprIaUe1r6Ib/D/txy7vPFAMwhTuMYAcwDyuf9N0
ejibwpoquuSGC6zRoXMN+uGTzdkeielYhwaTYB2MCORKZIvwQjGQB5Wq73gJJ4aAiuotXEReBu6+
jqXrjHTXngQJuISERNpBGHWQLPrM8mLjoJfn2bGcozWK6uLfiyrJGGrCqj++EtRR7zaH1cvV9X6W
xqbxcnIIhUzKNtTcfgBm1957s9Et/fynID2EtSFmMarzwxAoumW64hc81ec32c+5Ny5nk5jdt9pU
F5xqjQzXXJMQc14OJNspRxCe4NQXE3shPyQoC+ZJERtzSYrdNlPQkKz5wzPqSCGjkPyWx4MF857m
qFEVudu8j5JKbkilfSOJWICaM/qLzXPLXfTLyA5yOGKHwARQqWyKjyWk5ERI6QlLCJGZvyPehzkK
0N6RU3kG1en8ty2sxB/Squu+U66x2q8fqlBH0tyIQfevsTjjpeEw6gXp7swl/Gg0xbWixSZtIA+Q
VyMZLG/ZJWLEcvnDyXE/SHSFAfkXjODH243XL5UBGGW9D+k6lb8HqDaJ/5lz0r1Jf0KreqYXwgzP
Hh+t9zkIUwx81/cxGnvodmM3EhI9fMvhPMgl6b0Y+YTou7aHkXJq0ZTMvBzEBMEkctsc00d14H9/
FNWgAINeT3ibLyatAE90luvtBHy2yVbjcyuzv5lbNolwHWF20uufFOxHQpZaYeGw/1zymq9hSfgU
vd61qm8rWKGBEj0uOaCtvGPuP+SgbGCxEwdsxOiNZrihVSvu7aAPbjLy6vuSaHMiVXERLWh9KUz9
CTBaE6RY4QLgME29eDs01YGNGM5pyDzYUvzSrrA39cbBLCN1bN3FV0N/unVZUN5iIUv3ur39MNu6
WpR91d6rKMNVz5FGMLBdNDRpHSc43hhLbB8DmUTpFf36lfmNRTqSitXeWeR+GiGm5B/HtORgl2RW
IzE795zulhQuKWoNCnw6KIIQgg7A0CNyJf07oyWSb76q0RzSHLv4OO1HC2cOkioVH/y7hcpmXVXo
KkhW+BQdg5QwY8cv6TtIjAWwL1M2tz8JL6amDd2CgvaJ4zTQ9w0m4vz2C1Y+dZmfajC9pDhMcMyP
Uvie06d6Z+gNHDeGfdZEhqAKMunCnMmrcXOTRDtGZJs2h+MpcD6MiKGFHZ+DHHVm/5BfJ5kvk4CV
KWEsCwAKFBeVuBJrOzA+3Bm7X2lgzjbO6l/sHuNL1OgW8WktRtkJAVXe8GE4QKxcjkWceXrSuH/Q
PPbtj4IuEYW3KooJMXxLNjR2WXbq6Yu8FNhz07yI3TiFs7BG7jDqU6I19vRR5gK3CKPw7PxwwMj2
oM3jU3A135JfnuTF8dSr5ntFaml9BlULhtBVgqpjKhdsrvH3/pMVGQ9WYNbH90qnU/deI0GCG/0a
yfh6izCVwova+T2yknm5bterC8VdJDMzsvbX/xJXLUodYNTNUM5N5N7M4t1bMPgZmiEsXYZ4oUxL
RhogV2aCrpaOh2XEqC05l9mdbFR5RyAiEJx1ybj/ACzgCgaOUueGa4AWpaDUxBUs3GMBrDJcyEUp
TW+rbR11fa5j2ijNJnr5gYsvWQzsrcN1D7ohSj43a9VGA8tLP/e7VPHTPZsty2ZcqVeX+KbBtkQ3
dCTOuuaTmrfjM4vtlDyvGfli4xAA604bKHYmQu2lLyyH1HgOrAtdyLZeLb/EmCrnpnIE8+CnRf65
SCHZ+jnRIIVraCZ+FXltQ/SKb1wp32V2Bxa51EITfWWhk4gYLG2UZ/pq1CSUzs8COl6hGZXpDSkg
mWZTrkDLs2JcNsNkYONUfPPlryffokzw0l2atnAWVFGaFoTP34rkS2e1z7hG8r24Ng+6olAk6nGV
x8g7xs3xukjzZSaST5E8YYSUQmwN8+75E9re6Vq0GsofRpmmaP4L3+avDXJogNks169fjjI7gCdV
JYiH/fvYa3QfZEMdo8feM6vtTGw4irmyDYZghkJtgnD2cOfwq0WOaLsGVTh+wJHksGih3nVSfyq3
vYGpL4izQ4vFUxFvnPT4Voqow9mYD+bw749BKgtnZ5V6KLz7X/GxpvW5Ss1sjI7iOZhPUh72pw8z
wPnTx4f45QPaEG0tLIcxmmviIUOhCRgiHOTj93YkFzfk6kQ0Cl0fugJAxMuaIH99rS7LydovtmWY
/EzWzkvUQKYv1sc6Vd9fyb6SVf1/M/uAhzZDYCwsKLIrjhG37v1EwgaEpqMomcIyDNs5Vunqp/jk
av1lOQKRDXxsju6clYxpw5n4LkaR8IySmykBx339R5xQLtRwfjsy5LQj4Tha09Z6cBvVqtT3ne9w
i9mtx5rMfJHjEz/nYg3NJ7ZDej4pv2uL32nDIZc5/IFE64Nk4bD7djUkwjVHQi9n0pSXHCLidO3M
N2nkoE7azu8zarrxuBMo4u+5Yj+xdJpdF+pKEPP76nyICUgqxcr8G/AwU1/IEu6N7K9sxBQNxu9a
I/Ypq1rvw6Xfq/iNcqWu8kbA7bCsgOLRgAWI4s0SeuFhuSDbI8rC+IfHrlz9vUNPgC1pvU98d7rp
tGr0YALMyqaunIWEF6LMxdp78WyCL56h8ERmSgD7av40cxigopefnaeob0lm0fSBFJ5O38fqc6Xw
1e242kHE8Lcbgx5DiZ8/FMcoNzzkO+8GiKm1Mw7b5v+S+7oZesOWGU+z3SYAa1+ptNT2KHYleLzS
tWkh7QH0ZaeR3z3AOYNUnxQ5RSZsBdarblt3WBp9uDKIEvtxmhdHywBqlMBQkU+OYp+AO97ID8ro
CusqgoJ7vealnq6hebtCbwd6gNKHb+Zw8d9gbDAY+oKe2AWO/LBB49uauwS6boH3jSAlYSDaEEp9
IQNVzvJ4kkDmixwTT1QoiF9FmjKBN0+6r7ci/z3qYv2Rgk2SEO2jwjXYZVD0mtKyPtkCRaATABm8
PnsOVFdh3SnPaaoi6xyVrJrvVXls2BllxnVJ5YvV/FpS+s1N5UrEz4FC1RBri6+iHjA8MxUkFHTL
0kqW4Kl0P8tl3Dzq+aPzwdhrO0/++6Hbx6pdk3jFbGXZb7jFaoQqAvMYNu6Jlie/HSdPxW/gNv7v
11nml4urh5/zRgdTxKWnttARA1Noare0d3NjB3w/Nq9jrXKO1+gC55/VjWiLXaIqT4X62KbjEmLP
YYAI/nnFU4GmIWCeB6a6HXs+45smftuomlvvHuot8J0h2QMxNHOq10PJS6OFC5Cv+1vUlAb6D3dK
PVnstWcwZMwHsnmDXiV4WCKo/lsoNNmzuuO+t74d6+wRxMqhYcn0RNF5hjqCcAYz3oVE5pagzFW6
E/5ybcBXWfLQ5SAZxT3EF9owwrC0t/MK6AShoBClIUcegrvXxIG5PGn0SVOcrHzRNgH8M32LkDvh
2ngoGX/NJnyTfLVZtrZMh/Pte0vnAofpMs0BmbSIXhMZAxUmp6khVVh++OvcF8UwB4G8eM0nAFyS
r5ibbxphK3fd08GiL+LfdufSybWKjq3DxmrNf19ypu+SujdlFvI+hJus8/S0ifBwOEUNUna0jxVw
q52pTvKplLcobdKj3L0960+9qXoKdh2e4GAFKSS/JJdWisCw6K7ir3VACLkwl/qHUbxEnoJSdGwD
IJrd4PG5a1Bz3YZSjKEnZbyEoeTRizxrw7JWGjZwKLua0ZGyiuDX6SKxu31TeN/woPYLeSvnn+oP
+gqkOESjuQSRRl5rnq4E4yRLATpiCEScu7FRY2jIaMicyx2r9oyMcKIM5IbW92Onzd+sCH3YVw60
GEeBE40kxpDwHk7RNqjnWa6XgNb0ENu1GeiAsbs9TZFo2fE+9aYoTGxjyQnjkZM5K1xhQctBTKSY
m5UY3/R09aNJ1zOnQPxi0QdVat5nurs6Txp+Ip8tZ8A+9Q3UPWRJNn7h6TeuF1rH12EQuwse6ii3
KXQS9x8UrvxRnksHmdNdkz5RGGeOD3StjG+GvWjhp3nbsSFI+Ep6r6Gnamp7FrViiTJDuUiAMh+u
CVItPU0AvUEQoXSL2HEpidNnvywZXjbZmzAPKvOp0YlvJIu3/uNW5SHn1TueOG+WmaLC75Lh4DOf
jpntsnfr/OO7xFfGFtv7HcN5cipEf1Ey2LeaQEdoGJsWR4s+vM7wNPh4hAXyTha0iE6FzueiGY4t
PgE6SEp9CL0xoY2Y0GDx04DkrTBfKS7CgoM70SOGTJ8Wgr8cUHMaZ9R1k41fQjOSDbKdLCmic/ck
+7sFs/5pLA9sX+o0mdTnVKbJtnVuKh7Kf2d1854c6JWQW+nOqABOGPZWgcqUD0Gf71UilkjjZqBl
2OTBbKRlbasWK/xWCDCUAUH12Mk84vKmphOtrFAKgq+iiemuY0psp/JLfdojEKrVy55BsPzgvAfb
GVGjUhtPDlTHPJCULwJiag7JOZIYuSA8jLIP8vs97Je2oGzq3raoo/0H3bObWa3yWKILA9ChIrJa
BS/hU0q38elIy3VKU5Q4k4u8fxxr2KVQqVV1efS3zU8W5rY5XwSh8ityTcNlFd0gY8gHgfT2jhhQ
lUlzQ2og90hrVBsmc+oWomyHvQ/u5MNdpWPoOYl0pYIl/phJR1s7iXzSKBziwn7nZJVHNmhH1782
X+N37o3yPgWL1YgDvqk5TfSY5mt9O78TBGL0UgwJwdgKEskAAm3HsEBTZE+iyeMKIxsHE636cq/K
AT0oAQBjH8MF88HusUHJgZZ5WpTTVABDXLLep9+Q98XDUtc6kkb5g9V5ba1h76aOBR5j/cVxCEbh
FvIkQoUP6aflihACK8wLrtMIU6zm9MLUU03aLS+JXQbR/kH/kYj8AEC37+TX+F9irZgKayivgtTH
i7XfGoxyR3Lbg5IlXUtGBBAJARAQ4NClVGvuN+aD7B5IM4d1jXuVp8qRoosiEZfrcP/NAqtPLu4Z
iTGeYUuCx20n0AjJVnXJADSsEXzSI1ic6nyH2LR6mMs7/6Y+DaAaOyI6c/PLDkXfG1fmM1FC0xso
+nvmV11KbF+n66nKYWl2dJnrKtJcsZD4v8HVwMSj9u60d9rIuFmwviAy0oHJQENgHS6wAD/u64E+
ZRHrb+Lg675cui74YRHzNv0xx4NP/xrAFFvdI+lyeGl7E4B+NWCqR6P9COQXr1Z1+SDOzgqyY7iX
H1KR1kNJ2mZPOKhyywLmexJk1y3IhY2C+utEYzgpot/dYA/XNR//5ECx4pDWaaDpij0WoGVu3FA2
LQGr7RYxtYV6dqyaRrf4eTgnPfC92e+MB3Dh+ItVjRIhwknMWHael6fS/uzIQvuE9yShqWts4Mj5
+xgXmCtLpqt4H6LO01+vlXBEpNPo6V9ljMB96yyJA69ZwWPO6NAOrW+B4EfVo50PrG3JspjV6VQT
rKCcda0ljaRWji7TwMYgz4D0z0A3sycYs56f8deN9GgSVW3widLyhl9UMCzw67RPDP4DEUpenpis
Hm4mx3r4lQPp65VhKVFtTREsSqH0iDFh91AIW3WIJ2oKTELCOjkMolk1epNmEBsV9He4wcNsn7Hs
rRFLnV6dYiPPFKBcFJ9OOkTvcfyOaZmtBenJy69sp9oepJdae70jJlnNIQvmiOV46ASidfkwYR/x
pm11xFfL/ue71H3jxpzzsREoFg5DznRrqDr5BRfpEnKG2nTka7W6y6TRkdyqHOjuJj/p2G37kLhv
bcqamNV+0k4Gf5EV5U1wdE5wQGofVQcrinFH6iF52bQ2GMwSNh00cE9rUf8Q9HM4oQFYu26tAJBO
wYNQ7RKLtNpFVrJLPchka/5OuQolWdfXLZwkjdKo3hOVoeWZ1z7STS+ZtORdGeCb1K8MmJ1kyOac
ftxTtHo5u0g28cflHo/nwRMEh0ZNCD4//FU6h32ufN9OEbnNJa4kZdVHEa7QzErDjv4qgS26IqLk
XGYk9iNE5HZDd384QzH73M25PWep7cBoY5n4N55Jr5+Vp5Mo8wPKimxxkJ6jIf2jEi8A+hfs/lrt
QlhVR22amN22V0K5Dq6pE7tPVYwBlq313KI5JEM/jt+PbTwFnx9hu7ciMR5SSpnvLKpJpR84Kcph
8Ohuslf6MlZXMGzRm/Kyr+b5g7kd5+cKiH+rt9dpl5ALFqXuuORCHS1EBysGVq6DvA8HI55+5zv6
FGcJsZlQib/VpWfPy3YZYbBGHTNvIFiW3kZOQ0+0pAmlUKDnhAhMXtNbQx0Gwh17/sNo3qDSgwlp
+px6ckWJ+ynZfXe/D3zXXcNS+JwBbL32I2cK1XEMMEb+eb+R5IPf4vnmFAQxqq0+OSzHG7UjFL7w
v0JBfmh4y2mjMhMcDf3eKndItjouEt08oyXvwvTPjWODBxNBokKX2ztxSQQ8VNKv0M4fjbhtujlu
7Hb7X+QnXdNqOIR4XRkr+L92/85ewx2cxIZqW7LKi8ancsbevK6OjNhFyzPCCf0/Aj4OWyBTJYnY
1SjbCgmxgIrygPJ6Xsx4EZugEHpzMsl0oU+athHegZizMBVJNtoywCElLqbQo9JEB3Hc8BZOI6FF
VXPw5I7PmnqOKi/YQT94MgyfIwrejuTTv0Xw7E69bJhRjyKhWu+hsBPZsyOdxSGnTba91+EgHm6A
sFh2uYTU8EMywP+c71jYwEvN2X0soyOF/S0iNc7oJRuSsoVDcD24Aa4WEf6/j76O6Sg16QtGMiyO
2aVC8Rtb7Hn941sw2uWImMGjqdi1ofk8cbkfWv/6NKXxgiNwf3/Ity5pS9RN4fSWic0p7GAduzs3
se48DmcvSiRmCg2VhuM29C1XPRJNSMpX0QYCfspih+YWqNad4LkdTmQGZwDkI1jaubzwBV4Bwoig
6oT2RIfTLoRzLSD6f3E6g/bC0LMl3m9xckRSu+Ms9cMOIoLG0rtANrGBI7vjXvhlMEeslIyNLmQI
Dlw6TZ2+kjfg/emdfvGJ5rWScWhnnIayNw5g+V3kRiyDFyenO0ortTwCWPxlLU49MfCqWb5qR9wn
0XXY6G5IKCrOUcp4dj/oqQQ2sAM9EKLPxB/mIu2mgM017piJB07kjIctESycYCqlkxjOsNnw9Rpq
toEhHsBBt+sHv0t9ScyWRnjiTn4dJE7C8WTnfWOTV+0xhdFC9hlJC1X65fhf/tw8FghYznEh0m9A
qYZhCdt4PYsdhex6lDgA2bt1ugkAB5MYlXhzzLCDbbDT3Azv6NOv7gHEplWdO1+MSfIENRHMPYFA
d8K5L3886jG/jg8dC9DK8DhDisbwptFp63wDFBNoLyHh4naK2HqlMRAigqqqSXMzN15TjqlBk3x3
i73lRF9NgfDWvFj04isJW02LBZmPBkvcsy7QajgrFWIMCOHQpwgKZc8J2Z01Osh1/ReZMWKRbNae
Mz59HeWLTW2OUMphxsmS+RFEvdeuAUto4xYPVrC0pIBTgDRZUb6YUOia1x3ZNQYQ5pzeU6DlKLJ1
zGadXwq9O6ouZrnmMql53p37RTrUEotQfg27iwbwpm2ahUoDbwol17qch1Lzm0g1lxg7d6s2zvWa
9PIU5WAOxhp7ZcWmHa8G/uurtZHsUUAvlmB4llrkyjGp4NAACRaIupZFEdKWw29iTv6iQaxQMPb3
mB7b1pvDbdQU4TX9kHCAflneKDUIWKd8Yf3GFF5jFYQH64RF+cfD3fEDO97Z9m/w5wK/ceo8Cuf0
phhhKESDJZ66yAodQKkv9IIp4Vtz0N4QJVmZ7ARJBBDEvMhl0++woFFCaZZ+Qco/C504qrTXGjbg
nRzx/GViq0Ns+5UJFn4BpJxflzhPbM+px8wsPoZL8IWuMCsCo8AQTEAPKFEG3zuS3H8ND6YP4Eik
rw7EOYVp0+Ae/1m+V4eWiMngirziB/Bkxq153As67hqwlpfnZPUSScTBxiGsiPewV1+uJVnjNIcn
3UDskgwpEk2ql7N95Ml93O7JAoJQN6N+dU7FWX22rXWBSoq9aydxa0w4NLluihaxG5rzTS0Fd9Y/
pxOpnOMRInqNFX7j9+ih6i4T5p87dav6qGIv9E+623GeF7XUNOh+bLeVyz/FOPeqPIcp6Grv6Aex
sLuInxsk/GJVrZ60VBxG9UB1ydscWincWj5mUyJXBPPB574jawkl2WwdABRei8YnWRwZmpZ5+Wgf
lFY9IbLxtoRHc/DXPahiBxgp1c0AKKI3bNKjTUjhV3G5NVA21WWSeAfRY8NTt9iKsXIFWxAllqCS
9tWfYZrkS0icMb8KQn0xjeUiHILATYQTyBtqMGifu21cJpHDEzUR4/YFQIoyHxIOjRWbnIfkuHU0
i3fVskjGvQHOz7XSnTckEi9ReEPfXuEEu5zZush8HRxmFqdqerV9VZygZJZCwLvq8ROmMv+Edg5p
Hz4jwN56XUVUwS4EaboQlYeUF93+t5PDJCLqAarvrGAphPqRpCS4JufnpKScwDBcwR7vyoaqf/x1
xq2nKzFRZHenGF2BqeJtr80uj2ktnm4j+00vbeEdhwtho70iZTeG58xEgqC9hLtvTnBg29aegNz2
tQWYiFGSRLk1cNZ/ddYY3VCQFf2qylakcUs6rELUMHbIriTnYH09cVEuCoW2GYNuTIxq+mlEZjDw
qLqLN9fMgC0XXcan/GpKXiZO2gyKhbm62nGwD6Z32q0hqSqz5DJ0daXvxMg6d63rIMoTNUh/6QyT
GcbD6Wx2Kc8R1cs6+bPIEKAEQGjzpOzSyxGGZ1HxsFQMGsBYWjVchZkAqkaDCs4v7Ii8zsdeWwQ0
8Kbti7OcTo6VPHGpQx0qS40ATpP1octeFLD685yqbZIrRoxDoMtouRn0h9s3xDmELonhou1aEdqs
SW75m8RuYYlX8vWpZ+b2Zb08Lu0kaud4Cugx2LwGx6gNqPz2mcmXR6/bAOEX72mXYbh3byVwyoE2
e0Qbi9BE98z6n/bo9acxmygllWYIhFKZ+RyRJnmQaI4DKrCTz5ifiy8Z6NhRyk/w8lPsAjYKfEsp
it+rNaS/cOP61wAnggtsWf/VjoGw4ln/bX5Te01vrfoZpGNmvHZSc1xLw+xrPjqxs6JmvyyRZFuj
/oLdTuIDdIGde/H9O3tltL+EtiB+FHCmMdZcbB9NHfLrWSClqORn5c683pPvZ1fDtT3X86gOhMsd
qiwqIv7n3FzrzzT/qzGzVqublkRj3SmOmza/hhkAniJFsI7W2UmvUZmtXwLYNVjiu9Xy99mcQUsO
A56iORWmuzHijS1da1BOt92tyq6e19bsXl+CLrz1oCaZu/9fEDvt0SkwRx3POvhfivdYQ68wVhog
EeU8wzdVt2O/hWBJ9dqGeqoPmJJgZgeZ1udHqcwcvJuCJYFBuiZ4JJFjSw2ISE8mBTsATXhmt7UD
UzExnsTnuQRUhLVjki0iEmX4e3ydTnlt9kNFSEBNTYYl5CB/gN1spLTAAipzo2kmsRJRL9RM12jO
L9HcAQvNuvmFxBC67aw59HGsljoBaDy3noEXbvGWXn3DzwbH2hBFJAyAxU1XzFbZ/IjuJ9j3O58O
vI7MBeCW2KDDFtTRZifi9/V/P7ToivxiposE+zeRfwFqGp20Y5Ic3iJukmW3uh0DPzyMW9DaB/pH
VPW8KD9ZIuq6QBy7qeYAhJX2tGaz+/jfk4oD104lnAE0nRJJGu7xiVki3n2qwyF0ZckcTbF968rY
fdyW0xlNBQiXHYPnuJJ0R2dPgGvYPxZTRLHjlOJMUcZs252xBXrXiyCg4xgsXthRn4GRTRQyVL9x
FH7lF01Q3GIpZxZ/ofgbVc1f30cDccfiK7nU7SD9CsvxFd/xOTGnUCW64bAGTjAGElYuheGc8Fv5
aq++H6cMhWv/x8mRFqw9zAxeZ8MqEQSgkLVQFlAR1wDFVzqkBJbS+FGVAmpgg5hja/A/km44ZuLU
3V7tR3xhtl70mjncOhWISntznl8xsX9jwaiFg6er2uWZTH9YW60iG6ctQNnlLorIOtjAXjgiJkwt
Qs0YlZ3y4UOj5q0HI7eYQ+1NVTV7f+52TKfVYSl5edICpe5jxVk5gUaPuGY9jdnidmrWLsEQVxms
ULR5CcOcWs1Jj/7ADV1SBVJeD8B1jD1aB4Lu9ZFuvTCTR6A7k8jOZrYr6u/JajZukLN5AG1lBBSP
EyKufppPnaDKv1ahqlQO0IMs5Pn1SRjm5ftMMWppP0DcK1CC6liXQfehWXGlVwWwCxTu9PxEUbko
JDZ6lJjCeU+nT+CWOymd6KzOlMCWOszdPXAMQYYi133yMTuZPttXc6BuGa/ApS9NeGZ2zEBKF+Yw
MdnbNtDTK1VxaPNpA7GCrvgTltr5RnhTE46j26+x3GkRuzoRM7WiTuitIq6MRrkg+aFzo71KAqNT
Cz9UQG5K58ZWkg1wYjXLdfoxHgT3zYhr1EMQioNUFmhvkfun3TirRc+f7pzWD3nu5c8c3Fx8HIQC
MjVUdZdCAvp+axeznoHDnFTtKKXY/CQnnyFBRQqN757JzX0x7YuZ6DXsGW+Z2zT9QwvDBqodOes/
V64Y5FBa/fms21KZQ7rGeLb+iogJwUwVuX/W615zU06mKBeg80PQcQ3cv2vMJnnPDGmbcpERgold
guHCArnkcJBVzGhcsKxwD+NAe5WsSsHB5LMEsIPkRkkBZiuEBcvjck5Ez5BSBZq5Iwxhzmv4INw1
HwKwdYA44BTYZJtpTum8EqtN1kRncbtPmdbjnrT+hr3eD+Y5Kb550W8dPUMKOWP7RwW6KgIOISPy
5uTCR9CJqW/p69VbwyX3re0b+APK2X+ZUzMmpO2ojSS/pg5eEaJ8Bq+s3pm6vbMn7TSZnXJu4tgB
x4cxTSgpaa8JLPtdj+nY9CQh12Gz1GI/RNNWOf2HqoMJ6SQ8mJ2zThduPsuAMWK+EgBRPh46+7hf
yOtptpTglEcIAl2BitQZ6qJNycXj/yXqYnrJfxm1jaAft9puxIqkaSNDaUvJ3I367OC06j/YmhtT
Audwv6scu0tyPxUZONDnF9+5itz2tSZoqQ8k8fvkrZ2mEdBHz3AaDc66GHzIWo8W2lSfxMLCaZGJ
KMOYE/WPQMgIdwLcWx5DdzASpBDPqFEThRp8DaOKMwK4p/ndKbeqmkz+7zYgb8lxLfGcAZcf1oM5
kI76x8yCB8qik4akGnDbXJxMC9geHavAu4KAEgW/k5t0cB8BXgh+yw1Cai9hNNRFdQ683OU3tpEX
wvXtmFuCFXl+mJXsMGMX8VHDSwVHbaPpjI4i9dJUz9SDBpC63I7XtqviiosieE8ESnHy48Y4yeYI
B/7ES+XyG6ymAuUJKTBbUXHqulx0HaOT6B04JmvEMvJ7SmiKsTNowyb3XACqgMW/MrU+lTF+uVTK
6O/I5ndg+5XP8qj82TwmwLHCuVvj8R2/diu/l+I1PWsTXbHNjxyz/uSO3/Qwk4NAAnXwokrRsQx3
7srPxXpPqk2WLz+FWSTc6/OLnUmI/C6gzyPhwlA/NjdOqbIKyYonJSvCsK2g747oARHMFhiaTnDi
p4EWosRqzi3GjJoyliN16jKHR9MGDSLqZXKI2GaaJCCJFMPvpErLsneL3tl6bMNGMiZY+yqsCvda
9368Mu+09Vj+kLqv9O/I7XgiD3qfQ0T9rKdVZ5hM513ATyTxb9XSa31TYYRgfzlCzGqcjWIhYCxJ
Sku+S6rfxDD/LA/bkQ4NMTBm1ln18ndO4NxgJq+N49jJ1JOqmQEC1IGk5KGXI+j1AfT/Bsk6uawF
NHX+EZjmsDqBIlW60jNR08YSqhtKe1NNewKMJ7sgAzALl6KXa01rZqrDrTS+EGnuTtGoa1OgGJGH
TXf2cmu8nNePCYO6cxoF9qModmD46ze6OKN6iHEMaESq1G/1DC3Egkry5HoTe3GtNPHaUqXXsmf4
C0jfIM7CwcRZlzMk/+HW5MOMaJ/73TsbIoFYvGevv5Cxk1yXAGu0K9TOtqYNqRbUk5W0sFwSdtN6
GqTBnGxw4KombGq8asVGQpK+e1n+Ttm6EgpZ1Cba4OJFieEabeXLFbS8tDkMBvQA8aA+KKlBn0Av
Fm9jmtx6OA5EWx/NHRcgoZels2wL00OJ/tD/GJQfnF8xuLFScOiji2QUzQQyEV386DZI1DlmjAmC
7jmAGbqrGfJqjgLwjQaMn6JtVpbLpad7onCmQVLTVPqus3dDw7LA14rAjnfHh4YBoXGWsr0ghaPB
HSYPm4mkzODsIbYxhRcgRvDPLhwHBMj9zv3/VDIrKip6HKXl5KS3sMoLsR0vVez1P5Xkd9dgOW8I
hnzxr0huu9zAwAsblIAHGQO2rBX03D0a5OpRpcc4hiOBIuXrQIsBskx68fwLlHwBK7T7pYa7rOuM
OTaG9V21kqGLkfmkbj7Dotc+FzutnMDnBXgfcSJc6y2pakKZoNTZpMwXOc0EWuSFsp2mNKf4bHnn
1df42IF7JrgA/VSQTbQlA0yOdxoiboRJ4+TXwmBZoCHQdNvYK/U3CQ18FtV0xXsFrLAApQmupXtl
H3rHyyngNR+55gHDbMUQaW99FcPT8V/m2IX2/wzYtMxlhRkovk1IoltXrMq/MSF7sndqnEWAlo7/
OLLfMXyL2FDu0rCHHkmkXTAuatE3wwmqLIj3D8mBa6LJAgN3uD5LliXeUP7HMY1f6Fzdt61rWXZ2
A30a1KnjSoiDYsMLc36+9m0KFrhSmC+tSltyZb33Mc5Twp6NVYHAVkQ+W+vmiK3sjC85EkvK0WAz
leRHfvG12hqwMIbUmEpLmQ5ddMyNLuU5I3L9SewEt6OjnLTDUyex8tSrWX7QtZMLGRyGMVNILNFF
8tHLBpfwiaGVrctN8wxTd/k8iklWIF0LYgx3540J7FSE31FX5xfqNS4c7Rferrq+92UePOCplUbp
VGoE31hCqyFvBqEZPJPjqGkbiuEL5CedXvyzfkKvkvatCiLw/P5qNYXNLo1fubd99UfgkS+NyTA0
k5WZWxJmq3W1yeVlwthpNEImaOs/GxgPtlAH9qwgITphk2d8/79fi/RcpvqOZHvGyvRl8cDdyNiD
lSM+JB+OGYKy28HTYDkvX8eVJqOoEt6JVr343TpynOLMyqSOE4UzCDqlfMEqdRWEUg9M9r62eKME
Fme67B68VDZUMI1GPiB7sjud9W+s3MdzDzdi0v3XNTM/A4bHLLzSUWyAXFC8h6zyDRqdcbVnKPE4
nLSSojrTAaLOIH+WA57nm+9yT2zLz2tD8/zZvtVO82p/lLJ8WS4aDCokuxe8U1r8pqTKIaPPV5f6
9xRmb7S4h+qeUigvnt6kyJIEfiIZCyG+AUxCTFVcBUs9RKvOnrkYHgVvJmEK1YRl7gucR0jqA5xJ
AjhySm7V3ys94WtUCgp87ntJLEBjhbbYt1/tFMPUhPn6m4e0Booc2s97JLZOrGQEoe+P4NkETNzA
fc7yviVsF/JMwR3dVCe9+TjEasRyT6X+nWlKkKh3vwTRCbbykYVCOK0oiGqrBo1Q30yy/bs1TImd
hdsY2DjYCcpu/nHGphklHotuMb7D9qMopWNv0WZ9++Eo3d8wnRWWJBaguMxYRejDBoUMq3VqUN2M
hWd0497feMBiBFGS29HcPprAnAXXFilmRU+CAMwceLObSdVDY8zg9Qy+orvpWyNN+GMADZw/H2fe
x69bNI4nH+An4bpQbv32ZRqovvjvc3vnHcBqS01hjfAzQA/JKLUFwTQuMvIFpLyBU1MPlh8RNf0X
WKfAjoAhfJ5ALbFDsP/R4nH9+knF+TX5ytB88ugt692tQ4KX4Z6azoW/Di40kIpiDGDQlqkpsBNt
hsAoKnjoMXB7px6AWnbbXPK6vOpMOJqwshzjY9ZU0CcNyWLPMH+4hLbEDrOMMf/j3SeoodASWHTO
xqChfBlL3n7rZ9GAPwJrgnBaU6iBs8+s51IBfDji3eh3GG8EeHZTQhR87qkrfb3k0EPBrMvBuAHD
sHT1ar3QmLkACu2tVsARYQBHAv/7AxDXbxVn8CThEc7ipI6LDuybe3vXNCMtWZgx4tshR2vA9Fog
e/jpWKWSDsm7fzKP4ViyO9b1CQOgGxrM7nVAwmhwxvJckDGdm6p5KL8tgqMYXxfvKwtENAofxDfa
Z6/XugbHF35PpT1NY0onhB5/QBlsbr37NWBLG2DJ6mboX1tYEKRMhJHC07QR0O6dfXZi/Hh8UdAl
3fweTVi1JaCCm7Z6F1K1AgcwyNNPvnHwqHV8X2QV7/Ylyp4UbST5pFO5PXruKPqoBCe7Z1JX/YR6
VdPXhsn2ff/fZzr/avlMj+P1bRJyCgXMM5MSqqjwtAfx3RlnTR6CSGfBnwqTO6ggMDwSOdwBG2/v
wkk6DpGpyG8b0Nl5Zekrglf2FsbrH3Yikuuix0EPiYlkTZV5dm4m88VzzYENVr5wHPX2/vR6xtOi
1Q/rUh8p6QC9tXxPlV1N8AuGTQmLAtRb+THPJK1qKXyMiR/NMFbRXCW7RXEG0CbFJeNxQznvB6GR
pPgO1nkxxIF5isZMaQhKBdF5CDiuzFLXFGcCkzKXRJZODwj2+BRcWTWj/NfbakDGL9uhTMbTzfoN
M/8DXx0W0BQMN7niIJzz5vC1utikNmCc02l975dlfNhMBC91XYEhkQOefhp5AgiJJgRXX1kexwPz
OO9nbe5rj6hgGXNWOz50PiYX52MIGiK01X7kjd6/gmHxX4cf7qM185lQwTYUTotU7gFNSHJF13RV
7BX6kE+04avycc6ylouK5SIRWa5HDfpMWO3Rw4ExhqoG0VB/paQ4DgPuRcKaO0avmkBLD32fDtI4
Vw3kjKgU9PHhUyixn9bAcdve24R+HaS6gvzEKaISBZ2uwTbrmy2xjSeL0DG7kC6t8HDUPCUuO3iO
nW3GO75XDahkN0+dkp91Lir4k9OD6GA32upMlTfM/GFIgKKj6r8PLlRBXpyF9MRXDceu8vjYqw1n
E7i5HkgDoaQo0ZvpmKqnrVz/KvVq0Gr82Y0joyUBJPCOonFteTHVJk7XXBLEzTZ2uyjBrXhYzwbQ
dmcwGUWGs6dERbW1aJs+Ty6wa2EqgoGWbRtiQ+gMw09a4UqpI65zzkh1Klw/Cj1dIz3W9j1+W7S0
itUjAVC/vaaqhTUsCVkgGTPkyjIL6ecpvA4RB9/1k8gn5WjMxfkZYD6H81QTK/+nZ7n2XmvxMG7/
bVKgWQrE/qX25prGcjw0eaVLJcqLjfoNrmVJ2Ot2wCBULzR0ONhdPOyKkbGUDeMMQ3cN6txlzLux
e9Col5VyKpjhTZ8MDFGKh0UV92jqqvOOENi+a56bhLneY7TaS625OrnNA+q/MAo4k29qRr8iNiXP
czDqjHwlr4eZLUmrJe1x9o79f73cd2D5myXq66QyUOWhRO5jEWoElK6AsDessvP+GvMsK/okHSrM
QkBIlmbFVl6RFzGCWBIethqwOeMaWzjh2+EUyxdo1cRcSelsjxdkvRClFNtDL/Hrua/exB62fyxj
zSzDTm54gBdubPctRDkwbykDhoaeIekRe1i/fqMwnk//MWbVcaDHnTB+gYr0RsY2D6sXZ26ubFQ5
XERsuI82EWW0fK2EGr2iBVF53f1to/lcQyeyexb+bTku0CiA6X8cC6TQlz8J0UyjGHVxHrJitaWi
kg3aC83VqeHTiD3Z5A6t2+V83WJ0/dXMRJhGIcYbTyEHU4cecDv6EUkHyWftiPnepZNxzCwNc15w
GLSjKKLk3X9PVRqKYKKc5ARNyREIXKODEvn/MZ74jgLAkbFKBs+Ugt67VKfr1yEAjOM1qB13Tme+
FZ+lNlU8IFZAZmHhjVHnDxl7f/EZZv8Ii0Lcnl0zaslBoJ7+9qtvc5u3exNRAyaJIdr9RoyVsl7K
QNaNon8AZZpx4dy/vJMWy6mrWPxeDzE0xYI0T2XEJls+jdgPHDqJIrpuzR8Mpy51TLGNsq36ACq1
vCIEQR2oJmIa14O65Mvh2lmvAwMy1oRrTfKVtCAdPpVgDXLXGctEen65W3EcorQP1BAPT+9/OiEF
CmYaQT1lHEi36PfrQgViP11VbQZsHCTmV/2gp8BW7J7/QjkRgMqG36j29k6WQC13vkYCewKHFH40
kiCS+E95LKc91N8B8duP6lEWjTJRDCtyFISqNWckSfg/eyLSwjYuO0wy7Xq3OjTtG3zMX7/zwHNB
RJros81sNbNUFKCyv90j4g01AXfZn0dgp18uu+3UxaBHAHZueHkx1lsaiHzQZH4kKMrn9l2JDV5I
wdSRn9iOwE4TP6OJWr7aLMXofw98LYtpQ2UedR/Es0lElgKfkYze/TitW7MD1beHEt9K69uXBP+e
Ml69x4c1/4fiMU2DF5+jAPKgO3GOlTLDI8Eba5KgNQuh5F+x/NFMja4y0/YEOYtFmW2ye7+Phiu9
d62bEZ7QIkGYuIOlmXy3vl6Gj6zPSZCie+YUECGd6HTaFCeZFTRmfQGKt/QlmFY8d26jS4ASglNw
/MQ0TkiYsEQ1MDoOJwjKtp6s68fzDeJrBZyqKjkDRD4Q/5bF2GzC77DUkopbknSDJalSkylCq3Ps
SQNhS1sDe26l4Yc4MKifgLWxj+3aNmDPg4F/JC/Idq7OVGuvAPD1lB2SeJp9H21+zmQvk7Q+6C53
Po81LEWKRT+wmN9qLFuIdEAp3vHMexelUyks6mackjVhD5I9dA8MS5ke5XnqtRDcmi8jId4SWha6
INDqRTf6YoQrx+SrR6FF2WDmHQkJXszQNX6+pATMYd//f8Zi2NF6XYf2IXvWeshf+M7o3ROpmG/F
xW2LuYaykrUmrXcf4DJZmCpBikMLXIrXNLrzitijej8j6iVG2UYtpEFJQh576+EN3h5nqkHL2p1d
MoHLSaCGJ4NqqKWaoxmi5SWQAuQSHv7XKanfsvl2YRM5zIG2g3ThhZY/Kx8URl9ue4nFdR17bFoZ
jJ/mkcT1uhJyLi9ch8qbDGTLuYLVOJo7Ggyj7kpx4HR5WkdCK/AbSf6bZquYX4ie1hdwx/YllvPw
rkVsMG6G2AulqrYrD2bL7yo4DoEZp9KKvmEpKVVw8/0sOFVTJ0B3DGfBy6p0nWkRh23r/dkvBi4g
XdjuD1vReJM/Enzg/qpIGRMv1iBvolEx/aK6aDOJIwko40LeFnvQwgM23v0g0QemxauSWWUTYF5Z
fHwRZKJu0c1zEKRNExOVERL1VPPCCF7NtopvXQ+RB/hFpzi3DcXRte/yaZsZVL53B+s2w3lgkF/4
ZmVZVqCSVam+qpO9qaw1PEXMGS+gP3quoT2zYiiv3QoChqMjYl9/jDIbY0qp9t2mpLeWZExsmbFj
bTzQ3D/47DJkvrY7N1WUdSbgQ2LTQ9ZdwDwJB5Nx26O4U2zBeBAkxe0pSs2LKC4ipONSMEEWlWm8
pXHTYObpzPjuhpDh08djUi/D298CQ/D0n9WfANHIIs1ojPfAvgZsCRkRImouOK8pzg/I757gGLsM
vbkng+g2bCPqUiFUhGlE140/1yiHTMBZUscb2YUK6FKHIKi/T5VnGaglhARjA3DkRVJbMKXFnE01
Jo87U3mL+4WLn4Y4D/cYouZPF7U6/hm0gWKzLulm3LhHAXVh478FZWw/mckZ9yhsFgGwBxud5ctM
4JJajioNJXIItq3QYx7jsmHeIujsA3du4ReVfpbLLrU/QBFdh23DH2nCQ7HPHmCHyN4MEKqz1vl1
LFu6OQlEmiuz2LcLmBhw0yPyXjmJzSX9dIAw096cEE7gGFU/L6H28BEJhhk9lrcKjCx1sNZX6kwO
lcOwG4HQEjDgWck2Ay1AuAiXuIr4/Iopc1+3Z1Rfv8F+eWLldZgAFJw8EtkLFtALtO/3oRnHBSKz
ts71m9lTlzn9DGPCqA0Ps6+TVU4bHnrhAwsauGmPAEC1pCsxusKQI+gxoUWrLjd9XZO92mFvv2dO
j3L4s+49uQzNZmvel93r9x+aOQnVQL804FyP9OQymEI5pwqhhhY0LsUZqcWtl9d+wSB3bbgXTBbz
q+rBTG726y356dZrtfTYCGztRB09aIwunaKmWUl/QlM2VSg9jjEumT0BUYRqefWZL9IIABJ5VGge
Fi0n0dsyABlkMOGR4tMpgGJuDVvy8eD6/GnXYFv5Bc+mK3nHuy8/IRaO8lJWxk+txX+G5tkIeMww
iomdoSy8wNOU6Uh0WPQWm6g24TE1r0ENd/mohdCL0kMVWKyfJagmUXZBLweb8J73a6HP9STt6W1B
OpWZ6bDkTBXc4l/NR4OHOdOmFqPKWSpiLEIILj2ocep2QlH8n85X+QidTMDr7aoifEDSnawMocrT
6a2olSvwWhs7ahUVUzmE2uqKP0cKErdOFHERJsnA7RoI0ON33qTmrnHUP3Hmy/TEWNIUdGnOsQ0S
DBmCDjiFiJtmOq/Hg92q/YENGFfi8URyIrWikA1m3yPtvMwLhKaCMGkMM7rqAO02oAaloscq3NjY
HCSU8IvwiMh40izmQIEqfqbfbv7b3cqx9WsJo9PlvssK8RnMJ8tjahnsUzhktCVPuMJSxAnzGLzJ
yi15F0/aLnHB+fMxmK6RfC2HJ+1Xe2bqhartV3cUOufF2sJFDobEr5cDDk3JytQEqIQSVBzCwdlk
zU+YXK+0UIWlvfcy0nTGn1O/3fB6gYXtVwIO1iKZSHhWW/maLYlm4f4rA684/qt3hxydFar9TDZC
hS9pBT1La34uFMPgxzuJQsUKr/qEqQmUqae9fNIa2RZbbt95vkkRcCEs7VyP7lGVsWqSTye9o+KC
Ipt+Va8iTjSVV8Y5n/3alaZ4I5gxPOawFzn2YyPNcm/ehIR8Oy0oHXUj6cwhjLnnnX3z10wLA4SI
PM8ayLxRuiky1jAutoi4O+rj5FaHM1u8u7VdnCO0P1lHtNq4YU5lTfHKoxwRhDbXCiRYLkIe6q0Q
PqMeJNhMa5Mri+Yk6VVKrJpSoY7rCzrUex/AKq7kF79FoI5NiheHD1Hd5tEcgW+LSXAeNXnV75V8
wRddoa19+bL2NGsa+u+VJWtFaRMt8HtpeeGB8CkRf+fy/0fIdXqS5bM/3LQtq6nmaQ+F6UN+zGUf
qmW6S3bF9UtAcbsYwkv/rGwz1/U+LF2KBUwX+i1f6yf1u2ERbDCrVjK1GNtSU6UY0FIsX1JDKjR5
7Dfkj7OsPFKfIezyND6DHZHlRipaC8Qv3nCNX7hiOXJA77nwd/bc9c1WXqoSFqdB38sKwg5Ofn6i
gaMxnYWDb5at2Xc2a4HWqqRCli41y01KBzhk2Grdqep1gbSzglO3PLHFQ1MyO6TYl+AafkVt20LR
NrIIVjnJlPvA1FWj/pJeCmAwfADKFqf1097XsT4lTClx0P6ybka8gl+WFyRiLLeQjqLCN7W2Bddd
YDnC7xOZ9hU6wRUk4WjcTU8xdDVD+LcRHdfuGUJmvRhtDSUqVAFWmczs0etfu8Jb0J7OigPkuSDY
cAd2L2gP9XjDl9yniKUci5Anbbn5RYp7mA4jTlEynJ2MMXJ/tXqSCe8dvPbsqOVNlcH1ZZFpnGiV
u5QXyyP43tlfpdJjZGVNluJMESzW0/ZsPpOS0D4kfL/RkCvWWeS9kChOOQR7h50/vqz5UpUd+2rb
VyLHxC+LL5MNUOn4uMKhf56se2XaK3NIr9UyK/7iunh/4iBUUjLvGliuXgTrCfCUaEbS6k/aAbGi
Cuk0h47wFO8/VQcFGeskjl+9gkpdd3iHFy8QpSMT/of4pVotHh9IV689IzAvwX2Lr87W07EoPwOK
6YucwZN6urS5Yd1zJo9vbzdwdH0SI82K4CvNVaT2aCtxyfbZmozQ57ELDflDAiKDVix2EaAWIPYd
yLOVSFRvmUhf4TJNBCvKtjSm1WJNtm2IqAhowpOD3hGscHOP4vHA4QJyRGBfzTEkWxxgjD3Jmfu6
4718eLwJ2+4lxQLRgudiIhUJqEYpyVBzQ9ht3Otb9CxlWJKxy+N4TABCnbKMSPM4Y1Mw1AK7R/zL
uJzvJ+48hqOfjqO7ETdqQQYAjtZ83qFUGu9rPsld9g6w2u1ZKZCiVZgjCLV1RVrvl+8rmrTdFacd
4w3qxijhFWj3VyWUSDJ7CUK4xJefXW8C78+i4+NeUP7+A4DkFc3cDRFjhrwgcDF0hJdmqMlmiYmy
Bq1bIrJtEnuct7ri7/jL3MGJ2voHlshkFNxUeClbZyTQ7JDx3c0Kw+UulRe45xLkUikeE7/GXaOE
77OPL4NppNAQlPCWMSnCgVyoO87qKY8TGsnWBU+ASpwdD/nOU/eqi3jQR/rrBEyeNUgDUtiN+P8k
SbWtTgdxKe/WWaH4PEBdtfjTxhZJZcI5nzqp9ns1G+j0cdphUk1eQ3cb+kgAI3cEpv2un8qX36FF
d0uAYuFkSbAh397uGpykyYqD2s0jAnlSosB/19CkvbF2cXKvzOite1izd6YvR0nk0CH1FFUPfymC
VfclheA2dZs62iO1TW/eF/td5TLlJRELcKxx7ZopBUD5v/RTAAZljj75+5r/bhKHWpaFQ1DS9q27
0EEvIM0w1g99d5WS4FzMeHZ4t7x1XTptz3o6zB+92LGDt2gBDbo/+fwqtR4+XFyZuTZmKa8L0Bhk
RENAMk6Zu/w5DqgGABTqdq0YRc5CiVcn5qWSP6GoKFf/gpCpVr1IlEkrepjaIyA6ZFtXbuPLOKpu
0cWhh9Z+VseRD5xRUE22FiaKyMnA3Fm2eO82h1JBBP5onWbovqhHTSptErRyVu4S9xLeBE4lHWgH
VV6J5AFif1WNcswRhhS4j6vUSqkC2597uCbOpFclJ690cefDNGxQkmMnXUFl7w+NLvHS89OInfjf
dqC8Uk6v9vvZUTGFuxBK1l82yZ0mRI3/lthaAFmtlo1myrcqc5Vgt/LY6a6xhxXL73SnqIgMkU/i
UABrYeAH4x7DcWsAR5UeBv7PLZ86L8kDvmXZVfod07KqoMsRhovEjzUl4Tra9C5FLsLh68lOgqkL
A8EcM4+DSA0OfWKpPiA03rnybYbczHnXUq3gVdEKalHx2nx9BDSdTIe/5LJg0pF79iCHnDLM7Hn9
G4Wa1EnKRTQmwRQBpiOn8ZQM8CaEHso8s+qLanTV5Bo2Yh+SDhyoN43ZJPYgOdaFXmBEqm2mP3eQ
nSFSydFMup7ZslpH5HXFPNok+ONkFtEoxazjmMkpX/p8JJ1a3JXO3YhtowYHPme1chktSHN37kEF
+JWG0gxEeuiFr/CD7sm+2M6u1CrHhB5hb4sxXcIPJbEiDIF6EuXnIZ/HdOMECUEHWLYybAtrUif6
gHcxNkhJL+SF3TaY94IIbqezftmkNwlNUG6Il++dyO2E1GV2Ox9zdroN9JyojaVX7s0WViXM3oep
SeP+wc3CSZR/ccCwZmWf6TvDI3EqOqQj9gpSZ3IdYE+Y8h8UEzhXnJ11Kh7NZz9O3XdVsMpj7B+Y
M0tiuK/bOSfVWHbbgvJHmYCkySyHHou8ZbaCJcez+jhqorknD9h/nv62Y5dXve16FSri2f6TPwL2
JUEGnE3lsiOrHFUtK9VHEXSKbek4IInv4RHpTmVBU9i4KGTsSwNEX/SrU5/p8jU41JpSN0wdeUKN
kkwCWfNJ2CZhARMC5FapoJ4goNK5rsMUHL2ScysMb5xjY0OdgJcglmlCTckci88mEVZ2EC/kuPke
DyIsMJc0Ue7zUnke93QhxQd874+gSJMRYTq0h1mtnBzjtL42PtnAqpWooqiR6pRmmcFwuK6mbFbx
KFDzFZVgzAEMeWbslP3ss3JsDGZ2ZzZEmL2lhP/6Ny6flWaByunpFLHUWEK3ubfcZYJHq8uoClVj
4N+TrQEeItG/WbYGWIlEp4CdVgF97VwGtq329eIoumsZVMzNsHfW8JekomuPFk+VDTd2r28t9i6A
lHC/FqG86u8alIbwNZpSq+oysNcwS8qq3+oBvSfjgdtlZdF+YRJF3YZoFDEN+JK9ZyoSCNSSeD0u
wW7kynKUmZkYVQKxg0Rcc0/uJRJqDFsDrPbp8BVYwuoJ2r7yxFts8xCkGDQQIOOQLQIjPj/2VSOz
XbWIxOpgFGSKSWKfAgKlu9Gx6meT2Dg5aEydtO0UZDVMvg1UW4uFmo361AOttcuEk9CtqlN+worU
ggHCptnoU6rCufD6cA95sgesh+dKCwmoPyEP1iBcvx38S69hZ+zDiDX4WDN3d7LSt4gX6gpeXPYU
PuDFU6GOtCUddU4IHk96o8s1qJjxJIc7JAPV4Y+Ly1fHvKfzRGeUUpvDxAsuQqjI9o5i1VRbZ1wW
KP24FeWiP6GEHIbjY7F562X/qooGrE18rIglu2mnRlYoPUTULIqEtwqcb06afD25K17LZQl1bcAV
+bH2C/XAUllbfi1hbTv8Au6n+kbI2ygza/oopNuR9Ku7XkNAe51ucSji+7lunv9IZ/y4UfmFt5Dv
XZ2GeeMBovVFpIpLJlGzqaG+xS7lxICrZeJ1HRrD4dw/iuv68+15P2OMns3WZvSmSB0IuODOfqP4
LlKYgdplaq+GXNt0nRh6Qt/x4L+zduAruyKrEPM3gGc2u5luuPzV1DNDA2rad+WM+b4SbIrqyIqE
KPwDj7qrFHhzdZO1ZiOIZurUBlCXPpftihgDMKH1LlENbCloeindx4zXtREwsmOrjYZFIAFARo14
19NNAN/DU8KepJBAx8tvLfcTNMTBTi9G4s2uBBZopdyV0ztj7ivnKPgrYBLbgIQi8BOe4wkwU8rQ
RHo/zsHQ+zAmmMVldO5Dk95p8C6Nfvk6B3FwLuyp481utMHzyqCgCFJ51RxtOmGYUhDHX8CRjzH7
z/1AKDYLVfIsPRGUr3NZr0zmGnm2UFyI883dXqXbnAOs6v67XLNiE4m6dD8taO5KkVmcmHD0oZMw
vHEja/rk7dSSLLXf+SdcQEPCTt3X3fpWxGZBYLw8p/3hz52CITYqvmB9tKjHU8GswrIYNPobpu3M
QowOdvoCH8I8adTmHmuOK9chLiJI/UhHgmRL6WK1eJQyB1luVAYrUOMBkH+kloOXhjMSTKst7EWI
fTcmfSKLz6xG39S6ynitZUQfJOnP2Afga5MVX/icQMa/4YFJcwDg5sBFmOaToIjQ5D2GWROAw/AE
w2O/p5Ez6edLQZbMR5ocLbjP85fQtIjOlYPb0ViiYZHEjK2yE4sht0mrgxK7eryW4+PS57/4RHKH
IYOZjWkEun7UTye27lsN83nEtd/gyJU1RkxosvXN/7zLSV1KnG9DB+WpMZ0Z2j5F3XvdryIhirdX
E2rBSNin2scY/QYjUStN+6nMQth0L8tToalGn6ddUuoTIMWc2bKaYHvihSzzShZV1GeRorRQzxec
ooWnkdJQ2XnPf0CzZjckv76go1BDJmCvgAWMWJsMAFMZSFIh56NKyZ9tcUBpmR2ltoU/ZOZTSD19
VIarOqsVA2O1KROTWUm4tYdiD1iwA0So1lIdKbzQv15DS7qmP1mvPKKS85XdEqZPrNVb+mSZuHl7
TG3J0TypIMUQwGfuJ23tnFdMuV5xcX4Bep2akxSOs4mILmTf5QJ4U4BwokQ2vAIFkVTw+MmTYyq2
QoVmpnRr61LfCdGgVmeXJpHA9wiKDTxXEb8BWFHhcHJokdakXviy+G6gwLxQeDS2HYiuXRIRq5ug
70xgq05Z+Rf7C5xOOX5nDfHzM+3Aari/7P8CSKI4N4tIIowtqcYbyehKkcuRqOmyd66XwO32M6v+
DE4Zn9TKV3CgoJDhpRpBpz0kcTbS0wLMsKtyHkFEeqtUA2uv85H2fpOlrm8CTvReaMe9BuMQiwQ1
Z+Zrela4TY7anKCC3h3+Ohv1YT3NW8kUD5tqnN6Jh/7J9vdu5gWxoxsnVc7uVxI0hBMq0lBaGpn/
femyFIHzM92FBrqRkDesdrkeH0A/KAmYAhst/fwwe2MD//ytCRO953Wkp7vNqc1d0ifn5wCm5KXT
X7MIenqae2B4AoU1NRwx4oah34fzCwfW0hqVXMn5yzq9WTuOpQ3cbkhsrHObCO65Lu507hTMH+fb
8Oac/Y6gJICAr36PBvjWnGZUA4zwgn55W1IQ+FyCwHS7l4dG5XSlusahAD97YNSKq9OVLwSHS7PQ
r6cLWf82crrRZYQyyfAJk51o2Z3Z/wRv7mY9tWsNWb5iXRGhxDbfP0ztTDHu0kHcLgeZcb2rrPW8
C81sqUTxfJcOXPlR08AEPRHQfEbrxGA9YnEANr+o2dtTS9xHSZJFkp3BPPAIyc09/orrpHfDv8Kg
P+kRpuNiJgulnnOUNRkk8JX8WH7b/I/UTSpOruGKqPasqG6vsGBLxvEjoPu2RI5XPPAg0f5RymEZ
vmj6VVscnifvbWAGMT9pV36exb/uAdC6DWuD3kDlHu7EaeavB6MNXPoYmaNfI99aLQkoJrMqwVCk
kspyShcDjv183N9k0vCRGZ043ET6ihE2z2wAtkcAQcDlZr0bUpS34b25R/W/Qelfd1tlJrsKWOpH
ElQjjqRtWEycoyt4eGaa+F/YWKb16259qjSwq9nVwusMOPWORFg+lv2C0BHtqITLbMQS4syH8jCL
YAsXR/l7vgorOY1YNBFnH4eTo7XRAcmBqgKc76FJfIXouQhO+Kq33UmguqkzDXrp68yoqKbfdMGI
dTb/GXs158YFO6V1qOEGd10RvIBuL6UribsWvhD2rsFOMX8n68doGsfypK1X+kkWylj9pX/c18Gm
fV1O9QfCznc1mcNuWeCx79yUTaaKkpkVTVli/esG1onGgKPtf7ei9dcZkhA7IjTBbOD+gkQ1pTAo
iRfgLLSP1GD827rQJ0l63/G/X9fjnzhOr1l0ATwU3D4SypBXEgWtteaDCPDFGD6QbJk8lj5vaWQ9
vbE9p/CzJluKOrbLYNW5iAk3ueiiv+ArQiH/Si/7BFad3NumF4nIZ3eFF5Y4rs1hpqVHubd8dvrn
nddcYe6NSb2TSqFsZ3jdLptYzd5Hy+ad7EEu1TrEeH6AIogs3t2jP84L9EryinemqyTkmpNTHjvg
QIUcnY3bfrMumAmrRE30M08Pgcoawtqua5Wz81SSR+k66/wGV5EO0GEoL9mHmWUYAk5jUnB1TURs
msFskF26mI2wz0g8sHLngxGUMtyrFABETnLFGwBtz9BoZC6lZANSVFZCHuWs2W070PcGz1hhzihN
ZW08Az7dexwJtU/f2xG+6C5Ogc5OrdXZVqKU02G/Ejngukfiizzed+nGZzSYpdPom5sTPwBPG0j+
vdLFnbMqjcAA9K6+toLmAB3YJTqGwbc3sEmv9ZntP7KJue3XIBgbBrSGmBGTKyJDB0jOixY12zT5
Ajz8WX6zzEpYIygdBfNA9dM2b1k60Bm6M9wXEtBRt42CvoD76i1oJ1YIqptf2c4Og8QcJDlkdzho
dTWvkJB5OZM2Ftoopg/FjJ2kWEGMCJqJOBZlskx42Jr1cA/t5gATsbrRtaLf+xhGXx9NfqMy5Cql
C2KWBxGMsSkj6snkmWxhjN5JoQsK1guwMWCUWF0SrMW2zjB0z1zWnnUcMqFodFTOPmsSPM37dq4b
rn7c1DGvZOomWEPNidTjhBqInsrtIUukpscmnic9cBGLs5jfED9RRQa4t1Bh5htv9pZ+g2eNfYaH
QSnuN9Iamunk9hdvqRYBekS6ZRNWR67L+Qa0XRet8rVf3OTcFr4LfIFAeSSVsE5f27qlweq46dl4
2cnARkKBKblVxG08pmdfhTN3BUGNqxgI9Pmvj1gNRV/tcp7U0H0wknhmjwVxUA5r58ckFQwEo0t1
YNpwEBxmPve6VdjDNv74WxNFxOnDvm4gjKYCRZPm4oMaDBxFQBY3RP3I8XrerFNkeIvdXEPzPDtt
7pRrdJ7qLjes5kUuANNL32Duy6v8xDWkJj8nPC/+N7MBoOtuBCwNmXa3kx1628kZV7R2cu0SYfNc
M3Ytg06WzWGIbg+KD0UdyjIFKpkeBBSxAHjTlJbcpFObk5KA/C0hBUMpT3M8JtJlKJ360mw2cE27
Dke8dBFaAYI3RBRmhBbxGnFa86A1YCCREa0rhGOxHbKKMb0SyGn7yNl+y2d9Sow0SkujG1fYc1bP
7qiivvIhor4W9r4wH3qAibCf/oKBxEVoor3gHcnvW7gLoJOTzQ6HtCHdIl2w4DSVD7P+SM+sxK6h
Q6MFA7SqIFxcaulb8+AwAWBtZhURgvjMVAgN0o+wSJYOUDCInBKgzDQgGGmAPDsrBfMrdzPQezE+
dRN3UUP6xvDOulZFikvmU5qEgpi70iczEHBQUe5bCe9a1Y/TRQgJsl5rxTFck4uiv1VPjrgNYUpq
/1r4EAk/wXYIKlvXKG2UJSLQOM/rK/FM7r74i5N49Sbp5xtnScJyTYGsW2YUZ6lWtCfM0ab0ttFM
L9hx8Zre5Zc5iCaOXNqJIJxIYP9QWJDlm4O4g/S7+YdhHnQiyP31sH9DABbLqZXSxWd7bX2VmK/9
qL4uWqBtTJVxWn4ui3R/foOxdzIEPU2FbIsnBwF9KpyZYt8YMCgxPpgHb7TVYremGIgqyYWScZZt
wAwZWSApasI1bUu89UpXZJk2bMZx6EpD72eTpD78MZ5xYEHEZ3x2cBw9IczJzZaqQNdmEH3//3Ez
NvZYKlOOKX9/4D/IiTeJoMHiDEnGZphkms43qqABi9i/SAerrJjnd8cWsepSd91QbP5m6pHds1ku
vIpVjwgfo4DAetgE06cNOaqpDRSJzzTCqKDKdtVH+pwtP31FnhwPD/XcZl5/aG8/pd4bki+yqgUQ
HfP3c9IwvZGrYR3eWHheDEN9Cjci6lsqdyPZQ2I9C2daY4LbE8o4JfDsXHyvcDv9KEkdNwh6+5qQ
qfbXS5ec1Hcp3LVLpbFsjYsF7vJCVjuK416xo/V2t/q2c4RX3WjIHt56OmgJjEWw4VxUTvpJVCFr
y2JpW1vYixJfFcTY9oXzzpIKvVdn1jM84SJKSUzGm7VXPnaVlCm8tGppxPeW7Ypk+ZYM8XANci1c
9W5Wc3qzXPvrorjLxgzZF9sMuXzah/IziB2eq0H3s8d34J9sQusK4uiBMoeqyxTracVdW4XCbXT1
bCQsAGYAFkWgu2Rc4xsphRQotIZ6X1qNepEWmX9gIRyOWVp7PviJB0BZw0gUzdjWAAdzNL7sPmCt
/hMDWPrvGp0H1/sf2CWKYuJUWC8drCF3NGmbQWKvfwuNw0/JW8I4JNWCjr3NssJRiMnHIr2BjyB0
2HSArweX7BfK/ypAaH7ovzyiacCRM70fW1L/luhlb+wiGasxs287mkF6HQqMLqjXrJHJXsqrJEOC
29FbQxeNvn2D4mlv4fZZY0/DgWDrGys9XKDVwH3yEvVtEMqXDmYcN3QVtlpc2ue2uo2N/vtdxJ/+
Vxubm0Y84stWJSN/twJHc+HS9siw3eg8pBKF4FPb0UPLJpQtEJmvlsmlzh46eV49LtxY3If1xWut
dfKZC5EHYaM9SL5GzGftAb16i+2fFBPNaubmQ7oQK6RVvfFgqs+WcGiE8vorAbekTNkKHTWirjKe
wI2Yh43lGfe08dG8teqGN3THkeT0qRPLb23FLa1vvPDs2Z634j9bGOlELRDftr3OBiqMwVXgQbb6
xd+SIJlk2asJ6zKZ6KQ7r9KC3J/k/h6S8fjZcCJNAzE4TMwBUxDgIrp1O/KKcQ8ovhbHyFck/KGs
5+9FeQnj6y9nzeh+hH10HQ9i7RTkLuMVaHBQAkliYhaQ0QEXm7D29O7+FT+ZbPPaNbtjPejftqnm
Y5to786eSkh/WybQCJCH7tjxAlhcb+E42yeNJMfyiZMNWUyUvD9Dfp2jfY58SgvnhsRioyP+Ltnq
Pu8K+jV3cSlGE3nrsN293TRWB7gSBtKZhH+TyUCPPkVDcspxRuIHH09zCj94kwdctZCgGOHabWTV
zJB2WZkmv+A8JDd/V5pBI4/vHdIZsZBmHJNIy7ULove8bBO2N0hwH9eciYXTS2RnTErpqVlFC3vV
4rh0QZezhC6hfmCxB11HSC81GbqzgNoOzl7TT8hZsjtyNtTkuP51R1sNCrHjC9ug2mWGXVfAh8SV
b1bWtjjsFjyFkShWNKVt96jvqnEvt/+9fGQ/kghRNf6TbH9ZBT/DBaQUQ+dBKEftWx7JTay7ehAS
utdCFG/ztpKIuPIsAIW9yp1bsUDkFbi0fm1kKj1YRlU3jCXgXFJmsT5gRyyfLAx7+5VK+gb30UMT
IndOiSB0Y1VVEjIrL4BHwRJAYEAa97j7fmP026DHzwOziH/Zp0D+ZZtU0TqSUF1U/mCpQXXtIHO6
LgYMCI21E6uqxdiiokRUTgeNdstMJoOCSiK1tmi68jzdfp2gPNWw26krfzlKov2dAPKNaeiOhtOG
wpf6ZF3wYCn9Qy7rrEdWeycSHMrt0XdXmgw5jLpQzkBmgmPIXOcvNmqiKfmzDZJ0dPS12sgrseDW
I89D4CAiSH5hJdWeK7gc6UuLMN4T4Uzfcr1PIuKySIQNiXa4MQeD1HCsJR5E/LfrZywGa2yxW5I8
A+x+D8KF2xCXgycev8cYVmR+Pjc40XqRNSutWAfZLiGC6TDIMPUdWqElLANDpdGzKpKqEoiuwZRl
KCcrGIwDoKS0aLsxOsoEJW1Hy94EnRa7vMnRURLzMtTUiyFY60yyVMJzGI0kcXQIMT4ZkmQVg/Ja
T5+x3t68PX5HMMO1x5gkjLI+fC2evrNyBC9GskJ+JVHjs9QS5bdtFjKG8S4fhm/MB21Kxsv3QdS+
ozj6HVxNKp3JoNaYYlC7/3HkNm+z5TNkgVoAbMtWkVm9cIIiQkZtm0VBiJdvO24bxxu5OLeZCbU9
r07WsuFVI0G0qr3Zt4+KSzuLKLFUpUI5etaRI3itNg+llf6C0utZLmTnCFSEU0L09QNC9svpE724
wWlnDEjyN+hb9Y380RmFEJ3V2Y/J+Avf0Vz/5S/7egOUoi0VYXb8azy4mefeWpcIm7oQlbbTb8Cn
0iPEpsXoMXUQX1Ec5PzP9JTCtfHJ6Uz+gf/RS9r+v57aQ8yZDKMdFSzOVuwRershWYs3lx9O01Qf
9o9k4wmiZNyIIrSVPgnkRrpqJuZ1W+vfm1gs0sA5Z3kb59ip9ZjKmckj7WHoviRuvGJJcyuw3Y2j
Y06w4Qk6LWG9BVzXPChjYAd5I2kCA1nraCy8aR2gG0FBTRCiIdFhYg5GYl4YQVkvGQcpHyu+lqIT
oQZ1ORJiD1WSXfcFFu7r1JvxQtLkBl7+7pJym1pjJefPt/zAxbD4l6MKtAWcpnGDwww/TSlSsFjP
bDrB2aEncGB8Rd2PMV1Mq1vpVD430tliRfmYFz/+XnKqP/6NTBPKJ9o8DSbhazKQ5gmP7j+xyo59
x/rIPLYbw6McUYQYLYkZ2SJ1XsrRXWFe2XS8jxxjTienTAPz2TW9BDJ24uBHK11HheE7rBT/lWiM
9JPigvHzWNAMqqfuwlJ0BqtOoxfEliJHbf8fWb5a9IL9EEaO0cQ0UBIBK0SgREeN+hcU13PpvWqr
nLijdwWgna3ZPldaBL+ijilzxcz6+DTaz509OCle7hCIInWu8Df5AXnylShD9/C3p1G2bMskpAWJ
jwhzSurJh1uGd54faZFRU+Lfzso6+rdjS6OdD+Uw3YveGlbMRyekKLw9V6lu7DY4b7Q8QAVE4U1z
Bz6gsHP1IjENR1IG2z8SQF+bD2AcwuapjqxiZYXzM74UaCp1VtzAkCfqqkDOTSfKXi6+pANMOPO1
lCwgLe0X0+Zl0qvsw9MgGn9heJyJdQJpdAc1I2lSpXKpafq2UnG5ShX5h9tiK4BkSHcioWH89why
BsRRJMJjprMGHinnXu/2d13fETMq7+UH27ivkXHIn5BtPRPqROxMkdFBAGhH8JMDewsvIUbAheDA
ObESOGX3UzYhyd5fjruOrr8AFO7nDe/iDiiINsJFTSdwLMnfvBpcwqRZLimQH8QjRwSQFsurmlFj
hO0cE8IAhuErmwQC3Itooj87d0Ety4BeSR7eMvnwUasirN6zlYZAoc4Lp297lfKrXdQ0h8rDqGMu
nm2ueffb0ym6Do4mUsi2RmuL/OwdpMLMKX8fc7nY8Yo/BRnmFyDqWAGYKRV1CkBuf4KO1wieVgYt
mQ06o3js97TdSz+1GchSfK/tfMuoxwD85kicpIZo8fmrWId4Qj5VvUq/95SSfD/EJG+NiXwa3+kp
qLcXSZHH093LKnFKOhMrGQNdhxti+lFsr/Syn/e4JZOyAnCRqi1fEAncKzzV30jcFvBWcXAhIxtH
5AMQLmlgPcvCXm7kA9OTk54hu1Eq6Vg1Tq42/LRleNq5roRklqn5b0oNEQbjU+AekQS80IRZ6tVJ
7vIM/ydHWXdP7iSHNCQ4NHQ5HI6M/mD3eYy4U3qw+OSN1lTVFkAec2NOqEb/g2FL4mc7UST/Mb69
+8Io6/HBiG8d+WPZZhxSKgS3XQCcRltnT2Sx2iKLyzD9pNtBYYMGLFB1Tgm0D9At7z90ua9T+a5O
do6ssWoo0mf4/yFzZycpJmCX7Z3vmbpXS3Gah6lwo6AlD7ODbTw3ukcbFSTJnkeCAQWWnAuHR14z
DSqZvuar4X5TMEoFtxmZP9xB63LbXmBQeDeAa9YbzhjTYZXP1MzO+BWCuWeuTefyhliy78ochSNk
zCPUc6GQGalPSzA/aD+SBT9G1t/ARLXmtSmWQrCH3a5SxGORZhfvhfIaYtxVdKQ5yMRKmKIDBhMb
vKUOJaEvOZ97sO/7O57WeK5gXnYNIbHnJBEsMuR4C+ILCyPvgUPxVw18Gdbcg8GyiUjIybUgfhxZ
pqgkn0Qam8LekWn0QDHmsYlI9i8ulS11IOVt7YB24E4Y3E20JSD2S3B8ZjDFJ0KggcU+7nrc4uNL
3X907kVPq7IGGMD89G46pKjmpWvcJRDLbxyBIKkdLr4NxIpwfW0WffO8VNv0MXWsL438FK39KBZ4
STaIPG5r1HAtdhOqo+4WFEKGk0rwkvKtCjWg0R5d0D5XY9SqimjGydaB/Bpa350rQBBpS46XfWuu
uhxvhLq4p4dYrtz5stc5c0dn5NSaQmMuDXX3CsaJmcnH58mDGXd0p0RKBqESNQgUjz6n6MOIvuCY
9BNGCZkHli298f1gwLxjpejkXqX0basPfYlS8qeX5aZYK+Ji2UVHuCcFDNPnRSbGXcinFHUsO8Ec
01chPXena4/prLPGwP2SARvL2mPV6fb+Nu5H5YAdpTDK4Duf9OpiJj8MWSvYf/CKftrR5byPesCU
1hvog6iCFCqe7/CmkAcqGd5QTdn0k+6j6JWmGWnuNWuyXrSX+K2XU0K3/mlh+osu+K5zmlz4yrZk
Rykw8dZ3q6wfq55KrLdDCqpnFuM+4qRoQ6hHHC865sB6YWYnGY5Zracph9Qg2qSSLV5wFqQLFuu4
wrO+TkLb339ki7MOIlOOBKg+JOSmvsDMRy4YslMF+z2mNtzy5WwexUnkRye6c1bzq+Z5J+qQbOGU
WLpbBmpX4hFZ9i/6yqgB7pKmhs9OLs/ho9nN9hHPpwm2QC9EkiDzxCHhU9G89c9C1LqsOcsLWs3g
PKhQE/xmmslQKqRj47rcACO6pbSGZX8fEMS9ya/yObb/GZAHUrPOT7dYzfhYC3YgUuialFNeg2PB
g/uI4DpcI0FXSy/+bVm+F68KXkMdUTeDHtHnkd0cBK2t1i0i3fdho4f9dmx+iZW8gKoQeg85J4mA
tSQewAu5v0jp80iLFjuCYZhvsQXYPb1C3IFykp2/TGVraLnlE+vErOBJ7Zk0T7M1A5vi7EL98lvf
SmmYO5Tw8wPbK1Lz9yll4VKFO5NVrrTXsmr8aMLYF/nr+9bYjj46dyRM9ocWsldHlSsPN42vMFAD
tYrOGxn+IV1Hj60tlrF69Upy3DrspRkWRMA6DzgGng1dLC34k9J2zNoAh/Qf1o0mU+3oYVJ/k+7p
BsKbZWw5cQifojjBDvhV2AbsG5CoSjEivmPQJuGkVBL51N4/sso+sSWnHdD4YLhVH49rPkyRHbKO
SN3nxeDy5d0eonzQ8i8Lc19wV/6W1g39Q4Q8qQlGlQho2gfv59eLeFBsLnLlMDS5b0Yo69qt1VzG
aBlhUJ7tlTe41tkrYfYlT+VYcf+qqqbOY2tbKNFonb179YYKKwHpLv9vPE2fF5VGyqqwHakb7Off
QEuj/ms5blCU33U8j31wn6vU9gVx3C2D8VQ+DQVZNMd2skqnSRWfuB4V9EtigblaeUna2YCEv/Om
E1dDCrNc0SD0FklSj9yaVSfJXuTY/4H+ZCCWNj+lwkALStFlts0nnXMly0fu60zQi8ej4w7+x1YT
Cvn8E4I0sDJpP8KvCpnNizuoJTuXwOG1ohBUmHGtkIcRdUA3x/RSH8GbbS0La7ROL75ZNatMn2KE
TNiU0nlz/zhvedlZnaVxgEfT2v+Ua9r1mqFyAsQLalQ8+5ZgtNeemGGOQPvgXPsTWg09pJJY3szY
UJyE+e9/yA6ZqCMdl+oo+dLgpu/B6emQEl6hs7TBLisNo3rZwiP88G1TQMaQ63Mrlgo4tLDodAeP
BuSUwZVLBE3YIHHRbfMr7djG6/xU247qHTa9SgEgrHscjBzmvmwX6kGTrb65ikrjvsZyzgWE1kUR
8PuNQKnmD/MnIsantfKQ1ap4LTbddjNEiDINQaMGgK3CZE6LRqfhH+kgjm20t73DXu7f5zxFhXz9
NPisiP1aVZ40+t3TdrfHlAwioxTsu9hfuZEsKJpDmKD41URQ4HemgFw6xFNySu//Mp55HnGr+ldf
F53/Rytgfo5MExU/PHaqCcvvDMEyHQgPK13b4vV62dBX1y3jsvPKsnVfc88LGAIX1T4wPBmiw3ap
Oq6OpIQgRRFita2QQMTmrUgCjqczYDxYMTfvzMJva6LBzj6RuBdSoec2f+aoh7HUHKn9grrWn/nP
CfCs7IPIDLSHdWOXTxC8bykf5ph1sxTMb6QmnR6jqSVLySaOoHB9NqGBDjYnFPoLf0yqKdUuEry0
DtYhhnIb0ldZkgwT6TLuULGwTpmfqlmoXJ1Q+dvTRBVjqs9h4vwk68lvRHvFqFj2xzwDkKCAX1MW
0Y1y3X34B+831N6lHUbv+nquA5wKOrSyh3BGe9NSYy0tXFCU3ODGH+U056nU7p/aQCfM9yYbMCtO
bK/eWHy3pz04gIq/DgDh2o0TdfWTtc3OvPcBuNGP1TK/uwNx87q8kXblcAL9HpNfKrlDAQPh2qGI
dOfI+mUjheUEeBuLgkBkL646qMH6w4cJXtCrSASqEOoynZQzZuY6pdAeZ2RPb1Uo35FrTUjzBsyQ
wbhBZGsX6yeRJozrc63NphMvjYcAohvBhQn9SMiqcowwKTaFyqcTu16RzpC4dcasQUcfnvE8YF4w
fLUXPGpfqY7/odEKoVjKI52D2olAjj5nj6F/roxpkLc+O3DOQZebGuCNUwQ3164PWcmeqTsKBnKi
Ry1wgb1l2nAAtk77xT+HFPtlD2FlcBsH62v7caKl9rcdYw3FdVlM+R8ZXXgMkt/Sfa/2UQr+yL9K
XjqlKsW9Zb95jiUU19EN7M6dIcwErJZzUaIaF9L6KoGBL5oKg5wMDK0tl1qMCeAn9GriwAccC3Za
qPqe07ocGcWyoR3e87E9tzqmVeTI9zboGQfm7TAkG/L+O3NWy1r0IKM2WOytrQzfqDsMO+eX3uET
GFa2jArZnbgtRdpX7ztMi1pEdIGsQGpdVv+0U+e0zQWw4DHgWlGquKCPu+RgG2PmvkWwf/cy2p4Z
WjSW8CUP1TiNRlwb4FByveKT0VEXkNtKCHJDtl0AS1o3ZJ33ISYa5fZtMs3L61nMLJxukgiH5Qny
NyScwRrGO89CbyZ/86L8hAsZurzfeYs4tSzISE0jKQvxSSkqI0eiCyUOSLCIRIOQ+7JAr/WO5zWG
e0rU3tdfI7bL9C4sFSnh3f4lKAZE2NQYmfLeGizaAhTEUW7ewhDICkU1TDpGhsFUUUJbCCu6A+6z
GnQ+KdJOFXUy7AEjpYW2LZL1lF1ETP4eG/GGc0d2PfVad0rUPbo0vOrdG8ZEXW+3AnSJ3bKm9G/d
AuWmxF7EEffBDh2rrvAU6F1VKtFh+qIphfFX1Qv/JU2jMrF7gezzRreGUn+hwvnZxsM7sz2v/Ai4
W37/YYSveyCG2ywzHgN7OL/93OtKaEzeRjAZ37dw5BAjIbmXR8qMjmD8Z/N26qP3T2iKTZ5wu7b6
LO3ub/THZb+ViZ+shUX9fykVzPvhxOOS9qzQbADBXH8+7AYhuD/FsllQVTPWreYEEcXhOOjnFwNG
Gy+IEKsIVFBdPAK1Pp1tF3Kr1pN6GnC2M72wnHjyw5s/2JxWxt4rQraNWSq0KWUFiCm+AvDCTJWm
sMutCJz53fZ7tSQKmxxtty1vfveDuthmHrkl4JJBYH+NsfT2jpCf2FiIbs6gSKx0WB/RtP6oX7o0
cJZkwQVigeC+cSXHEPtKC8+AfMR5EQ7lG4Dbdr9eHPurBQ+DMlvg55iQcjivfdGV9PNxfvT1yx4R
UbcIOEMtNGt17pPpWhbZ88HYLkns8sHlz3dgXo2pYZqmITj5Wg736AEamQemxpb0tJiHk4fgvTUT
Tk7FJA5mnrmfl6xkT4QRTXkiuQrMTf/sOosy+OeaXx+aPYGBsZ2xG11hQChbeLERec8DiRg0kHXO
WUNZLrzHeb22yGoaElDHaDeuci1ajHlVY7Hx01ty0+vUFhSRg0pNt4Ix5nsDf7cT9KWjbXM4/KF3
pO4AxLpzglX6vZBLCIdXaVRiJ0MZXjPH7HeExiSSWgxY9lcS0+/3En1aA2vo9XPbvUuXgv9AGfZU
ww7w31O/WgvcNzSUuvhrmQxeXgQi+qUEVKtP9LGk6FIVTyxjWMgaQO3QuOkp0bHLv/ncbc9VPKxH
wPAav1neHdxlgDr7GJ8qhMtN3GXQbgJ5ZiWRsYj8JMzZks4BMGkQZrZklJPqUSfGhZvtV4sUtNcA
7Y+y1bT6AHeXua7I3A0nldLc0zcrtGj0uAImVka1P1GKVpf2vHIkftr6MZwx+HQ4B+yEn0iWVFcF
K/lc96jLxB4BIKKq8RLCUZb3QtuGBEjlLHd+gWR8XVRRfPGWOviSvsiwQCjh8Pq59wQ3Ea1Hxmt+
gBfJwSg1e4WuirFYVxUPc2vqhhamauKMQ8tSmpSgDXQgURHpULdjWkjYwJkaonHJFIfl2pgKIKvw
mLDaEIGkMLbCSMrRkYzFZsaSWGKuRRr1EdPurte+IVq+DlJc0gJoQlywSm4v8OcNm4YaFzH30gYd
1M/DEyQc6Uc4NSmGUPzhBFuXyyOGhGCm7fk4YIiU/fBFGzeTIM0bpwuGwOWOHT+X63DaGzm+qGp3
ZawUZE89nxT3vNG8kWiB9gJWbMZuFQwOZE+d1QFE2z2cBhqhogA3UoFltv7JOLqvZdclONCzexF1
LbceNLzYDtbUFKxjklHA4NURVLkGVP3hNgL9aU7JhDuk+4KUWl809wYTDRv8hlo5V6G5CIwPb4rA
Dy+iiRUoZ6mQCvLLWrgeIlMBN7mkh9Eb2IAeLAoAnwMt/rVS9AJmkCLlzpWOpDeSfXS6SXN+bV6v
vyrmtE85xU69ioeFMrMpR+UHOZMYH9J01DsEE1osWxcVw8FTPGNl3ti+rR/VrcWkftYLA+c6YgYg
ZIicMAjgvBaXR0ikbrO4QN7CQhZIKGtrAvsC8vcjtXE1QdG3XOI7G+Mzuv+eizdpmPIuT/NiT8ok
X2KXwLE+H4+LlfWGuPjsyOcgUi1pLWLnxJBJ8lOYB0m2r6DcqEuBGpjRKyAXPGKeOcQVMFWyjqrD
2u5/x8Yus/Wx1DWW5tWNzBTRjsDYrusJy04vfLq/cO4N+EWPbD341OKB6o8jFkWzKLKkjRuBzwvn
rToKpYmPQJV3zdGA5RZmKeTLJ6BJM5FjQtq1Ez9z+F+r+Wc5DpJdwXGdvH2EPgFDG7lSRdr1evK9
rcC/fcMy8uAjjAOaOTYPjGKi7EyBrF1CG0cS/dt8bqxRF4la2TyPKgDxu/HJk7ZcK1wOwab07hEI
YN3c9sOKdhYAuoPlS7r/OSv2GeuPmslMJIGH13YUxv9nWw5QWY9Aopf08r9O+O5NbGZlI2gOXOlP
cA+I7qN8AkdGOkDOMWHTlTbBMA0Xeyt34QaR3zFIVyZKFEhNHPNyyxHMdqx/xT65q9DiW33RWsoo
V3JSvXvuKuI5ym5ndeiPwoKRC8emDjpEhUR8u0rLfK0nua7rlzhIivKdRChTFnxwQDMWrqXPtRvA
LdpNSkYfLulSQueO5mbDUXzadKTsOMNmwe/PkeiGs7FtD/jAOOaJcRWUCUqypGYB71MECOQ8R4GM
ruZm1oyAEBxxVtfs9MUrYx/2l5i+hTM6H2y/679opid7hQrziOZvEOmPML4CEupaopMzR+qIxOjD
wwgeV0f/nEVl66VVfndPvIy7ThInlTaNiRMClGn9ITspH/j7XnJ4wXGE196jsb5vipxvPriBr9vJ
6GDoMxdO+IhTqqvbamEYNb0es7mCfK5t98aIgCFYSB3xzQb6XJayS+bvOUOuEGLbshuq8eOr7tjr
MFvAG3z0EWxRL37i1TVXlAtv79BIHJvweuaGzZtETUm/eGnRcV3tEzqX9ZC4rU7o0BE0eMSACxz9
d7XTP863alEe3bW3DKNVTjsmxl8+lsEc4zD2m6zI+Y1M/E49KcF7w7crpF3l1PRc+8jCKYb/SEVF
nrzuTQTsDpuk8QrTkE3fsNtHvWKcaD2cWpOZnZXLtF1nSP+oZlmwC+bIfjISBeqgS7ViXrTotaIu
nbDVYGQh4tPyVAtSgD5V8JnO3mswuxNCumQGCGHfgk7uiCt/LnMRJ8AZTha8n1MnuJjzoqit9E05
TaiLSPm3+klXY8FqBtNhoIbUp5hq5/+XcFa0/3HZXWvsizUdBCq6UXgg0yyPQFT1ReI42ZjuMRez
K2yM8Il0dXn4k4M8/zwdAhIRxhhdePwvVnafF0odxDmhuOLkFFyVKm4KSp08zNPowkWRfW2Js1hu
0KWXXkrLSb1PX8TQVuUg7yzT2YTSEk3Yv3Gr/9SjRujae7t0Kux2AiweAt1S4vskPcoHSUVOeslp
YwJXMLexJFV7H1iA1cAb44Y2qt6VWv0IMK6DQ6tp+i961epkTIMqexR6RTx81kPymtf6FCd45Nca
7vz0mmklBD4C3sDB88FrXvUgefjegCmQi4ZKx5xN+pIDAekp73DnVVMezqKkPKLf59SfKDYkONNn
l2ssOBS9+TIY9bYRkTem6ug2Zj80XDYpOIirkdMLejsvKp1mDPfTXf0B7vi7WJ1XDBJLFM8cIHGH
FCdFfjZ8XtRWDuu7q45Wxl4mU0kZSAq/G9qmVLOM+vs8l75kl5bD3ZerfdRMlUvXa93TLeW6P8rv
svJcog0qwPZCr5/45tid+5eH4/RQjwlpXSu/x+eVpmqdMnWTWu1ko/uRu3YojZtM5Cq93K1r89ko
K/JCnjSgLjWmm3K8ERXUHrNBvGcrk8j2sLMpF3cT5weGWYVymz5LUs8ONHbNRU2tefJECPPr7fqX
89MX7XjWLP3eDZ0ZdbRTwdpWS1HfhwE6JGx25wzK6GE8yLfaqIHed22227T5VB8/NDbKTtRNDAEY
9tfktqFOAgKVpjujw0q7zWQfnUKXQlVUEBv2f/j/Gv3lOSYtWcTHCE7swbAC7G8iHLuneiIYEWQH
AvxZgj2m+kM7slwIWzHcOWwKZt8+vorHiRdNxfmFhnosJoeE2JMfwyyQ5XSETK36yuTGcaJkGYpH
Ny7b8kmY3ldBXtddMQH+4B6lkCYS6gA/Q8g3S0P4NUWYaV8gH8uIOqJb1Fo9lVugXcqQp3dOR38z
RPhIoWDwyAf8dKI/aWrphhp8iKeHceu/X8FHdOGDfjgnLJN6VsBKbBXX0Lfossahiwbq7JeAD7/8
boygxdODy8raFPqrDK1z4XN+NlW5V/rWhiNDDwo97RNSJToqOioFm7WR9l6ucip2w25Ye6ff1Ds7
HNlcG4VfmFX59p6CJ/WEvujasqRR6HaUPMEv53Nvr1iSBxsi9GfzhKilYk3k73aPyWFZt5VSu3ov
diSd5XQZUnqVcQ3uwT0R792x59dyz+Z52J2BXyNSs8emivubAcIK0dHNreoJee+izie9og6xLJ5L
pwbqNisoVQtWZZyl1+0gUZiOHNraT0yF0nOoYdVUg/y8qdEA8b2OEKUlS3+XK1jPtRpslDV7/Dqo
/VtgPGg8+GBsGLo6iyyScDi2K+emSe3cE2jzeRubpQOIsiMFIW07TDY4OCdwPzgiRtfoJ7TQ+RqZ
fHEQJtv/dPe8B83F9nSBCOgSEVvZSfWVdHc0BQd76UJk8pX3gea8kryau+VSg+XVcUfOYsz9E0Fo
GZ16/xPQ2jk2lcuxEnH/RMTxHFc0SbyR0+TfdNk20HjlKWMuQqNoCqOMpLLfONBL9W3I0rONF+qG
QuENSELfNAdD6WTjM+Zsp4ccSonQlMpZDB12IbkCcHusiKVCWAlOmVuCna2iBBokwGVFBkEU8YdT
iw20CR7dWmVjdT+JWoiTtdGMqCyIrhADu3CGkg/hB3nLZPaDKrT6eiB08RuC5Y8tuClJcKxUCljY
msie/9nMSAiJ4hxf9BH6xvGnqx2GcleOuJQ7XsTP2YW3T5VFnLkYy5nblUGs/9W9VkY6GlBhB8CY
uTK5bNxXBuC+5poL+7ssyjzv/3nnIUsHI+VLslPcoItzI+8nh1yK3C7NiQpWSI6T039q1EeYnh6d
gZTxVKQBz1Quo+BYzFM+jqsmW37y2CAI9VbRApDbxm/r+VIDMNVZtbUrguIXkqHvDglRyiYcKY8c
nGXhQCni5D2uIYv85M7/UeV8CvaNHbCjL3DvhXaEJSSSoYwQcUdmGOKKQYWrROuL9gTvzzr4WV+w
pyKFOurGh4fCXPKc1fTXef86uwk/NaSJMKZefL9pLSrmWVe6ZXcxGcRV5nPo1X9uBVHxI0LwluhR
4p8szo+QJE9eiFh5mVIx17pUEKb89TGVhGmol72Gq+JH+nmrLsL3vNFUk9WZCNcecPGReTlgnthN
RPix2Tc5wUQ5THl8vIG02wTX5djb07jYBNh9kRRWFT5o2Kx3YlECMmJ2arTONkrCpzsWDQyvv2X6
sXehiL9xvaG7ys5tyOjzGktmmYaC+ESfIVj+4ZETJ/0Aj9sVzt8u2D476Ky6U/IKTn/ziTYpbiOT
GNs3q3iME71SPMPj+FBPMPwLUTPrNvsNPMSbuPCu8JLGymiywqtMUfeedfyMNfP/zZ4HSB1FVYK6
hR8gcx68lxpjEaet7xDvBNEX/hsejnFm1+9rd/wqnUqLez9HeAe2q7WQYNmoAeDIAmhTXFamrD/m
gzpDYMen3F7WqSDEt++8vFBD0WMP41yQYulALftHCgIVDPPv+S+STff8vxFApk0QSzPxSqTjY14i
h7X/QhI7zM7nJkAtedMxP9ocCeyQJCBxSNAoGcbc96KJKKYTZge8Qa7zR3RYBiuinfajhwR+rkB/
NoLf3VEte6OKt6a3XdJRD6F9/9goyaPNqzS3ooaOaox4dsrGWTBQ85AqrVXz+10dOamDMxipLXQk
gK/7qRlfoFDsuOO1tm8qzFwL1Dk3GWr/IVOwbl/lorzcAA6sqKSiOGvE4mS9cdMQtPpL1J8hfHMG
uOsQTgrkIKAtEje2TNzCTohiMq74ZUNISC6+0ah4AE6QZQ8qy53uUMepeTllyYDWPtypYNjekFEO
DcQMYH56AFPmDKqlrf0p/a4FpHEuBPQAC5Yv1gXLFGBjDM8EdFbyRziBVy18qPKCaOPKt9lbIyFu
/1k06BBKEzlhFS4f6m08jUQ/kmUWDt90nEVmx/S/D689H2JYLFgZt/sNo7w1MJd1o956WbNTGrzx
dWxHqWDaHXoDen1/FrcrbVz0Cj6qfiKysrnq5nA6+Dlvbm0rkJrUpgFwa13/+aSQTNgJpjDcO9Nt
QLit5Q/4Fl7LGdfAdr5H22Wd9VEKDi2ihCWacoroESMKCBEfxeV5z7h6i42je7yHUq3qrfZs/A9L
0c4w8UQpC7TckhXRuYe3uaWqyzFMkiepmUQWUAYb5cWMwCyiq5977yDPJM1ulBinypgh/eA98G8P
xWakVVs2F5zK3v5gn0ZIySCCb+nZjP4T7Dg6fyJIcmqwUTo0BLStHBOCrBBLDvIas6qV1GFpdefu
5qJbp04TVNSCM4JZh9u/Jo98gLylEsSw02NzymiWLP/OEUlMs5VKITluYMm5rNvbSs5EaIEn0Tsj
c5leVewTCANPlDf8WK2aYMW931+1mtFdzggm/NJ+6ZR3ANwtOa36/cWR7gOMoxAyzOIqRZtddM1L
sFd+N/OKHkUcwhcOCi+HWgHfpFXs436IX4PkzNDSh9ByyDBMuqjuSAfgvpGdPaey6+eFRdlGLOAY
EGtandgVc/upFsOIGLTi8WW8zECJTf4AH6d2cro1dFLSytJ3TUxt5b64vQbw+qUVq6XhtbbR07zH
EDZ1ahgqe6/XPrMlw6WVjiVtkZw//M6W/Ksy6mAuzHBFRfn1z1wRIMVNBhmXUbtYe1vPstX9HTYc
Bx/F5a5GG7imLr8tXBCnspGm/uB89FycvuioEJkRV/hd8PII+64YnUvDbaXLHFZvcmxSnelUiKDt
ApwEycekA9QvWS9nb1p6/AdCzWL+kmPk8oawY/wFmQX1k5XgbMQ/NbmduDWioOsFWWs1TMCDw1l8
NNGOHrDdKXzEYkBaWQ5Yq+ulpEVnhJmYL4lcG0Xan24JsRTr5vUvnrJNwM8L2cZ3/YvXWhomMewI
55ppC5d49kwalVcCe4zqYyLn7oT4/RDI10Mxp/yqJyXyiapNrbWDxsd+hHGFj4u0BoP9rwGKgIfs
YH87wG4MhseYl/rAqeXmrfX2Be/72DzsA0q8iekq02i9OpIlKolqOMh7ylEciIoETLjFIKH8Mflu
a6UJoaVXg6fitpaNx87movWS7XcNVidvyE3EHmMP509FlFp8meRMUnhGLNGhcVob/YvR+viFNj8v
SJUxsdTayN1iUng1aZkF1RKDmfZ5swX4TAgfl9LkUpuZPMQRLkUPubyvN4kLd8PUSp/9r6iIxjga
0vkvkc4TZeFlJtsybf4eONPmmITmNzDrnkqAHodD/9cD4maT5svR/iNgwj0ONL9Hz+oLUvkH01AR
ByJyhREVtwhISrzlkzTL9caB/BK9Af37KRi6MwUo3+jrr6XSHlfqj3SyurauYX4UusWUJvUoVA1+
X3JosNQMr4Oak9usoznNLnBNsyuIvX1+oC31WPmM99svkkmvm7LnqYYlp4h1M++xhbUaRHORUGRh
Qw3H08xAYnU1Ou+suK04qegdC8xEOiZnR2ZFj+lDFse9xpjdqRGV60dfE9/vPgLaoVKpkpRBg1TU
yVQcQ3HFutSwIb2TNs6qEIkhNYUng/DP2DhHlQMs5hSGXNRqMmAPDT/22IquqgzRVzWUXruT+wBB
25XZB99QEaJEjvRkuSoqhPxAFFh2Sb8bf/iC0IVv2O0LgmC+BLP8arQxNAK3hCIKNmqc5zLSAVAx
mTvhmTO5MhyZizxxKM9WGsxuJtML65pX1XzVY92EPQ3bul1bNneQel/eFcUwpWK42NJXS16139rJ
DpKEJfjBkTGyknLQaGlOClUYPVMct223PT51qIdbQAiG5GWKKa41Gsq28SDE8BEhdL26K6I6DB6+
aTfQ/dALBYHgu971NcD9l44XdTdDeWwWtaUm3uurefOx73jLH+Zs+ljVVduevnbnnkAIfV4XxGpI
CQ1+FdRcDiFPTd/tfIEAbEq6LQsZQuJEPWz2uZW5dSOH4kSE6yl8vdsMTXY4aQWT9qaVtB+Qm5B7
mYBMc1HLQbHUJUCY85MVQukl2qrbmUITAOSCkJkcrgf6Mrv6zlaHms1sJVxqTddf/jp4wrNyn0Yo
Z0i8GPpQu5XbUjHw4Chgk77z3RyHz7YsjMmVFg5lbwm9D3eIneJBY5BKQjTgMqX7NT/ddvXF3AjN
LTMgI5rfkfL28/nUUg3DW2ISuhtajd4k200Bi+C+nx2MD8q0wIm/qVKKEIt7UMZ6PuRqHU9irNlj
uTJiLS+agKxPJB/WdhtqZ4JXIKGn4cdq8s1pkyJUM6V6ljqd3SWVKa3rEupGueD1YpkELjf0FGpy
1mpmnHHxlsqLHw+mtHQbQ1ThhOIroTBoMRo/WIHtMksNcqes2jSMbr8xXruIFh7icbaWHopaK/cz
D0sr3j6fM9iEq19OSZ6sh8eERtYO4bd/fTkKoQ+DiP5eExhMQEldmqecKiAVdA9u7K+bUJ6hdrpH
xWcHvQ7QXy7ZGqEdlXgScCKdNVUGNMwee6BdRTf0V4133koGFAspHCrYfKq9OOFzd7rAiCHO6BWb
e8cVHqfekgBcIErs2v9iN098eVBxrSgOWGaHNfT1sl4IBAegAJE9VMqu6+pBmE3RWmBXmtgkxk5d
8okh+DSX+PzGgJJ+O38+1rsP2EEdjSiJ1vyTp7hn219FVmBH7fkyaD6JkorrWQu8Nd0PgYRcwmST
Uuzlud2AMgzUmnNqtE2OM3OcuHtPA41HtS5x9CakZp8aVXk5euOecz2OL4xFxKAQJHIos3KxtNBc
QW/B9/tZLvRGFqUDNSOwPzI4W+8bvHDpbAM+ulc7IOPJZZZZdvZJIsbtTCOBxxXXdmDj5Wfvhhro
0KowN52UCOq+ReKnrvc4xGBlfFliXJ+YO78y1HsM1lepgbSEdO3Tp3UJ2wUIU0M77NsgHthcWHTu
6WKB9QfbvIx/1hd1f8YSOEDyOJVVIXjksXpi/lqm1vmwZSR0ITYGU0Yd8Hsbv3mkj7jxL4QVG1wo
hp4oIoI+JQAVpeNSH3dHsgui7XtaMFmZD/LERSLsFCzJY3sklGGNOKzJm1Wxwr1NgeKUw5g9u+v8
ZUCaAP5YxfxwPLSZ2eoew7aUn8xjCLv8s8Okb//msHhO0IfbeVMMA0D4jWJihVbWaL516p+C+7uu
iBo01n3mAPG6/2X9yEw0UDzqO1s7kkTauw+inIlcqMMCGre3zU6lkaRqAuG4AnIA0JA21kE2uiMZ
u+ahn9kCNz4+VbnAtnM3UPo6rzz6JSziEAFEk4vpChfQqugBkL24j6T9yFtrk10U9oFF25wTvvZf
xUVDSfK5erWw/Kw5mdk70AoY7VnZGeyWHNnqDtz/5r7GvmRr9Zzg4CVGQ9z5o4EHoFx8J5s9gXbk
rni8wgrPiHy0L/s+IGHHhnoArXaaWiYXTYNAVFz/32Sq5isY3mljIyGzfGNjOm+aXmDMARKO71GG
gIYTWor8M7XdaS/UfE7JZlZ2bpAGu4NysHoCJT0jUY6pbJEOqxO47s8qQL1+tOYpXgcXnf6N2grM
KJL6eKOIhhOGRv1lg0Tf0UlHwmlvF6Vh3ap3UHDyO8+WlONSsta1W8nTelSMv1jp5AJcH0yEW0Kd
V8Yez5ehyyhjbcWn3+LaSUCk2voKpNpomtqI5+L3xW6jXJSQPMUolzl4rA7ZxXI6b7xAo0EflRwO
IHwcNx6YhAxXqIbcXbJA4b74tWgw8OBxezbTA3TvxyzyQM/mPHBrmkjcW25jTbCAO37OcXj4elQU
YHi/KzdXOziZhVAVf4cWcDbrEpC6AywguZUUulLNzldGbZQdqwbooYlmTWInGAAr0f6v5jWnwsep
IhWeZVmaBU7UH2hl8qw/4rmFkQpRNppDiEt3Uqv5QD3fV7qtWXHN2BiKApr9Kwpwh1v5DmDzN9WS
vR7mYVT8qMMoIcJeKdikwXgeGlgB1IJhGefwTMN+qSx/keRDhW+5EKkyi4bmraHiGsixMOkgPA42
R0HFzfl+jvFiu1Z51lxwaXWisejSc/R1FKNS9z1hsE5yVbtKhHpPc9wl9vkFd95y2psdF2UXVO5y
FEYg0A35ym+sZ4tWZedi0GcNAecOg4ZMtE7k/zOvMhW055NRW8k9uH74aFFPITiU7OtQQmkiMSds
QroLdrtEBBRVnfxBY69BnTgzUzqufPwF+3rvPdIf7Ch3a5a14qP+s7yUB4e0Oi0+iY3BXlsRTxtw
g1l+8nmq1sNN0OmnA/yuX+WYU7BrJwvG5SuQ5gr7lxbXTSp/Pc95Xa+S16Gz3KDCOYUQM2U3bSvf
MthHIv3S5n05ybqietXOvRLkeVkyydktpSWB5+gxsOPIlnia2XzzlMp81aA1AUnIDcRn3B+eo5zO
9v4SbRGcoXrMVJoQ/xXKW5Xc9uoqv8uBRBp88Ng1Ek8XMfAdW74bNorzDG5fhiOvRJu3kuJIcmg4
ZazvaTuPivaUGnrvmn5Hm76DO4cZ/HyY0Hcc/FZqyCVMje6eDIqiZ1Ta3jpibMkBaWDVDQpKcc+N
YJoOjG08cs5fyPkculkq3TaRpzjtxTEcjVpcsr8R9vxoaGD8JDfz2IQVmYE+ZBMP76M/KAkF89Ab
ipLEKEyF0m7lK67dSDw/ReQQcI+z9HuiAYX4O4lKsxY2k1ouxwiwlymqLtPzmDjHFLrq+tTgcqmk
Zc7XHccgkQquiwCLhPEzwrdUBxMahfvoPOJcWjatfoF2BHp8y/m14n+tmq4cFamINHLOj42JD4Y/
RtzHLBSwHImFZrfg8DGTgWiV/BqInxaJXU5Mfkh/y68CvWNAX0sk4mgOSpfuqQVWRUMl9sslj/Qi
ZwGRdQaaqcR7XLo17sqbAvXNNCEuEke6z7PQUsSVwmAjbonInB+lDEaik3JIu0zgeNg+MxJ+aIyq
UQesNrd02Or0hCTCs7ER9cAGhdlx1Kxb6xppedFB5ZkWbFT509De1M0UKmD8UYhhHgn5d6Vv08Qj
w8ZJKmC0L9+ZWMPT56bXja4SmQ+sX9JQwWDLhJMbBrXe0czVO3DR2DV5539vCPlMksljamolELCO
Uks9InXhxO8kk0cQmT2hrP2EZcbNaLobeJj1FRtFbE4w7Gkayz6jmx8s2uqkwvAof8xcjgdlW72o
k+26t4aQhd5K+cnyeksCZIH9VH3Me8ET7hlCM3X47BfTWWkM3KSsp6UI8tW/VJ0TLUDFgg8ETmEC
2e8pC07hseBxLLrlMc9haQZZ6ymWDYsFOGgsM2p6j+sTKu0DFL/aPzo5gi4zg+3p5IbaF0FvPNkN
yS4Z7AqRPqnzn7BbK1eoeQcun4stGtrWS2c7mm470mbMJ+bJlL574gj/YJXTPdZtkCr+9FmSODPo
VkKoNeKl4TXbK22mKt5ovixfuc2oPEfUhAeH4cVLuLkgBNZekwApR0qsHg5slFDQ1DT6vsoEO2xY
EmaLxY42pk3gSolGqTVh3lrVsEQ6+f4JkTyCzYMvzA3z9wmrm0dBAoiODjQrMO9s+SAU8HdKKdvm
mRmK/1ziLTuvs3V0XOESvJXI6+UxqOaPkFPRTM1O6A0exSjI418xQTNXv4PA5CHQmdYEkARmEnrf
ROooHh1WpDPcXLu4pxbeyGCU7GW0J80NRGJTMAlKDUZS0LgBhwChG3ig36GPGwCaz70IgUsXN6bz
FD10ihfjh64Affl3VXta9gOv4nHvi7eCzzTaC1C5p6m3Us9BpbDz5snypcGlLmP5eBE6alZY+7H3
Nj3lv4wsp0BXSOt/Vsm28zUdW9XGkE2Xvci5EnaqlQ3FCAZKE9sJJrqm+rBx4Y5FWw9lLlWwtOru
3gBfgz5mlIapnmSk8XIKq1KYTywT1nO3xscLMtcnj93OPwJN+q+B9WGd2387nRSsFyD6iUhR4bFZ
5TnnzOfydkOEHHtwxq7ICf50CGCSAKRUcgwUJinH1nIy2q3zXUJ/155st6MeCbwtC6YYpCbznhyB
MnpGMayn4LHS0OMGXg0/NITzmpOwYb+ulkTWNounyW+dYsPzvEiHenlP3eqVFxcFYoIejaNFoGnY
le1kP2ByjuIZ8s/rGkVm6szhTfIBaOjrXZIL9rS3pyh8ZY+YSZk9rfpzwS84SqxqJG7UKYJmZwyp
UegeVSVJg9tV2a4Y7S+1QIZR+4jO3nBXknmBiyip96H7X2MZcTO57SE4vjEyGj6pfuZ8SeCoqWTc
MIJ7KCeYJL9w701TjXOk63m4FYTJgPOA4Hyr/S3eMjIjM2CUznUzbZdgdh0UTn864yDAc7JQVG1u
ERM8SqVjnY5IUI5J+Rl1yi8dFpgmK6az5Hk1ezVpey8Dz+1xojLzWMx1Ezn50b4GqCqdk4G/cVr8
7CGvQQwzB3Qiw8QdNU/DMoL4EJSBJK8pqAeHqsxWf1ct5VYpf33QznUcimCSNnWP9ZP+pSKyLNXQ
cBKWSpRpogO7VzRgIfed7aW/HB3A6UopD4OUmC28RSu2hxP7/yBNWHOSLOPtxoUn30GAxlR3vde9
rU8gePRL8b1jsrEc8lylczlScsSm7CZ/HtnzEPO6Bz110odF31Pkud8daH6D/D/qXAD1oRJweqvP
GhNK88bLEvWEFCQFUpcWK5D2vEeZHFJbT8eCNIhyz6UGVuM4zmFbmVptoEUIfi/zAvVF+tImhhLd
gX9iHHmG3Nx3pEZ/pze0/EdHZ4Hmo1hsQJsVDdZd5ldpyBHxur5D4rhsqvCHnjKXJXmLM1pcAlPL
M3b6+Qzw7xB0O1xNMxK7+PbfXxjylM6UbZpAfmw/fSSeAfdG5uFBMgmOA/qS8GS35k2i81bNrilQ
cyP4eIBNslMxI4XmVu7ZBJQHVcLv3ntGe8xbxy0MMVBd6/UioGN9zT4kfuI5iuRLkkWa7B9guGt1
YcdfV9rTvP1GnJQd8HM5H+NBfcd5MEWmnn8Edp9ds+LdEdfax4W6x1gq7QHaB/JlKGieul7bnDb6
EVejulDX6mFud+2nmzyrn9yZLkEFP/KIvNsO/zFy86vtI7RLlPFipVHsISr3YwZPyU6C5Egpx3x2
jZLSdqPlm7/dh5xsfDOUvthRooCIlHttiS4ZsmKKsazsH2mhsRSkekPAOpj84I1V4xKkWhlSO2bp
gS5xnUp+EuUDNlyu8lsdKJpfcfKEbpt5QwhkVOIlou3d2Hwhab2eZcC707MinRWvq16KrdJd8PnI
RxIlTnuD+2/2ox56aM4/G2zOxQAxMQVDeU8lXrnhN/mchhFfa2/PWW2z6hXbRCw3WxfP1QM0it68
QDupp97gKvjEHiDP0iF+b1FXGQBkHrnnLEAzXnECoc0QJvMlqzYDJQNdATN3CJ4niNEmnIMAhsSF
HO7OWL+71ZYEpiUsOuRfGqxAY+8YiOqKtdemMYsCF/7hYfBP2oAOrq1RyY3TlaTlFsgeYeuVUoKQ
v7H6zE2uaR0IhzLaHo/2NPfvJj2X+Bwh3NhMbK5xAMiRAKVYVQh9WTzn45EfL0f+O7pt7hH/y7gl
54pvmKA4WnldVnKbw5l/uNVBfTV2oN8Aa82TOrf4jEFQ65j88CkhZq9Me0GS30xgTCeDotVhtH2t
0w0HzDEZajUU0UFiauhVAcKDxYS3rtFjDV2SacnRNH6grfLZbuSce2A2jedsDHpCuGF4swpiNWpT
pzHDbfJ7auMwAWsw7mTxTuuQl30lKu0zHbWZzpcysWqFzK5gvguq9CASbsXkuO+wK9Bj0/lfeR8h
7pJ+gDfRFfdFpUy1HYDGNkJer7C/nvrchLoGrfZFF47nctpXqS+7Fi4P9azjgMApiMbZweYRUcYF
mUFANFrB7rSyFjHpdwAzIgrzLG4ZaaZ2hvF/HoYA0d4vM5aUYRoUY736rRv1ylEzCD1WZUTVUhax
CwAMYcYzcVxIkO+oAdsTHunfFu7NQ+sBorHCMiHZyG0RpkIT3KcGkCjgThPB9JzzKJf7W4dx25z7
7fm0rnBD1IZFv691yQop22/OO7DoQXdm9SkbsPmI7yOQONcynhK+ndSFDHrGHPWYjISxaX5bSG1U
se64vCludPeaFYjHpaz6R37Q2GdNNct3cDmQ8zlQa4cV9sUvbpnN4nTSpTkLyp5S3wvab20H6m9s
TBWsx4xaqkIVaH3BDxgslrTuq8WVyPMwFri7PHKTkGAx6DkOViq8sbpqH7m8wZdfsn9Cjrt+mbaT
N4BvDdpbGmIHbauzB1cPUu9IAeQdcZtP4Wrc2TC6OfDbXjNr+9Q+AgntrelzG3dX1KZxtL2/Rnl/
9b4f7iFEuIVPVL+yIZWZ1prvoEpfrOeyya12j/dhwE4NpLOaqBdnavCn3p9qI9X7lUpGbn0SgH63
lH0R3t/tLiQpJsQMviz4fbz8Gad7mMfhwFS3BsdUt580DtifB1kGnGagc1sxr+X1+UcHxJFrrIkp
Dxt1Em02P6HYhlzhzVFhXU/IyKl4DgOWjKdY/OY1/Nxad528020kvIa89GZ+l1bIWui8+61vA7XK
mzTklY9s1gQ2pU4g+1dtUdLe/X2mB7EIMMSGcMVbUgSoT29Irw+VPsa0f+lgN1GLpQYgbA/E3jFD
dvxS3XOmE248bNkSeTRAXXj7d0/xVgQHRtdBDYn4LI9dzZ6q+GiKwxigwyeDoPX8wCfvTbQihjsu
ddLRy9zfQK0V5nNJOOY3SEgm+zBOS0fRTDyZqstCcJmybJzNGOtFhv3XcdAoSI0MLMvm9D3SJrx9
8iFZhsns8lBBp/8jryVsF2OWVIPW1qYyE3ablzTYUFq+sDOID+sYKOWBCRcWfUFdxJEiPXtykp8h
L1pw5C9G29EKDnHA3FlCrTOQSAXCNss6A0lYK0Rv4ITYNp8XnLmfMZufR1kqQAnf74R8tGnR9jTv
JhCQjqW1FrxAptL71G7ZTU/+OoJ0PPqAYr5g35cHFFiOCyoTkOvuI89BHQPYmW8sPnkHAVhY4iDD
zaJqFdRx7EGpvEK12yoULX47GywPEtA7A3KbYvSaMdwOPXj/rLHpoSWwx6JFAJpBmHSQyd3fUzDI
F8Dl1NMg/FQfOVqaFmu0CsCUvUMjondK7GvWO7xMskb/dPHQSgXoxUXA/TYoSqJdrd/zvQaxZRFe
L5qq5PIz2TzbTKhNyU412JUjLMeKgX2v88j4ofVMr2JPqUnR7xwv34EQfLo9gEToIZThOKsdF3Mb
iD1WAlc0Il2FEYO/09RT4Gus/dwBvlCH9U46j/OPVTMKXJNqxp58KDvhVRx9ULhZ6Q9PO3hTj20G
Cv3Yu3zgD8MHN45iZXQGhHFqvZTHuqo2mxsJ6aDP9dUGAF4fLkeB+gsuseDLQZeNZiYYeB2/p5jQ
5P6qSthuEEYrKolFQb70xUS3AZQQMiKX2PdhDzLX9E7vpPSVBDYkkpVrZi9wb4wRLa/L4PP9T1xu
11z1eB7AcHtLSzPZZVBqLWLRlGIZIOExn0woWoj2JTh7L0Wo9urp1NOTeVfEWrgR9cyonqARdC+E
dY7nkhIpV019L9ch/h79tScyhmLhQuLQx4cjQkAQ1ZwiWE6eHylsHwwp2a2auqnkIVTWqcF9r32s
mApYpnlljJOGoLc30P9bnGP4qbbijhYkonl1SHNXI5fEwvu4cbc+H3tEKhTeYUkqoyGbIuqvBYOg
KKVhJBwgblcC9PzM2Z5VrhI2tB1PlVzJWpJKpXy/GwaVgEz43Ow2uuNPG9/MnJCQXIGPMzG1DHa+
riHQkMOOnZiI9TuJAvg5CVKzFKIpuUUg8+KqksXHP6OgGbV0pm37IEGMDts5u8Yhag4DJqp9RDEQ
2owi2jP+EjQbtuhkLkC0U91MaQSHrZ6pTH+N4Xu4nLDwaGJvI6Oi1qwWSg2u1c9kAZGF2Wt4bz84
7nDAASUOfXuScTQ4j+stLoDigeUM3+PYYD4IidYjONYRouodMeSDWZAj+x8pjoW36708RzCjJYJ5
FTcRqyBsFFO/pvkz6Hbg5Rd1qB14Cih1cZNyGJwYOEadREnP8sr7x9du6RO3xx76ZUUx+fEscoW6
qirnbEewaPO8C4zuOkMrrktV2H3tvWExVSHE/iehjl2xfq2mjivulfhg0lvZVmOD1H7Hz7oaf7KG
Hm1B+WeDF3BZj9YcUn0fePMwvamwb0H5gltIR3EPBu9WKjL1KBE4HPCqaHZFwmIoP1+hZQNJpljv
tteFaCIHqy+60pa/36CnGY9j6SC7D8fM5IFImkYdCWFV1O5DRRHIN0rAvdNbeniVcZRElkOgeKbx
w9MTvFpIlKRZegcJRJsm/RGyz+Qg4sS3QTyJKV/xs69+MfG/JGLLDdiCqYTb93Ty2xkZGB4lw860
g+5LR9VDvNkjIAsboZlGzDa/r4wk4Njm9agRY8dH0z3yuq/tFJx+sAC+gial1mAxUkZQc61GMepK
Yww16z1uxZhNpdkEmrXg0AfKJprVzTE3ILTi05BBP2hTa8xL3OWoN1mHrfk4NymI2wDEGTXyoIVG
e+azad6T+lC0M3FXmXm7FhOJdL0q26TepJSaF2ii24IKNRAOvJLQY8CU1JSxepawOMdgmwPsmhfW
0+WBK0mswEiWwHQWP/PQT4DpoRIFBh1BKFCGGEP8EJa5yNAy4aGEHJgR4E1+uB9y4E991oX5gFLF
dDdD5vcIFEBEWkInHLXl0F2X8HMKVZ4uZFViIwfAz7nSrYbF3edwu2o5MqvVbo6xcqeTIi1Djn5X
I8cWipjWku/qwnAEtHEB0geyoR8izz0UkEGhHfgEk2Zc8oiVNQyWYDZoNIwZrOUfc2zdeDMRu33b
AHgR5uuhFnGY/6qeRKz5x88PeeB3Ixm1bTXe+HC5NByHev4WKDFiS0kTsZVQ+2n2sofiPtf0SUln
RnyNxRQKAM70YsA5jkrBnyirmJ1rBMJh5t8IiBHjIV33/V/QzMtzoMRINkTt1uu/rWNUqkfuLGQc
VcgiWoS4mJzLmCzVsgAszn5lCoBERoKOFaIFljegHidEYw8XlsoMR54ZVoh6NJYGHImDAPCBE70b
mQKk/xLiWGHeXf4qLWJzMaoIMJeLaVJdfSMCU7Onoax/wUD5/43i1+SUW7n2Byzzkgd1G0q5YlVO
gv6rPX5FnUMvNeZQIdUzSQpO6Jj8KaiNFD05mmNwaCTOxtQqQYUtc+Fwug6aC9NgKGpyvpj0EkrX
b5FGRwXVp7Fsy29cWA1DWrLiyclvVeo3AnM6LjLZlcCgzvsMojup/Lbw82VTW9g9T1ZPtBp7zZls
jcZhXvy1fCxzCPcmTspyMmbZNNX7GxG9MtLR05KgF1AgdRs3kIlJCG4PFvMwschKollOaUDL8N93
0VfUy0haLcravaCh83byypXddEav6t7mlhmYYSaX16TS1+irpvYJ+G/D98zSlFLHrWYJMRUxyP+D
0+rMpPZYJbE4Xy3RCQpMDSqrzPqyuAGb3nojftnFNJQNK1F3tDZh3uHPd2h+c6RQ1Lqv5ul0U79o
5DmGmdvr24zgTN4RBp6Oaq1PfaYsLKGVz+uOakQwhqzcnXFaeET7WCU0AUT5kayz6xhsngK+71g/
TY/HGHGHTMRvsPZIUsmPki/DEnZ3zhTT9C81ILYSWuUad9gk+9z9hnoceEgEHDr+Bu23SSQ99fqE
NxOS8NDoKwqmo33vOLHM5Zlvg4AjEg5woMazwjtz4sc5FG91vYpTiSY6/x4bmW/isPddnAvPFNb/
wmVKNeOlY6UjTqfgF9C1ZqyRhhoadLGEGZAqKCYzhYrWGeL43F8RFPzkA/LstGal9Wh18LAqal2D
MDQUDntHS0hi+Gsle1lGf9NBgiedKZ+L0oSmTJq4aPlThq95SkLYD1hGLYkPdKa2aFJbm4nYTLYW
E9JFOlCdKr+8x2xtZTnO86a+pWPtWdZoVTt30YjwMFTNMaddOuw8GQZZ4qFCQQnEAgf7MnkP8142
tTT800PAbAUm9eMJWGxUZvfpy6aI85qaDzxVt+9yPuO0333x5GOZ7WsRh2yZNuEjL8V0Rzk1LAu0
U+Auf5becsmbSqo12bora1HSuw5DAS1dYc1U0BBJfop+4Tk2Rc3JC/GzyGpVAQAG7pkwhZP15wW+
h9vxjSWkPFsxAjnNpyt1yGTVVr6c0+BkzElh0OGq86bNIXNUyOi0k35UAVu5hamQzbWLYdjvj+OA
GwMGonmPTAa0vcPMr0Dy+7ouJ8dnp8un00DM7dyOeCqUZCUF2877m3waaRvnIY4cG7f4FtEqA46Q
8fyWP19GWQc4SYYwC7DsXQDef2rmYyirM39MHQPnEFz/7gLUc5f8jSB7bvvIX71BK2XGXEQ6EKs1
P6Q6/CK/s/QwPY2472eTyvGBreoPIHbboKTUMboQHmQF+YWmuvrYcwIZt6u0TALBOhe/UzAk0d2O
MuWXA/OwgITQBZVXtO95IgWk96MWHJDL3GA9j9J7OedCa+C/Vj9hVqNl7GhCTjv2ghebMWoG7ol7
k2LU341snQyaoTtxaoyxwjrLBgFth+BTtaZlFUxQ3DiC0wyAjg81qMWAaBH1npR63Yni5a+iYA3m
wRtTKyelwdfzCRAheGDwih3Ilj97YQ3pdHUE1zSUxYw65dI3hZrkvYw9nNl5ZNy783JNDeSo9/Xw
i5C3RR/L7aAGVpOHWVcKqYobukyckLmiQvbkhN0GBeTTouPLJortwFCQbyi6HZapr8Y+0SrF0jGN
lxkjn6K6RLCnlV81LxX7wV38k8Vj4aw+67K+TTQ6NXF4Nt85+yIC9ESxGsSPdBVvtmgnVsXPOeB1
NuN8u9yU1krsPddHU22avn+/mYKel4s9Pu0soFWbH89Io2shALnHPHMk7MRvP8hzzVMLq0Gr4BsV
6hbbWXUwFydrKhIjW6mmaxplceF5xOWYVNvDJ9GP4VFffXIapFq+n4IGCSrwW/XeUsDjnIVjIdvD
6TLtii9xZZtS8rmSIFkl/HA6SDzg6f0he4Y7n3+ylvxv47fFr6aUEqGuR0pp82hrIcwjFM77pzDu
wIuD4FPN9yN/urwyrgLjn5j9Oif8U4WtdiIMPRlD0nWCpqztLIEBNoujc+XjMFEuPjjW8SFPplEi
nhw+gS6/0yeWwAfICG099vL2gslcwrrNtvcAUW/UpW03DS/YHGDCoThz5RcVTACHHteepoW4DJul
vhDT5r0mOV3/HfZkQhX3JgX/i74iZBrk4olYYWg4CywWt31rFsbRS3MkmfQn7bWPk0wL5Vys00af
NxCPf4LmYD/ghTtFCSyZoPTO+CwLLNHwW8qPDqeEvgRRhZvq0by7RVtVMoF/N3sjs+rQj0gLSq1w
xoBXFk1pQe+3sDePJrJiFV0VzrTD5C9kG6wdN0UQqlUc0Tw2dYAdkmC0sPttSI3kKkYTLnFlkEMc
7NeZwznKCaAHriQNDdOk6MPBof8xGgplq7+FYdm/PFG2nLMO9K+pM7u9sZePZBQrbXNCoL6bxpod
XEqB1yO26zD8CAacQmhtvUnhu2W+8GIUlfq+QOsCfcZsuJYvkZFMKs2qMQRuBClIQp471N6XsdZM
U1uOkS+/hqKDVohzoOlnrrJWgDmjEkoGIE2/a+Ig8nZRZr2ekCNM/BeXYSRNtN3d+d96WUtUPzQZ
/n6GywdO+96eG+DDG1e5VaF7m8mOdssUu5mBGaHDTr6Q2Ij4at66fVdx5Sqd2Ze5NNIoUmBIcapv
wH99mjar4mnaUr7ikpxfnRq5POdPyoca4ltQm4BV/pUt4coQdUsu0dH/CirXtUxrHBIoI/sqYJlA
mpa2V6bLpPSi2ZMeWJYMIluTfCEHx/ICWhM3X+QIqr6G//mye1A6q15mt7YNPeBK4HfF9XYX4DuZ
9glFoMB3g61vUmvvYj4e5BdCUH/ChPMKoBSyEHZJwwnXHtteDmid69RS4UUJAv1V7M0WWfJONAuQ
J8iPIQcDIu7jTapY04Dxza+KkXfP6PQdtN0SihCujBSE1EXa6itddyrxUAjygFFgY/E1EUMg8H9r
Ic3c46lxbGTcR4tyl7ecuZ//IYca40wjqVLVA8JhVZIhH9qKte4D0E6aIan/f5roEWqsVbXmhqpu
pp3F4aUc7oSkaTwXgYEoTN0I5xg6qpX+bB4joPX98gAXw8CGaklEQieKiSJEfloL1V1IilOpKIq7
fGcuOGayuljFsQiO210p11f6a9xmoh68y+rw1FN1jpCpNDWWUO4twpHXAWg2gIsPcKF+l6rbsrYE
aGhAi9eOkv5uPP5OSYZg8LSAj9Qf3gy1eP4G6zFmjN+wX9E/yk+lBsXze5iXPUAKoYTSzdKzLSUx
aIwfNa7uLsooNLvMjQu8AgYv4NEGE8ptQCaz+I+qCg70G8L4dimyml4dm4GwOEVNOoVt4oSrGzat
lmNQ3vJFBbC+JAelH9XJG0bZu5nU2wznD1DWuuRNosQGJOorF6thi5p+Hp1y9n6xkNkAke30BqLU
66mzWl6sSJ229v1Atzis0g/xKwgcjoJM0g+/Ux1bqo3Pi/NLWl+TzgnHBw8pk9YIt/m1bSTJIqfp
f1lbWPBgnH04rrquA33MrDzWXSQwopOGovuOz/R3iqY/gZB/d9D/u5PpqPrbSw9xAvcgSwTgPWh8
qTbgAwWi6RGScp6dT9OeGrDhN/wuj+3ntLqEmrXTB3Vr1nb6zAaLyqXXXzaQJXlmqK2/kHfL/4Rq
POFtEHfCrG7XX2g20UlM/gwmFeN60L6hNNFP6+SYvlF6Q4JkEAcGxPZFdmFbeKs7Rpl8qcVVqRnf
Tf0rSAmdvigJp0F5wDNQbgQpJltuLDcjuYfbEcUiwrOketxT35s0k0iFDaec69X9fX8N1iIlkM6q
wkm1RJ+yoiliOMpwgtrqtNsnBdzVX0IInOHKjsxTvLB61lqTlFm0f5bKpWZnrMq/p3ajli5ZsVOv
5POUKpJFyBPmY4UozWkBTTyC0aCdumCUWrdViYPEXjrCBNONAHuZ6qGRiVjQpuV2zg8CsiBsOulK
Sg+RWbfAkGOnAxMYWVv4htVMUg/E7qVy5xC3BB3U85Gushs49v02bG2NyPuJcjOvs6DvAjlG8lLD
y/8yTbjBRldYjXfo388Ldw8xjyltRkh3Y4quuUBcTWRQyO3eHOyM1Nm0+DE2LI5VjWhjPMRjmIUM
0bvVsLfwhd3GW5DG/0FNj8Ig86bkvfa8nxNG+tbgNP7SsKPlKa8TPaxu3HPPtNQ/+T4TCQWrWeTB
BylLxh1y5sEXVZZmFj+ycL7pAQkwqHEttDH/F2urddb++LABjgKT4PkGpkIUKKzZXizY+cGKvT/e
QcLBrck0RZ556MZQ1CyByDQhjH0fCMYM/lGMrkZeuk45Oova8M/V2XBzIFU15/Krt3gQWrKc8VQv
dvk4cXNZOaB85wr5fGU7uq2csF03j0HLrCV8ML1vJ9sDdWAxTgIvfv9Jbr0zUPRmqmgn5ah/Fo4P
hmhsmG1mjXhwaTim4Ibl0Bg6jNigmpOaJLgbuQ3Gd1Bfe2/nt5WYMf4HGPwgwEraLX4ygrDtZ6Qe
2FpFCbMs56r+qxr9kPifMwsTRH1tqdsMQccEj9RM2xjUI+K9U/knGk5zSAtXxdklZPd0g9lxf/PB
l7yjDStI607DSjufud5g3QrfKKd6Yow24mJYVQGuPd6kYGo5eGUe9V2d5/OsF/xSHRQ6Mf9e5dBu
tMUssu8A7Qclbz2o81Yvl4b8Z24AR/K5lEtjwWH4H/oyS9J/NXCgDtAOLhg6becEICF+BG2XXLKK
ahdGvn0gZLlVxTIi02kfLgv0rlIdeQvBJrEDx+1YGtDjvMrfGfUrDNEvx8lNbM8r5TNH1XpbwcZe
nmUa1ZxRvZ5dAqS7qMzW4BUnZPzYAyxBwJqnLvUQxlbk/1srZMdzu+wJlgORVtc5jC+A1XJYieIu
/vzKKhnI6tFepYDWvEGMD/ZipPyWF8vSguko7EBc2A6pbRxPeWzTfhthJelHX/9HpPOOgsPkNVeR
t38Eu6oKMUV62aUHYiYVCmJa7O3A+KvjBXxrnHGCtf98I9LOMVmev1iIpoFnX1Oj9ssmEnefqqwQ
Nqqb1lUchuzyC23C9CQlYJF5lWKeRcNRYKz8+GAxjSnnm4lBcgnJu0t012PDU5+xJulQJiN3z4mV
OX/pTR2FX06KEMYOJM0BV2w9PPrsG2FbLfOOSGpQAQ8EEBjQGF/paWZq8Hp0YILAKSisypuRCOIn
816mQxFp9dlkYzrmvFw7FTD590pVPp48yw1S5KAgAPvNHrga5PYkuJUeW2YVbbr2KVkODyZEpU82
vWCkQ5sIsZS5U2/MiaQqq3risskrZP89HykwWhkBozHk1bdLjwnov1MnK1eCYxEfi4SriZDtM/NG
HCrTiebTY/pjJ1zOXwHFYNtEJX/r+8lhopQNFMl+zRNUQ91jGXFLgXgwRhfhJIBD2xnrgy6/b1Lf
V8g5axfmktXK+UrR9++XnybBoRY9HZR8dIOdlXvNt9ldFLlTCeeJN2atDQcVtbRjsGKWbXCihzH2
v1X9x1KhWjNfK51sio047f6VxqRh+CrBLSurUDH8nmomvuP+6jOezqUGdqyNXKaqnct142LVEdwq
yB4ojHEFkRacT9yjH8AMDBc1KiuFTUne/Ra053qxYUdYJtR/eKgPTuN3VO0vSjzNkSldbs/KaFF9
gfA0PQZCD2QrzmwYnDR1WW5RSErZQZbgZydhHT5mdOC9pXrseDAn1bRZF3v3q6KyaYCmd+7AcmBM
oNXdskZFyoL7wuDqeS+e8a6pZ1aHYaJ+lB1vbAWMDd4DqXhdcYkiBg0Qq5sziZeEnq6lPcteA0ry
2HrRbWlvdKdrAcFfq9xotFsNofzoB1BEXrB0LZMmo1xoArLEmjJQqj8ubEH7EG1GHpEDq+49z7vp
botI3WYRTK69ByjRsfG4/pjBeiZEwZHaydp93suLMMzpIM8P5GdHl2tKo/tF7cJsoPb+RbdzAtRB
XGL13OP7bc/cs3wu4ADpmgBO3GE7pV+b+09dNnwYof+4fzTMTEKebXGDRnomC+B6wIICsgP6SHhD
0AbFq+UOvVKl48ipGp/sRed0ajEyCumprG+Rvba43muEnDUmJziKyHCHOnpPYjNDStHU0msR3PmJ
NvIGhWiR2CVWrYhV+/IbB0IGnYsiN/69aO3AFQ+0vqlj+o1MjVjc3NqTzqVJlgP0WaBysiJv1kPT
c9bOftl1wk3iOBqIKmByKqLJHjoY7B9wUFBVNXcgfGK6AH6JY4HP3d/m5har55OqRpqtis6CjJcw
XHTDpdPinfZyY2FUWEmo/eYBUfXhsDW00hyrgRHUqoow1I09CPhv+IhaBSVowOai/lOU4Kfp/kWo
DUv46YRxTc9bkKVkMUftytSTr+Ds1WWasW++ryo3li67QCyxvtWwFVihVJhmMH5f/1y57tHiinse
nV8wYX4oiuKasC3heNfTVLy2dM7FLv0RjHZ3nbOdh9PS/9lDgFDHvzmrWuJJBCdEzoJUWiNapNhg
+hhhMvZ/uVRunQEzuDLMAJ1qrVKV0HgbATZSqJmlP3g4vX4Yipaw5DKsH9ZtfiDbME4yFyFL6SVW
pHOzr/hlWxy8StjMCztkIPId8ilcC+gcW6GJNTW7/4v9mkd1X5gpTh2AZeUURQBzWdISZmhUUljf
x+h6/Kz6fqiOQ2n5C/dUPAIQt3iogmXrSW300jTiY3OzFwpF4DaJf6fGVDLEHJBTb5JevgqAE562
9Ery6fLiAubevkREU0zjjmNH1bNfCXPpscJLYKgzztllGLPM5tCAFhvVNRyxWk28aekyufjOETxf
oH+/cmju0oSXT+XTEH9ONdURN1vil5CZrZJQ/hiHtQ60vfP/TNUazBFCIxSB3fZClZzpHB/Hk7bN
0Q6OV/dM+HNDDte7IwKW3Li5ZmjjaEGbEdy1QlUZ/idKAnR9qgnNku+Av9SLvWuirrFOPpB7jG+m
ecmx9pgkfILDgvv+SHm4Ifa6U4VyNUme1ksA6oVReSG21PYCVhPVqbDJdG99Xq9k0Dt6bo0RG4tK
yyZQd8mL/6aQIKLpmDysnt72RxseJWHbYxS1O5QVoJ4oLuj1VuHIP2x1qwNhchr/BZ/fI564Pn4U
aBwo8P9HCjMJ3Gv1LsVPkwNGcsVFrtYJnZ28y225ywdqg/E8uAiKoWH5gVAvL9Xw0D2s6XiTb0zh
1uOrCV/B9AKSeSG0gwizonBVAJofNBfGxnZJXZ5enH+sW864GIgd7nqi2f8cYMqSxaUzUmGNbRw5
U6mDsZpFWBxfCQjXhAgFQBJeikDKMjz/F/E1SpTlTs1KxHduo4/TuPb0xlJElBMpg8dyxL94gjC8
pbdOC5orgK3lEI2yuyYIQ+oz/7BaryBiOQPWBwXrv29yAzQ7z6PbXddlGjdG56hPd7A8TA7avzWg
m5BAjsDMx2x/vW235/W6jqW6DD7ZOr1YQ90IJeg+8TdRh2HergWOvVCJt9Rl5oBstO5Y42Eo5bNE
qALQImZZDIpM8PTBUDZodNFS2wQ/mm5xQs9O/IMMbw8R18IAA7Ysi8P+xk5bnqCb95QLNeaSMc7Q
A3As3GyVuMURSISWnqkmrkPDQsWjrZ7qKl6xmSP2ErvrH0C5JGzbWr9oCfF0S5vZJoubpwCeLcH+
Q5GlmFcWOy4+DVJyEuFYhj/70dzrj5YJp4fmIBpBIA6Y8Cb4bJ4lcs/VPcM65LyEegU7MLiEWiDW
BVwsretU9VbEs4XHdCxbwwVThlWHPqe1LpP6l50sE9Qr4dvozIWEpkPl0IalFprvYwgchLAhE5ZI
p0Rhi0MRy1hTXZJKbxET2QorN+DYvvVpZRDRx0cNdbymg3BoD6RnNABX2HowcGCKRabokMu61s1+
RhgQwsV6u+p4oGFS0qzOJMG1ah4fNi5/HLeMJHyUw3eAi1Z4mb2FbPZqh2COnp0yZ1vWZdFNI4ao
jwFIwkPV6EieFoG9claQQyrU/JGIVlzd+BEKSSIuTzoNayZkH2UrsS7PHjp7+LnEM8RD/9zj9zya
zjHX0zXT8eEiRviItFVRTPrzIFvxhULFwVwiteT1WgYzlMqRx8WYKTO3REzWFkl5fhBca+H15lbW
2/Z/r3PoF1y14qcKAoEQdWT/cTIHsLgTzhS5chImOVfPTwaw5AnUNfS0G81BBTt7F9vQwsgiih6b
yMERZrEaI15lOMGgIVIbcK6x8wcgeIOQXjWSNH3vETZONwhwz4Efn78CBta3NWfAgMCiiVe+CWN3
hv+I0Y0Cwzk2pO0KhAxwucbTQaz85tMzxBOXXby62VbeQEvJAuquzoLI0JrEU3ug0m3uzHdh10Zv
1xCelmtR8fkjAz37UKBkdqe2t+8TY3+WoTwr3Hlat28uFUo6H80sIVTghhnZJ7fhy9M3PY3ei5Sv
ghRsPs1Z4UmscIKA7VkbkWRb0j1+tcZ9BamcmYb4YZh9ZPz5G6/K4TT19jqZVAsZVRsfG3KQGbln
4/y8W/v3hZK1A46M9U8ooq2c79y1XrhfKi8UdF7cM3c+fWJE160ZcmRJ6jQDbXOM2vyDPo8owo+r
c+L7yCWDfdrnXwbQQe+OuSjpP9NrSwF/5cdLhcNeWW2/Zgnu6xmbJaU9vtYr7FeNzPKelyxie/uM
vnSQqzmAYzHgbflT3PpAC/FvjnHTCpisdUqf/6WiMnBIEyPcOz02NpTr/OmUsPx1YM78PZk2bBbh
CJ5U55/Ki8DKVkAEMmAEorOxLT4J8fvPPliYxmm1+mRlgw57qBDL5EkdkoUVXO7n8O6vCz6xK36r
3pHRhRgpLWAl/yC51nuSKXKg7vLgHljAQAHxKQtMQB8jToMPEZYsBlEVr5DCPOcBTm/7LPEIzFCj
CU+CZ4POkUF/+zFx5lQLftQapbyjfP83RQ+S7ZRzuPJHgxJTX6rfQoxURuOg+64Gd8lQu+3c8vi1
VyOogComG1G3rf5NU8vY3RLP2ZcEVvoJqJAfM50yzliQwfJ8u1/RDkGjCpZJRHol/1zpFhC25ZSl
P7W8pz0qgKEF9L7VpODCe9Rop6DaApnyfQ1WQRLkN0TClH9AZ/FYM3y1kWuswjM72BxbL3XEOGK4
OSJibC8Jp9cx2u+xFxCi+WB/it4meQBKtARF0YjSHS1AF8wykrBRcF3ywJI7dU9XziOQYKdJblwN
gDaMDdoIFkNiN0uflncT1PaPZIJGdzvmJuyZccfIw0O5sfM+4l+ULKnDgDOfICzsFpKXom6FgpGK
577DBFjH0NpILwLLFKqawk9kqeSfo3M3EMQ6SncxtJORUPHjG60dUgijjwUcTpB5WTLdCqQEVM+T
mbSc7mLJuV49xqu/vod554vA45DVPuoCW4/y88mns3jlsEyOU1OLaUalmhByfN3H9nlS6pgNVOWa
v5zRUl2SUq0XOw5e8GoSAY4tgQ+MPyYUxwhle6vkkv5/+16wVxvW1zHqbRmvU6JCBvFxZqJ03FR6
Tkbv5Ltf7KsHr59C+02ixdmMrZm2ITuKrwDReRcZb5KXr31Hc5mF2xqvb+0LYxgU63Ji36Nj/hTe
henbTIDEFezccisIAqBhtd/9llRlb8t1FAD/8qKQ1U7sHv5hlzwvkTRTeG8NgdVBT0JpDQkxntNQ
Md+LV4jrbQol6x8w4z7moBSUaIMty1Snu7XwwPKL+IaAjZkIqaHzb8neHuFfijZzVS3Bm2Yp2MoP
cb0TG51R4YdBq3x+triPZkQW5tsjzRK18vTX4ku1RiLMy4uZBbZEObma/ikFeGJBRW3tavlva+7+
fD9suqwDP6y4Vz8N5SrCpHlkHnf1BwDRfa2nr6FLW9Pu61VWFwzvAEqiN/LnGNcb5XLUq0wRRsT2
AiOCuCDMlIjhfC2KQipVwG4pFq6f/E7kquSwDFutITynPWpQvFUUQaJHaYOIHzNGxL2Zp2ADYBnJ
w3lxny3cgyWhperq8Gbpv25X0LAj+lhykX/NSKWVe649Gq349n0Gd5UtmYyp7yGJXenoqoqZbDpM
F/Ty2OeOXyp6LrpvAVIGNLuyDyWmm63PpGVHEzq8ulj5mHdDa53M/Je+3tmPEkXfIN1NOegJcP2Z
Qbhd8P17PRLodhCECkGEQIzfd4uLi132F5i8019Ml4YZfvkxEwTNGBAR0TvtBIfdvTpFHHflmhgI
xuA6/1+/ouOWLxCBqQKFk2Fcl7ytHwcRMEKBdHyJCoKDsNz/cfcm08p3AlGj8yCr8GPjVB9yGQAK
AbUmg3o7NwkEjKYSN7LrBlpKdsZCqzIS2o0GhjtnkofbNAU8UoyN4O2LXlErTxgsoBGeCb3aWbD5
Y7X7UlSxDkZGus17Dh8wgW6twd8cfm2bz/UYdGPxflVN6UyrYC2Iu38K80udmvDyx1PMbOSln91E
kzPfp0ueh8YXmwfubDeWIeXD/ISOpW6ZwBSEPH0zUhNjQMfEF5n/OpiQP9S6wCFk579HySzueD7Y
Txm49XQsKsGKxD6Mp2O3B2F55R1YS7aKdn4EEF0H8LXvRO8BYFfQOwoUdlageInkldhwv6CMqtLz
HpDmNSatVAw85yNhJvrBRhQtj0gmH3ek8NOVy9h1vv1l5l4QCRq6ar4Z1yoc31OqhEJ0cp4SW+wk
pO3SvY/qeWVlEEAlTZ1wH6mlX1GiHi0nkxxSx9aTlU5Sr319hSm0MtTrydKvYa9TK1/KXJiIEqP5
rByH5bmoIYISCD392zvOHYxk7AgxYMSlDIs9RGId0ymvoD//7eKLCQ08DFFPi9GBhjzjqLhv+Ys8
F/SqZXYBe957TD2JuCsM6wYq/1NKYF78KB5dCBgohz1jpIKSyWWSbniOCpLW+KCHvktGT3R7Cv/j
H0qdYZt0OhDUOmVefwWNAWsA0bAnsa4pyyh2Z4HPAGKIjnJK9tN88XK2QQqZhsl3gWSc0pd7IW87
ix4hPxayowD1SXT9dmM8vr18TSC9SKh8+KLm0YHAjca39fspaYRU3TGEANeNHa+puGx/+IS05Kyw
Van/HNge4VPZpwEu490v/Jqv6rrl3GqZqjvsDYQ64QC1FsvakQh+j2z0gxQYRgP973n0uP8qM9hy
ubJeZwcI47i/2EjpdawK6sTe8nWkGPJ3u0lO0PVy2XRuMYH7IelOxQTOJInX77xAw+kYppYAMcCX
twOJ/716g1sFdagCoPUIztpeW6dOnH0wYsySihEzZYMh+Fge32LCT9efIMge0VZlVeeFm2vbVh/K
qHWCoLQk9a2V1lVH5IezymTLamcgN1Isj1jebywpymOdv6swMVxrdFP1iII8bFJYv86E9/fgrjmN
jFMDLS0pCCYWLl21H5DBOxnwBvpZzRl80lxiFrkw3j2QOlpSLj40tkV6ffPcUQ8lzTHhCK7S187l
v1b1LlXWxuRvMOvmKjBsjWutBIjxosHWfxgRLPgttLt3Wmo4ZqN9h06GYJw9Z5HVL8MEcQyKn5Qk
9wJm/qIV93ZlUgCzmjWTIcHRR0jwDOtY9efpxHbckxo9RWYQQxjobweH5Sc6jRg1c5BpR4d7EIdy
OWzqG5MmsBj2QbQif1NHXTujFIZzCR6yFB/aonRd+qYdIzO5mzFOfv5HBf4pgkNBVw499dOpN9AA
sCtLhFx6Gld0ZVKbyQA+uT303gcVP+lcLaZnNt1ao4vI9Y5KnvPM1HsBE1p/eNaKsHb0CcuhqsNu
skiv6cmCAAVTTF+SIYmX4tq/Rl88Wt7M2qEgvfUKEOfhPewe/GUUajetrWk1Mzcu7grYDyKrr4Y0
VNSKKkf/ykqF54oQ5HRGH9PDpMGrKrba9YP4WzIpjWJuUYRQMd3/ADGM4QE5c4Xh5GKkHyyhB2qr
dwYwFtWo4OXSFMVyZxMyQsbQjFmoFbeuZqBxQfjFWVy5lzIyzsSgAppeThG/zGArmIZcnzAIqCpV
A6eT6IDipW6qkRBltr5GX5ZvJw9//9R79uV5f7EXYTFP1JSoiQ2KF8W40+zdEMWNAO3+kFn9g/C1
piHdG/nKLdojnDhvBD95TAcYucMY1uj0hCS/789k95eymIPKRu0Rad0VKKCqMvbIIWduHJ5IYDwh
v1IDEHKZsyZugXmE/v+jUL5P3XpH6w5E8IBX8F0BEMXFxyghrJOwujoJ7s2FjuP07+D11wyCmthZ
igCeGqm5lmBIuWOdxl/V3J+n9r1AOliU8Z9gRaSUqjjfKbadiX/NfDAD9efEuxCpQKtpmJmGIEx3
Otx/G2HBL++okeA5TgMFDKfkulRKECiUa759z1lRYYSwW1ophj85e3z6JDuV6/NHJrKzR6Ii9hgU
pKc0+tOwaDQO2df73bAgAU22Ov4tXcDL38T+xgTimM7Dg4puTdlJkzTt2EZJCaW5UdG2ARCPedId
sJ5Fho/x3KMEaZUkvyKAhcn7mxuXY0cDj75HqVB3nW1wLmtRn/V7hzPb1N9X9uRdAC1uCeeVHVE9
wwBy/6sPEKYN5cCkiG2inlyouKG2wepiMk8ghlS2Dgb0TQeICdlvi8Qd3st3I3p89TOcFEHHPGwp
ISchNcKYqEek6siW8OZQk10/S2UoMw5pBvt7dWqq3hbd0le14O/ZIKWmofmCWouM0V9Jk/k4Kr4Z
L3zjD8sfbu9pE15LkSl9Ltb45EDCaHp1sgBfaCjybp2n/vWvUvghjAxxiwXRJ75HBd5OGL74elbj
0HfllSrymrahrgC16YWcF2oqybOxYTk0VMCPtpjr0TpZDasJLqOHoyitvVwZauqGnLMLzYifKALY
E/e9B0/f8gzGnlJtZ6+Z56vd+rOIYcmJs8BxYQwQTKEzYo08IblcDtB47cDlRRWiekwqo6O9IDBW
dLvqnipHGzKrqAHnYy6VzCHvBuMd2XkEqxhr9/z9BH1l0SG7sPzIHGLCL2U0TJGh7HGt8jBfk0Zs
mXD0pMHdZpGovmq/vvc3oWl3ePpVrab7xOMtkdaIS7TZXxGCIheFei7UY8HE54GBEiMA1eFe2Zto
0Lwv28Ulu8fwnbhKuAoF5kCx/uMqYPGDQEbSHKd7bGW6JZJwAFV1N8/+qawBTdaYNSw2qK+wky/n
JDBcD0vow0uApFQQXcx90MEqw0LMns3dZ+sxmPRvISDe1nrdTqgnUecfmXaslrRtJf4QBsVO3kFZ
1EJrdhn2FzNtkuvGsft/bLSGsVbwSvi6h5faETLeLcSQoaHWFKtBgTlV0r/CvNgehXcZNITBrZe8
5fE54jni9iZVOjMGOgxql8/EwgdTkHK9+5mjexLkJ/kYNSp5Z+SU9MaWVIajEnsrv9FTHFPXc0O1
Ksqqu7Qzea8fylTRPIT8cX1eXN5w1O4YoI6DpalJ/XZokKtV09jwamehMBWNLqLQGex7PIMQyPf2
+iclR+ZfD7Y6Q1a2Unv6fbqj9F/HbiMrCSkFxZakLiwW3tc6LHcgKPgSl3fc7t+HU0QEMtfwAvEg
X+FC8tRR4YUrIoeABZjsKqh3Zd6MckNDJnPUjuTfT+4kGyTsqUA8ibPFFKf+zF1U15FFo1SICgyr
PCwPwMhbPiyFmzCj24YNJX7qIGJe6l16jrrMoc/xPevBf+1lA/g7wBQkOk3i/0Y/sJy96Q5UKtdG
5ekT8/3HgEk2k1n8K2ldHYMwPq10BGwabAzwgbaikMPuouvOJPubTte2ux34rXIQoq1UiJ+QlEoY
/I6Ie7HshTZCfr7rZCB3kTGs6qRH5zYmIa9rvTEqpzAPWFqJW2m+yIqGlGI45UxLLq65aBKLPW+L
QxqbeV33SuXz6nTC99EMymPjivY0f17mJlQjzU3HTjdVY5yT02M+woo1MxXTgi8WLrBp5QCkKKrY
DjoC5akCq6NbLu4/PSjWCDzf+OrwVXgK8e8oHz5HSVUH76zPn0VqCaMP/ZJu6JJQ3mRjjPi8sZHB
FtyJS0fo9FMAzl2uJ0w6pPEdQw6SkWwlrC0wTay9XRZIVt0ntrmaAWuwqDvEvqBYY3hTd69LWSoa
w6kPNg42ZKiI/4mjS8tgXxTQyGZgeYhei5NQMAmiRcXrtIlLsoriuxSqmZIiVTcPoPI+BUQdggem
m6IzvOcDryaLYOlOlgsq6ZbjADd1IKv2nYYcAambN//vIpZJh9tBIZNJUW++EwDQGb9TOO8xS1rY
N2p/Bp5Tohim7F9glfHFhFgmcxsE3TUnYV/RggQmtT7ynOzuVdK/l2R7KzYW5bNhilXTB7Fuk8Ra
CfzSRVz83bNc4KG6aifOM1EpIBh3dExoljFvNDYazaAk9jvFv2duRQ9aFyDM58aSZ0Q/RdEWErE8
93L4LveJ+aUpoQ8xPBHB5ZmVqZwHIDtqZM1E8eniVSBz0MTlJ0BUyNr1NalJj2xvDrEko2mTzv47
EhhjG8Xa//9gSSww/noxUXP50+sZbQJuDmceqVhwFWIKgpSTvpQVXotcSn3S+gLC6lcWtTYB8ytF
iy8B63F+YTWBz9yhCdsxHUu30iQuppOFYtSMt71YNKSDD7C22PFYLnHOF/vjOPKhY1mccwqpzW/f
BxrvubXU26fgTkr8Snx6VZPRr9DEOJ6ZMVmZxGDELZ8QCgngAS8NeeRnfQoCX4BTSsvTAhX+H8Oj
3TWYs7ZiR9ORsspwbnyjZm2YtKkwxhD4rQKT4dVmv0ZRtLpk9jay4w044Iuhd2XDwK/E+59U15KT
atH9V+HXG0pv+KMUtaZBHDRRs2jto1aBacSNT7qRv978l0mG50Hfbbwoegx/BIJIgaxx8xmq0Oos
oADrusQhwI6z+rTnm9CyAXmoqoIgHvyD8iJxeGXNFP70px1P0QEg5YQxKgcfv0+foPWNRgMoXopP
M7eLqcVZPMFgr8z1v41lzQsFuT/qUNmpAril8AiFGgAqGfMElbtsUL82hbFkOYzwP657fCYiXEWC
DI31X/+sAwkSZ1DpzPG6j4AJFcHonDk+FiDqjDxE4YAudpowcOJxs4rMcQ6PtiCpTUMRx32S6P1R
YZziW8nOiUzaHRbRmYIQREGP0x5ETUHrBH+V/tq9Xhig1Py3B/kOZuTVmBkjWyqI+Pv2+J780n6z
1yQNKw90wcEHaqGnogl5vZZBW4Nqh4bZ16mdY62Tu8o9x0EC7WXFSTc3NwOu5gXqsnfPetzVL34p
3DUbpe7uFwfmYYYb4zNQdraLbMR00KOZOK7sosD/lbN0fay2f/9iYaGZbW6AjvtA9vK54CcOK+4L
B5+VxeO/pdxNV/M1pj93pjUfi4cZStHD4ASBUsRCFWnXfjqLE5fXmHbpUblmQzt/z0MZDvqBryIW
epIPdlGdNBGocWveCswpXbSEEJ6GY10n1dAazDkHR8RdPRlase2dPXiDhBv1ChPAAR9qwJxeNwKF
OacT/yiwirQ+pecnIFj8jvrsEYBlxT3mpNKOAPr1kORYOLtnQj0O6tkx/ruOFR7m/tw5uVLMzDKz
7RpcQGZgr23WrLQXt9a0jm/k733XkUiI5LgQRNDpR6y2n5cCnXV4wS1pZi+xN2nNPF64PUA82HnK
B4UcVyrqsvmns4x0CkaNlN5BSh9LSXIdzxfzFSCETLuUD7g6Bg8xTMKpMT2INKvvDTPn27hZB9Si
B9QqvWMVvJsEkd+Ku5qH151IhyvGLed6Aqtie5hbeW1YkMbToOCON1mkfgaG2JpbYHssEjhesfLE
iRFLR0QPpyhs5wx+ptvHZBCf3J5hMVvJkGlMQR2hiPIR6B+HuMY21QRds+Ux50yRhlUnURBrGIoS
Z7bf7RCYeBnZikX0lGosxHZa9jSocqNMHJrylx8hBGs23Vo4PAOq6P7NmjzTMg39ho6jEc9CS/F1
TsGmADQoneXHehtLOLQB0SaLyn5yUWGjK4CdrAJMRkTPANb+doQx6Xiv1MKcOMOtujJJCofflZ5D
goMe2ujpy922V0sKYu6d0pqjKyAjA6Vo33D14oimqEmXhOmZDbL04vAlrSJKUuNkLWCkyzy6a9jT
x69ivJkm5Eskzo4ybqOdZ1pctmbdr8EZAuQm/AyQrLewVG++2dhbx4O3MxcnujgGuwto2BYyJ+Tb
05RP1X6XIA45BZtK/wvaz+T9aahXP1NJlJDGn05NdvzamcB1EXhtrN3O8nL+watuXFJ2AVQYdwbZ
Y6QqFC4NbtEIDeCBc6Vo8arITuI7KzOLRqnFcXfGW8S45Do8yCoNXr6CuxMxya/8JTOxjCNov5XT
zgF1rc3wF+BnYSxC/Ky51LQa4sLsQHElMBDhH1cZdJM5/WmLBedOePWNbCezhl8CNvvBZ7nn2iCJ
lsYga9YGD8TVipG8n2t0Y+Te6Y+iCm7OYJ59JWYXvmPVcqSn5jg1Rul0ZVLAdd/NoOQrfzJgwNEv
LvufUiWHGeM5v1YTPcBWvES0uANPj7lSsQxtymA+CeacAqle+Wx5vwnHcSE9SB6oi+9X18O7kxgZ
wADg62Y6NUziT6Mgxiyu4P7ICx3Z9NmmEmlPPnSc8t9LX+Eaz9d73M7yYctPbq29+J88p73t1kPU
V2CerbsXLqMy5EZtkfeoRCSUVCjxCH1Y42M/2T6EyE0+ux4YmL7ivw4dMYccgT666dPuOZIhxum6
gXiTaRSaoogBJFN6Y6IMisinM6i2R4TFgmF0uO0Fi3fbNVe0a3Jpi1Gq+z5YupXfETCPxpO4u1ag
/pzvjLG/ZfO95x7w/+XwqIS6lD+L7BqKvUwyWXl7CAuhS4216ylEFEfaIL5m8Dtwm6Ln1TPDm9zv
av224YIkkCftp6X/iFSF5Y1+y1xbH6XhpzSLSdmu/X/IgpwVZoQho6+VYNSL4q1QrMcXqclGuCq2
JvWPonvWfE1tl6FJFE2k5hN5j8VH9G9tURYzMCQVVi+B9McAXlLFGmkDDfNbnUHiw+f4RRXCEMOH
vK4p3DQFR6I4I/inenDm9lEtzGsKgnyvm50GT/f3iZFu5ImRwQlqJDeSseGjroIJs7f3wfgbuFEt
fNsyuWBjRHcW9GGgAuO/3aOYx+L2NEXM0A5X/P/KeRIovtzsNtwuvYaQmion76wTUMIKmcJ3VmuU
zL6Y96nLCxL5cmk6z2lTyOCbUjXP1UITg9fI1aIU7JT/dfd6U2+41vD5hb5eoPCR6nIGnLMEzIlq
HQuGp3MlCsuDArr5iguxQEPqlpubE+/T5I+UuhwOOW0Uw5WPoCzA2F/g3NiFeOkcP/Vr9ho4sZQa
UIQk6SlVWi8QjB8+LRak84qI0bwOr5DF4DV4TWqc12eg3rp/piur8Fhq2OPTX93ShZooHWqFuz/i
jmdEjnTHjzP3gkX/xkbQTugsW/M3XkIN4Mmx34skrxSmoPaYysZYlFz+IHxRTAe9EFqEdgwlVitK
SOgWLKPxhkAQxs7u9XGiqIikWzEZoxKXz0qrORHeLS1hNHE5AeB1evp7PtMhXwTvODqPKC9vQwBw
byBEldxeFKeWN6vVGAvj/SeYnZh9CF3YQHcO0XpMvigNEZKDxG5mPbPiZVM7YSVw7gjKUcqCkkQG
9/HA3kB+kezXMJ/dy3jkcwnfE42yULq5iAaTmJU8ViJEeYkbTbRdVJ5ueUeUKKr92syGm+R9aouz
y0dI0iUvx28l9umeCzkyH6GU/2LQyn/08J/7B7/+MFrIxZS2LS67+eo5luJNxtRknpbM4EqpcgWD
Sugpjanf6AgOdFAFMBLS026ZQcA1xmkP3rfrLxcLqfcSr900+jlHK30YDYCQLQk4l22z/lL5oHam
hgNacrOZFBkH3KdmkP9Av6Ke/9gu6BmJQpVc98qEeAh6ycnJRdrDUKiNJ1yBaQxZzJLCiA8grwN8
okkKklDKt6Io5l5Y6gXMvJabSPLDpXLClDkx8ujpRXPL9kw+a36dmArUdUEVBQF6sa7GD8Frjt0Y
A8m4hPKL3vAUAJ12DGthq37f3dFxmgcHc+3MNj+iR4E5iu1mnmtQE+sF2M82Wm0N4Vn6gp75ni4m
CcllxiqHH3jYy3ImGjMga/g0wH79PBlmSQa6qCalyKh7yokwHpT/DO1iDKpnzJYcHUNDEaIQ2QOt
PhgZjb8si+j0fA8ARbQEq1mGytD4+r9yrvj9WgkP8uU8ZJ2tMedgD3J1/G677PgKyr+TdU90GCQx
A//8x6skSMyADUVPHgN0iFTVNobpbYg9vlUAAFUFH5zK4sfhxs9vZPAFh3gjGbzos2hhEOPun1KP
IaIT4sbCcJoc7x3weVd5XJaAQKxkl0HKaB4pj9CLjFFHuf8dVCzND2lHduvtOOl/lhCfLs668QgL
MjJzW4uVa0His46H44vmvR0goFJfKob4Tk/PcYYgbTAtLIZrymVtUUmjdrKDezrFZIDN/R8pb4i8
pnfkJ1AZTuhXi/NxDcoTEGSK1UDFdYRcStB5ZwpEhL8mZpdXk+N87YbFefKTWCvkn27LpNM1g31Q
Ze+Z0fqlgkgYGk3ERkIeEDsKJP58GuzSGN0L0KDJP6BGbT8FYkhOtJ7f1GIf/lGkesD8KujfSbTT
xZZT02UMeh0cpbBglO0MGYKTok+fbMjlvg6t6J2fNwwYQllv/IzoA8u4cZQLvzKdPDXtQqnQ4LPV
MbXCnTzTnQ8gPO0VJZWxLjGfvYtWF2zfwzA6W/dPSrlkQv5szSWGHm1JWL08WszHLOFOZgUpPceC
NwfB87nZaJpcq47NyUh4WmNiAsXPxC4oK6dNxZA1zBkJVgaGLjMB/2guIkFC/D/usUowDVyoChsW
QoO2qNdHzttGZofCv376VILVLsl47erz5qeJxA1IaQC+XlExyZCHYsddNyZeD9pGOD7329LbdeWB
5RJ+vfeN+kY02yTSfequRHQIDB2vEdRbwQvS2Lw8wAKtlUf6NMpg3lekhv7Xr5ISwQAQMfleC2zw
otU/kKrZlnGM/CB/hW1VICn7kSG9EMwQ+Mz1brKyFIMf6QsUCMACf9R/G9W6vB3ooi+ZI29QCNTQ
NFmy2p3SSj93F7F0930Z4mPwURhz3Fmu9rorS5+of6ijVbgQklIYyJYgiP+XwpaLgpZI/h66ESbU
hRMN5ChBdJ7RPZCnx1VTuq8DYhGCuhDzh/REVwxr5qrfwHoOAIe5jemIdzmzJmtB7FKLTmi+u8GW
YM50UMAiURznGCNG7q3la/JxaTz+cwfI+D7+JXcHRODEqJYzuvcSKf4T6jcUnmZsy+LT9nntQrtI
/gobrpR1N/60ttQgPJJWEy8vfdNabfDZYs44FmK4f0Wtbz8Dtfg2aPuPusR4Q33P+5hn/p7fRAmc
aQvyFQgVdirYgBEZTeFIJY/uVfom0Rdb5Hp9OB3jYMKYek0m87v0PzdbU4UiQ5YbH7f+ov6to94k
wcSR+eWcfFDpe8bapllJWzFOtZWMw6CoHnEQTMHTBskO9F6pfSSPNLxe3HFG1gIZ8FB7n0NPbmYO
j1yHW1hvCs4cr76o6P5BqGkXOjadzX8sXVjIX0pBloY+guuAeLltLZfcEXES8a7IHwXHSHCmqUDn
nOBYfuBBrc8Oq4N3X7gt1QicqCyW95Pf0cLuq26kBsrTb9Qe1IE0PbS0qxfuzP4zqdeteaKeZbSp
kREUenSrB7GVr70Wt2iPvHYU7A7sdVUbXsCmqDTzqUmOGuWpVe7wEKdLdJnABZ+Cqpsx9MfSt+kO
3uFugXvoNgOBzn/wj7/Aw+/xQx0IKqMK4j6x3tjhiaWvoctEtvIDTbEr/ISmdHNbU/BXCRxDlCj7
lkIsxdP4m8ot05XKjm23vnwRJsHTtJJX+g7sQ+vpR6NEqB8KOgVAYo/iIcpymzjtQjgHLLebBqWc
oXVRaPXIPJCRx7MMOthQQUuPKtJ4aoPozqVQkqrIiqDwgo3rV5oTFjKOS8osSoDvhw0AxrhR6Ss9
m2V2HjkQ1/yXkmnFSuoo4WTYFyoDOgW1aXQsHik/xNPqB4QsFCbXYoa2es4MDv68x1pK6uW7nbvB
BnJ1yzkVwBVNFxK24D7pWskzr/F6VwNfxra/It8P29w319JIpig5vzupzoM6WqfFuarXHZgOHs4L
D7ZTRVe0KRS2s4SxnYKLq18DCBiEK2EB+O02k6sRgYt0Sm7vpN1CfO+XfOXz38RSmBNs7HvmbXOn
kkUpJ9v9OMQHxgma11YnjtxaVWw+yE85rv98fCa6Ps2mm1Ymwcm2X/I3gmjKonYD9TOR+QdXRTOZ
PXN1RdYPUz686dAahzZciU13bFskLhrltpmOPWjMFS9+qAtevFsb9ylGOJQQ7xCg9owV+xHsm9jy
AC4UitUkg9ylDZMNDftRA6h6s49FfAsKU4YZUKq4Pg9tEThFEVBLnviVtMNvdlIX63SUOE7n/ciQ
PfujDenuQ1S0z2hoB6ESQOcfODocpXnQyxpgFtDaTpc7OHZWdCP4kaRyCFru2rTRwk380kREhzLr
bdrnh7zZEGU1gOMyp/vWYW8VPp0ws+HnzkChJynRUf397DJ7y7gMFTuPyJFRpzCEkG9M1Ci7N1uz
6w48Rz2YpGxsRrdDrgfeO2P3RXqRt/xqezFqgrrAcZriTQctUzKg69bhuAyNm0MYZUxIJGYoGsJl
k4cjEnqDSyYZnNv1W6AIVmCfQiVbkt+iLgm+mLd8SNvNDAqJM6hYGZtQ6uLJFIGXJWi7RG9vTLn0
bvmaL1ih8wdMHKZA5FR2ypfLRH/xwEmTZSh3IObQ2vcjao1Uqp5zyLoobced/COBSS5Vs9JVpHbm
08fHW/CS+6CPYG1I/bAXwT82oY/H7Ga7VBqN7b5Lochwe4RtsL/GAFlblPBGpIGoawy4Hfa0MCY9
pO/Z3sqdrbDyMS/T/VRqbnK+ch3mvGGdqIPOROdgX4UlzmlVWMQgIx2eZvuNryDe1vaWwGeKhU2c
IJ5lwU9el5sNgw05m5Le4pUSClW18iS5eMsBURcQOOGQ+1/+hpYcKniL921S807TQ5sh/E49Mwrh
dj1jJPEZf6YKHlQvfLSxKpIguuXGQ+UR8BhsUyfTliTEaMBnBYobuooUeCSrQEGb+MjaNxrT6rA5
ror/7ILVegPABRTYjnm02w7/jsq4fbax7GfMIXNR37o/lOqAJGALGBrtA+8rnNqat4ysn3t/sWXj
FaR6X+rDegcKG1V0Ee3xT5na2KfZAMMXcpe5XKNHUFvb1RKDsW7bW6brhOAAB4QuBSBr7dD3OG7X
Lk2spIod+P3yusjQdz718+41JLebgnD+4Vgoevg2uE0aAPTXInl4LhflT2WZ+MImoTs/rgi5+ZHF
kdy1k6DSX4fEjNRZ1z9NpeWmfzN7L+OY/pD9daXcCkIPScllAWTo5/D+3O3UHcVTVmeVSQTaoX50
5EBKfabXtjZHYy2/SDAOkz4SOZYwZDr76Fy7RLHL1Kr/TgDLCkSnxiU7R1gClO1xnarnclxVImRS
qLoLjFjNzlRJ2Qx6/smj9wT8VdPZ2NtLOPSbVvNuRnuInBA2UDP7z0Hf8yO0HohZW4HUOlQRjfSc
JEWSmriels0QBX53wE4ciw34fPbMTs9Y9Pr2WCwbxB3iGlAHtiglnPe5Qku8gFOjAIlFcG4RrVOK
m78MqKm7ejYcIujUKkkRNKxDEQe4T4Mgnu0N1JYQIP8YoYBjKzmRLz4BFHuBPvcOb6ZdqMFrnDYa
yqdVpmXmIGAQx8tWKCZrsF7AiY2VG1nnGYk5Hp8A2gJpo/d6vhO4x7revkVJjlzcsAA+BErawbih
80lWA8npWWquNtHITEm+JZiE0awtzRi3RzSr6O9cI0WcEA1E6F8qtgJ1Qp0szxzQVnet3Rh0WX0Q
FJoxevpoHJBzRf+QhMFjAJSYGksTAynVsf5RECruld4vXJb61i2toBlkMjD4cRAq5vt26OLulbXq
adF7jdkGnbhTSSSoyCPCiABEPJOElmqxasZAsiJffYTtSBbfohzDW3tevFT3PMmuickDeSKIrry2
h6uO3gzu5Vj2Oy+0uGSPb1j9Ew92VJnAfPvAVblFgHDn1JQgu/Ji4a1yMucQNL4Ve+V01Q5j7dp7
zQsXd9B9jPcB7lHstOnN0ZxvIVluKIVSVMKes2RLjA9GyDR7xu8pmbbso6D+Jb9Qm1M+LhdPQYOR
BLILE/ERBt6R11wWB3OC94ashbYHaFXy/toYQiYL5wIHOA3kDue8vMTwfIV94JJVOdnUYcPR7/dx
XL7EI6YJLjUiWfhwDXQclZoPKEcY6ITbV8JySUGU8ngOl+NHs+wQ0/ParMDTR/PpazPBZOJYfokY
9A/Pe2Il2oBk4ZOM4aE/6Hel/CFMZLHKigT899jPdM7vN6OmPx5sfxJUEjH4bDmlkXi9WMoP7Chi
7YXR1n5sigJb0nl5FoLlSeWKBJSm1q7bA72zE5wSty7qij3/I8EjmhK0qLX4soSfibpMXN8Bc77j
Pxafv5I8WjOliFYAHM0SOmTt4ra4HmYTColAz9+gQygG268mfhealvOe59Kf1X+6z8NX4IhFkN2E
oskdQhgTHwJgCNgKjuXFJlnqC6n+sxGPv3Wjx4XO4KmsCNoYmbSJ5c67+hH2d1eDRJTUR/qyGqV2
Ta4Ip9opf0XWnGNLggrTXAY0KJZp0m4HJdq5VYOV+X1E+hbPbn+NxUsUzHn56x47ExEoEViU4wo0
GU7Qu4ATVZuYagEOxRnDIFlEThlDpMdiNttziNZKp02uKOrsQvIK7GDl9sYUn7fGno0+8/pu6Xq5
YcRkPLyNHFywgPU/JTs4Tl8cXwHjbtv8fyUW0TZ6gP6VZEenvevaUGsvLbMcYutQ/FQKKxpEDvkO
PH8SGKNObwtmTd8yspgq08mQki2H+4YgRippWOmI7/RV4xhYuZh6kPv7FyfmFp1XT/hgSrIQByrq
auyQSN36hHk/SScUezaa2FVT7GWLq3VgR4PcLAXVNse1ICBf1nC41PBafVgwuNvdoB2bt5uNL8In
E3NQto/88qmZGXwHBloBherTEbceYfm2+dKkjyRpDQWazF/tmZggpGwPb8I4FVlzmNhqDEhb/NwQ
fBK2sF0GNtNPqCJzFzi0EFSnExXxArQmwev3S+aXL2rlM6VrivVhl0v9fYOFGr4ht6nscFrBdRmF
7Vmv2mfpoYRhxfdqGrEbcE+Gfr5vFW/eH98SUTAfockQ2f+eFG5ruGmxVzZ22YSRwiDPkXxcMuRM
ZisYUv1aXt9m0BQ3aRSyxDd/I2s/bE/tD4p8XF64xkIGtgN4YWXJK2xeu1Q14uuFknlcUm+hlIAt
ZEju63RCvTZ5evqOZ34lD6tGw9uxX3JdNZV78TUZGxWaky3Mb6H/uFoD5C/lh5e0L9Qj6xJr3cQ6
zYoM2sZm2iBhTcIie0Lmk/gn7Y+VrJjOagVpOuV66eXq7/LH2amKifDVT9yIzaU8NaNPLJtfizeQ
0zxDZyfojjlvi1puHR9IBFg8O//HCuw2YMEPPi4GKBlUWEVT57UlbA+R74OY13BfgEU6aE+A5nS0
T2r6I0Evw0KNaLhT+361/2o7cW4NegVqYnEIvIaoUThvBzStC1l9bGLPYS65Lpx4BO8mTc5jRv0Z
MKRAdVpyF4d0aMFd+JeuTV7onbzmA5T1l4DKcrBJMvyvdjb5gtJ1bTvRJKia8U0qMixndZvm0K0K
CR3XPt9hztQ3VeicEnEEZfg0JmMAYQiYaEmZSEvs+05NayGFoiCe/IfERDkEO7YjjNl1JA0HR5ab
6NPMVh++8o04dO0+nawm8hvnQAQGZOAKJoUw6+oBUsNVqDIieQDSgY7q5CtWpG55/LXdeLdm96o9
9b/Oi9eJnkI8AwvL7yfgHvkXi12Pd1DEBBG+4LjtxLPhuDhwISZzH56PD5OQ1hwRO/l6mbwlCRi7
+hZtBB8Sse1NJYn0orFITSBBhDR9DotbXSq+gBSdOYajm4tQijCu3dG5JP10go6UvYLwDUIySxwv
e8RQ18b8HE+ozIlvGykPce3Gj1iGVWJgfQBwm71SAodBy5j/k54sGjOZcz7zmlWphpKB6wqkB9l2
zI98v8/KUX8f0bYqWZNwJCO3uac106muTivjVyn9ICGu2plVUamlmwiIWLWx0BahS39/JNHIrW8I
Cb3MGWZy+p6AmCB39rfPO+K0uZyiZ5omEorsdi5/2CpAFZcb3+IbOtuc3FsqPpc3FJ7SMRANrMo3
Zh8kRFrmNWM9u+YBKNzHQo3m2S6CpRl26YAvyYXiUCuVcqlSX4Y66K3MEOciHQEP8KGzIDxax8Vl
NLUNge2HO/5peGOIEFI2qJXCoAp7Mz8pSoX+wrlAeWF3b5aE7MV+dCrnuYYaqNdY3pRBRBaO/zgF
laS1PiOvDwInU8mnDb2BudyWy+90TIB6xw4zWF9Zo1Nqzk63JdQlJgdHmLpcywvM2nULlG1z4UaP
6As8lORZNora8wy21Kj74SD67eLXGfZMn5sy/AZFJ/BixRVccBwoDoxKtcoXHrJNfT3tqUuIwTAT
C8zCt82h8XOkqpgqVPYRhmwUq2qjhP7ln1OfRk2uN79lG8p2HlOHADTqIJBq4L9NMDyhn04ymKAv
gUYsK5FkGQ5oIk84Bs4TlTltGOOQQ8thxQkFuN0kGkjt/s9ZBq3Rj+eXTvVFEUw6bkUkxwUP+E+2
gy5i3DK+/aZT5LMXlggRjo6rnwKWtx1uFhuwGZr1hLqox3dL/BBm2doDGYeNDDlfsJdhOIA/85Zw
k8xiUQ7qgBvRDnDrkbWnLqAU1t3ZnFluNnfzzlbZE9r3FfzewNVyOVaEOwtOW/jc70DkMllGbOX2
161rt1zms4YAgTiOVdsruTIufvuo4JLJfczKFgeJlAfNp3fQfFsVqF1DT0HaAQLcHqiYrbui6VLV
85YpHmParyNPKYapWhvbrZChYQzKgnUDYl2LjsmV7VJWfzPusCiOUMTBZ9FLpeFtjx+uM0kQCeyB
Yt6CiQx4KF6f2iJ3hCDDGkxCtW28YqzXi+LQBQINRQ3a9XjOoJZ4ARGH7XrKGphBZHUruboP5LrF
CsJYISvl2JBg2zlSDv7Tdg0yMxl+4aIhXnwdCqXJaTcytftuGmVcXTSyrr+gZS6W09Z/FAROD4Xl
gHGBa86cidIUtWkDeSjO7QISR20lMpz1sYsrnpGJFNKQjWKytqxgk4oh+IT57GDZXtt/bZ7RmHt+
5HrANcMqpWqL23SpLPPxm7Eig13F8NenCmtwxKzvgMcipyptxolbvXvAzNVxX86tcscbRTmM7Ei6
iV6ZOP3B12MSBpg2DFNxFldy9nEFTx8CA5bsqAv4xcViU6j+7B2kgpjNs9pWFLv9lP0mKgEckVRr
O/QRkLKEwFui5ufnvSk5sdGfMDog8q1Dho20Y/tDHjBl/k3GRaXsk1Jpr2PL3xNcjjX/Pf1vtSRS
YcLSvq4W5S58m4ktCVr86lGJiyvLhsTwJDlQiPXC/SaG3tgdIeIMVcpFxYHPnpjEn04D/AVwx8Rz
RDnDpw82EGm38DTUHK6X2pZ6hqgeNKRzT0f5kXNCAaqx9Ts1vALzQZAeZH30QOfTbCN+LJYihhEa
TBSr7CR/U7gRDuaF+Mxrf0frKh4N7V1//oZjVefaJgXijnWpFCiJmhefGrb8CB1lIfUJ3YuXIfR2
IjUhEA4MCIWW4xolR0Sj8Tn4dPhVe5o8k85esGS0/wzwYtxncWVuq1pivpBVxL4axSWsBpk49ZQc
TA3gQ/Ug7127fKXph5p99aHaNaNhQSCyTUS9cq3R+lsejfMNy3fsadHAXvH0opASmmRQ0qsgBM6t
ZubsT3QxVriXNM876icVxkSWcd3j81FGOUaa83p6PpUO92dhqhvtX8n2kE2QsEcDIH9L+XMHRePT
TmqgslbGY1cXfx3Q5UuQvNjM3o1+Vfd47FTzWaJOpzlmS9aOmviGtqwwvVd5YgEF/cWAjEPse02J
QbSwykaUcZeXXlUuZ5dcziLym7PAsrHeU6IvkRcKY1HkK/CJN6SyjbnpzbARXOJgkH5+eONCMMhJ
aOgpM+13da7ugxOw/xVjl+m58spBnoFULSRiQ1ae0gy8iPLAQLm81L/iCUGxBZv3g5aXki4KiQKg
hNf9I+hs9VmDJk6Jr/N+cFo6RxRsEoeAqCEXn6wEbhjUF+dDNIAayjDlEip3AFNzsqwQfDn6Lu/P
7WUniUDzMce4+/XVm/Dkvk6oYerxHExyI9zaWHzXSJDLivkdZe4vqCAbixrPDsOEIhU2aF861pnQ
NiB6c/oRPjnG/rY/fwMhpSchiQaQznF00b44Yd6/aZ2sCYjIbI4EsJmH3HmEl8zaJ0fKVrodTXax
lzc6R+uvPbSS2Q88ucCQQxlN6JUzZkviBhgu5apa/agVJo5skZ5ponDtxAF4CXsTfacppm0puTlS
TCoLUnfIBY/g8SLQRyIedbC5gfvSwfQobZh6kmYLH8tov4EQFqQE9FryzfO6cnBkWpqStidWv7r6
BPvor4ybtEtkerGZ3fnefLakOoCt8Qwh1wVho9BpTK5ZDHoA/vX+PzWKuyyFQH+ru+oDju9zkHx1
pDNQAT57DDXfqXDj8c2zBUL1nIkEYRGvS1be4qnlTHv1PQV0ec68FVN++PAjEb1SBp7OIV1aut+i
q8pMHKVDySZePql1KTD725WSS4QlZ9salxDmO3z7x5C7kl53+cjW4vCXVJ0uenJgBbfpFBg8H9y/
G5oynmIECDkmjg7w7x872yxWy+s0rRRE2McogTgSPxIZefPLhO42g/x0TnTL8of1+fH1RjfnsK71
mH2+aDU/mseJCvS5I5trDWK+jgGycWbYX2slnBgF9Dne+aTM1H6Rr6as3wQ0u2eyi8vjoS54xwod
Fui9p92RJMnjbt4jBZCv85loAZ+LVb3vWhYq8/6a6jhvezewRimbDBMQ4/sj4sq0ENTemlja2+G8
hCtBMmdM2xmsI6XmYVTZ/yIeTSrZT3Lv8g0zsQn50Gapp9NAX23RpyO9RNXRy4yVmEjwQZz3fu3s
LDslLAg4o5M1t6EkVtjauMJ9CQ9BJmFvVz4KNew5KhPB+oxI3TEjVxSTOYLcW5gx5RwB4N/6l5Qg
ZhOvBJoGQ68Qm0U9zYywxGh5fwHE4AppEnCGqkJphz/jSsLBGBh41Gsg5nB68ONBQaYKNtFshUbc
BP97y/1uyK+cBTuRdTZHpwI6SnOO9zFzIXsHIEYY5/qTbcGndvW+hPkvmOxUMKL97QEYBRdYgOe7
UJDrHqJbzy8izXzoOEofMoK+sYxiwALRfN09hGrc5MECAjoLDuYT2WQybGtokNgs0k166PK/lY0u
F6MOiiEGCZ2fRTSLQZ0K4S2AvkK1df5Jy5o2FCV0YGecfTuEQRfErBRpk+k2jF8srvgvxKGJYCbM
Mo9QqNNlD8aifjl5uT5u/nCDF9cFAeSz5HDUH0I+KxFsmF6/fJ1GX5jHcgbyOvpK4FUP1ZBgLf6g
b3tyw0ILXz6xhL1giKdB83ofj7cLU4wzhudumsDlrSokKXI0IRBa9HtwbT8MAJ9z4nNawDp4dIty
Rrc6/anyO9oO1sKibVZCr0bbXpTHulArHh9xHaU/ZgYtWiD6JcdehB+W5DHwWfV7iuqhwJVa1P68
xwNjc64wM3yXP+neLdkGe71eAJjumVZWm5V7BuGA86ZhDLiFTp7+RV0qhz90OrMfjuLkNfCa2S1g
PXk9FTKS/YrTnM0IPW8wQ/sh98NIum6PVCypUX5BLXsye8Qx/0iz8uEK9QT5cPurWcopKpaVkCuK
W3faLNNJWy2B0QoYxwyGCP7KLGGRlwgsn6aU/fCq41cIpqcWRwSZhYsH47KNwKixafu4CG2tngmZ
gznoloZdAS0/0HvXqx+yIam2IateKX46vfb/5U3nHm1LJQ1heUVPq+fjsEj1hzg/5u4FAzsYj36j
F6r/vuoAp9BKlQIv9c+8JJu8CSF1630IBkknQPzcX1SBJo/VnKid1OZ4prB/oyIM73uZeL5KE1ms
LQHTfJ3sQo/f8s7MuH+WVl31h5n24VwfqURoe79fkF/rtjp7lQUf4DREpdqWfqM78UuYC8Hclavw
F0mRO51MsMB1QdHBh+wfE7kIj9KueHIaLZlOds1SLCqDzr6TPiIiYUYzFoaTcSjMAeIxw/IzA+55
DPLUBKA+fTiF0SH85UHjzVnmeDgct6eQjJ2ZCY3hrLvI5UI+w0txxrcce6uMOp/HR4lQX5xIDYrR
oYT4meX9dhEW5o8D9XfM7fXDrMdvnuV0kYiuLeRxkYcQ7olVc5bZMVHj4VhdkJU5HQQtOfOHHkVh
7MBFCfkTbu8s3FGuAvzHhcTcXR/fW6lCg2kJ5BD1rqOxyuo7Z/XrMS4Lpt38euRvbFKe5KlE9PLT
nbNloYhH6QAEG8Tbsr8QkbvjpB5EitE7LaM3NGur/IIZ55A/7lSVaTxjQH5FMsTcY8vRlThlnP87
DSNlM9kmUrBzXMW1tpK8dBt8U6ESCF1zUlQpUDPEzvAbfvBo+tMQoDCc/qAQUsk8VkVCq435duxG
/zLTAywiwQIdzkneNlxpYjM98vIj5CEc7TLKlZRB0yrBrg16A71l6OSP2fiBChHIyLndHFQW+K3J
lS0Jw4Fiv1tFkaSXV3lyPubCgP1VSVF7oW0iyBOULEwg1ZNLCJH44hRvyvvRZUwXEaZhAj2fBwfM
2aZJNDBld4HSiYXVkv4sC5tFPRcYAJmJsZWkxPKkPQCQU16tGHYfgI2gyVV67jVdBaM31X4dwq8j
bZKBRj2bSv5QkrEZLPZzrOtmgpPgyhjhKe5GcyphCafciXEnC4VPqf8hg+q8HpYz5JrYKGdWzSGv
8XuLfmJcwEB+XFjxWlxauFq1B/tuh+hvb3kEENon0gplOJcQpvKDUDXnPvU8/+UvexdpdjxDpacn
2LlTOhdUAsdFuwArVcbxj3H/opQeGtXP5o/5Qng0nB/aXbhETTXGizu7HybQDBIfSbgQq4hZ3h48
R8DuBYQXRNoIssPoOOr2gZXoDci7zgAoed5vOHXpYLFM0NZ1M3hzCXNXuFpsitDer9wapOpHZi4v
7YxVgag+UggJeRf+e7Wjktz/pXyexBfuYhpBKfvKMNEOBhc9q7DpwGmPDBboc3MaWKQDzspHuSMI
tj+NocKOu4NaxvDCiN//9W/e8ehC1/VxKlm2C5tE3Mx6rFWXJtimaPoVN7XpPOnRWJOQ5m8l+voP
wiDZtN0sv8r2XdPXZ+FZ2hFaZJFe/tFjWJF8GF581A2l5SPvdvEesFwjPQzGHfjt81Aq/qGHv5qk
rrvehk70xhRjJbzwkJTpP/z8KwGUnyBfHEjWKxcCMe5UOT+y06SyuGALLeERCElPeclSPh5jD2fS
oRLnGIlIxHH8RXVlYR596CbE8Z2VddJ5ozUfFLyvXRddLd9oQ1mr4CdWuEIkL6SgM8GAqm0hpHQ0
Dkdd6kFztVevneLcLiB/Q5akEnOSR6x0/GlWEY04/uZclXtHNTGQfrq9+4wMKbKBkNm+gxzJy8A6
MsM1mCXFTyasTrFLkhQ6GFuoC7zjyjKj0BzEaQMgIFt+cC1mDR/DhO06qgabr1zxplrBtVS+WKFA
4fLjSp1u8TQbe3UzzW9egS6kA/M7f6pdn0HH++QWCzNAW7vuWOOX8Ae+6SU/UNJAs0AIhZ5KBr7X
nomDsY0Y8/gm2ItyvFRvZCchQV2l6CrTs0YMh/evdxqLkanB26WhFqKfeuDH5XdVCIC0uCPJQlG4
Rmd7BwXumBwggW+gnCG8Uwb9D/TEwE9IlfA4oNZXvWtkb48DHDIRdlRcZkg87HDiLr281OTauwef
EZxpn3KK0oAj5kx+oCRqzKjzHIySRNILJi/xHDWu9NSo4m4D2Beb1CGoPsF5g9qX/j476Ru6zbFO
Vf8r7DuDOv8aWts9DRU3WwmHJtAfM5MWfVziOnplKGWm1TiWXUW8dAoAlK0A7jHOKCW8aGRW3sTv
lHxE6fHd+h9+WypbxKLs/kcZ7pO3w1qalyhIk+WNoaNGPjOcsuxTziXXd5qfW0u4w7Me9WxRU0pL
EaYHkVYvNK+fW7YvcJoZ/fZf6PKJC8efM3cCsyz/66r7ruHTJlPN28ylJE4EFQcHR1n3/bbeSMeA
ZAP1fdbovpokJq97tMcfeuDPwqtDgbF06ziy6vDV6j5PBINKCmLlm19v6b/Dglj2zxLw/vPbbn9v
uCvuzHXOVMLx6Fr6lawndEB9NwT0uYDhF4sNbO7LEw8W4E9yrsrvMcFwavHndn+oqVJcmYG86fNw
DKrkq/SOngEOrDfLEQxi8XWHaDpKh5fWFudOHyrvIKP8LEVi+eXN1mK5hNkeL90+wPcMXRpcSUvU
lxjKj4YogbH9+wAJ3lkXVzKQbLc2ndI3PsIZ7Ibpa7603B8VtrlCitwK8XBMTKrppxGImuFjfG0n
5pFM0aIFj34nsO+oB71/sBMngwvRxml+SYtdPxS5lK2s3FSa4vUgmoqyePIFGtRiBp5FKwPgl6hG
20Pl4YVREUiV3HHxvfg+/Dkf1vzdSrvX9qg6QIHcuUkVVC2F3gUASDXhsyrEyn+Dt5SiiesiCZvQ
0wJrC/18GDP1H5YzembjeFUUjKw+ayj+7RF9GjP9EwtNsTAjNe8Q6tRsD0FKUFNZhOv/0Ea5DwBF
BPcMXCFUOurESrhMgFOuowm9ou/Yo2WBtcuVnGOjgoFsruZyMkVniqH3g/NDBJtVdOUGA/ua3n9G
qjcJ1vkYxMgh07JkPcsWtAOs4sdtFufhMmFAfWklF+NfeTjK/u97RomTHPv1WhJfAjbOAZY9EIfG
BzuMZUs8Aguiue49KKvLBwQ5HMUqv8P+diThJlH3xGtIcshAtqGsk6fW3sb0o4po1gFDoNILD3DI
ffkfMa5F/Dw+uMg0b3g3FlROWiPCsFIoGBKPswq+JYYzvH21k6eYuMtcYYKLxuE4lFT/XcgL+VnF
WeCzCJG5+SnDjz42q6e0Sfrdti1nhcgfnuCqR81CMkC2mMznFO+i51v1y9cXYb6tstQMaZRhlc4j
LZVIDeGdtai6miTFQRq1frSJhko+6skcoi2Mk69xKXtAow2xHRRdqZpfXM9A2Hmufn8V9AE4Il/r
+pjCsPNPBAgjUkUG5+9CMyX08bVp/PnrDPGUYwPrFVR7/2INavls1MRfLWk2t2HqaVdDQBur8z7w
8qKmkNmjN3EaPqnjCeQo9KjnExmd8bGYJxhABHnC6JoBRmysri+XTRKwmHVyUP4QUpvSzf32ephR
0VbwibGw3NmsJIl0i/KdqZyvvfr+eAsLJWfpsapgUFHONAzhlt6ECOnjQXtObYE2rF+iTA7i4OhI
1MHdFVYGHFWfAedK7Dd6usomNss5e2LWj6Yz5VMzZ31Z/+KHaj2BMcv5+cWr/GEFvd2t7+lUur4W
dsKPUjdURHcGvXzoSPfOSK0f4nCja6e5Yhuftlm9ydLzGUByCP3hckQpBXfNot5yHdyNuXfJSS+q
fjUoAhwooeeJUOFetD2lPUTR6YfDVV507EJCVpiNFGqUSPMJESGW7e4pj2xPCbXUgPBumB94ZWNN
BuB+ibOeMtJ0WCJS4+9JdzcwyaMR9Y7l2hJEkpaKYU9uQl1FIgCHLqJK9S3XaxArd5guK1oOVW2M
n+uM7iWHteQGAdOYTUGh2OyFKvNS/EN5SXfo1jOIelM0w5aVi21WRI7uCkWiS/NF83S1IhnaK7aR
7mpax5woj9LUPFUdOj5qW7hzVuwJaba0rSN1F58bChdenE8zCAgoD44mAo0rPmGjhf4QpTBQrgqn
IV/1DrojBN8gAlaZe2TdMbiXEWob06zJblAhIBuCoXzCCS47uY96KZjUCbLRcrmUC3DyiAEDl95k
4wr9cThMqv2KpE1AFVjXPuvoyu0jU4CDAz8bQnRVGYqzqcAxPHNdNwREDIltudAMLd1eF5BjeheN
45IMCtZn2Y74aynvPbfD3N5YsynwcmobZXswTNZ1/fl+b0v10CSxigaNdy+4FLCe1v4cys+2Iia0
KibdaQsHrzStTYqoSPgPj6RuU8aXgptz1o+yIXGy0ansthw3iu3G3DDcfTD3KgC9+pUW/zBiO7+E
Go4lE/UdkQO+RfZboLiROLiQZ1hAZYvgR6z0T5PyFJT/x1A2tIaZYDYwh8vneDOu9pUz/01AXU+j
3hlO6vOCOKUsRzCrrvdS68bS1tSntMySb31tKUZAlQ26swbV7XnUClH3dXmQAo2f7ZNJ+jtkGN/G
hlxfb8prQbV87Zka0OuJbtdX4yJiOV3nkh0Ldy42rGDuiXNzlQ7rxjhKbu81fp4CQ1EC4Vz214sp
im2TSfFVMRVDJjmE40LMK2MeNAluMTIIGWFX/Qyl1roviyB9PpewwPlmcgpJIclThY9KluQTZNzT
Hb1oh8CFMlt3+V0L2Xi0JrbxP4eydPEXUNRwUGvHz7PrVL6hwUvrYXj+zMpDxwkBpNR6btHZdyrw
Gxn2czWx5LHe6UHV+S43267rkvLKs9vB9sZgOZ0LOApEoO6cOlSov7m9V+Q+ZrH1NDoZ2cRFLOQU
ujA9Tk+klrT9T+yOcN/HGOpAzooL+uE/NnmV8w4HV87MMxuNzCoCI9DLmu7rcE+d2zMQEUHx4RDO
6kaoHuA4IDuvzTJQWn0O999vNAwLtuwS5F0+KPlOKdMM7QPdhLpRGY/Ysl2QhLjd//vYgkMSrcG2
hKQL3fzpuFce4vE8gytdcyS/71kGYXZQJhh3mWPn4ZLJAzghpZV5ytz553D/M0j/3qq+NBawP+T2
QuxSjb2qCemZXSg+t4tHhTLgpNv9+MrgVGgFYIXh91GPqQmghQay//9p4P/uxypBojOOSJZR5S3D
2bqL7NZwCMH6eYtgUPw/n1Ss/5R/w5UrmoQhvBuxrWk8Z3D0I7KNfEdA4/T+RHg+w8gwFTeu+wjH
fo6rK+DdSBNfVaJOk6MmQuPWpiiyLFcLUS1HQMmhWQWiBixOax3rG3FOWtpuFoZSnRH4ehg+/j7k
jmVzy61ILYpvC2OUWFsoxigvSXe0OSWGXOLPKvvrfpL1/qGZp4YyvaYMX4ERLWQkU8HvZVNV0kFF
VEinU56Xq7Jke45hAaBqB4idN34HEFoOW5ZlTRQ7kChSu0PdGjFSKOmcRRHWQb43lew5U1IOhzKQ
WWPgglH0kGRLabybyRdf4a2BlHpKUrJHRs3MAKiw0YEgA6JfXRHZrDP18apcCYGnZ/GXdn8q/Q6c
5HkfKhJF4ThwU7/qN5labFckvn8bDZl/6o2T6PKINdWo6DMsEdbC2WMGDYzhoIZqkPgSjg9nTLoO
UppZoq+7se5JRkSEl8Ky4J135Vk2WS2R2SiijdrheCaKk70GEcP7tXswaU31Hx6OIuJZjtgZbQlf
iNCdy1c90ri0amm9/rbSXDERmNmDbPRlKjIITgpSgmRNaKTTMjmHQRz6PPBeA6xRefSqBvi2mpy3
qJHJzISZZS7YxdkEeYFWt+DAOhW1igqq/EZPTZZ/+eOodahtfKdvCEtUrecWGCM7QFPygszcpoxE
Ahlhxe5pGnFYH0r1h6nEL4EpE8XWKhFVOATjoQ8vztdpy9ss/+/t1mHvMF9rqo+Z4CPJZtAkdNwx
2r9NX6IHUUNMeaDHdsfZm8uQDCyW7uyGJxNVZwjPhjWH5psz+tPmTFbBSDY8gAJrRhkB70iqoTx4
0OE2G9HJeHwahLavTBZWGPdEq1LhzXbms0X1Ayx9SEsnuoaULqcByYASYUg+h39oVvnICgf/hK8K
la6l+IysS2BPpnkElIQ5mjMCJkz8jDHN6zEq93u7ijqahTxbBsQQgbqu0otveXq4GoZuxyRWBs9y
ZffiYW7pKS+LyOpINRtTnKQ0qeQXKmTOKEZEt9TK3d5d8LmyLpda4B/IwmJ5OLdNvydmlvL+M200
RYS8t/5/TcIcBug3Bjz4x5jvACVpfZADnyzt/yZyS312a22CQr2+D59N2OCWwiieWepoWLcpBkMx
r/otkJPyIUnvjMDOF6PiZ+OhMneZd4AivrPvFHvdlt9S/MycrV1hgGdFIVVuP+UYnXFrYdghT60v
0vM4q8GhuObjS7m+hQLj5L/dXNyVrr9vKJMeYugHXybwVil6VEtXYzfV6vtQdtZ/SEkd8hrW1Fzz
8GoRy/Lmp32uDl29Tb89Vy0AMM0qOjeDg9H+632Io+UDqHB0PvI86KtqJMjlig11Q4PrvIN75RcP
63ouBjAZoy7A6FM6zhToAPKNxaj3v3KK0XNEsqvRhyhcn4dO3bisOfudTyd0wb8VhFWp8a+Y2cTr
MBSqPumr/W9moYdC3wIuihwdYwBTeeTclNM2uD9+4lfc1mvKpXuZGpy6/0AV9Wc4D7g4yFOPcmmU
sqqwmBgRQby3ONVGgBfaIVvve9D2huVX+RwpUkmcbM+bTUcQs5l84mvm2ky+4IWySN8tUaGlRtZO
yQqkUICshOWjz6OZRABcCbvBke4QGekPZzvOPHMpJakkxhXghIZs/xwm/JTCq8OM33cUiA9jbQaX
Vj9ri/+jz+t8aLs0OazWifrgGpGPXL8ASdgC9ECUd23bF0GgnZCdNDB1jvcRYwgAwRpYck6rCQve
TWnSoz9NLW/V5j+84wOOZHHfL4MoW88+1rbUt1ni09ScuxM8fhE1QalamyWHqGzprRzMPuXcuFiw
aU9eHHEUtjCoLKdJI3SZ1HDJiLZA5cNNkwlthLoUIvhZOUxTUcNXogzDXjndpbV21bIR9BVvXtHV
ZA9JHfIJ3RMotB9wQAO+tsIXxnp67HzKMHRdU0Yb6Y1iWEevCC6j5+N0znYMD8dh4XKqKjGzaEPW
/mGfof/5/UXkfhkFG33WtoZhhpTMp/TqnfYvbnu+1TufVBadwEXA/BFIR40JBw+t34oxeFREiPU2
5ttwcw6Fr+Wo2R0pu4DUG/5lBSbo2OuMZkH2Aiv3UycgbXarOhJSSmXC6cBkJPXTg/BbdY90H9yH
tpJZHyn14A+uNmorSjRlXdAlUIvpM88LcU0rkRsw2grx0PFULrXNBTSZ7or6HGWctt2y0Lq3Ky63
M+ULnblj14N3YUtXPzsmFL07F+bj9qGrMjtyEt2Ny+/D6uc3cnHxhx2DuW/vcbMzJo6rSP3CDrxQ
0W08rGpPhZmJeyqHgGcTSdvCFY4bTQrUuy4GpY8JUSYYelybiuZ51PeK6C6s2bF27OxeOtkgYvfP
JVWgmB1/lMSFxOPfZAB/4wFj/5liZ6LMqPKBq97e2GGJ8EmqjSvBquZeZYDMWwJ9A7aTadVcWPPX
lKMlF9SZX027pQYfSKGwAvwGXra/bjMsFkiRxrZF30ou2oo+TJSdtwYnnakutobbDAEFq3mHQXbm
H2dWOdyDV59y6iJSnyQmuxcJaDorex8CA6J5yEjaIiL1Z6JoCLYSxoUAO8pzwVSdOaDcxLKvpjVy
CAIEjJh6fHyLzwwyAmCC6z1DSRdwA7pd1MdRrAc/0IKi99GAoy2lfG79GRV3iFJmjzbRJPh03PZA
o6pBe6PBBmhA7lD5C1XjeJSgE0KZJhmW0s99LLKjHyzBfZ2PoXwzKbdLjcikPcbV8OtRhKev3Eug
ZyW5cptwkuby56uWV4E/MxuQbNoOElyUd0eRYVD9V8snKy0J5jQnQl8jfI8/YXgr+HIQW9HB5mnt
a76LIMTDg6RZKzKjg4RucINKATs3ECb7vT7NIQ5M7h+98JjJ6aK+9JPxF82qZvVsrmMM/40IOmTN
T45h71P3i95gDibFFYL2UgPjeHczp1Z2LgfCvEHpRfTSD/4M71TcyYFBSzYVzUNY99GPF/2GdShO
H13TlFNXf4txX+66XPMC2bm8D/rkDK8Pu4TNz0poQzXPn+e3L8NW8vqcOip/gZlI6B6UQtd10Mat
1B4KwmIbV4trs6ipEQa3lP3uOCyZ/k/PBkVEcoi3I03WzWXHTnDZ8Q2mZ3v/eqjEAkYS6sVjVckk
L1AWhvMR1aLqqah6SyoxOjSnFtNmHmj6cT1YbuyXjFuRFZIeVi0fvgy4gljFm2n5KpyVRIXauIS+
5ShSKvXq/InNtIEs2/OqEunAUdSbTsAHCGrPwc+6I1e/n2MMqjS4yP6Z7tJFqvVFOWxzS/VyWj2p
TOBWz+AV08JULNYRVaqOkiQ2Xttmmh83qM3hzC2q8fobHga8Ub6i5v/q8rfRr2SHeQHoJsyxx3uG
SOtarkAR5/fhbmetwd5F5yK8Iunvcd5M3UWKyH9Xgq7xs7ICD/mHeXwXefzQvI6uxLurFtykBnZR
cD6sFzN42Pc3QQLrkY9A4KYH9GzB0+pNxYx6bVR0dD6vTaVC/c1di0LRkwzlvIsF+7tqfleRWpFW
pqUGIfiqjmb5D67AYEMQsPNLovDeNJ8s5G8jdQaQbnQBfehOAK4gE4qZQIZJHhgaLsQ8rXt+nWfc
/ERLM3F+AQD9IPFmCryzv30Gq5B9UIo3TjjjlnMTIiQhhrmF1xyBGQ8Er2AZt/n0GFf6Vtn8sjg0
oCDf9eeikS9tCmnn6GA+PFvvp4ltKW2mo0Tax5jqwLMn1T//OiWBYw71fnQ1gdyNsl+MEMP/AgBs
xncUdT1OyGhTYVCa52rboDRu0fDusQX7jiOIScVQEh/oMEXM2tmXjuExFSQbJzdoU9FlAI97WJnP
2/xX4OUMAzGSKgFUA6kv3j97ESSLBVa81SeO/obfnT3FlDwHCCFYv5YezHy+JFJP3RPRRKM5Umyh
wl9EScFotYTLs94Ku07F9xd79ZJlQIAg2vyLPCZnsCu94JSkp11yJdQyniQoMkD4QNf25IPMGyjF
5xf/F+AZWe8Wb24ISWCEsd5egy35AAuvIp1XP9DoaZZiP2c9uuvuUXq79bdIdskLi9vFmYwhUxcm
wYIgXZMd8VB/B5LD2PM/fFryt4zVZ6E8MggYSkRfdC2hdZUUKFeWMDoYGsuYQ1FQu07IbQGFy5D5
z42nRjq4wE11xRHeHRauysYH3lumGsg0yJibXXD0q/BK3j+ULg7yMmacU6BzilPs5kqYOpU9JnUC
5iGJcpACJw7JFlU2jSZcD7ov8fZ4ycXvv1QeVBs803pDR0tB2g/3P4++9CptRmehYHVM0+1QDUwG
J0jIUTQp45QWux0nf4Q7zWOV+dDNttbRznhFRuwF5V09Lg3CXJbjxw1tV5tsJ/+9yiuvBDCYG9sw
o7MlhGES7QsfB8+TJWw7OMk9Ws3l37Nr2VkoohSABCoJMlXSZJhxdI8bsteLoRvag8EPpW/hoLh0
L5YwwJC1lH24LEwgVnZJ0ZN8aTgeBINQnqxnDbM2juUV+LRVY9S0jPc9h9P+blPCm8fxpx09qMLH
HVmVX8G9Ou6Ay2mQiN7PzTcinu32NHX1iAe2FrJZVyoah4ppZ6aBsMU4JOcO5bw0ixE2Wqjz+bqM
b6ukc41NOwHQLT7/i4ADI5SF5Cw/3+FW/b4g8enl2Ftf87muEIuh5XQytWZ7RPcgubbC8mLxCBC+
iPvxh02j+IGmz+ESq6SA+m0aKSrK8FtHND5bUCicD3XW9ydFoa6QrCVcmpvWj7Vb5yV3Ldussha5
VHHnqBTcFd6f+XOaDs7mZRPNGswgEuyGpscc0XDa80vxWiwyHIB6YKcdHZs1MBaDxJ/tYlTniLpt
RvKa7ijL5QGk9C8cQbST/e+5kQHHRrr7ZQoZWYxsy+awAu3YIFBB9zsLOOcsCsPT5hxfRBzS+eNv
yqwShW9fMpF+I98+AQ1CsLI2jzxbyo5uWw41/z5S5MuQbrMMaOPkq4ZV1u5N7LqBlqvb4tu4JFU+
eW86kXzVqA388J+x9UZabl0w5azM3/lymm7FDw2KTC1WlNRoq01cAhX7o61mrIxbfOrCWI65C8j7
4OjtOmCi7rwOmseyPPtROM1V73pOf85A77TS3a/bPVk/4mJIBbIa6zdw2yL+jSyIIiwkLhkfsPhF
OQCbhvtY0p/GU/wWuXXapP0nH1650V1Wp8kIM5ToxRj4UAVMws+GlEbfXpxez9T72P/tsBkakqsM
5i48EDJc2NcxferhzJ4OI4LR/vwsPsxC2KgjO23/D7O6nyOYrfMGEROdaEbKtqRF3dHnkRGUuXeX
trRSU4obK4BNQp3+Be1QPH8LWLWeWAiCyBqUhMW91RDlohZNNB+ZNZH0ZPyRgTYBc3OveBo8cFJ1
VvFHPPmPpsXUi/RkOwbWMyPCV9X28JDuwPlp92LGMIReZ982VO35o+vr2fGBv0rK9EOZYZ53b+yY
vGxdWpYjyeiFFoBKSwG1ymX80cZ9YZFYfM6NtIiyA7CpKODBYFv8ia96TI1P3Nmzu54z7kaUGs/u
NyuZ6Yg3eK4O5qSv7YUANxo3hUOiHEV7J0cpG3amamiGZJbDTe8rB6BqkAiE95HtTYvl/SVg4lgo
rB2Qr7/mIRB1EXxQaQHUEbTujZzvvle+MwKlC++qggIGF6dActtg0u2ix2k55lbj2TeDaUxcQghx
EUerCaKRqNNFK2CpkP/c2s04UgzMYYWvI1sbw3XBRncfQxKMmq5ZxOKAS9BtPnLSD5KQleuZwPNg
+kkcxi5CvwalwTR10Zi12Rnl7kFk0YGRU4Wc6e4CibGm76bBfXF+/BFKQZrDwzjhBUk9nvuz5gSQ
yKmQbHycOM6YlcI4ku19/jFyGfqPzKxLNKuWnR6QgnXAWjIROR3vL/oLt04E9XnRMqV9HMm4p1/R
QZc8hR0UPmZIpymlEr0MS0979HS/ar0YrlevLIMSuPi1agZ/RgxlosLHq9EGpDD1Yogmy5TpzLBV
4gIHyGb76E+Sp6IvmlKg9ts3OoEMH4Yoa9AZXp8LbqP/nY8lWSVVxAb2ANrSqi0gIKhZVBG7o9PZ
b4+W2NtkxrzT5QuKSoo7v3cmEFxaIPQLheDr6fR2HgmoqHLHpZeGzfRC9INgzqqRTDxqgeuCCYsn
vbOkmdy2HVV9yl7zqcnH2O/tWly4k7iVm2P+WxW/16Xat0YVV9foiBL+zNqi3TGlmsjcdxM1Nq7x
FzY3vEZ/Sxyk9DfNOMbSQ68EerJj4AYZ+j92Secgoj1fiJbsZFNDlwHi1ge2bIWDnSagkqZ0aGOW
EfczcOo/HQxcOjjRd412OSOI7QE+720ryQbzDxCHW1dA62X1BamtEP42cI4AqHydEXapREpf3v8b
UXlETlwGHp4cbLkR7gLtuwLA6n/jd9DTTpwo1AMxxapbT7Gji9HXIiXVABuVqXAiy/Kggx0YRxyy
81tCvyNm1NJhLNI4tFcaKiLOPcp55H0N/JNhf9QsqZ2x5YQE/hfKGR88zvwYJzJMfQgTmtuwNz/k
OZFdMP8DEx83woWdZG8XO3pkjnIb7fQBToXRWM8y6okqEaUrizgVHjZlCzAQqnvEOnuwpkdS2+Ln
cL2jHfOAejJa1+piVLEWhxPNsdsmBXiPQ4DHzbKcYDjT3PZLuO85/6hQAUSLcujeClquNn7ie/u5
Z2EbqptehCcDGaI/Vljbs0uHjTrwuFOW8m8ybDDw1sotAIdFyI6WcGIMto2M9VnQn9v3ubOJpY22
CYIOtckyiG27j6O3qPMFRR2R2P6kk/Ln07fcE1Cx9h7RMhUooR9LSnB0xp4C7wMDlib4Shd67RkE
LCEYVEAsOi6hZ9iGyNh0v3z4wT/c6U37PyC5mU6vk1fwkaZC2S5RsrCzyNueJBvq8x3EDWV2tcPm
0tBBd64eMazB5XMKSSrfQQBMauCqWsH7aP4XmsPegroqLTlANnbLvQxkPCA7x1X/HYbNkn8HDcYe
0GEq5eiGAWEc5wlzaMwj6A8VfGDaa9RhcppWTp/59/8jHka7D5WFWaSjCzrj994KVL4qVCLHB/9U
U+5Xa+f+vqbam0BcWUSlsUrql94Nb/QUHx7JOC7bj/6TS6ITo1HG2YRFgwSqiTVahGcPGPNHrU1s
AgZPgtGcOo2sUHI5xq95bODJCNHGWIEHHyXp4FyQ9zofPOXuB6dWfApuVnScRvwvdMh+jQVTa8tF
nWloq1kvkTen1nNY0JspT9/Jxs9ytH03XeqEggPESkbw6loXnHqeApBqlEzQrSi+QDRoYmMDOb4K
tpRh1e8Rezj95KPeRlHtHPglx4AIrRiyZJOM1s+JpDyzJa1blz+qog8Ia3OYiky3xazOymkV3+rt
uoj3m169U8L4dW04SorpMN+sXqpIcxpN+sjnWRvg1Wz+xG5seFmU3sUl/zBBzMTH3CRE7ZiuO9nh
BPOLRkDnmMQ+g22iyPA3qvezZxmhYdHD6nJD6D7W+X7XyZtDbq56SfN1rD/a2W+mw6BErk6T4TpA
xpGGUBuxxijiXjPjW8lvg9b9nXuvhA8pbNfmU0eouRkz9nCFBy5MQWA5+C+13iVUd9JFECm9B/H2
nxufeDkbY26/INxTRt75X+dfvAu7aReK2BQnjwh7e0fNTAQKrWWfqU/oCMDsgWcMtxGPRvkbhbCc
VzgBI5gr9JyM4LLvtTzNuV/p1GQ1qtiFBODUEavlfaANk9NQuFyaJrnkZnkWXNh54/wKGCjBxzoV
OqIES5qXnMhCRvDhMzjiJJbbErhUAYznxzbGLoHpyolQAXXetaqAbJrUDCsT4mSr8DvNoOknUY0k
KseTPL7eSjbo6kRt9qMqvpOFhKwIqwYQO/RyRZfy8XAJga58vT448J9oXYLR9erE1iYev+qGkvEZ
eLt5/K+gkBg74FvY8tv7oTXU6Mc4m/7FQPvYgtw4uQaS8r/ONKTKamIs8eOyN32rEH12X7RI+ZPI
B/KK5iOm+aOJSRrCG60z3rIvcBE6fcukq5ng+utYNK/cQsJmVcCJtV4+f1qwgmO5HJVF0LNWMUZe
6QMdgwtDnllBES5xEevqCrnzKc2YaA49rH+Z9BMQ+lo7QKH/8wwmtRiOLN0tlNU3kvaABUYhg/fp
MU0TqjbDbKNQMeIEK1rf7LjeGa2YvTcH4YrnbHihCcIsyLMlT/R3rzQoKCdmLPlsnW0yV5sJ0Ima
aD3P7l+E9BD0dQJpFAVcTlu36g3xSN2et8OnuwO+HGqovRE8FNI7rjKUqlDGmDr5Ca22TbCdGdUm
NvMSHF6CbwV+qYZPlVBUYCbt1Rqx1pxIhGvRG5u2ZSPlL6OvwuCNmRL7TcDKYJsWhV5Bzdr6P04j
4RpQlLgTizbqZPbnp4YfxkQlbJ/inAxde1V+vbyH5CJOmkr1NQe5vRAG7eppjN5ZbeytkihDwtGm
jvMZENBsNwWRs+j6hsCkz6vyKiqQFitb93ajF7v6d47QZBNTZgRJd+Ywyzlvn4a+xX55iRNaK0qF
7YjM1DnlfRwyWZ8cvi9qPp4FFgW/NibSCtzMQIMxzjiyualWCEegvKxB+pS82PM4/JAGWTEtJzna
6yzFVYm0flhjTNSosfLzYVeGDGms6WAsAjDDEoc4iYzZTBi2f6ebdFGOB5razxqY9+P45bajHD79
dxOMmboJioF/CORMVvVVbMD+PZfY/OTp+4qqjVbqmMC9dTPU6VugQF3XQyTcWLC2yn70/mOcaZe2
5kEGNnku0RQ26f38rhY65FSba0kaoqNiZwAJNBX95wJSqmPSfWQXCC/JG5dD9SBBqCeyJtq4MuBl
PGH0k/db0OTcUEua2aUVoRFQepWAvR/wio9LayexON1MuqXOXwHCjwpPs0vnC9GSjesMpv0KWndK
cag3IQhZ7LhN3a4sXseIajKwEtXeZaEwh3ZXY9lwjRts4UyMyBvWEeVKIZY4pOC/2xDrbuRqRgEX
qD8LGyenSLrpPi7Hh4Yg/FEkp9zaPk8yzGHobMx1hVKSgpayfL3UfXAKkoL7WadbrcSpYT7xjH9L
Y37emr8AGyJDuXh86XvTlhq39NGQh38VfE0rsaytkZ03DLW67j+OLBjV3XpJmJMUWI+ahPCvfg83
Hx0d3tfbzPdjn7in1GMm+9jomKWH8Xh1KMDhaWQLErdfWnF84wELpUY8bodVFyCvxOk0CEiYt+BL
grT8eej5L1LKEzMZmFTGgo7TVFtkxBwVKHPnxuwAk4Db5V6I72POl1ZhJLcnxPb+tBlUPUtLq+K3
QTrP08PjgDD95tHmIzLVmKziAvQtXiPusoV7LaApQE4ZGUUMXZuFHLqqn5H4iAWrq4tyVM6emZla
xv13a86543GJ0WLjASGk1EqGe0HZxqnYbtORmUGfb2YgnC3VnQuMcpXquYDBu7Jz8dH9vhQi4ZpF
mKrpJGpKGhcDaYmO8VKDAsOChZpfV7x3ZJkyjzs3QgvoFyd2mO183FmZa+5EuvWIiNy0S8O17q31
vAknJNLQnZy/seA6aRNbJAhdOIZ8E679nHT6HjkUzhJTBYeBc4ahS2k8Uzf9p988eJJYLY90Sdtz
P0LzVW9KHi/syl4QkNyTi3WUtP7H7FFolsDkoFrh5LTbzm1Eg+h5ce2dHJlau76Jgi/WFzV9bFKJ
Mq8pK/D6AjF8JqP39FEsTR71408PFvR6x8AaC+Ape8bF/oUksGqmwd22cyqxIA9k6aQMkmQY/I5p
dDCsT58BOwM7GG1KOqIQuheiajTyVMalXudvQLIcfurxzEucoKG2vIccMTYY+mQ37maIfymkpv9P
uKhctZZCwaX9DaPa4I14LkwMtAxGkjW4K6LWlo/dyx1IGAs2FEl5S6sfcdMAd/dj1K69pOUVCNKa
5EKhSEmpjW5E5DtO1gGMnVM9ifXftlsIRB5X/2o29EeUiRtIJfBFULPrUB7CmS0vC1FPa4P6izjc
Nil00S0s7E0gXXAhPUWKKz0PwuJytOPbv7EK0njpPolpoSVAEQM5UaUV1oRzlzm55xd4KauTr0QH
pcVilPBQ4oNIqO0eWQWbkbg46RZbG67/D/N5kJnEaKy7EBm9wpetfvaTAhO8sTCtZuKzZAsWq8TE
bumXlKxYY322dahY4dZY8f70g2h4j5eWxo5Rb0srU3ohc3FYmt1nwTYJJYIBVis0Cczqqqxg3BQD
N0+1weuO/PVXjAtPISK6T8ABmvC51LQFKU/W4TY8xXhX9E+qY64g2phEF5KEKsEwqzfNTCuQxrii
d77msqvhmfW8Sq7hOEXkv+WGH7F2vM4XbcZW5yWRBr5HJBzFKnx9GVOeNEP7L6tPHHWnuQOO+baf
gCeHlTQ49QfJQ6NOA2IL/wSuxeqcKcs6N1dtjbbRkbGdWnc4WPr6KkLlw+IHylovbhngk+159i6G
kQHxCQdK76KAsgvBPL3g/7787adR6jOj6DFKryFsdueg1qbQHlUi2r7r3YVd1jdRtcIFQDFn+UQj
g+cRj8DpBci509YcuDWONmsw/CmUWT901SdsX4FcyZF1HEhh0JUps6Tw5x76ernagvuXT5/4c/CB
kYMw5PPvPb9/CyGk044OYlb7XkJByTKUlSlRDkYUl5dkSaskgftHcwLGiXgMiLsT3d1f8IP5m3IE
ydLL42rX3xLbfEQGKQlawZ7zvV2apHT/YQG5EkpMMbKDegCG0D8WgEKkPrYktBRdQ2eV8E0Jyo6x
1RF4tvpwrNp/frJyJ5oo6v6MFa6HAFkmXHVe6agIovQX3q1yMkU6YcUzwNn6gdHC5h1M/keWZS/R
6ILd/Fjbzq52KuDn8LNHIwsizUFhdlGB6+vkyOSkYDFMbsOUnBNI7OnrBeR/LgnDa+5XbfP6wU8O
sMaSEG+jmctX1k/vpo317pQNwgEmYDv7/nwnWURCL84JaM9WzlxmnGy1Wkn8lq05SUX0ucyfTzEp
kWDYdQ18bWqjdx71Kq+1MNl+RP84cKbhKY7pQKgZGSNcONWCUudrDA3cYqxbPyiicmuXLm0wSlxe
7CuScvVa8YGGCuCo9Mpfc2L6LXiKIVyC0egewq4aiRM83MjnUPIzMgD2pJv9iKHA8p64OKieYjJM
7n08hXeAitjuXYzNDgRpEGH7n0CzswiKBKq7DRZo5nTPqbGn3JCE1Mgk5j5LAjKMjWt4ytEqCFkT
gYDRAJJFxOV6XscnH8dW6r8t2JQeRZsMMPhwIFCNWsne3Luu0Lmxz+P3QJkybk2s224mgYL5D4TA
MDx6f1XrAHmaR8OEUWYLKsRUrjF58xTAvdGDZwewWh+PdNFmslEFbZvGlV/ouGjv3MekQpJoIJfx
Hi5kjw7CflNM+v17J20wrd+3ev8Rv+ubbROmx8I3uPGWOxBdZaCFgR+Oe1DnBBEKVapOGBa73cso
Mk+p/lisGhq+nrhvhjN7jd4ZnehKp4myAa9agPahdgCGE9KFESj225u2tf4bzjbqZrM1hO27CJtF
YGaTYw4M5B0nnIZX96IgEFQblFCgjfUz1kyiGnX/cXy0y7j1Ezq5c9V0v4ATV9rjItj7b3HRgl9c
SEOy3tsPK8OFCWFgdCGfbnMpfZUq7baYS9v5F3QNvAekQ6hIfibshOU1yNLRMBmSEKlZASPU8aub
ME7i2E0skn66M+73zJRo30JMLuSoW1xZv+E8CGlTlVlXb8+WL8CAh8bW/gj4t+6sMSpCoMY83pJ4
NOTdn0o491xtEKvOtKlP9CVC27VR5tXVCAfkxjaDwhfkjdb1bi+PSLlINWWlKhyIZmBYcXd2bbGf
tHSg/zFizZ0CSiF2PuAFJEFU57h/FA6w4zt4B2lVkU0mJB+CeGoX2ULHOKDAV7AxVjX0j6IxFRLl
Y/ZFqSZFieNJrzEOkjYUn12lAftXBq0gBKSrvkqvWzqETH5PC8kVsuquPGZaC6zitZ4iMUOcWfQu
1OW4GhXVT5Ve1Uo/DSJ5ejCUMumL7BJkfnLS33Y8oTuvxdIFaPt1+CcQy3e+iNyND3rqdncg6xRX
LLlDnjs6gYEeVdolBmu/akV8XnuD9R4F6TJDlCApXEvf9KV1tBViWgNgtRZV6Ma2Z+494K2EJBdn
65ELL5/M00VSrZUKLgbyCpr0xcSnWJWiWF1ghCeKu4D3BXekK4QJn1NYXG36IC8tNLRI7E0kzD10
VExQtr5iVNYf+xB2P9H+ojuQu+SqBMIvOE0OhBdpZ3OzTA3rQv9Hi2E35lpHn1GpOkLcJWD1cnlQ
3U8M7Plk2VKtJ6BhmK/o801pCFVty/h3qr8k+V1c+Y80r4LJAPKPklBv95scQmUKZghbMW7RXyMU
1KAa9h7O4aa+sX6AqDvDv1F2axEwmBEhtMzQW2nu8xKd2ivoqAvnTvay9aMkxysVWapgikPiPdSz
JoskmBgXDFlf35uiiliVBlKHiQfBY8YmQQK8f/qjpZmBGTl0zDCeF7hCVCIXTsNATuS3dH6KgUWW
AKDRsFAIgoJVlFbOXDiPbJQ8tvtinCMqfevMYDLq/6YpBsETxJISuAAOrrTHysDaCMXYrV0Jd2x0
Bmnz8uh1Zk+H8i+ujdHWqQ7NEL0wxUzOCnvhYvF1MLIGDIBVI3fWzFeFf4QjZ3v2n7APa9VPh7zX
IfQUCHSxuyJwguhZ9iexeAtKmW5UB/tsdCT1kJxni8n67DYKV/DZmwISgXYhHFV0lrWr77KusDxa
b5Pj54nO/LnOEvmeDrjU71PSCtltv5oyDrAhtIVGp4xsKj2XQots5LYRwrQNbNNtpl/WbDxd1wPw
DjaPioxynjENqJPsQ1+1cjavNjqYNUmtX1vvzPOUvzQigbmeM8+TW3EtEzn/7f7nF852cc/2I+06
B2mMt06vDu3lRli29WoU3YI+Bt6goRhLzu8JhvjijbgGfk1hCP4cA2SZ0/QAP8+kNo0GBRrZkchO
91rCRfeY5I8jCQJmRUVZk142Key8gQ+XPOWiqXkF1AlF63f29AcBYsyfdAx3uxTBI6+eRC0ktAVh
YQySRLcKtpSFTKj8YeTsnp3BPF9Pk57eg5DjRCeXBnh6Apx+HED7NssdXyCHoN5yelaLi8Peh3DQ
YGdWDLvOsRO8q1ucTGg+FdaybWBuadkqTlzD1XJd+Rsv4Ui/Ja+jfdhJy4CtlmiwqUiQPpfXWue2
1z67r3QCZRNzfIQzwQUOIQl6QwWB2K+cfkY6I4Hu4RfzdoUGzWU9jKi0uNvl30BdxMpEfV9wpneZ
dGhTDsEhNJv1lyfoBV8S7uR6nWb/CPEKjxc9MpkipL7Pv9jl9VQ/fwlUoZ2RVBlHSUZzJ407f10X
WNPF3hyZrP3c/6zaFGIWCmJoGZK0HoDzMOaQLz5xZ17+9d9z2jEsMHxf5lswD+M0aGxQ8fF92Bu3
MeopJajL+QAPrKGc0m3RTn1A19MsGqEg+9WAKyT1cas8C9JvJXya/bfYOJGiVK6zqYSXmGQYBJWL
HNbdEDUf0TPZsU5kEZ16uF1aHqMTDAmTMcHEGsgUn9488H91BhCASIonUEeLTJ2wd9gwvsgV/RAs
dlC1vfDQxr1F6pPWuBezsze5bFHTVoqN5vzYltB6DtQm0B9mX69QX6z9/zOp8O4/LSDTndIhTCEY
WtXjvDbrtU3tYaU67TNfz/U5lLBXydCc0MIeGl3n3ZlOBo4sA3jBPsNYlXS8jBovHJ8Xti+8O04d
yJCAZ1xyVI2Zmn7zvtKRnTlVD+0F5E1qBqBlOwdwaruL1b0INX+Hy9U2/RaEMpET533aL0Chmucv
gpdzfXAzTja9R3PzxhZcOr+OZ5S5s0IsZmUoiyTokkud7fUYloptI66xVzri90Dw+JL2czmaRbNF
D3a/OYnwaAv10EmgLGfZR+lGPxS+V6dasahC4SlX2bHV2De3nY8/xgCEIVPsk9wCqjm7qnnwrRwR
60lgNAu/cPZ/42Sm3cyHTmKtn3Z6LbfGO09ukZFl4oFRF6M8mqpvSzvzqTj6t8j0bE1XVmlj3PbE
g9LgpK86udRQEeoJSHcuZQjbakRYPx18Ek/dH039m0CRKWi5pcRcXF7vvou2UjliC2e9Nt9dLp1d
v6xmfgT/jANVTr0yvVPkxg8uMn1EnH7GLRk4QK4M0Y1OHKtn/0Tn3QSZbs2dFGyDjpElAXW3AXMi
Olm5NzlLOc7NhPr5fr0UnRh54DUg5334rOKJJADaP6mIGKSqv3/WN46sUMGMyynI0tt2Kn5+6Ktd
XRfETvJpExUfCnKvWSjl7h+Oxc0USe4H1ife08xNGy5jDS1YwnvbWLbJjky7d21Vw0h/FEhU5N9y
6dNan8NZsS0YET9lKe8sLYfqPOYBk0ZGfHatJJ/vdEBgsGadXiMAeOe97wJRNIKxp3t8lwSZZhZB
aPDTRb7R+PJRMmreZPMGwRf2sL8F/7nWSOpfjLJ/ODvYSktBAGuPQwn4HdpLt8rkQUUBmCGZI+u+
3O60nFfp5DEKGVBTrVjfh8edn9NGTSHKBcFKZIysx1zGbuRADfyHKdcu/0cXT3Qyf5C1a7ICwfdV
ZwmzkJTmbLxY37a4whRNpqG4sohp5ZgC+mFpAoOy41WFqCSeiaHe9tNzubkf4ooeib2Jln545Ils
8zYHezOzkyoSOAUfvAMtofZuWFyY3fGPwCOT+o92K/hjXFdSwU2tmWmrHOCFuUbaAtDunk4elsp/
PqbJxXgvvfjc38gpIjiO2o5eu6wrsJraUF+Rn/qpI9bm0wL+woILTlZVvFbXWIp+dWQ+JpZ1Hsc4
LiqbO5bHqy8kxMas2TVhig40JTWYTuUn0WPZ1n5rWkpiXwuIGRMaKxEmAf+XYwW5QJNvHNAX8lPQ
yyVJB2ppV2BrajXD3GqAFjhyhlYddOLf8gfyzEBDDcWeP7T1q7ng5FD+udfqZBZw14dT0+UbxF/5
jyVGw1wC4HbGbkve81ufLzga13RcyGfb6XRzc/TW07wHU6bjTL1IZ1Iq0TkNGz5EX4NSkGQd3Svz
5KQDTl38Wm5PmQPdRq08mAA9vjBoevacmT2bT0nyGMJd1nWzRtViqjdak/mW88Y93dHmcBsAPM8b
CqHAwyhkrv38ul2KU48lnn24CRvHLHb0wngsY4xUFU7oExV7KrarHMe6hC/4ORUZUmmz/0YUCHLU
PPXMOyBDU86xeNBUrnOYvml1q/94JKbSNpEBPf7D8O5Rqop97Ph6mkIGrrkFxj31jotpLvCBkgju
1sPxYWsSgUXhmchjo7V5Y/jALH/iTUCO2nANvC28m7HmbtFNyBKdwMHcRSh6BF/7iJ885Nm6wJh6
T+ssXj95oOZDXisfV5+4tzuGj0c+6pl5+0PzMmkhdfrdVyy69sCk6ooxtQz6IXQDv2mWd2YFBZUj
HNOWjFPCjTNE1XjttBLet6lgFWmLYAjhw9+coZ1wIiDN/ybHwzLZBF4ETVCr0p50M+7245w8mEg4
vJ4aW6RVqvxuBGfni+R3o6CqH4bgnrYXD4TT36UI7Z72AAnJHXbxZv5HS72Fh9fc8gfs0RTaqp61
XToeMbz4dKGzR8t9zpFcbadJIE1GkKd5v6V7YmBObR3i1nHsxt94SCRK+f/di7kEhCebFAl+c7XJ
ZqU1P2Yy/ij+yvHIui8PzrRIzheoeYzzmf65dbFnAsEfDf1EvNIeKy8AnJjcTfbjWwm3AT1TbKEM
xG1V804p3npVlDS7o7LfDdkoQuw/UFrN1gtrMfskYNS3fKTgGopSBiPHMc0kcDn7tyc0XaCDvjrY
USBah669qkYFJKytss4fY1ogfNTvYc0cNBPGlZ5bSw/1qYjT/UEgIf2UMbtXBT8r9joVlQYP2LDb
iwF53Z8REQ9USbEAGLCCKmyvfZ++rBXNVbioxA7FGRVw9m8Cv8MKKwapJMynmYlo784DtsN/Z+g/
RocdfFwwwT5wIii6BqpqOjsFbj9g8qtiI9tBqbv2st7SSkcruNyFIXTbrebC8yX1bjsIr8i6f7ru
Thud48Pib5lZkXyqaGzyShGmX9wDs39NMPskSGAINDPoRWktYGn17TesMaqJXDRV4BH13DEAJyol
idzzPKyWVsLqn45UHNh2mIaNyQrCFxHFtxt/M0uwo/ceGWGU/793Rse8PSvg7TAxE1wthH5tF/5Y
CsrfHC/V/OJf2Xqi7mXMbQ266GwsT/s40Wf4CDIN3Nr0n2HQfeF5zmAsS5c53Rf5k+g+95gU4lJT
8fcK/rR31SEq3z1q4+z9jp2WEvFMQXoRVzvc7X/L+1bKvOpp1qGbxp4LBtg+/CtcCD+m2OV1qHxX
roNWcryLlzisYhkky8fL0oTIUwdud+6Yxrm0lJ0SHKC+FeZ56iu90YWaC8rw7UJWiVHezsRDHupy
viqjL+6IVfkrr5ix8zUsrc5RX6zduhb4P+dj2lbBXYUyWoJH8EqHYSrrdnfhcAyq804qEd5TPXMJ
E6ymJplOrsEUw1bu2VfKZqyJrZEYx3GdhgG8hr9Lrz7TrVT1MHtX7jMooSh1qKdjv7KzowKUhTP7
fR52E2tFqx4derkcO60if9S2UVhYRe3y1ib3/Q2b4OObjTorVPhUc4fIviM7j7nfUby6xSWl8clL
P5sv8QIJ1r05eaKksL3w9Pew8E5QtoX4VHJERJGz3lO7Q9nkych8zznd4634Lyd2ABtfiGTitaGC
DqMXk8vVhS9mzvq/TdMTlU6DkIsOmjGbut6A0OcCx8toKMZ5WS3A0CQ3EBuEjKYsKNwmEUi/5v/V
1YhZ3ACIqL2z9If48U8+LxZnVo4o0mZ+k3iq1IeSlsg5qNXHlFovWrfgAf74cxFR4YGGH0p6PJEf
CjrJbJTco7AlN5Uu+ktb3L+/xVlq2kVY30tG9fjuuBM+ww3/i4IOk5hOGRoUWIxR7HrIVReJMjkI
/zko4zMJUX9G5OIf0rF40EA34R7Q98T+Mhn1dv5/27/CI7ZfpGyTr7C7pGn98CND2YPj0RD7+I4t
vyAtQxIe6l6asK4BT4Wi0sH0pUFtqC4PAWrmeCpGyE1pxFuQsvtErFIvGY507SioGhBZknHGX/HX
3wbF3+zbpx2HSAMiz6RmUHGCKA5Qda0ozDgwsqpxPKG1kAfeWeL1tmDMG19wGOZqewZR1XMMPFgs
T6FbnvT9tmiZ9033knENbooVrkconVHVO62tdVWVYvNrceBxraUnEgg9bp0laEXJRKrDZGMQG/9T
I1N+3ZmfLdEaGn1MEIurOb1BOWaI5FLm5RECxlxkWXcUlo+83gzeZFhFCPMlD5Jj9Ayh7yJPEsD5
aVgoHXWjqSZpUhPSDumec+w2XE6rW+0tC1ejjvFRFTBAKpmVEbn+DiljfduAOmgtscHu1mizV31+
AXQDNbHv7vVx7Ykyau6z+iCWQLD0do2k+JSIihPW5VtgIsYqcFL5c29x78rkUpB5J9L1CUa8IRYh
3alUN88FOcK7+lWqI4rjGxCbkIj+/NNjrJcyexn9zsoj4Zg5FBMUGN9HAMKNJ1ODfoqSWmk2Ozg0
ZD7uPSnDU5hVLTeba2Z5Ck4gzImmDiYqTWs73fsdU8r3oEJ5yD/RtgG7A3kVu6bSKlDNGxHGLrxK
ixxF00jU8rpI4qQq6W9qsFQFY94Gz7ud4Owi5aSlLD0KrVDfRx4cbn6yF6mFKunFXIDJ1PKaaHQP
DdHgIsrQj+nalXxTgdeyH/PNg/QYyyGY7wlvLQEaouP7yU323RNXuoRuS00/I/+GbT84Rn+I+4d5
JBigB6AmKorPzdPT2OHNRBVQhD+PvmxgIotaIb1plGSRWxUx3meZAr/fQ4qtC7VJAGMgUgkrAV6/
/O4AlL5gK5RJfqs/o6XkET/I3gxLxby1tMzEIGURONnE7/9iOKzJEvoPAwINhK6VGXTp9wWfp2YW
/8D7YZH+so6IBGy8fTa9E5K3jpOBeHmrtChvWrj+MvyHY9pQJ0Fa3VKz5W1vuzx0v8cUaRqPAHet
szqUMWusVvUrFLbqB+/O5jb+DW9z7Aor3OuMtXUBkaPSnrhjFX6trkRp42Ctw8hC9Hq+EtJQCZls
sM+ANyNlZGCK7qDo4ntWeW3/JqOtLaeCdMElVi4ztWwGfap2IKbU52Hdb8/w8aUhXtnFgkgiZQSz
/3GJMjkrSqf6JwbvZ1HbgUciBj6G10HbKzBL/GHNHsY5s4L9vMoh4vl9RqkJOJj19vT4O4yIzH8h
FouNRCsoHgtkKQsxXIQbhTbITnfNgcErzSGv2Y8co3OYmvfAHJNgeg5gNi/lantmvCqBB1uFngWL
GeHm4ZLjYWkSklusTwgogtbGqwCLTf/vnlyeiGU1eErmZT4HI42quBQvJ4bh+DNXJwyJ6Xz77rEy
iIOyXLRWsewrWmgjQu7izAU86uJtIBkplcqEpB5swEXn+8QL28tMwI5RwKiVh7Hd+soHMR1N7fRP
bDi/B3Ayuc5V7/JOGoxNgRixbHGD/NRXZnRuAUD2ygfUE9xtQy5ojU7AZpMLeuBRaiv06419Gu5K
2nIGGP6kL8g+UE6KRKJcm3UCGp10lPNzf0bG7b5OTFjO1VRd2sasp/wa1v9LnvkRPXG77CYO1Uhp
u8Ra+DZ+VnyIRCUaUoXNsDSpR+aVG8dnnnhJKmh0yAQcDGpFvY8hqItHdmvkzbrkM7GzkPux1Kpu
dIS72nYQmpSD/p2wdqGuyaBt0mcG9/3eq8vi7/wOwAoGGSNQcK1gv5/obdI369uc8xvwjQSalXgg
X7t3ZxgXaWuf0PFSdLZH1WbHEQhHiFMaBGUFVqtgHdUC/sElF6QbfVxmQBgXDRm2KK90wUnXXLim
PRGf5uv+J+9uBUvt2yhj8DPdLQyi6HEiKkZRealQjKihuJT68JtneMhhYKpV/ubCfvYVMoxjOKZm
cZrnvAGx1L/AK708hBA/F4I6J6VSpanNR6Qe+1rg5qvpRsKJ/7JnZ5a0hJmLwXwzw4HFeKE98T/j
RlnjYQ1TxqpeBk+AdzF2riQ2k3z+CHsUbD8zsRLGumiI4R82aW3WHm05H7wIqrcSIX+GdiMGQtMX
iGDx0e45x0wx+22+Mj7EXE0YKJoFwQMdLLtXB1fuqbKGtaqSAtbKPXJWBJ29+Mp1wWl+1wiBSGYp
BLfAYew9UzbE4OclPjVXRj2ExNKMueR8RrjVfbk/sfm4j4GvjsVaxw0tbutP01f3xPND02srRqtj
sYBtHupN1BSKMKVlYJTbR8fDRRlVbNTNT/MyhWIczMgsriBQOoCQy7lZkx4Kiw4Ahu0SOeSIyYuH
Df6cfWzxTrP4Aa6ebNg9Hbf5APrKKbENF/F4GRL+H2fIZti9/x97LJSPWBkE8rziuueXVGy8jUbI
3UTfw46Bz+ymU+4wJ6sOnG/IXdgoaHizNh4Yi0SakUhbU96OxSsCXXnQWwS8bWmVrdQtge6zFljd
Mu0Yf5MxlbpPKaoT8kfJi4pbu5Ss9Ruj9rgfRHF6leuo9z/Pzyc74Hp9mYCDsJ3bqADlOc+72GWR
xfsDS35gLxrFE5HFk1rUlqz53SmXrFN0C3vBs8DhkmjfEEbU17ufSv3J5Q67n8lmfTfHoz6G/wrK
DFy5qf9MsD5OWVjLbaiuFGGzdcGBnZ4y0B46RXIj0GZXHd/U2P/SpNF5xDWIMmzgnEeJaALlGHCM
rpHDsiQTTCbZM/QPMzQIGapTe+HCJ2btjkYFP6yaLt7lrY1OeLUeIWJfRCsEG3/sWl3S9xQN4lxv
QVt63emBskDUXMoaj49mEe2zAhYXywFjxR7+lrjqHIRKFyP+hYpIGQUHwgfN5KlGyY9LHlb2mCT9
G6v1zdMoPOmNJxcGwSrqNg59XC+CADkuN9S/5OLTrlwQJXoJmb0b9KB+005OH5Xd0xvhgt/P5NXg
E3VHYL47f0OsSmgoVBgZnI5V19+Vf1FfZLzbrnCeGKTb3yDektkV0zl3L5NW/VggKszd8QagSxuv
5cC6wPac4Z7+yj5BorLHjuOUcF0u8Gl6XBHyI27ctvnl9sSD0qivQf9bOnLiG45pL+J06aChbO9n
xTDczgHkAaWGsI0FkVk0n43OxE8ULeh2ymXAu83FixyGYJy9PrkDKLsG7gjz9gM3QSfmh1YUzMDQ
kRpDAnUZ/qHgiwxDh18YHfTnj1PeeJtMBF/PbQQuRWTa8mAEmL/tiihY7Xa46GuwMwNj7tOJ0Nxc
5JUQ4ke8FUDQM4PyL1O2jQ08Hgs0nm47oDJAlVHNHfXOzlu34lihg6dvzO6w0/8QxXz2IFnOyH+C
DBCOyzeEmIfTEyGmeFTFEprXGAh6uuHAY0WE/Lhv4kjCf/23WLEp+ChPFtk50xmB/DFvhUMc6qMv
IBeMVgGiQv/ue+MscpL8fLGBLiXrU/lK05fllGIw2Ln9NDbuA16MrabwlnkM/S0SBeNH/1vl77L3
GFLqL+UEsXjqU6eL26T60cdi2UzxAGofxGVf07RTVvPISeoUuqYnWYlmipRAgwMKeXzeNL2IiLSE
IXD1QIUnjnBu77/qzZC4MbQG8PK2v6mo3elJFkIkKI4WUmkzrhSH/HNqK+tmUT0kDEdENlGIiuOU
6oVF+3A6SWuQcZrCQO59KAVW+uSmG0urJ7IlUFJRgPFguG18SAYSXivOrP69x24+JSmCxYbXIGd1
ZPP76VPVNpZAwLHMkziHElA1NqrG1IvfTNk2Oh8Kp57gW/JooBSBpMeiktNtes4lBEM4h0umcMHA
ZsN0QZ0moLbDEzsZZVXpzER83dX946HzzqW4QqTtFN+pm9T+da2y3qBl25/5gzDyb/pmM5i+bDjB
G6PDC7+0V1xKiBkw30Huy7hMnjCSjH6s3fjj7BAtUna/u7jNIOD9xugkcyRJeUOS9jrv1m9FS798
Lxn0uptKw/S3g6N/pyCB1kK4cS/PfONuiGmPprfg1oZVnsfXrtF+agebXgm3AAb+CgH/2IM60l47
mAEVRGKVOTT/2cF5y0w5GFCVFN0j1CYeTYr/gR5WGQ124KSrIhy6elQbQY0jW8HiheMaRI9LWLPS
U58I1HNi835JdwGywKS6wGNfTGkxefEYxMCL1GXoXZgkZ0BAPbm45uvrJxLvdCOK0nKu8CqOqawh
rRgYcu0SdB5ucT6AajiitKQOO7z3Ji9EnlspwQphAzKfQh4PE+GxjEtLl2p1pd0KMw0xpLVciQcu
mFtbOq+RKP3iwmragZDZecYrwkkvlZqIvitbGHBaM5zEFrnIXWgd4TLtDPOYh0rRcbwGK8SArVtO
8ihnGKlgjSw+xVse8yILAIfl1yvjMBkgVGWH86BGSKYYOe2JAbPpcrmOMYAOp8womIXZEF49y4I+
zYj08xiMmqeMXtVUTyZv9DjdPeCH2UwO9TGAmCmsRb+ndeQbjQXwsNo7+SuccBruCISFt4B/C+PD
9YyHekQY6vb07XygCab9cgk6R8S+vd6S6yPP8YKm3gzSixcZixQlCEMmRcgUPefYR4s93ThnKL9V
iB7B83PhQe9PrzXgJ7nWDlTMdQQGJfm2skMTo4tVFxfNzeSKxdU/q69eJ9VVtRTBncD96y7k1deC
K6AQZgn2XexFzdK4voODr77mDKV7s/N5tlgmaAvJaP5FPcv2tcqdNoPnkK06kpTeIdyY8eJorMvm
ZnB/wSqkowXybHciiQuy5/heG4qdUeVUgarMi6YNrxGr6a/EC7XkVy4hVP7Kcn0ux6tTMb1JTECX
MwLo+8PDw1/claQsvtB6Dj5USNkoNmidFhGK/wMFNIvEvWBS9su+6VRtBxtnJu70fcwNI/M4Uc6l
v3Q+5rZuP8QifO9/nG5NKuhG4kyTwJ+HuvvH/MSHhSJYvvqxXei0z9fmntIMY9pxJg7KR132wX/t
8mOaLIVcaBJvzg1Ywgi8ucbf+Yr74FpxC/+OhUvXzWTJLuW6tWN4oiBhxqEglby4ncY/taEaJ6t1
ox5cjpTUHAdxoxWy8w7l+SXJYEKuneL2dp8t8ePRA3Z8r2M7Nr6qveimPgZpancDeyQfv43wQidH
f3H5khAtqvHSwVpTt6d+qa8VR6HPFbMrbc8csBweWACf5NEx7UzYzLECPFUvHpjofJnnl6OWGPDx
VahtrXgsEhwgdZ0kC3qJivPJ6aQMdHLlDFVnqhukQ8Mp/nYH2ELsAQdHrM2lclq1cHf34gv5qPUd
7/RVSWUntshuBrLFBtYc4EruY9mfrLFfC19/uEPNqqXOkgStvlmgL9raYCquyh5dn6GIGsOHKmE3
PnnQJZuD2txsInTydkqv8ztZ0QsxDw+Vuvo20Us2syZIJab/xveXzWMr1PxRvsv/IMezSnZGUouG
aBLpu3NPY6xjQdli16dgdWMsRB7cpLatoJc1W1TRpevKuiXbTGXYbveAbGeOE8nKhLdbWnf46gQz
SmmywJC4dzY8zrp4Ag4nrTsYWoDaXC64DNbX+fNE4ZlxoCmPh5JQYcAygy8LJZSD1txuMxl7hLHX
JSI6+Z5NewT9AyhEymb+TLEDFVa4ruYXK9N0k2RQPpkiSN53I0IKFSrrRLwbYxbcIRgNPR195ULq
UaXLG0jpb9aOqg8kNwtbNFPjF2jr8xzdCVfgDMzSDVKZWwFCT931/KjDVvt1FO1aW3Rx619WvGcn
iAAUzuy6KDbEM3Xxvg7F7xu8wL9cKHlDJvWMRwZ08+44XP1AeJW79OYUlBNsvo6nUn5eXKPdl5j3
A2IpWSGl3jAKP/90Ztp0swfxZbyOO3rznd7thwMxPEH5Oo0brSTBDiweucb/+qUIX+QlpRe+BrF9
yc7SaDs+N+Os+k9Vlw8qdtmzI/GMXWngpNyd1iDCxSdlOjWPDQVruQegnyLN+mMoyznHzv6VoCDy
tg2G7uQKUDmPgto/Vb71Xxg9yq8VExuqmJ5hlrlxwxBl4U2hn5ojczQTWhL4k2HZbETO8W3IrDrr
AsfUcVpCqF5/5Kw/HGsYEbRz6qCSTFxD3oH4gBxuGXyitLadyTqHsuGaQlYmj6RIeRYzyoh9ABPt
QprsxTw3hadLCbMW9QtOL9QZwG+d+SS08XtVQAcJNgS807oKJkGWx4dw+mTNczAQTWNFYGMv+Dx6
ate9dpzJ89tbpxznDGhQ3SR+ixbeG62A0+apuWJCPrSeNU+cgsAmqNyL1T3CuK4OQZYsXCy3wJTJ
fQMpvqCnBDsxgD1UW1T/oJZlNcYsp/sKH6R7mJeFisHQ9A6mKDkkXMZ73ct7zJYj5GoczJsguU85
uUzj7UKDdFrfnRXfuTqRlyUWrEAt07B6WjgTqCysnKvC9zf9vX0JYF2ScQWDa16BmPrWUUQ+ERAz
5yVX0Ejh5tomn9cu43030KqnSp8o4qBasCC97+vU4dE2yIM3ObKSuQPS8HvPVS1liMqkhzPAt+yX
zW1F1AZwQCuDmCvJZ3XSPDhi8ypiAKq0ylNiDDoQ41+LSje+thv+wNy+7d9cQ9xdg47bXrcQlUZo
7+RK7G6t4O1FO8LvmKi6xAHvFVXsIQ19uTXydBAIp4zwEoPIBdR03ZDIU6Yso4ou1faIwkQSlLRj
7Ek3eKleuAY/DvSGVB1kQjiG5Kb2+HkTyK9faerwcqu5VcCutycA/MocVOFqALsu/oFEwjmJBN4x
LKzk77GPrTBJp+NNBQNsQjd4kh4/EMu4TWT35JQKpEIIlH+fhIBnlcHtzk8OcdCBSpDbKW/cyQic
FLCopUEtXC6tAoSiGtCQjE1NMjsUZs+EU8/LeDKJPjJWCpyP1D4DHSJP+YIq+6vrNMOwe0IBHwl7
8Hm85HL21iSwZnDiDwu65StfImWX26p52G095BXDIaeYYYbFj4sYMzXbWqpOnynxip6uldogCIRF
iPUQaH/SEojvVfPOErKbZFubST5vX9477WHWTmPVIgyJA/62SHswJmGbM6CB7bhLY93nbRwSjM07
kvEysI2FT7Htq7Nv65Z0ab3O45DPRJmGDWwEIQkXSqiNBcg+mWxib16uU/tD70XXgA78OwxiXeXu
inxpUI+xkB63+X9nosFz24UHz0MEcSjx++p88itvEdmpsCtJljHSn7GZy1y+PyrlHzD81IHoHdN2
mIEanr34HTi/sOcIrIrw+bvAwYttmOj6Znl5K/ZQnAx4LC7mFBiOr/lu/St8SXyHVt67ogfJLJyN
1eVO90uTn6O7JIvg0JOJly1OuBp4Xvd4r66WVm5zZ8vzBLrUPKthwxYF6DRD3VIA0CDIvucq7dc/
v7v6goKVLcMs23rqN1VrkWkeR5kkEYKZ5ifPGQPqbBFNAuDEb6igNEIMGdeO6pfjojdygBfGuWbY
VCh0CitfF9psBo/JHpnZFOk+Gt069gSB8swL+H67K2EUUCpXQk+UlEx85hbDGM6rOnvVvZqg1PTq
21AhpfPAZN6REOyr1tXrOUpFrJbvaH9HdI3OrgVUaj5Ti+JfMsiSvuEfj6tgkx8+hBaHMw2s3/K2
EbUFyJ1Me4ZnK4qZnrZLIhw5kQuS1Tx82zOZiffgOz9rPFzYg+/ug9WFKgkT212DjuKBp1z6yfHH
KgbV6u/hXDj0MdHgwoEsMP2Kl9EQi7KFeJv1YwaH04XbhG3rYC0zfvqlK4VffDP/8MK8Zy/zbbai
yhCZHyhCIihDREGhQjqoqK2Qp6fSj1MAvP9SNsYtfDQKiEvkG3ej/6bsN2NH/0gD1AIzIw3e+Y8c
gtfxXSl/iWjTBSq92OblqHhm7S3F1SZ1Uvu2KEfMzY/Xk+hBvEvZUHKmjliJzj8TmbXFG8diIPXZ
w5EMRCJdhKBjimhExdtc0/36yBDkfCh+AlQlVtBZRauNbrBb067L4LgyPhZMnb+0yDmigrrqFUP6
1hNQxQtjZNSx6ekiA1mBs3l2t8djmmgTF6Wy30dxulrH/KuQPRW0uOmwhUDLnGTeenewQW+ixVky
7zvAPHptl6UzLOG8NKMZh3xplgOF1GESaHTRaMNE0BbPtcIBYvRtQcywpZnjYwMAfXFl/VMHI9Lw
tR+dUtOP+GLp0aKuRFL9TG78SiNGDpPaWRlBvPsx1P7qno3txdTlZw+Hmpvf1Wgwnww1DRCFjKgR
wEn3QX/EmswStdQL/oXN6iQvX4QsVDy492o2J264I9ISpBGbLbNJGYiMckWc94pxMcdaBBU2GrMC
7umlwUJliRxFdZa0TmY4Rr+VRrxCoGv4xXq30q7+JZSmXRSMQHXW1jM7BdBoWyts1Ypz8WOFR53D
8BwTLGy4DGilD2VgjyloIFbZoLh9TDCB3cYgYHXgmOegzQgUy/5UgSuuVNCMfHMQChJDDJ5v87dk
QUQ2008SGzS1mOVOMEO9FUq96qDqeeVkof4AIX0BA45dhjvDSr8TKItF6waOiCpB9EeUEgQaJSUt
fl82BNQPwDZp7sO+gcq28fw5T+mGc2A8YCF+qhWRMJYvd5t+t2+xRbWH+YA5JitMY45vf6r8sMVm
1ebUg7lEmxX4X6O6+i+kT2L/32fmHabkldRQbQuifVgp98sbFqLrvIxefQIxWyC7uamHOurbhjpW
ETx4uF6nIKfY/1NMNxHgTRYHUHOfe0Rt8cLa0u5nW2vHkYJpROH+eEm0Of+BPnjg55gSqbK4APNi
49mr6CFaVGfnsliBciloLGLeUiiyA2cAe5A1+Max+5zpBd/bkwKHkd3iqJ0FdQHWSCBj15gxBKOl
XFP+vRpOvmfvyULIRN9vzzq9gXC0zM/BjETT+Ie9/NTsrGpoitjsdrmBiTZcb72NURjrTnE1oMtE
neFYEI79N95KzG2DkoEBWnR7GU9l7E/O0cc0FCA3nKJ0RzRxNpPDTDrSgl18WERmw4ch1uwD4i1I
gGTtTCS5I52uMjiYASsiyYLYmmVgeUoIDTavCm5sTbJT7CrUPya5m8dUInYv3J2CTEGS52L7iQN0
oc3RFKFz06zDTkDImeIvDu2UR32t4KI0Q6YspaQWSW91rE0L3+XMMokF7aU50oQSGyKH+WkUR9w0
jBVPMuxTP05A6aciBQK7CoCCYHoUmnPh5HeDrBSoAxHdwPa5K7IMvSe12pRkMV8OkBXgZsUWL8OU
0YBDgGCffhRhSowXWvBceGDK4lRjZD18pTWj7n/0/RzaYf4LXvcPHkjiiPMjH4HoQTO77ExKZMz0
R6XI4qm+XBWTRdiUWI6b+LFmXziXPVJ9bckCl9N7GM0dQogP/qqbBEqG2wkylYCDO978w0Z8CPEj
iVf2MqctyXG0aFzRjydR4d+7L4qH3BTaWrXNWk9dgXbuPObVKrfq4kl7MZvsmwWJKQExrYiL4xng
2gUhe2HSBGIBuqvA873iqekhTCecSDvQYi/5ZhLUXB5sR9qTe2KkcyzoXxmm49PRO9miNeeZlw9C
p2mUSCfr5vrYRNDmbZ78+EEynuAfYanTrXAyZXWebxwic/JU4ytT1GocYcFlv0/1YtLucG0Vfuzk
oYtWdFidDpSoBPL3+p7PiMYZ2rnS3wh99VP9GW8M9O9PNdG7YFlhm1afEzknITDuvgmORQLKjMmP
WT0cAi91dtptzyx0CiDkqzk4O1UH+MsIdm7bn/K2qh5GeHLFMDacSpeKTXOGCeKgbVJBTtEJL4NG
HTbRPS36v46JDrNp8IlGQ6E7mAtFf8Q8uv0ugxRI/PNy90Anu1yjAakra3HhydA94OSQhavFoQWw
QG9RJBrj3XJwBkqGllRmcx95iwS7OuvvDmi8WlupkkpRO0t4goINVmK6Dv4AkJ+o3IjDQd6AXLnF
SIdRZ7Z54vwP0w+zEPkwOhicEX1/nbMM5YvH2YQATTnnPhVz8gmmA6CFZQvK4npqwirt17VLvgkO
E+SzVSFFCzyl5J/TVjAJr26zggrt203RntMaMxf7aFn2QNlts3n57p/sliY9sQwwcKP1UbQ76GR0
MehPA1xtsfz5Phuqr34U7CjbXo0N8KjXJcZxCEMxTGJBV41G9VeSPL4f2C3d97Nu/bEYGu57BZSE
VFARjxETsKwm+OV4E4xuPzeccMbN53eJAf1TDt5XhF+hykvmBQle7EFd/tbYUE5VMPOEVj5p2Lmr
QJ63W1qS61Pv/hQ8vUlDJ8+cM4hl1DfBIRTMKWQPQ69tzpDe34RE0VMq5TqRyAMqk+bXYer+yPdA
18pnKd8FXk6/uwNTomOH6qgSOGAQEjeN/T05hRo8IgxgLnHukaowA1jezEUId728X2U3nNqSlzJs
4c8XEmSua27IFWlQY7/A73VYEyBzdUY8dl1bMICPXaB8APWuliHksKDiwrHjjBbcrs4D3Hr+RlPG
vgtRDsPFGaIzhPVVhonuj1CVdQJTOpXGJNE16LMS80Fesou1ITRVMTZXlScoiob/+moJmC63csuz
F3IomtbmBeL5lZOQb0GrRfL8NGKCRPOKlPOIbHbu2N5cwf7CwdDMojiZMSTKlHjZ/mYGxuMyDT0Y
KRN+DBuYnthUwnAFGkVRo274eCmqjj/kpwOMGosZnL78YEPC2l28wFgUdBvUmHgo9qsT60eH3Jx+
33rOvV4s3I3NrQ23yHmU2D+66FGcCR4fWFBSUJvOyMzn/4MRtpSIH3e6sNV6dfStJyYCjIb848OX
/1oWVJAFLdWD+VW42zgfcOretL9XDuCnxgb4Zo1hDo+qXQqDqmAJNoZ9FgCr2fp9j7+94+6aiZOB
nRR93Uq2l37ZE6tqJ5aKftzQ382JCQWpS1nkpNsyn7idtAXllSYUwFKvRERgmJh6pqN8i6iB9b9Z
R6zdmRbtcu+e/LKtEeXoDDvTdkJmqiyF0rDLN1MMhBAO4rRk+LGsz+IkKW1xtm7MauGBormFTfIG
zMOC7Tgdwk0/7cwRBbKVVHjHaN8/RFTL4wLyXxqKnqu7lJxQdRZdvEr6vucaXPUw0AqpdneN9YNE
ACHMzU0nPU8+Vro+LS1l/r6vV83mUgCQecG9efpU82d5rajccfVDrt4dHvbwtXXpIwR/kqcXSHU9
tMNvywsB2CPv/JT03fYiNJ1f2RBKl6K/mLZ+ks+6WK7Sx1IFOExLlT2671PeKxeR4GrnCfLivWpw
GeYHVLjRWb3eSPtlAENukD7NnZhq0LZqiKZB92sJJnxsyD/Ikv6TaBPfqYHBWdxEkqiaeNF4qunp
uNxJUPeoDJoPw+VK8ZTQokgRgSdQ9I6CBRQZL1lqwWglbV5hNrYEgwfUCCNbsoZTiSKKmaEFQJow
+w6wtsy0St8izECPmBffaB9Sq89bBKU9GHEpWEbqaz00uBMFyaIJbywbCeempJLVvvLhZFLx6R4E
qWdxSm7ViQBT5gjZ0S4LfXPHi7CXADgpCfoB47WxvtTp0DI83sgpR/xjSMBPV/HJrQ1yHyZrTIdN
rzqScfpbeMWNI0RCUdZYCbI7hvtXdjBurwVziMq3+/w/Rvg/TCEMnFPTJjpwBizMmLlomoOuuXyF
nlRQPmgXG+Broci8c4qSyMmmIVNlAsQwFYdOE5oGx4HPkMOdBNMqWwQsnhcnjxalpbOGR6Lx3Dul
B9zCfdC/f0Jc2aMzGgvPidfYcw7HioGwJJSWHPCB8OlmWjX1RbhQ8K9mAJ4bj8TJxdDv1oKS/apj
8Tp9zBf0Dcni/wG69+GLT62zVMmKucjB1oR7iN5+O5lY4mMjKiY81J2wMIpwdP2m/86aJTeqZ1Vm
Z92IfHmkLwqPIK8+PiKR/ouPTmF88JlmVhRufYmT6Y2LSciBRqKJJn+jo5HG974TOCLlPoVBS/y/
Z369ZB9f2Offb2VXwjkDFEoAFqKywOCh6dvB2dagDyvu3LyOFAiFKKuNyTCewxXBTMcgl1HDZKZE
zxoBXieWWEN2TGoA83dSOwVosNJGbuebgFcGjAAZsX47pbNDMt1+8+rzWi89zjpkReAzvjFCPKr8
9nY+5UhHUUMXEeM5Ec3xQXJB0bpod5TI7EdRwmL/Ccgc6ZXG7OdB68sdQFCj211yF95ai/O4sbGF
Wtl2vJlLODqqk6H/VKj4706ejwhBVZkGYwrhJnUwURJxNMAnjsa9zp/FduZ+oie2KDayzY/7z0w4
uCuFaBZ3SAjcDWBWnBLNV/Y4IB19ZyE+AvUjB4Y2SckCIjLccjiHqsW5cAZlg79Kb/ZgoeUyN/26
Zw6ZOnksUzirfX03e+WhTfqy5PKqyF5EEGa20wZXbpBaqlOjXfuRhbj1BXqx0n541Z+W/Ey4G6bA
dKtlRD1uLFCB0pAlWGZT/URFIn3IsS5mUd2oZ4mRZzC7n1ccMt21b7lvB4gqgpzcmFJ6qOkc58uj
MEXC0tXIBa3vdI+lFOJBQS2WFXudabbBv7HOujaQEZs4rljJv9IyZQ0xqEEu/IatYOase4E5PBpq
p3xCv3YMoDY9tjVkyWBGCKePGmwwAQ7oTrlzUSzodVEzGIaS3XCRabUHdSrbLyMMwBoRS/4dI/tW
CilissV+IIT2g+ffA0lsbltiSZ74tuObkprX6z6pWNd4VAl54IMHKQvLrxrKS3Hs0oZv6yivnSpE
6RuVRm0gXRP0Z3kLPL8Bz/jNx2jCfDlQl8blr6xxrlrUr4FG9DFsw384jouQ9O7OZFJkfNW2g9Xa
OBRDM46lvASmIdLn1UCWJG+HfHAu0SQ2zWs49ko/i0VH7ZtXnP21U/QH0Nnho2mOpVYAIDNmFXgx
YYl8gWQeFwEYFwXEJ8Voir1hpAVevfAl1ogCdjJZT3KWCzVNge6aLY6N4t4VJDRZtvSaasMsQE16
Aw10MRAjTDnvFKao7eaqAEOkiE5WFdAvwDrXBxyX1gUqdzePl+VLUxhEL35pzUMLIUzQIo0s/M/G
J3up72S3rs9UZ6PcwVLC/DvM21xs0aCEL8/v4iTAwsbCS5gOqPozYbuzSj0zrrvk7XjC1xFU4mkJ
MCgYx/tuq8qNjO1flyhPFg0g5yAY/UctVLlWwb2s5LRAX5PsELuwM0kQmCK06ynsAi3hgHYMEztd
27QUoOatLhvTYVUxyrHoeHDB5plmPq7iN7seLADO91MGzUj0e6fA2rQs0hcCDIPppj7WkeOHRnEO
2pDxP74grlz4punDnudbep6xhKpvp7ffIPKL3us2Yl3VHkgYm8CMVxAO1i2pPWSID37UMC9BpROC
jak1YxJ1cn4gAyUGDU9wMEkrUzFfzOI1wVjHaLlTOzpT6Sh3sa4EvVj5gfdYyhT4FBggjMfvLkYI
WB2tIXQUFEk1/zkx7IGQA7jacCJpz04rUt6VYDuuj475GGFauu0whJ6kM49AnY34A7QQ6Kq+v+c5
S2nJM+rQJiPuWSRqrfYpZMxy1c4dZ1eyjOv4lEwBRzaGf8O2gRdERrnoXPg97obs3wVQt8S8lD0B
K+GvnR7hBCYE5FBLfVYHjGXoW141tJD2SVFCHwzhH0nycuxOB50dw1nJT1y55yF9PNwzujdvLBcv
fD+dCEIJ3iZsUDRhKa709cDWIr6fz42D6tSR30SUyFHPrX5UQ9qLxPsbVqvXesbSbpDZ3csGaYC5
+bsDglGMtisSVxf+0FTJFpAHB0AbAW9dGtISxygoY+MtlMCJIszDRYfsEpLfu6w7dcFDro1YVw8W
3v0xiw0IByAmtb/kUI+zr/qQeNk2tM8gJTZRuNiFHPdBmFpKs/J2y8L/aXGAv+ZbDtFzHps4yJxQ
q+nbMYBiBgjoeM9nC4JK1DR8xBqIrYw17qAEbSJ/5cfGfJsqDOaKO8sfa/7LqnHb6L3jSBIaUAZE
D1Zo9NxniCBzjNA/o0dO7DEHHBlCE1GvlICTCkrNqCPlYBEcNCe9/yeKHzKtqpQA7eTI4/zgD1Tm
oxl4j1kxhotDYhc0TQfJ4sZX0ZOQVblvI09530li72EY4JQafpF85I+rPwiBdnbAC2WqEI0KIsww
2Dvi3BKPKfql9nEeKHd0er5IqPTj+cf0zZaptTHPyIINFAewoHjHig78He0QZYO5i+W6ZIbyTuqu
txSyFOa2J8G28r70DaZeIVCjo50usY3F6hWL0uu8TJ1y+KG0tH13JsT051LUWJf/mn2fIhCM+Avv
ECjJy6+JT5e9Urw4WbiTesjeVlXWW69pCADwt4M8jFpbfJn+0bnlo7/Ye2lQeDEcv7Eol62xmVQA
7UkmiKaMGlTP/xlcmF6I6jyy4GzrGLdwWDEK4u4q0gfT4wgf4ap3yfg0b5gsc9BqzqPkCfiSoQ6j
cy9H48aQkMJTTDRZo3uhdBFgymHIrR1HYkn2V2z7ZSUda9bgT5g8ZUMcFZWoQ+AU+jvHPcpXwdpT
UdPWGDE4qkYCHWHtojr/e5YbDw/5oiqTJvojI+N7WI7MHYPIhj1Qgv74iIPKqhe5dcyFplBFJXyh
NmMQPVJMS5Ji1ooH+MLDVwv7DV/ByQmF/x7PS0EplpE9TP6cA+TTCAiTCkZoCOTGxBQHVsLGP1PT
ufc2lFbX5Vl4E6pibUZNy7YTrk8MMAsJ0mYPHsgBBR8/ZVtHoA+6AqtrSbr2eFJZHzVICdm6GvO5
uLr+gxpmvtBgDTRP5ek6MJQmdUNkMYTH4J4sE5FdolWDgco3b27W/lDCih+VIMOc5DhwU+KWYX4e
OwDCj+g6MjPXAzbdGH/aEzOIeGB/y2JZ85FRqoLHLQNQyfsjeA+BCh6niP5SpwyFFQDvG0IEexia
PtqeokIqlHw3O4pn4s1FhCn02ss+ZNETt1DISM7qQH29Ad9QdSNVjtBUsp+PAT0qtrO/BJ3TCrgl
03vJcS36ibYpaoInm7mZvQEIsRKxJORTKqUdkkEfQAMGwaFFyRnW7xZXRl8s0vKfgYOebj6+RMKd
+Ht1E+zkNZEMuvoGOY39Gd3rxRlsTnr5yPSTXm6qvmyskWoeqMGq9Z4syoa8QJvKLtjJuWiI+Y6j
HW2g70yxDTVYEI9zG/Ytbe8SsUl0anJ/lAlFvTtABo7BPu9NJ9YsyzleOqaDARCQxMnPedLO80PG
7TLy6XMu13fHcB/jHxANvLREesEgRJW8ZOASeChB69od3OvgGjGKqWweG7uqAF8QbWEDaZqbxHns
VpPy7rZHOI6Gtn1o30FQVcYKZdp9LwPIMaei3ff+wWTqQBjEpCoZKFXC62iKyj9cFhI4JQbZ1BFs
udMtOQpXnD4nrhLacrd+mWMcIKo1zeDa6upARq/qJ+NaVXzlzpxh0BUll24mEcoFRyVlNyD6nXvB
Ys7UPIYW376HHhu32PQ4JFfu6NzH/7sbg/5AlEYmuJA8WQjFgQo+gVSO3kDWBjc8Ej162F986Nqy
/1oCGEHJDjXomJ685Oc3kaJPMGnZcvNN4+273XkWxMIAxXq731fsoEU6D3/U2lyAuBlPinXmFjxm
P+aBrcwBy7P5wWIKFbJMc5jU4Vr1cYAugK1uSmuWweKIdRn3w+69fMkamKx0vmF77maM0icxUk8G
XAlrV2CQEpem2iKhsBU6C/Z7n4kVbvpi8COyicZDGU0igY5LX2MCPOO55w7Dnwf6mkrt7QeSK771
mVZOS40X4dAyyIqRA7LMRMaDyg19J4BG3JXUccEznUnsy3cS8wM3FrQu712A7c68p2pyAc2zIf5r
/FgRRrla94HceJaDVLCNo+EVY7ln/hLLjmmYDxy03saYCrDb4s30ctarGbfPCqRNloMTp4tS4+a2
NKv6qUNmvXmaCHCZ22z4y6lCQgIZt6fRCVyRTP4SBrxm5tCchRjMGV9X4Y5OQdPgYJxreaoHyiXC
k8YFNSdeHJOsbpL1dLeTylcDF2TutCAC7wYAHlFnUgc/ok2gcAKWifZ7f1fwSDzFhQsJXJunA1oN
aSWiDw3c7iLCz7vseXNdVN0S/EPAJrlhr/GBOqvGwhncsnzwKSYPS8/deKxm+Ij5IneHo57kI9qr
BxMye478hms1okAL4My2AW953KjlUiDmQPomCzXK6fZ41BsoOXvwjMp6tprKqT3cj3K0U1MCr+CC
wRBMgT1fYmLEsth/5I+j1jwUU8MfEXWwzSmOts1aoO6yZRGHn+HbrgqORLURePeAaQoUrQEVvLtI
x0EUzbgBQDvqY/rC9BNu9nJnB4WcZlxFeke3PYkLsRwl6I2CyM75h1UxwWoE8oV6DmxF60a9qdXC
tTl+18myrNYVWTDaN3T+6aFtZ1zLwa69xszsGEOEKxyQ2DDsadrTr92uUGX/1UhdqekPkiFNTY1C
ivM2Ns0AGYqqp8fkVKJbKQjzfuM9Cq7p3ojo/1oH6Gvfe6fBvxmftans6F8BC1g926vKgShc7UAc
RwJmi4JdzXNWpcAb/KWNmtsF9HvOHj44a9eHbCJXgdN6XAsCpSbAi7pRAfKqmv9g0YqaX4M25NVQ
w54zu0culSUQgL97cX22580bAIBGZ1SyY+vcdjp/xQm6f9ttBQ07liVhIPBKYb0/OssH4x5ADbf7
QshLCA86CZinZcPmTPfU311FjdfRH9xCc8RG+P/erySsdNPJfOU/wjyGgw+Ic+BGe/hLQsVJdN+M
DOeMtWiP0VLhySkY1WfuKHoog8rWIM1bHfBaFRk/kpmwelHYvfKDdvUxcfegYZ94hXCddykFjOVe
9tNqxDlMsPL2PtirXj/AZ1yUQ3cLSormLuiQDxrWNnvoLhsrqCZpRcLUeTEwq+G1JIsT+a72Yr8x
CPsTVlw0Oby31JJInPMgyTYBOrOX+es/0DJprVn2FqhJtHktrrsWt59PZPWgESJ57Wsim1hYzpQb
e8hcB879L1Plj1OxhllfQHlBdckH7HuzxGbAnrMRsYQywAWlII9JX3ljXDspA7/cShWpCALcZq1R
89+swClBivynRv0pwRN0WeeEVIxzjmwAWyJUOBAXyWUWmnbqKsHWutzUPoFJBgdZKLEHKfvSL3nM
5kiTdbgVpkiJRxtw+uTCfbYOcIAinVW0cPE9uT93TN58G9X0wIt8kV4qV/cqlJ3v/xVfP/mkYvqN
WINTCnc/2Gj/mqcEcvU8oPEweSN+l32/JWRrIHVwhPCiFWB6dDikfCEbPP3d0UUoLzJBMIuwhp+O
txaKLezA/S6YPfApn+Wo+34QgZlJuOz6EMaR8AyCK9l3bJlEmPkILn3byEnhctLklyOQF+y3bhZg
JjC244wK6mhdp3Rfoyjx/mAVj7odEMk15Zsz+maz0TqYUUB89Pg8pg9JBBjjqRWSQMVR5MRk8txf
T+2LjqrW9d6lvktm+oPFz/a//wVs85d5uEANpT81NLz5oZgGZ/7PA9dLS+z7h0NVei1zfMvE/kIw
SdBnC6Preidl12j+UKDTdOwIJ0S7Ce+g88iJChAnTivEzrJapNT4JhNa0BOP0SRMw6hgwAowbLND
mciqWziY7zrkr02G1J1/XAObHb80WsO8ECHg7uLTyMhB1a8FPU+bw/xgRmhrKwdHWbX5WUiI5DAs
Od1MwMVf9JVDrqDaBVdFkUMIbGNyvJtaUWDClzIPAzvtx6jgg2S7LI8CaYseOHQf5MTwMzyGRrQA
X9lzM/SnRIHgj1HSW7WIAY5VsJeubpd3mWcxv6EZ03tjAEsd99uKqlcQfgElMh+o9/H+0lS8mbga
qKY3ucgwl2q1m2I0E4Ywpd/hjGWCcd2OhtnrjogMizQCOtKwo2A1IYwN8oxo/TozOkuqceqqYv4E
oIBmy+sQE7sNhNzeUOlEKO0oF0t9yOfeIMjgaQMBOhfvCdS5yAKzBZb21nDIARQCD8uyNoUtclgx
+dAEX4G+7vCImL1kH95pKqrGiQUU/nL0hZNefYgekc4VgqgIaoLCObrjP8oqM4Ss5evQ6jDkeWJe
VTfttWnvwpvnlSXjWIDBk2MqQkJoCmDF0PyMqJ5200v2yoMqR16W+KpJbIH6JqeB4/q2wJw7VdO4
TFjTpFB7Vejbj5RT681j9lV87j/uESKz0Kp9L6wWP7GXnaunStmtqHjEMGvzCegkXnrJm7Uu4obx
n9BSM1Zf1uDBk8VacoBpPPoh3aH3Ntgmfsjy85CMRlJDfrQsUsUtswMpVRsFC1Y+Stbln1Ntc228
3PsKOLD1ePfBIB3ABSGii4umjKMLnVRg6oRrmXDxm5/A/+Hx2tr9D/hBh/Y12qpaPF/+yuSFNO1C
y0tfA67y0JJXDsadYV+Jx5xA2p8og9SV8uqikz4ocNk3XQ+swKXz1jG/xaOpW3MzSvNE5GkOullT
roxOdxq6H74zBvEDzkLykO4Ptz9F6JphKdPcRQlpIzoQBSIkTdhrqG/w48opZEQgIB8dwamyZBPm
3dEZFIOYboOgnXebsXEFihzhos3ayLcLGmgVWfnGI1PR+JX1HGePd8GSvDIysv4kO/bUyxiDAR6Z
7flmCq2wPiTVwkRXGOg4eH+/fVJUzhYDDwAsl2hZPB5j4/kRWygUlSMclLmgIxjQmW86mVdo8dzd
1uG8RNMxv6gGSvbfi3YukQ83BDMnC7+GAKdef0dpdpFnLBWcC6a3R3tUGGHncawYjJK+PQ23aiPb
PfZ1rN5PCQjvCpSZ7iDG9mftPFj6tebcUVhWSFD6J6sn6azYs1w7CHh7Ttmr+pOrNmuw889RX4w4
v0elGqzrkHY7bW8IXIRzNkSEzJaPdFMfFgB5hh92bnlwhAkO3n81SXZ5bXnuNiCfkXEKwNhPuhRW
WHwAFwsagyEwJpu7EOsyXLbsh3TacZjbmyZNWSwOqrCq4lpoaCoGfmgyDL6c/LC0fpV8lPopP5wo
8TluOqOM4C5UxeDXABDaia4ngKZruc97mz2PKhUFuR7C6b7QW7dMxX9cWdcDc2AYwGvGTBS9Xp0/
0jFeQT/sveuweAt/yiThqAN558es87P3/4TZ3GzSwpb+nxuZr901RswTu5/Wp05d5wk9vA3bxz03
JGJMuw6tUG+cbxCX/lIZxUfcH37KemZr52omQQ2dA2E4aJ5F7p86VVWs3Hb1O8OzhhTEONMhTXHQ
3bFlgC/CkE/GiGhERwkGFPLl/vARN1ZiMjM30zdMYTb6QvqDVN3FE7mzwMIxyx/xKN49PrJsREqy
nnSLjdBRGikfEeQoHw55RI9s2tYwOhxeX7oIjuvmNdz50A4ScSCAyGh9ZDN0REIwJFTmYRf3B5KQ
KqJIXeeyC04vW3CQsaE93TgqgLFVLYSeTu/xV3Y0d69uHkV3fhSrQuD2ngxiP26gzjJCocbEGAsz
+siDrdsq8bppUx9olc8wPk0f3JNwPlme871KIkNAlX6Hb50vDMTbKDfH9otkBcaW7wvkUC82A0UL
7bo783jzZdaiIwYwQKCdZqYrBCy2gw9+UXU5mVe3PQrAtZuNUOWGy5AnQZcQ5WBq5KKHR8NYLora
KoeYV7bhfPK7nL9CnMulJDhG8z0PgaJ+JBOHatsUE6DPsfkMahvToh7A8K4IiC20zxnsC+2vd5V0
jry/T1xgfSUa7L4gnKXS0QQloy43rnzGGJXEu1Ehz7zOsyRdJGiV4+IxF2oo5yybM3/p0eR5geKk
gw4jsUL5g8l6fL6/t92Z6Fr4n+5U52ym2hxmp1+XNkcCJZw7jY7q5M629ZaJ8q3Ptd/9RZeq/ohf
3F4M3GRM1ZLLUZAqB0c9vajibyVNXQrOLK8AtKBHS1kuWZoWBeJLdzts/wLW0eGnJBvDSJsUqTxG
CmCKZ4NVqWEsK4cyZ8LTBbOQsFW65GL73e047WdLg+7sA+Isr1Of/Z84gJswBz8P/IAC1hiJweEH
SxWG096B3D5qwbgZZJNx9FPA3fFwcUjhCUj0VtDmcHvBtlpWkE2JwhX7MuGIURUGG4peoWK6jXqh
ll5/Ob4hWd/sPtou3XU7fBlpUMKD6kr68j3nkyg34JwAVvWjSV2v2IaAiLhcXZAL51dkiQDt/ka2
ar9xNLXYLbKCMXQ4nDKgwh7vkOrYCDOrrtFpmmFt60kCroojJaYFAnySAuxY72xK/5Gon5oUfNdG
dRUS0IKV7MNjVOsdWuUuEZC+ITQtdDwX7E5P1qibyDoGKBJUk4TnqVAAmtszRQ+sMnoqpXWwt/Bx
ST+HVEzQQmtZhnRtFlI3ETfaMbgVPAvcfXRXmkKk1rHOfIdiupJrr2u4wDiwVfc3OPYNVGq2Hi+T
AMXpbi+NiWA9/Cu9KpC8G/pKU5cr2xCuozMGrrCqbloUPUPXT+uRW3oILVOEJMSRfspdo76CPYM+
W/DJFsxquj155uU7a/1wQ10JWNZYU1Oq2FenjxHFVxde3oXRQm41qBMa4dWOufFY/KTkE4cSsur5
Gq06VTwiKhCpTyJH0tCs/1Xfs8jMZX3P01x+k76HJfONK+BVkTfu63CH7j2AdVZJAl1WljFufE4D
dGUavdZjpPz2pvj840M9kDBSREr9+x/WXBzvuQ3C+bWJQzU5NpuaDZhry5Qwyxp03lEM+dmop+7K
g6CIWlaF9ZHTQybT0NR1wTRh/wVNUGDWIfPX3ZRMS4WnSZvaAOEa5fZeY8kwqdCEzuYUadqXa6W3
bIwLsmLk50PXaljPQI0NAOorwhOerODMYL0TuixSP4Ugs0qRl/doeo8IcaRRtOhFX6D48nN6fIH4
0fKbiyGcgIWfNdLW/QOndaHVg7LPmk6x4GmWHhDoTRYjAXPl8ZmsFwCtljxdR7gTi5LPxBn06yi1
lYMhTn7v6ufIV4xoN6WnGWVdXtKzi0kyBySTRYY7IAjDzX75W8fML3xa2xVO/Y9LFTwEKH22lgME
tIFqSt1lyt2uVcIrk5NlXVxc3syALEm07dIPRGQ6/DTLDTJ5voV9VSArgGYM7+2NtaSwS7ihcLFx
yx8N7I/T/AR9udKdz7xym7iUW6+hQeMYq8s9iEvjcTu0j5CGdfh1GYIbjjG+hVrTt0sPkMjwI/WF
QP4xrdOYp74zFkoZPDXkoiOBcw1ujJ+UkFVAVSeOBJwFbD39gJc0mUYM94BSS2axnlJiAqNoGlKJ
osJjo2l/VSZR2mXrXYNlL9NMboRz+hmfw6dErpE07NxDJNpMDaO2G8HXMBJP15Qmlz2EgSUpsqoV
tlHAYQB3HrmYXRvXMKIzxCC/+VeExjccHX67b6XP1U/Ns5EM6MRjYfC1ku9Xkg6HAYsdBkZesDDh
y/aqpNWiPIBUaSYQBg+VOaA/S4ryvFe7OeO8AG+OkHw/Pl31RWK+Lb2HJYJB0hJpL1cX4ySm52l1
IRnucZyU5I0h9c5P1uSm5agZMXcK+60flgOj48XbtJDcHTqJp3oPZw9puUKptXi8mSiC9qijBY1v
VpJadUW6InV8alK5Jv1KNNd4LDiC1mBWYs+uEWwmRgkP66YGMNCK7FNcb18rhZmIdNq8rFq03064
teueuAOMSeA1nTm8I3wbPrzpIvjZKN591L+WNfQgGUSctI71sV6fg6PtYfJPsMDsIh7OmOAaOSUc
l3tLAyRAhekfOxHAOEDqwRHB3LI7LtxgFA3tWXKxES0ugD8CxL2BF+iCRUVr0Z70mUlfDJ5H1pDN
6Wmzyv+LrVNHCzyOGdURMfurXbl8b16iHH1l5uL+zucZB160GNG8nduNI7j9rib0FNxY7AlM6y/o
TfPpNWj7yDvv3lusa0C7Q7wpX8uqfe5M+35qkcBdY8vtNYIgYC/UVwULI2vsKj0Wvvx1mT1y4aNz
hfdNWFoPe/8YPetlFfC/MYdgwfg7W7vBlGfSP8xdv72WB8bruZz/fWg43qd0Q+DLFd5C2C6r4jpL
lUixuZaxwJmUBmymy/d3mu7kmI/hW35pQ5RSlMEzOPcROdHpB+tpM8fDPc68AIfXd76k51sLKEwL
bIhSdrh8XcKXFo3lPhPZGszJM8CzEsIRxzcdtjgY4tDmEHw0JsB+R8gRTYPsG6B1GCWuxYpxQjWq
f2a+4h+43ANxoT1aCRSKckWS3fddQfD3joLrG7xSFa0UuDVzBhxS0Q5lkTPgwT7YP0rfMjtBgmG2
wPVDoTXq190JiP0XKuSFfiz4XvehrifaUQDJR50RmUFGzpbyPsNsJrisAR8MlQWpJ+orS4fgh+sI
lEvXxBCMrf2jvLVofM0xafqWxpNfGS85SLBwhfxS8UqtmzkPuhn+h161OkGsKZCjUCTEGS8oiTei
H10lvlTXVrm/VDjpkDkOLGqHLOVnGa7hA7HtTqveK7a8y4YTUblF49rypSqmq8r9hum3mYvCo+BR
h2r5Q1w0vYJ9UuVMufUNlkGsD4iHQ6na0sskzo7DUBpb8LRohzzQVaQHY+Iv3xgMQB8J8S+yAyHO
vn1povMXwRUEtID/Ph/8zTY0PgNHwIQ+GcZPwhLl4ZAUn1jBRDq+zbt7iGQ5m0gp3Y6vD3KsR5s4
rzNklD4J7ibCl3b74WHZYl/bVhaHzCILj3ar1ehLneWu+RYCbhfITgSUdA8BL7FpuUkOVaSY6IS2
3h8ruba7/AtspN0aU5r3tuo3jzs/CkYIh0dLeR1tQ57kazMSGG0F1fsX0ubQtKyHGoJnTFgiCMlp
JUuOccZKzwyKhIRAY104Z1YNr55zbfMyxAVwpcVnF43Znwag6MDKTaBe5nGT87qTT/el6O0NxS7h
f0tgdTLlE/qUIPEZDcCjC31pJUQ9U0rGPR/rPNNSYwBsi0MYRymY3kG14z5htdhesgTfH7DVs0xr
pHxDxAzSTpNgrZn1Zd2GJStiiEmgIR3jxB0vE0BO/dGoNPtHQbJQrlUEL2RBTz4wuN+5oqoqi9Ht
NgFIdpjoo93p9k0CDHvyhCCv1/t4SaSJSJRqdensB3wMknViWrhr15/8GAHZBxUIVMk0B3Ukt6OF
MJ0svzdDcNKyeC2bCx2ifHpZt8I07KNFr6SqWyNU6Qp4FVsSWsCwUQP6QLH+wWN5VXKiITkUCL6j
8kFkbydpZOW91c117rCHi7IpvaYOObSH+907k0AOuVsdpK5yexwp0W9WtI1J8pR+VpAGCBgpY3E9
iwVWXVTQhq7gsh7EYn+gLqpqlsA76czClBZhXbwgPjq/Gjx5fLS9oN7C2m34mMupokVjRS0Xe1Xa
+lOj65fe3UYM4CdiIOyagotlT+HHPIBZqQ58HACXoJqhy5Y0R2moDUHfDzIZ2q/3+PVCRX+TLc84
HzyGKrLUjSyemnZoXuGOOIxjnjUbVXr2r547hE1kEwGdrZ6OT9RFi5+CWGmvozjOVrA0L3xRD6wU
q2bdisWuNICsyGP6pUoPhGWkKQYeQBYSSbQpbFOKT+RgracNxa5RBoJwJx7SivW3xgWBRe1Zoggb
x53YFFhNOwc/bURy6rI/0f+zs1XsFy6oWj4mH++M2Q6QeBdQY3GHUF3DqjuC6D9ey3Uo/IwJkUBU
I4e+NPSwHiNdgfV/K7tv5zPEyV6gQqN0QxJ54jdhIV8WYGO0FWCbuBH9nHGJqOD4h5ResjEoU0xP
xa4j0Imw/tEH5msPpjBPx8VGwGrJr5IunCKlsToh+Ly8IY1pITvbszhmSgbYCOe037ysHEPHMLno
xIPXAV5sSzcBqWZ215LpsKbsPMimztZpwZy92FVZXkJcv+W1ImMcUKxWN5rG1ZhhgquHb7mZg7BC
5Rh1xgy3da7+1SmnGFkwpMsP1J5HddBb3gmDwTf5PHKQ+mYRxKu/fv15cdRWTJoPO7mMAIL4Pfz8
GAEbY+AFYLedRtYh2GL+9e2EDhEynSmGHBdryevmmeIGQIssdsPZoCtkPT+P/qCdGNESIEcojk2A
8s35DWFmO9p48j46ITpqVwRa3aUQZhVnHnuMNsxwJ267l9J4bQLjngSZWD8f2WBDdZg3MXPNRzb/
WWslRxcL11CA8kh97rP5EGSKmYzOEUlXMqG18yoy2gLA65rUzaihrw06Bq4H37w6/EjD0aYIu7Cc
hnIvx/GMCuchV7C3Y2ALm5i/5nZX76VyHu8RQnUJw5xbGMwdj5tNJhIXJtEUK59FRg6iKPjvBawM
jeaj5bX+R/vf7v1WVlJAHiUQb3kNE3mCjrYimSktSbPY43KDF4FRf5irQeTaj0Vc7rGKZzl/e+lu
bSyobfWuxWGaCqbSDg/Vtg/l0vAbg6CGiirR7Emj4CWL+3LaiOMofwzugzwrvNdM/D7yMiCbFE9p
/R5ymsKbYfEx/t7b20lVuUDVoZOVBCWt4mZ0xt4CNAT8YweklEKSPZ5HHRo8zyJIVu4tTz2X1rC5
yoCJK1HzRenVu48u58jpPBEvCEid5iaANvic/TtDbS2GayEZ13ld1AaHYFYN02VqPJCI9p6LNZVy
4sSCjnIRllQSSQ0lAbvYKM7YktzraaO/mhqeyY0bF+ael58xgznbgSp+qRI/Cb4GY+8L3lFORtRR
3zEqH2eFX813kc5zvGHGWv4vlhWXwxtMXz5O59dWSair9x48mlm5F7UFBOzXG7FLdAGjKcaSDlF6
7wXa6Gef7jtZTrI5+jY+4e+o+Hvk9nbBFS7b/N3IB8/NB0HaPTp16Dhnzn6r1iMgKNPYIGMesSsc
e6L3gVbB7YIGWOOse9Nn1UStk3c75+abk8PAKKyIveddeX0jrF8PLEvym9t5Ye8dr/TEcBVsB/ZM
fshC14qCmps27wCIwtHx4iR/F7+kxoJYNyYAa4U4VMda0b4ZnBG7rn8nEr0lu0QwhQkJrD5ESqIz
oi9Ds0lUmPCr1jI2tlfAyWsXy8I5INdryU9TUL/V0DQIOnBM/avoZ9kTt4xqsnwAX4Y6Qhvh5HPh
9cG7atKmklP2cjN32ceo4VuIy+Ys/w6S0rY4/C+HIRyWOPC2z2CNSdUyV64wLTdESYXz3+ZxEUYu
1fHRK9FQHVW/nqCXxbwEaU6yU66pFSu3twpJW4WZFAov3L8KAipGnzJ65bhKtpj1X/ugIocdtMUX
sHyToKu0pwt8/ByMjg+/5W3xFBpyLfsfN5TCGuEhGOV1Sirco9SvVE4NuCEHwhrVbG1SMM0qi8KK
RXEAm1yFGwBrms0LXgS6bKNUSDFeH+cAKdox8Px76rT0ouyDYFIFvEFw9bf9h13YLwutpgyGqz4u
DxbcBR5Xjs8G7iyH1oWWzKn9l2f0jjq3oNLU2mc2aYa8gn2OfssZmkcsUy18pnuxnxUt59St8wpr
9lNhUQJH14T1YJPayjGcQsXY8pYDTXfklhFe9iOAm91JarTf07GVQbF+swXOoK1zIeSeZc1eD/Al
nh/k0t5fwchfgRfXShfTgy+x+3UK5eKxwbfLBtOX1ooUEVqy/Aj0YECIy+HxFzSrkEoHz5X0atE9
xX0mXFR5y7cQYC/2U5DFgqOKjJi5xZM+o4HG5mg7Yx2qm1CDUlFjINsHG4TjvT5rhSIo/MRsqHzb
b7H4mhDzWES0bKzoHPgPLOFps1iAsK0fE2L9lNfyIL1/E4N+zyo+Bb2pbVTcEo28AqR/1/ppgdCD
a2kqriIavH8Mju+4BXtarNCqxHYTFZB5OFRegQr4DPyITL1eIYoa4w2GSs71ghNd3R9weKfL367M
efiehn1Roj8l98DU7Af0IbGpL+WUs21y4ygQQfi5D1D0itwIhgmuTLsOCRhSZKhof8wK0ZUFuKmc
LrJw5NpYunPZdh05xQeSfHE6p8FPY7XFnu9xAajzBC/WQOibF3K/10Uw2kufqJ6rW5Hry8SEomLg
WpBnKCrbynWflxrHMCJHkv2zlDPAoIs9Sk1CLYbJrUcoPYrh316qCbUWv+gpGnvXCbGIam/p+doZ
ReAdGJy1juJb4PVMWc2/2ZjMRT7a1FteHPRrj2WRfCxSkCGBOnBAMrwUijHm6+Jh1+Aagp9GrsCM
Zc+TUoT874APCsG05yj7qCmU0AVFy72+z5yyKQ1YQ0KbvfHl2hHLeCj/n+dLjyk38XnYNiuksC4k
9n/zdmqIk0fty+TiSGuXBg8pEKMjhmsQMyo9OfRYVbY9sasZcN/T7jKsiikdmTJK36J6QDweVcIc
7tIIoLskqsIAsm2ZTvjBiy40WHiNN9HLEO80/nC4JPF5cy53DbM9aa2I5teqBSJKONenPRSMweII
3Fh2J1Z4sk48OTkROcbPCAL788zR6wTMepWGjNntBdmfren2DrcxDemn5R5WK/NWj55hIoJyHlI0
ORqk8xys+y6psTpAyhX+YWK6K9GRCecDXW7DeeOXBLyPKDIhv/MIpnLpo735uWCCvnn90FbMeA+Q
UlEZRQziTPAWC/f9fPNRFU8wB8tSK8zC/OeQI2hnzCEypxxmjQ9mORCqqKV76xmSn+exD3RfBiU8
nyWwptSBBPS+IkIlGKOKXvSb1uE5u0Mr2+htnKM08M3f24geReVxpN7r6DMWV6h1CEEZumTD9dQj
naVM2SoWE0nGiURqDascgn3DMjiSaAJGz6eQM+UZn2RW1KwV/DgLtuWQzFdo4akwqx84XpGM2kM1
1R6M4ndGB3G1di1PuRY9eyn5eVpFsN/MEw4X4BnIbSDqdNK06HqMGV4MWUwWskHcif9KEiAQ7Ppt
8Rok/Cy/r2ulRMUQFXReWs4ssvXZ7kssgDqwIlAh2kfW8dhldQRd61JrpDfKfkL9asN2OqD7WUzM
9w4/XqL+jdBMuss06EXbj3j32/MtvXKNR6gDiqd9PAu386rN+Oqm/ssKDkmmD/+BliPGl/fYnDV+
F2ZtU19jjnW1Kl71tIcMmCaK/5YlvcdARloCSdGGOMZDP9Xn76Jnpi9zERMmukWUqxzzbmp75hiC
Zh1E5k1oq0ZsBa20wo8OkZUCHmZNXw9TvXFyc78Am9GBgSaN7tJSh6808J//lXSvjEHW8kXDFyrK
VjcL/heOr4fQqX8vwrak8jxuOgnscwJTeTINHMXu2jNstpOG+9ybLRp0o7pV88Dc19HJjKeuCvD2
tL+f2QhMc1OFBYpv7CNzEo0aoh26TSWCQI0Sh9OzLgD5sr5vwXErpSng1kYZhk9v0P7gxbuSsnYn
y3/J5hAXWyCpfwMm1BwCblAsfekg/uzfYNv1q+qJAA3cntc9Z0IM26Tsj5PhHgukFU7Eog6ntawK
/8aGyZ33CxoL5AQRbJRnux3iCn27mReSbxyZjIwfh6eqxa3wvSJSIH9nyFgSkoTfw86tvzKlaqAJ
lNVatmNjKCq46SAWzeqk+huq+JDZ3LMCh8MVc2mnCke5X96ZU1lKNf4/6M0K00njkNiGaHfxpzvv
IaaTcuRGo+wEZX0h7nlVIBEcgw9SPqss3bDgeV51EUuVQw5r7YFkxnUH8v67xRYORbSGYgTfz4Jg
XAVePgkvazCw6/OTSseioMH1AR93NfztjAuL0QqIPiRqHz2pxWh/1k5a9FSFtQxdlJ9tOGCmCCqo
pEMUrnswaWE/01uHDqIFZe2wWuB63WUUrBbVTmROIS3cB7x6x752/TOcJH42wYNnFPjk9hoAwMGo
OpNlnc40cEyNwqqNl1GsixBAqzw5NaE7P15kfYGUL5Vlqx6f8iwPVF4BV4fqC3w8y1KsHOuVZiNb
sXSkd5jcGlTgH625TkgnRGcgPMdKjc70WeiRjYRBQORFYZcPg/PlW+/Ic2LWQnRuyGxfG+z3f61g
nP6Juc+rzVZxKl8drf8wR6twU6m2Bo6DaF8VHLw3aKizD+W/rpTfV/VBw40OqSdF9vtIX0dOds3r
8WEFu3P+t4CimjMJI/sKjM3FXEK4KR+uYeOMbleWytbLw5EcpkA1qEsKGqv2qyGMnmkkPpK65rA4
0domhrxJ+ICgydkYxQn8e+MEbCnW8W4AlODnHGRkCGf7r1LkRxLr5DRZjcpRsawHyppMrnGnHoIM
F024M3QQNbGFkszKacv7o3a6k2UHDT4N5CtSeqGuwJEqYWzQ2rZxZa5foCxv5gOETD+Pvdkt8Sc8
Ox87LzGHV7FkMEwqc1DAt4YGaSTKGak5CnMgHQKB8MsVLe+xfA0kSvzswE6an5n21Y2YNFBinfcd
52xYkzTBWLBZf3j5Su/yROFa1AYc3/Vr5IF4swRQdwJFsyfs/lXt9IfcGsGHDW3P39nYgKOmFvyS
Vqrx5zsGOOyp2qbyTRydwdtLcgg0mUqqyRgMbVwGYD8puxVlYjoXZZum7b4sok3/RECE2yiyVsJO
3IRFV3Nd5+gTo4SzGjz+Iww0Z/GJxiuYtvpsJbYjhpzPNcPrqczNtlbbdeqqzKX4ipn82M2RgcGS
Xx8C/DRaow5l79UxwwMaHoqmSDltbhX0QQKfTmxhc0ukoBVjje7P3eSxaun8Rm/Azsd11o1b06qH
1qQjzn9xqGi2tNsTiu3sZDMB4w0rdyWL1gqrF8VpHwpWtBm5XyO/8M3Xa4iECvOTQb+8FTj+AiuN
o+7Pj79+eEeqNeN67PNtJ/+kjEmQBv6y4rFaLnYeC38GuRL2yPsgeW6u6XhKUTA8uxYsgWH0gmUw
obD6QAepnfYlYyXo+9r/nx5a3io3N/ksRUfCzYhulqdAa0HlN/YwWVE26bkecsJruaExA6oefCxZ
d0I3wX+nT9MbHtpzXVwjkb5F+8d+ilyS7pM/oiTa7DWbQoe8/Xf528vQ1m8nnlDOEQw2R7YXzgN5
g7d43i4pCEyXVMZ9dsTydlUuMdWh8CBMx+a4vpxjLxBOq/mAJ/3bZF1JFmC2Umfs0Kskl+qiYtHv
Z9qEMGqPX0NHoI8INRH6L1mFWThQxSycqCvS6GSkPNudGLfhp7LM0k4T5xULpFr2eFFeJQQLW/dl
s1EXnH8Fa2Kw47MOSaiqw4yyNh+pQmqwaoQJrT1tAq9cRO4ykVr+ccRsD25vRpBBSOrfSIs15qPz
EGY/fG0hGFmFXqcn28wGEaQslnGVTR4RPtYe4IiHXb0QG1ZwNVcRer6v3tyIQvMIHHo2x857wDbU
Ne7vS/073EsgANiSzEmkJyy6CddF/yUnq1t1qGBfIDo8V35ooBamSe09e18246ye1ny0XYrjkzDX
vtacG5Q1Ojsd3OYQ+0wJG8wk9QnFs+skB5MtlvE1qeU7coa659zK5HoOtOuKHZ8YoBkmZNVcA1E8
QoBx5GJ79KkNH5SMNE4XuUuW0KPzy92xbkdeg1uQvBPrlE0OtfjuRs9TN186fdXZIf9UKrVLNcyx
EYHbJtWRM8XpMUu4MUyB/AemH/PcrmtWOrdPamLhV0YLMdQOdUjkKSrX+qofawDEEIGEjSWSiyk6
Ftq389Aqt+EVO6BvB8/l5CAmDVEMNHMvRJo4+yU0eZjvRnecflIOrKjLG1D2Gsoo3/KtDS4ba1iV
MdbN2IuqOlXzjfOwsHvhRDeUJyrbBgQ772bX8Q5FnOM9/hBlVVS7Eksh7Fwac5OR2PG+wB1l3V+y
/YgRKFO+Q7bgT92MPuZCSsUTUBqX5XPm8H+shvnG/RwUYLS/Drambwm7p4BuZC/kxL0+MOb2RfYc
6StkMRGIFldLY2iE9mus5W1koUPPO5DzkPsZmEwx/VmcN5g2zyLZzTJhdDH8pmpcYsc5oGaL4XKy
IZ7+5lreFJqaUC3qrOdyv2BSGYG6bhaGlbhC0GW+DAK6cNnBvPSnmS9pgqwO3Y7i26VOdt5l52ks
9gJ3iiGG39PG8oFDbryGekgLxrV1sVc19Nges1hWp9VUeUpwXO4JGZjpju+FvGyi6OrW1L3pUvQg
oPgcZQjdQJeggRuyyrcAlhYYK+bzgrI/JifQyieplB83Pr2SjMIqRT9ozqjSEfGzwiZxUHArl1Md
hxVGpomY5w2z6GqyTjMitmOqGUFjTSsYwfJCJtWUhtPd1DxNidr1HU1t/ckqHyMn1gZEJavAGjt7
FgCoqffGmKmT5hfIV4FmIE/JKXeyI0eCfT6xPdhxpdDgkgtTx2vEGdUs448TBtswzLLfgy6R2QR2
7vuU89dfsJYZlDQMvJMILgLodgqGqlC+ZvUNTPhd01VZ1lPVxw48MeYEqOJj6xBDEMs1lC36cb6f
wxbQb3ao/zDHV6W4LU9i4XEYVIuhmyVtWiVzQgc3fa+nfJNzkS/ZNLqUh2O0D3ktsdg/sVMuRoef
emCvtXguIxW+Au0S8BMVXh6kMn6aVizdGSRW5v0/YD6mwthPRa/Zj5OmiQlVszu5YfSFROQILiTN
P4fwTqaYQ1KObYmZEMJ+L512fpTE7o01fNsLlC0cGhjiD8QQsjN6335E1mNSfLKJmLoov3Bg0kAM
thRmv9TAEWFCiVnFJ4TW2r5SGp0vhFcBZkn1htBrLD0P/ALTKBexgCDPRuy5l8w98F0g3xB6JZvP
7Ua/KQiC7S6FJq8BNlGeEmH0ZwNPTgTlve3/My6vELQjJ8qWHa85rs21urYOIMrPhDrtn0MIi8Ob
dWgRd8BAyqOUrHkTIbMa36kL84NtK2sUyVVTdXB+zjHgK7UXYZhK4NK6Hqx1z5FE9KHgGqT80tB3
nbXNdCoe4m7wRdB1OUYhPnnUn1mwEj+2fqZPTiZ0G2C9yQ9rMgbf5GatVsAl5kSgav+fCJogeWN8
UinvuaU83GB+irL5VZSH0Jd3YTmcN7YjHoQ5a8I1bn6CdVC+xA8l6kDplKSbnXycWIkqMfnhKVsI
wdqn9V9m5J1kh2CdjaHIyyq/l9BlrxaSI4DKtS11YN9g8G9ohABljMvvvNLbLpHHJegK8/ohzBu9
XCC87UZWm0CpiseF2x2TVW5mzIjqiJ+fvVGSzb0dh1x/5dSiwHtjIdoPFHI6io7UWO2mCEJHiIYG
JBemxVs7Q9yun00U5qHQRtYTyDSeDx+zlcItU6C9M2noyWGYNobp4iD0TkTTEIMl1C52qEVyH7Tm
kUuHHZVjM49xTWGgFOciu69CGAjVymFVaL2UCXU7P2tv+d8URv9q2q0cJtdhpVqh2lwyiwLGlL3d
hPMhViH0+/M1EcK7BNOqZc2kplIlsqaqctMHFW6JDYUNFqwmAbGNTKEu/pYm4mFHswsF3Nr4DOrp
SOrjEENSFIQWcQRLy8Y2KKWPQTk2vMXVqSQcwhVlu0mUFqfcw+uK/FQbRkyiC7Grxz9zCzsTzJy/
SxiOsQsaQ3GCFOzPoRQIYeRzJ+cKQEHFQT/pjXz4JsdhCx32BM+yq40YbErJFyWSE/xV75B51XK8
qwXRyqlV3K40ZoTPjGw4iIfwfDYfwpoKi8j+GW6g7fuDvanhbyF1qnarqAC1J3puqF0MzjLU4rKF
X8hY4JAe4TgU8zapa9cubjTVz2fWEJ/hvipKftKS3OWZeQ3umo8vfOfFv/pNGr1AlPpNztfE0dId
LcSRwt+1nJ+IQSm8Dwh7j3qOxN305rNDn0kcLCchuAItbXvP3dQr8C5ZriOBVlezw/XrWbASViJi
26W+2ocUk7IyiYbFHmvcWdjHahPl14kyT0ogXHc3dizD3Y0LHYOCMU9xg4zRJ9Lp4qiMOUnGgR+R
RPvvmq49fTVF+KkzOI3HxdyP7Xc47EtCb8Aob+f4WHzsNuKws+f+idx4uy4EeNKh2JxrX4MVK8md
MxlaSh9z3pJuYeinVLkKr/6X1ItsRq1kKpMOIQY5sFpuCZqsYcO5diWEgSDULEIViBIlBdQ5g6LR
lNc4lYzrXOD1vQ8clNRXO4bMJL2qp6SpqOZ7qiHV3tZA7zQ1qqffI/Oe4MorcnOWU9cbsTC+uNOa
bLv9eMYlI2FelLa2C7kGIuWVivht6/55Xf81RaohTlqsPMcI5QR2JhjIdAF5ADjRGASRr9aJDNaB
FtdCY8M/6LtwDBoh+0Bw3uk4agB7jH054jjovFA7XLoebiuYEDM1KhFOTT/NRQOJLhENBno27+WJ
9uOU+KvoDHQNqQeVlHI9L27MjPi8jU6N/intqhOqjH3+8Qu5KRrksDP4cOGLZ1Dc8Rbfx2/v1fH7
1EJ0xv2yfLPyggT8Pk07+Kk1/hE+PAaYcPdA6O54AH5eBuWv6I7bSetCQlfDppeCFdSYK28QCuPy
jwTDLCgojlAKIGeqyjBTGt2ALWQQ0axwwRIaLe6jBSkBlD9sKIXmzUOfQpEsu2+5jLA9mSuctTS7
t0skGXVc4GHx9NHKq57+DdowiQk+bZCbaJLHE7FtCFW9cWWyC7a48En0g8rZZFyShhBB099Gy2/j
CB5Xy8PY4/95nZUpKTn2QMJ76tKpZ/xMUO5dGLRPhtOJWnUixhMirG3TFPW7XpYz5ztuke4NNphv
KVnAEZAnrt9aVqrJ3X1yNo5K1RDI90sFgyGHggBL8kEHZDDjihOWDzeVAmGy9n6st2vXjreyBKmM
kFn5enDCdKWz6adX9e0aa39KAvFOOjigIDKxR6MAUiBekwk3g/v24OxTinBscUhY0116lWntpo3t
52dzO2UTf5hvVcKesillPKHWoOGj7L/PI59Aej6CNRRj5PG2y5nkFn2ajd0cx56k2B6JyPEg5JWt
H+qhsR7YZzVmLn915eCUtlSU5NLkapm7ISATmj6OxeXc7wDEZcwusj56+9DtO8fqHL+vwivG9mhy
3dnVPTadWU1SdBR4/IefDIM2jLdFRbAsQa/0lxcdAIHmlPXuBBHqPoEuKGpHu3l4YehLiPDyk5iL
u3G3yHNHhYwoSYOxqZhpo9HjoO1swhAPGE2JaF8pGlBp/NjS4mlCauX3jb7dmhDn9LtZ1bLjZ6le
wVOJZF3VDIYD9/AmMvscpFZ/waH/KaA/76jnEPTuIIzew9m9jCzHABOAblQ66ts2XDi3HaKIIipy
QyC2neXVDbm+icXmKVvksm1/m1GvjXkvk0CE7QxfZQTlV9a0dsYpp3a3dbAzpHQ4pMsD4McA7yur
DurdSUtif77M+0RRqxgrmzVi58E9PZ7yk0+nc40BtfZ9i+BIEYdUgw6F6pVVEko/b9ulFM/YlC86
4yOVj+BEXMh36Rlbot6JFPoV2+lukZZFJhb7UcdR0xAzFWsN4e2OcGvNIQROhs2P/0tgoew0/vwy
2pnn2Uc/mgsVf/ADq/ISpb+P20C2Z8agPXnsxstDro1zsOy9hIN3LSdh9+EKOwaTzHjEwS/8s71J
kdNbhDFU0z3xKFdstVMrKXzDew/CqlSvMCrUjBoSZgf10zS/ppFsAC2SFHRI121vZS9SHnDrk+lS
NuysGs6LmPFD4swkkTWPn0zL+BaOV9sujLI7kQZicHibIlnMUn1g1rjAoBKDVwCBYyHQyAmJHl3j
W2p5EQSoZQelepFx+tL8W6KofbCyjWsDqnh16bKujUqiSa8AAHl38lcHHFQGGz91deIRu9R3X3Nc
fHJ0DPDeCIs1GT9Q/MsyDooJf0WSG4q5iqS22vJv8rjMva+ZuOUwbO5kBrmy5rH5RladTP0HqQp3
V9hnQL64oKtNh2Qb89xEu4F74FUVawY2aOWyvZ37vq7Q93AtI2NO7GXRQiI3aCP8JMCph2l1/c/Q
wokieU6zmJwerRAENiOXHhIo43rlXCIZxO+uhPwRv9it01H/qfPjBt3TK2W5J+oIJwWXymIV+v28
QKdESC1nOZDmoiHKqgZSuJHBitYRxc6iynfKEm0/rRqiANvwgFPTX9pnjC9deyGsTpf3g9zSApJY
yZNYNEUBeFETyiTbxDOx/lotW2jnLi2HdXxudcGlcInvuwMJ0tzvHhMqwkRVD6UwyOoAFOMZmWnn
XzRkGLkzyaFZKgcBtmhgxYRHapVtVYTlyGo22d5TlEBh7j8IfMcoNca32b/fqm64UHfOuYmSL2cE
sR4qJgshh3cw5RBZLbnXzd171AgSwrwmJmtITr2MJJepsGR5qenASzXfLzVXe/HeEjqHrz+AeeFI
XPByf72vtZwUNP18mRPi5yToY0Rh/vZrbe6ZWGdrsdyEkpTozaIou44kl/5HXSjtLyQfICDP1Pn2
XNBj9eC832TeI04drW3HCC6lrpyPxecaRf8miinS8h3ZF5lpMXCLgWrydXw/sgAaBkyF0zXVBorE
my0F+Nuc6zk37llwJQJCDKtTS2Arbnh66snZk0Xz946hwqAi+GxKUuluIEoMwEsPXXXEOZHgL2jM
6D+ygCJJBkAPshCa3iSQfQn1VF1OIuTkQijENUsXhwojvYcu77VsN4QbO07KtXxBB3AdC1TbgyZC
3vwADMe/trzxOI4pVGxwgxG5yad+AzPLglCqtvKhHdPUgO7HsbqQd4t/xhygGR1ragPqxF2p1tGp
fesjzPSZgHEacIa6t0/Wu+ggrhwGHHIveFnqCP+XfZ9LvcBcOPkjwYk5VkrgVqUib7jlPfD9rAqq
1hMi4GQEv0+2Nn8AOn8LAoiVQd4zKylkUL2Ml5uyH0uuli/RWymNDVpHWbRaISMvCGFayE0mbnXf
tpioh5KiMprNsMKfLoxHzY0HqpgS97pJ5A0Yi8B12R4xHZi2XgFdzbdP6VfcTvJDkOdKR1WWMcK3
NbIr9/5kT0N/YjcMDjpijcsdk1iJdwubanUkrnNhHIjgP8nrt5T4E2QI0omS6fafegxYV+132OF5
gr643nur68JRabPzaWoPizLqqPf6Wk92eP6hi8bSFI/K4SUNer0ncctWFSgM5oSPgefiRsdakHvq
r+CQYKIDhmY3v6eqohL0CzXU9z1ZLo1ywpIOTPu6CbkVL4A2cHv/SZw7gvK7Pm5Tv+JY1dLMyDyD
nE/PIk/IyD67gZc98BDBPtrBg4qylBxJUPDuc7cOImQMCdtiHn4IEFTuf/Iggt/bvWEmlzu0NtJn
3uoq5jIKpjI0PD2+Gv4t+Nb99bQhfDnGbpEZGecWj1VRAvOmvKYq5inBa361Zav/GNxTqNEgl7el
R3gVJf8s2E/az79sxUIQUZl31+svzmUoJkn08yLXe6Cd2Sja935KI786ANdGgO6bGyx5Z3pygsBD
+t88fiHlNX2Gc5wZ9d48IlQV5S5Sm1wLlutUNMDO0eREPaVWoXTwChbTzMIKlXai3LhChVWhX9JL
0D6mK0TFSSZzRxaGhsgrRMUPEIxHBLxvbAJIdELwh15OQNxaXcQx12Giu4y6KVDP2Tmqc9MmFJ3Q
tgmGwoWhEyD/bd5Qh7fiCKI6WAEdL30LTNKKGWDNlP8Z8OE9O5F2LpFaLEizkZdCuV6cBf+lLDOV
uOkeR7aJTr50ygmABQb1+GTLTPHaJXjA554b4pc+eOksxqk+9k7A89m8/klraEuY0Mr7sOYfyQND
NeLW8c5+2nDbAPDD/tgHf3Df4wFnlmd3T/E96fm3mjC74fbHrWethezzXdaHPF0MUlSooyBHn3DH
MTUYLJg9sha+PG653nYbCJgd5e7H3c7PDHdNS0+LieeJhzWx02n3M/GmUCiDvNymVA25Q7zjF4bD
hnEJtn5q2VCtye7imjSaJboH2Zyn3ecFl4LjTWcsBfrjBRyQ3bofekB5z0VnOehnPqMPz+woQERK
BwmwQMMz6HuMoX159jfWLV6fQCG0hrdJMIDdA0lAPc9AnmIi/mBmRK+A+pzW0Fg0ZNfHwv4GG8Lh
aAT8WJ1m8reH8zzj+We/Zs0ECyBLnGhJH5yUcpQxLoHlpniL6NheyfMc6EYIGSb9QYhk0KDfZILm
mrCw03KxLqb/MTAEtLNcQ4sPzrOItjMYUYs2sNNPl1nz99hdDj0ARjlaU0HGOG+7/1ISOBa3FWy0
BUkMIBbNixMpYNAcjCkc63hphM63sjttsfZdgJHuU8B0BWxjn66Ut80r3qfYg1qtKhp6WSYnB1Zm
wpHri98xWDsdoXsXjlZsPoeWZqbeb7wkfV5ly9U/KSezZYBXxRwyt8ahRBDA+KSFfxkPMuyj0tkg
okhJvxV4Kl6ZCHDFCnIeWAFJ/jZWXs6+7takt3f3UyNBUSJfXLQVPyWo6QTbDrhkMQOJwwDcCzDd
YZruINgRyvvPvDdR+0wOyLbw1Em6gVa8IBzqHE6nRsYPVcMchLgNa7mIXT3r29S+mPo2DP1heH6N
5l/FIwGAPGLTJF22ksS12WayRhr5f9U6SYuoHSNbbK9w96uz74caZ4nUwVwKWWAaFYRzQsigbZhX
5kpaUkVW0z61mQSGOOfDKc7H1M+ljCZOICUPH8RorTJUX6El9ixvh62o/Elu8ZWgYpqhOJ7k6hpB
dr+u8V75YDtKAW/j3bsnOCI0f5jA8oViVf8Vkta6vkQPujSN7uqZZM1fduDCzH2Dv2jRyTplaMk4
V8hNi2SV3vNzavuDoHgdbIMz1hqUEKJqntapYqewtWs3iDSPcsyZYAk64OxHul58mB/myNhSdOxk
3vzhACd2iKx5GcKvc1VoZTaxWNCtxY0ijIXuToVA8njByni7imJsYZvfygPASeWq+DqJaINKQaXf
nK9CD+FxOul6CGw1260ilZ3EanNOKyeHypqnhUHIqVTuXR8AMybFpVcG7u1NLZnfImednEV2zMzd
N2a0gtF9ZKlOvceUGYmb4rc63O9Kp8cBZhtrVv4Ke0xDYkPp5C+kWLHO8yVeoIprQQJRID4GopA6
ATpeHPckRdsfO2lUi4bb6Em2iQCuS9LFjtUwYBjuF7zsti54Tvxvu7EM/JSknxAAj8C2tScIIX1t
xjNsfr7UT5duB+voY/IGBH5CVJYs+TzjmxZgsyrmwynPQzlWRuUb7wxBygTAUW31lQc81xjwSgWg
SldlGVdInJWzV9huR/WSVubTSeqtUdFPuICzmNGOgJmgf+rTc0Z5H7nvvzUdvqjZ9oqfYBN4f2Ee
D8gOqTUAzbpt55H755QzTYkJ7nuBHWnhYAcRDHOZX543qJAB13GOYxd428fdguAo9wyeJDGSDlKX
H/VCZwUGIeHl89nC42A7Fm9m9ddno4ZhZmMNIb0/htgZAZHMBk4wbDxY/fxOLxRl3oCPvyNrvlZH
J6AyN17l0ZQ20fXze9H1LxdcG64zBRprX7fffDHgn1lLDhMJ8qJm8vCoqMwatGJogoZEMOpROJfe
gMa1y/MzJnprxqkke6GxJuI4tVd/VeG1nxAYjXjRbpT5fwEie5sueowpclFFeR+yZUGKux1c3l5d
wobOEWt7CdTWprR//UXUTq0z3CxjBfFF6HC9qYt/DDeHSBsSPv4TS4jlR2ZUe+Ib6bGumcucgZYU
rIXwIiNIXcwaNqFY7Zax4xRp9844COGVbN3YkJOO5L+umgN5drvkPGJNNzJNfs2/R/TGjDP4GIG4
/XBrK9hS4jm5iZmXmql7qtN1yVUV7Ht0mpUppg6NUqR68GZI6r2bOfsPI5AXZO8v9nRwxggdqLgm
sTNK312r0w1W4LsEZBsjCXaTFJsX21S6XEKwGCJeB6jC/TN4JWF8gVT+lczCHh6WVc2eURkaIh9c
VIeQacdw6h4eiAcO4ejNtKHhd1XBEeiN7jUPuB6FKfRjC8itCZp8fhZHz6zwvwx5ak/jCaYaz0mJ
XkwGXwHQh3Cb7sk+vMXtfXhKtm+ajOEXl0WJeuBH/gI/9GB14fiZCaZVW5EVrnGrEWzFXJzm6P9z
PbzGqtSYkbpdu4KcT439NzaKLgk4klOOgl78tQICwT1q47S63udEZpcRJjmBILAw/4M6y4lRMN5S
MsuPtaz6QAhC2A0v9sMawZuLxuhCm/9YHuybwSLIkFXq33FWqNRuW5JEkXxUg+ftowAFtnXIGK8K
MImxH61C7BRjcbflm0LRj5s/0YjHzlfmYnxnug+NmhjkuIIB8ugEs+/QuVoL3LjlZFME5dfx4+R5
P+GO02VhuawmGWCE1xyknNgZp5jhFxpbgUsK35UXE2K8e6QzY5093J+ehEllmi9RdoIkUuriC+gH
wqgBydGyjMetTd8DCqkzDmM9CEhY70DPCuCrupkXTc6YpnuEefSn8RPlLoUJjjsdWg4QmcspJjYm
YPWcxYr+U0cwxJiNH8KZYHmNBWVzPcOMxPV7yuyxdYFo7yv5mDCsXg2OQNMtWAuyfiZrG730pA6n
qO48MGkwVeyJwH2Sv3ikp0zEm1UzwVi3jRxLdUhmdbTOVjA35apYYgsonTYowCGQidHsE7//HNAt
hTkoGQ2/Ok5t+AfmemM6juImssnjQqUMlOItpVHTg/lQrbvzWDQys7lYcWUsQjdidoqT/wuNYvrM
xR6V66+5pWOrwnNTC33FmhMbeGqwMwG0xm8xvc4JksF1hCDwkFgn2DSEPuKJs7IZ/QKsJOFVwRft
6sB/1kE+U48AjaYKbkFP9zDIINXD+Pq+g44jYjfNjYl65CSAkSQkNcU7MWTVG+H6Ab+0n2Hsa5FC
ymtqS9AnOkqQjw+pule9w8t3BDjANGCrWggtFw6FHH4Fn+Mc3nUtE8UA9DQNQBcQzjNJinEM74Wf
z41lsKPZgVdu2OJaT3cwpaVjnXSg7S4g7Kah534yfFtOK8Mrsi63+sONMDvMqXhb6WMrfcTsVeLY
XXLj583FEkwN1pImnmGwcYa9awtulKTGgE8DIVQjEb6JTalG60MM03TQwB4qFd58EZlsL96TYzGL
SM9rmdFgFBflD8ugz6LIWFOyHry7qLBHvVBEZLpEE7dzzRWxtzyU50NW5TyZxF1CC20Tvl0eDbBg
bPYUzAVRWg4KfuW5qexQRSeGgGn419Klg40xeBLN9FnxZPB/bk1hVtVjugzv34cDoi2xgn3Ipe2U
DJEsQq3p5H7hKbZ9V15nCxZXtc3kUcIUxzc3iXBcEcYLzJfcWIwHCTy3ijiaUfqsjFrIsxsrZu1s
f/ampd9lj16DzSygZzmwgrLVxn4oiJNhikiuvrmNz84Xwvoze6t6nHYYYvWHuEK/K/RS9GQtFYIm
ouCJ/x0S91vD1mGE3LPQ3WzFp8bo6NfP7EgEYL+Ml+ocSWndzYmGsY9qEYbc3qwrofzX51yquqE2
z7xZqHGT+IuzQe0rU/vRCVQhYqK1McFDE8DkQllbQ5Qp2NErlgY3o0OKbbP4GKz5vctbB6pgmFX1
M4aGD8STB3q936EbjL4DsRrxuDbror+jzM542O/p1GV5K6yX27BET2308ejNZiHQNbfPrdpG6psk
lBxTlUVaKnZmWdCsX76WqeWmn/6C7trqSFftXLp93suoIm4TQAYfN35HlWrQiPoGIurbFTaJOvm1
nUfHsCdckGMeEQSzPZ3UE/BlHfrv2GiEZCSHlNf6tkqIEH2NNxXIouPc6vh/qSc9xKwXzjPgVKaM
xiw2nwv2fDZhlxANwXUm7YmdFp1D1wCWoA2bZ8Wz4UYTH9NYKcialZZy87hVlRr2GSSmDGI1+dLe
OJmFTrgSkEtXfCU+eFksPzi8u/ta3OxVwwKyClygsfVp5SfWRwKAaQPJCOTA2uBOwfgUwpeQsH67
Ysmm/x6XrjWSAspvLPRsoSE/jet0nVJO8IJusCeUpApnS32SakkKzAYMi3XNGL66/NFcw5gc3dKn
v0wqaAUlDwnRFKuLxQ2PBdrOlBEEyGQi3gFLk+bTi4jDFcN/shu8sWFXMsHWmGKHz/rP1WTsGwkK
UnTbnpy30ouoQuQMLWEtZMCmfEMYDK17AbJXalK+9828v0GTQzdl0vOt4Y+RkIAlBlUuYwnyYMW8
AjOLPbvq9zrKkTj2d7UH6y//mKLjPrRwk7jfvrx7JH/UHxxKKkIPf9R8btV+3FOI03L6a9NRqBPg
JYyL7aGd/1wwGwtowancrx1ywALb79aBputY0XHdP5+15BeRPY/FeXqjGyBD50Q5j28i4qIyP0MI
TbR4WJ2jdYcZpFyzuk2rljXxAQx7WeGJvn3WtKXa1fAKSffFBf5MDkZyBGFhauU8xipDiI8YRrtd
AqLrA3lN9Whh5z+RjSibESPCBGzORO/k6w7Ed8RwFhD5v5LI6YlN9CN0N7GtStjtVUYSpjIJMi3I
2WGRrlGN3xBZmS229EHNzjz+e3lYjdD+iizRxmOlwK8T2UtdLdXxYBRh6VjeMZz+m3MGy5ADRSND
VRPlmgPPD0qOKBwjZTeH9MUvOzyCClxQJ5NvbwgnlWaBhWW9U0JN+ip9UkWZZl8/403SSdYtCSCs
wRPnShNy1QVRIZiYp+ctUmKnWk0j0tu8y0BXcBSOM9g/DUq2D+1lYzo2Hv4Txj5IuqodKpcg9OuW
GWRhg/8p6+4iXLEc3RcdrFm73BSmk+oPxTY4cQfavJDqENP3FM45X7WDU0Evil/olxhXvfAvJA2K
fbVPFeelLpJxTkLwWqhgRBurb9tGMk3C2sTm2nlBdI65ixaoAb1FvV9d/gh9joU7Oy7rGABKCxQo
9N4EFbMNcys+hSmCqapxdN3lCbsuxnbjM6e6t9QWKsqgjHCIYayhRouTHy4bInEdAbKhTffuPjvD
DL1kD72PstFWagRsgc3NXnJ1mORfv8DJb37nG5XJj0jgiPbeOkPYWjbD2wtOmZgLM4zQpphUUoef
5HO+ByFYTtfteGi6QSkEHFXyXNzn1iyV9YQAurR3pQo7ookuCmOvB49dAiWU2cpJSN+ojenWbYVE
j9sqdQZm3DkJKSOaci11KOst9U7xX1OXeqdzA6b3RRGvqcqjnMTMPh2YiMCMTNGTV8Sj9pmll8Ot
ppRyUfjfo5ClI4stus2h4JIOC6aZJC9OA+KzFOlbER7xYaTLlO10GtW9/fNALUNVEAYCJL1MxLV6
Vck4O7js8vBuHV7wIo06TTrmwhklMynpZOHl7cGAsFwMPdgHVdSalvi73fqNV9ajQFxRbFmGnEkT
QcNSuaWccPM62WdQ22qGMSEMKkpefvTQLjs5+Zm4z4cQSpL+jOAMbnT5NT2P2wc627EZuPlrzDUI
99WLsCppQRjJL3YOW7B8oOqcHnxfaMkiRdXnMOjo2AegExtulkZ7pBRhM7HlMYWm8Zjfi3m6BhYc
cOnKRnIut9uWxzTwBA1MTtBlKO7uJSSeF0yX6gw+A23d63G+JITldfVI/pXeKqBPO80+Lt8wgmB3
6a2CZRw2EYM9z3/oK0kR8ztCM+BRpd/8xP92pfO+29iOtOSxqDGJ0xIjiRHUUWcBXLb7I+yPoyby
njeQweb7kpTe2njl8Vk/YxskU+tCLp+qEuXwPSpjKdPIw8bGjQY8u6ju9C/FHNrtBD15Cf0BLtX8
+Hb/Qyg2Gw/pbiR0jUzx6QG5aH7+Srao12IU1kUWkbTvmK1gLohoPs/NMLINljOyVnL7B2jl1i1n
fI7c6H8XL3h4gM1Z9q2fs7KUxkryZHB7ZamD1n/tINw7AYnT5iE5yiPfuya3ZUQvwRHQe7g05or1
Vj86wQuGKmol3RCXmmNUs2vjzu+HAIPXCl9e/YekgKHVhJ9k37c28YL+DTHZrw5WtJ26B3YkXVOu
anS9DtN39AQyAsHtn3nM3O1v21fYdvwWnNx+oQFRC/e2nyygKbOjrbsPQaJVJHkEv2+rpJNycl98
IQ1MMbxqA6TJwXbDiolK/IrGwClmbpGUl32cWbb1G7eoh45jzJQJ5t7NdsDBwHedaOdbLor99Da8
vD5XRpxgKMyIf53sYyCfnu+rrdpeMx/b6/7verE2FZDiwfj6Y975uRKUE+Q/kAbFTqSKE9Qbc84e
r441z03tvEhMqls8Xl7NRJSutFW0VGku8/gG/j4e2H5IT26RCrXkWlpkgDcZjkKxObbl2EJBg8kd
+tn3m6r/i/sO3A6GBEDKrUWdOyNgc/0VAI+BvWtYgopA6++V4lcEU1JpdnQejplGEOl/S3ADgmlB
RPad1UJwCJ1MUG36rAXQne2djocjv6FF/aDDeYNKEVnlIvzH6jS6Xv3zPVeeeKgPcnr4gOF6QuxS
drcl/kb0VpF0ccD4oSi0CC3+U7ubJ1+UgmDq2wJOKXKF2iv0fNX6/0WCnGG6qFj0he0CN/Y6Z8fO
m0NvccJeBSt1Zh7FZA0K/c+0xFKbwasAQYGBrW4duD/iO4nPxPRysuDlO0NRYjzMV+5EN0vl2/wA
fvpkuv6/neFoTHe836wThi6A5w3J8/ygTz+j+1UMLrQHo+QBAEMrje3eIrsBd6jKCLknM9lzH/pV
trul9XN0CkIRI7eaFu85maXftAp6TRPdZIjFDYKb/aIw7WGh6fjwOOnbt8Blfqz0V0kYQY6JprgQ
U5yOUSGtMqxTZj3/g/c24kQTW+jvSKpjR/4/Uzll0pUih0tjYhL26GQFD+ipb3JwXMKChL+qKfJG
FWL1OPLzRlTO7Gi/5aMKAPah8o60IkiLLJPNGTR1OG0WvsUuGxH9GfjVZNnj9BjMi10mD424FeVJ
+wL0octSmFUFbBBZxXTTd2IKZ3jzySl38eUEAnODyTRxuyDc9M6jRpyFTEzR+MOHqwIz/klY4EwQ
nvyQuBadn8vwdw80gG3oSxpXt2+r21L3jAMICJIeAzdRaLoHtv4paYSDK+3D0XRN6okOrpeWSRT6
f4r4YydTsUIRQg8bvEkidZOF3eFudhxa2AoNr+Bi0z6VNpI8Ucs5NhIOtedX6NGT7UmDwYpA8W75
gH9oXJU8luuMdirPsq9fRBGJtdL69wBnFxsZX3VE2UXqQ6bZqh8n+OOnxSqI3s6AiRj2iNA6Ufgc
IGThCDkj1m9J+3baA5sMnNTjtFHV+DsqqNCqqg0fBcQZaExXK2yiL/twjx7cS/C94X8jycRwYyFg
XJqv5ihHv8Zib5F0PmHm6W9rfyZveRLcMjBWzersv/reFPEjCUw4q6n7oPqca2STqq+5gUbWREJU
eC33ufOURl/crfIcmOfJyvYmw2wQ4hueEjoHr8iatetc7M2w5uL0dDrek+S2vR3OhERopcXDRAan
9Zfcxvi60kuMVbHOedrEuXohVD61wK1LMUOfdemNRvd84hnqkefuXwU1RaOJenesQRh18BbygWdF
2o/r1gTnpT+B+vyWEHVlNjS48X8tl/Ba1EqG3VduOlbEAfOAgX7rM5/7c/H6udk/X0C1IGnjHUMh
QR4xwN5C4kYmi2IT52HGOOj8GojxIYa46NawBjOYUv9rQ7s2gIERJjYj7vjm1iHhMTeW/NtQRsDX
BEdOjXo5jq8ngMFNDsb0mSD3lT7EdYIZfR6EtOgcR+6JvyYMTDAziYeYfI83hRcSpAQXU0stp5ko
LDPApJbQ9I/BrWPO+3Tr/L6W03gQVZCQsssL9QyvYs6lhrSctsLlR5wvASUYnOgbDL64RfuxEjnh
vTukzV2o0b27i5HEqzPDeUk54ntoLmTZ7XbrIvk4EP9rUVEZK0fOUbbRCz9S5Ef4uc7o/d5BoOxe
kYASgXlb3vVBmVrPdbaAGYDowTu2lriMk/7tgqH5A3vdKdY0g4Tu6zYNOzIX5xq1lPbCuh3IRGq5
MsFnfeIjeJneS4g7PpoXgbK26Svwwmu34GpiHMjJfUWh2iPA/vnKbVmUaAxZWmaNkwnqcaOY/6H2
mzZx/EdAM/G85raj7F00x9jkmOZpkRYjMgxk73hjmdnU9sHxedy9/qHwISgC5+HRnZk1VimUrlC5
4wXU/uxP4dyyCfLvBk+mQa1YZnW9uuKDa6ObJ2ZnrI77AJTSIVI3jBs6FwIXI/51/+x/ZaQpzlq3
EpxRk91kjRzrO91NLdmv1UzzlnwzP+3vNHmi7CKxqyFMapegr2Hc8+EZ35GG5AX+q9TxKxZwkzar
SXK8VABb5vMW8zKzludJvHMYB4/zXdurw2nX0+jus9WuhJ9t6QM/DrNt8lFhiVZIjADJZe9U7O9s
UG6D/Yur+SUmCzBeUYOktnAPvu3XxbITEWIJBrlO2RgDmpkQOhUw2bFfnPtfQ+YIZzXM7j45nC32
u6E+1n41bI7CdcwnSRjRC7yVfngZS5nAcvW3NiF9yzTPBnxrtzBjfV/xI0wIKQvFf5kL4Ygpk8MB
Ple4djYS7oJp2tdxnGoLCzPelSA0cPuWaFVYg5/oLb3+7691pCATnRhvq5VX9MXEQMLaVMofVTrB
xslLw5hAIBZYr0QN6MODxYpBwmtetyT1aeSzNtMhhxj/Ll59hMdammfcVjUDuyVdKci4ElMpG8OH
DWJuYGE9lGtU6XCEw2s4hL6UQ4h6RQkpAS7qn1IZbo6kpfx8PpDWFYBZ3ZdqhkHVM9N6TQHBXl2Q
7g+srTDtMzPrHOZsuhvOc3WtubpEJloOdMjZ8Mm61RGvIoqi/PASoBo0LKVSqJNDnMkij7FhIr94
3CoaQr+TeAnO2F6TWHe1T9BBO98SfJnLZie9a0wsm4Qu7WtD9Py7PWK0l9LepWrxI4Cf7RZnkVOj
sR8STvgk6Q7YAoAv5kB79rVFD+Rl3Jfb11Rb1xqTfyagAmNZl2479NXfyGG4MH1zsxtiNaHjDLsU
quU2Ji0Y7qRAvEaLDNEhy+0sFsC6QYCZ+LDtEje7fkRLvnBN1QwkI+tVbjveDkol5WxQyxJFN0NV
EqkufNMYBAnC4/6VGRPaUYpGMgRxFvHGacrbyRuNh/Pbk3bhZabb3S6Rzz2se0owMcd8dg4embT9
xWmebsMnDZ4cOwHjYrR0YATcQxtSBgU5qemajegWVNv4ZzJiT8wF27LBQMFMHCxVNtRVbG6P1QnA
xBaCdl6ilPbjz07i7+W6DDkL/iazQfcufsvdGBZ+tgkiD3TUzKqQXCdu/wm6y9gG0VH/bN1mSY6m
B3MsKRIR6rZO+n3AIUrRbLkKletpU10yYnnr9pPixmT8eIlM9kv+3Jw5RhCHHxiMPCGS+s4ogi85
ylK9AoB1x/ndZgW8Z+pmHUm5C/4CeSPzi14NQAo+rG++JgA356eKPPhS0fyJJIpOmOuTNxgcZfbH
6OeGu4iLUxXNFT9l29N5QBRNRkUd045Q2gGD60TV/s+QnrWSl0OQuz+BAql35OAQmqxYtADqYJJv
cqMnMm8bY5Xyfkz5vjNTOKtZtheaH8OVXkjTIQ1eLHzsjFr5cR/bQm5sM+CPIDDikts8CbZEV5wg
AUgyl9Dpa5WPexQXRjyM2ebz/KTAeBWz328t5Q29+Ynm1U9tkal8sSgN4joyyp3ySbn18gCGhmTu
i4ADC67uFLIf3ulKobcFY8grx8T7oJeKSomO0BnMaCpxFcP7RisH6ZIFBrzQE9mUTHq+NMZ9zArH
b6ygOrPEBPAsp4aMlberD5dnON3HWPUIsdWcTxTmELgznB9EcxW3P1ahGSZb7hov18jXofRNK8CQ
Xp2BBpESAKEzTJdLCvFDd7cC4NVVmI8rqrYcF+4w7sbLrqs/dDNJY4yeInl/yqVGDy0b1rhKuy6c
EIBp17DyA/1putTOE6N/uNEC87txfrDdvZ6BJhPS8dkFlqHRxtjaAsoqAgmaFXbiHiAKjH7YRRQq
8HLrHz2JaABFw9/ssnfSztCoTtF/3rbs+VLV/Hfy+MABVq7RFOvCRHb7pGt1vLA/86wVA76jkLz7
z7XU7pv79rHDPEaFl8k0krrlKTv7SJh9f/OlSOytpg1JwGHE3/1QJeq20x8mL/RIafe/9uWaPGT8
y0vf0RvqFq3WsbH2qJcx/0/3HACHSkkjXr0aIq2esGa5J0aInDQs/Ah8u4IRDxalRQcFE1jIp8c8
EwsgYIwUGw58fGujJaxzULTzgrNbUBH+weetFdO8ZwNv6b1MzDfi7VzGrJhKdFnm1t0FWq2RAOsJ
1HrTcgTZGbpapUl0NWDaArormQKkXAu+JumiaDXzEUgQpz5x0+N1waOG2MZOcGdksjsPmKBMnAEQ
LavCXC+7mwyqEL6HKCENEXn9YUoYTY+cg5g9cXB48/lLDKtlmXw459YirNrzROlq76NQtabas4eI
WeuoYDvWdb7ohBE646Ruo0OPtGgTH8UwQG8A3/orcegoatglZ966KHsWfYerRiImqILlD1GH8V1l
PPQuRf0DKKKilwSiDy/pWI20Mn8MSj0F9faO7e1OhuvKWKQHZb/mfn+4GCtMO1fA7G/Ji+FoZahv
4NxIphL1WI+xac5nZvd24GE5N9uSzOMpyCtKeJleDmNdEHfbEhgD7Ro3/mMXEuCEEsN8zjObjVYD
hGTMDH2BK7lXpPZZoI2tttCx8BQ3+ERY1c/1qOoGHQiWYgrFzScXIL7lav+ldGj1dIiH74xWU4Ij
Yx0+32KexGrrv+0fda7B0OYmQag6E1IS8tg3vn9XGuRLJqUbXxfg7Q2QoZSCSNZxYZrtVZLz89qb
u4/5xcnxbMl1ZHXm/DSghzcU2v1H2lgy5NYLYl0K6l/p48pepBV64PcOn7wPRi7rdq63eqdkC676
tFOz9eVIXi3MWDQmfeBV3BeTg3wZ6sAL1BrtYbAcMura2ychw45CPhTfeCm97qSgLmOFtkbWo+QG
XiuWLrMpw2w289pvxItWjPPwhpQKlS67FnrOsk6kfow9ZP37dorwGM6S/pP3LxPmpuwEnnuOvSaq
T2BURjzEvf9FjCPjsLmp6gornJN78yqaZstDbf8Nn6NziqYUD/07XyDQ/fOegtJAicOwewApDL84
mDsycIGl3P1Kfl6xRo1DadnqR7/Kp0b4VS17l22bBEOxSz9Rwp8vLYieg4bhlMeSVWFokE278H8c
Urp4XPXKGZ5TuAaefqshV9xxkJlSuxTE9KHWMvSfJzGXnSArL62krkrs12n4rQlEI/3ndpGATQ8y
z7UdASQkcHuMgNCAEk9LUXJfds6hre12tbe0jTkHAvdiz7Mfkvkh3/ojUhPutYtxKp684uAKzbKJ
pkn8bgSzkoSpRepQkuy5qHvyF9EXsF3l7okU9n2n4G9akIeD8zkTgWv/ZTtXUPzHIhcY7t2GZVWV
NdjDBtGDAAFQPT9gh4gvde/ka5l5Vpuhg8eMZqr+AksfEzWg0q5Gq8XXeIOenmU+3YVNlVOQ6Ank
Ikvl50E0S+XfXg7NFm0egcEHV7L6/RgkiWyzXaDShzzUAzHxGsW02v3c4jSriV5Z9GvKvjTfMKVq
66ul5PY3S2Y4M9ktOM3wVM3dJ+yZ/WtBHng4dluJQBjbhdj6VzJnZ+strn4lXVa7LyCV2HEeDlAs
MlBn1+b/jmnCDHIK6l9tkrYz4ODhH2NF9j9QnEDDvzzT1kdxzR4B7B/xIFp66k7YProM8e2QDO8Z
M0nfDIdRjH5pGHbfmnslALu/OHUvoDJTMw6zFvITSal7H9p0Xa0XNfNitzECmJj/Wxu6qY5OyOc/
WgSRzkf6Kd48N76g5UEaYhovAcM7U4Cpo4ggfmi+Px0yMJjupP9ehQfLylpNmcf4fpCOtRt2hY/w
4AefOX7SD9iroyFNit8qRjglzDl4mbTJ5GRcEkff0fsaCPufOvcKqduLRJiIYDoffCDb+ru1/URB
uLPfPjqAHEn2sGwnthmKssJqcW5pa4SbzMokN94uEKnXGBGfQKlRzQ3wLnShTFlQPhGAestPbuxH
jLYzpaTcksDJ4C4w0JGjAkaPf6KeC3o06MGr/nXly8/wtqXAn+VZDv5WgREC7e4S5o/V4YvDHoVQ
tJr7NBuOtNUif3T0S2JLkdx4RXcXeFn3G7I7jYxUKJ1or8oj3ytoQn4oIkXw6DwnlGG+jEt5ANR7
EeOzNlMvUr8KXT+dMT58XgMhNcSTPkjJX5h2193Ise9bbUU4aynCsflQ0ajE3a7StaV9TpPactW2
yyXCmtn/fNX8V+j/J0SGpMTCP50H2kJuES0VDaZvGAGhJJVjh3mOdQ4HdhPlg/913yrezzREXzTN
jttalDEKu4vHbweuuH3AhtXUuTeGQU3omkThme9sgJLL80knM1e4XKsVT39shSkIhIFsixeJrce/
JbbBcgBkn8Ydn6myc1vRxge+PdighLWhV5jKixnPhNj1UJ0mgtS5VvHoNgC5cnbCPrS10DMjiUMk
TwqyWbX45FKcs5CPcvSp0M5avmlXLwhJk6t6Vtlf3pw7LsI/qgNQ4t2zqwpQQcEFs5TnZUzUsBQk
St5OpKUuGl91Tn3ns4rQJY8g3mBfoVMSOM5NdqDCl+EyrnIWuY5p41+BoB3u9ea2ccderuy7B9wv
/fCmMtI4mPaKBI7IfDSROlQjCta0v+jgX+rd6HoZUmbaeQ0OEizxgH3Y6zDOtOhPGHEhetdFPy9k
0xSXRP4UIGm2WUrMYg+YADv6xcRWIVHw4RTfe65trIjdS2CtCwppCYZs4BCPpnwQKaAOfme78b7F
dUR3zuRTWpMddgRymifmzqPRDN+pNSrJUIK+JitpS/Z6AFX1cFgeHmNxZL5fk8IiVaD3Cg9/PloK
sAiNKxWHGVTGf/ZdxfAvksUaQb0WsMof4/peUC848aSz2u7fy6Haz99M9cDfVR8JUSJKrPMuyyhw
yti0hM9c0sCtHnFYD+cPB4B5dor+kH+9r4sRDgysux1SnvY0yv5yNJvqyZyTojLXu7rj7lGIJBps
0Jd58HKyd3h9kT/igpS7BnOLPlXp/wT/k3KIUE/r6UT8nbDoEI18Rj7sFDXPZwQcbVZPEWnNeiXx
9HAEKeCZjOnBALBPulnNr/hKfTP52CDBhJs0jzC+tD/ib+T9XjAhVuVMWsazgA3/yXcTtkUZcnAl
y/psEWwTOLkktgRjZcBN9EKMWaSLqrupTFr3kURaj+s2pEJjVhIaksIUGk+BFu2OamiMwFBuos1Q
o2HBoWZiNZXljWlpvML7Oqo7Bx4sfkJh2a+498OnYmT9ZIeLtG5cCV4AdfzWm26FH8XAKF39VfOg
qIe3HigCTy2XHtFdstZj+mdR0QSmaoWG5oYOy5lg11Fj8zhPV89LEnlzXp9NlPxIOWDef9IDR5Jr
qKG8dn2gz71HjAiqgSOmiU0iS11QgvskhoZzaADf+CL1MhP2b1GoH0g3FCmfsdJUnFy3TfX0cORJ
EYEiVlwCoWeQs8YGj96jv7OHuj/4JLa0UcCt2RP1hx22yQrPnnYroLNq8gHcq+xpcL1gdwPrmETf
4f/LPVkTzbqkiBaeaX01zs6qi205lMYku5l8zEQwwMu1uLkvl0f3gOor6gSJ7scBEqfixRodxwA4
ByRSrrVc1sj+Qrd1+FszzL11LWs+yicdN/x5cXDvXy23Tjrgw2BLIbOjydXa46yUVtnErF9yGFWg
fTMqG6Z8biMHNvjl8LNENFGMBf/bGJgZOQJYtzmJg8pXs5c1IKVuqDvL1wPheBTq9jTvCFALY1Eu
VwmNLUwq1EyuaCIAg4SBQqf4A2PJvV4YhOKt9zeItAahAKTJARLiZk4hi9D9xfzqSAYSDvnMulta
huLLH124JDD0aavCto81B1fc2D5+ZXc6sxU1LYCuORpVTXNXMYlbBZyDPNdkddrrYTYu1IBTaP6l
X2SMrpN5zYWx5OSjuu5q/z0oiInrKE7Pj/J0NGHcGX5pxIYVA2Wd9tOsjTuMlJDNDtblQ/c69C2x
GjRwgVas8HVnRhOI89J3ymFOwC07WOjmZVtZnxCZgPW4HEbHcoTsNNYEqxP3JQn2KSWrfo2kN7z9
gZu/e52xK1oLi9R1pmlrsS8hSVWirSdbW/h1uHzRY9wQrUvJt4T/Kb9hL/3piY9F9XDcP2jHaJMf
/5gT9FuHozUDzDhBklIh8l6EZ0Kq7MiN4/kLhpyocDSbzzu0m0eeaLC31OdJkj0oY9Iw6feR/mjR
mKANuKqIR5Btpz2zdd8pWP4+9l7GuTx2W+XYuByfUpJdXQ2ZLkY0hseG+U+OTB1ERcVe8fD5xW2q
Wn3DKlW+a6bcbKwdoXCXvMq/Pv+qmZdYek6SnT4xN1wO/Q1CoSscCyJ6trBlL6U+wYsHL+p3FULf
Y0P1PtHzgong77Ccx6xD6BK03t61FdmmWLQkSynvMEusfL6TQni1eOa4e17E7stm454MBEO7/ZYj
ITMgtdwjd8C06DDYNEszgll0Shc9hAyl53kTovVqSnAclrGIorOVp0gA0IAlSBGK5ubXBj+qzWrE
JElror7jaVnkDnanlPVlbq+CysDK+Jduk+zuMluK+ZJI8WgP4Tt43+/sPt1tJOXhceOeqKZb/X/1
9nO/Kbz1rBDlzeZ+/+OTm1cK0nik/6FRlLVJiOsmRljQPDcgVG6fW4TUnIBh5jzn8dGXRfEwmh6W
ICRGR+u0PZ57D0D7i1gCULQbllvbVW7KT8cmaPPREYGeDxL5ER0B81Sx50CFBU+IvIZnbKnEaD7M
2BacrTQqlq2Uw5Wp9DiYBXLW6jdFbaz/TsNBAZeedjfA1+UAgzMLLEAo7RfOg4ZFMbKuBuZxfijX
iAOPvv7J2Fbo0ornQP6blWLGN2tMfzj71zR44KLpTo2vKiiGcFtY+Z3BKMh3JXrQ5zd2rq5vmB39
hjD6ZMrdH/vj/5o3QqhVChs9NCJ2GHo/I97vJUKYAwb9CzVG7WZ+wKEpMd8ULN/z/cKoUzPhapfP
GFtjnoacry64066XqHJCII+EIKfVOUS+FPiFzdgX4COZ1YD6TDGofe2KthVhzP9uF75lpdxLD7Nd
43AJgiqad8/xCWiUk4kkwwZxtG426CBfoEFeif4GmI9KevJn8uVP9/gL+KiuLXyFsHvW5L+2Y7tG
nWfsFSMuDlyTmpFEVIX29tAzcDCRjwi8gMds5w3xRS5eauCqmaJ0hPNwltVVh+Act8uD9ys8IYJh
9OuC1fXjE5ZGn1KYWrcu3a3aAn6Z9dTbREYW14JpX4MIZzd5FAyJ/aySsN/QF3bGx5eg2yYS632s
g8vdJuDX49dCPdY8ZrMMgfozEodfvT4crgI+/zBa/4cua2P7lOvrKUQHWbeg/+Cch0oXvjC1RfxF
O2SUwDJj1rQLGruXPkd7EUnrpLjpmVMq1HIG/lVmp38SDgJ4w/r2QYNP4LVREqC6tKkj8tczGYr8
TTfuSh6pJRw0JR0Vlu9Df828AeAX0QtYqbR3KdwG46U9T7CNLfY1S7+H2xqmxllmZ0qCKx262Rmr
Y0QUiMhe66e24Tds2iKXhZuxTvUwUu0z4Y3Rn6pD7la42gPK2K/Yyipi6YkELo/xlPLnyw4og4BF
UMyWWDTOGZzW73rARqe61a1zdK9YSS/cTa/YzZbW7tAEgsBhisRwpr7fNsethP712EjeHEI3mgFq
8bhZTK4vEZJUiyT/xGRzeNxSTYIdXY4SigedGDmDDmPh4fBWqo5hCH34slOQPBwJg9ZQQVQyk7g+
Ya1/eBaToBkivQGnE70kR6Nnav5142HCiP1yD08PBoImuUaZT1SdiJNja5PphEpqET6POcesKL09
OvneB/DjntfUOM6z6pidZUNdDkENz9vdBN/kGqp2o41w4VJ1Z2FQF+EvPHKgh4PvRuufgyzl7QRl
dsPHS4O1e2oeXrL/pbidDOmPFsbBO+qmHJI646YUEriIeAm21WhSpmk0PgUruqPmiIGTCqQKqqzJ
x1GxXkTeEYRjucWEYpgE4NcAdZKrnWWMD36WcnCjJ9P8mXTpx+Dwd683pnyxnL1+R6CAYYm3nvnH
qWBB4C8rnjsBitbUHw7XmOl9uERyFysX7U6BBKZQCPQf8iye63YS/9lwTarOkJ7AWr6mqiH1narx
fxBi6BaDtKfK1CkisHjvhifm2YcryZjjv9fUE/A3Dx41hfyX5WisL0dx3KJtynuywUIiTbth1K/A
oG4AS9vT9Sqmj9CCpQeVCWdCdyNEKc646trkZpLs19ksKJXF16AGIbnclTS+zfi00W74UrgtYbIB
Fp+TdP6exnAjsVgRoSqDvNsFoGxlW/o78+dWrMgUXI0xMFGImfntFL4wCoKh5ZvQeJuJRivt7NwV
ckSLScKZ5YFtk1xYnL+lsMVp1SjWk04OAIaE6kp1meFkk/dZjZvBjsFCvKco8eMh6nyd7iY+ejbc
lH+V1BDNACFqlk1ZWvjRGVkEAdJp7uFVUU8DaUrm0mr9xaspbPTAqS3UjI/+QIVavxUl0KMxyJbE
lPeqZu+YW9y2QvPwm8C6PLHDoAxxr+NW3aieD1N+1CslZauiolvo+hDrPZ5jISZf385j8hEjn5tf
w4cm4F/rcuI/sdmbeH+bXh77OP2A7AYc06jYx517uK42XX3Jqa62YzzGMZboQ4stqYi3jtI7wVeo
8tVDwjIa47v16tpKIR5AzOxXrnyPEmdArpeu3uD/xkN5UaWJf8PK3/r3JrihWqDkAOmGCKzEOUIL
wZZ9OJvUTIjywbYHfXSV77NmocVq4qfAdI9zdgA8a3M1LgRzDl3PxCN4vFc9rbm1mP4U0h1KfzFb
a/6VaCrEaLcS9D/HdfoC0Et/EHFYfPgyeCMc8+gYhPa4yhzmiShEWsA9OwAbzwKy+LnGp4pj28s0
WbNEK2zYjH6WfxJ4zmal1QPvzEXR9KPjxpWWRPwM1ta2xI0fKeMgrAJ6d248/FB5cpxoDCS9w4Mb
Ybf0CAXccCRjOSBg4B6vghFtw6CYNYP+yKmncxR46h+vI0QXELMfFwDRwpPev/UpxSLkicK0yKlK
QsQBKBwwn+Tpq/WbdLXXpYLllJCu2fRM+HhhrmybozrhX6AIodbZo3a3/YvNoL8spydFniHuMRrB
UR06F566Tk5UTj8y2yyGSqTQqprvKRKs8WlY56JSchP/7+ZpGbnmtcRTKgb4UbwJVyGNl1ScCXY2
YtnOX0EC1ED7UV+Rmgzkp9vBzfWB7IHDFDK9+252F6Uno7T17IOHy16HQkPACfxAcD3hJZpnQZYX
/NUTaZtPEttlnEgb8RhhNsl5wqmSXKAaASZDQjuKRVCAfEkyWaeVUjmbDs662ofnUYGlIk8fidPV
4XKCbKMgmYMiDDq0SWycaEZb+qtGXrM7I/Q4BVyf6ZP/UnTySl+S9DgDD2WhCPVOO6LGYoon2Ezi
Ndn2nzGqMIoKPPym6Tcvnyv9vkBCj02eqipVnJbtFde/Gzs/tC7S0X5NdqZw4ngZLpkDSJxyVl/o
D9kfGZc1/7aL9L6Q0KmhQX5HYPccOVJH2RQFekf/dkDUCWFtMQZCPuz8esuHRDTrGbbkWeQsooWS
a1jgq/f3MzQmqeRetETcHScEm5Gn+3LWkxToxDAIhCKWcCFWzV1jp5GLJT1DBRyyfqXqfvAfqD3i
Px1e+IQy0+4vufUSxYC+qomYdQIyEJ85RvudJ1qdJOw5KbcjBPCEY5Kzp1rfjZ/pdk/+wVDlEg55
UgaSp+4ZLYdzOF3gMhHw7geKJ8/lFEh8UEpW/g7sYcMJQqYOCt8WRDtJxNWN1BZkMdj27FKgSKB7
YTmdpIA838XaE8bfOs8ToipZVpOYL6mkfYOZUEt1fqYxrIl/Qmn5Bp+VL9YiVWUTgTvKlra8j5SR
wxNVPEU9KX2T64N0qcl7wzgBcc/WOn9IOjHT3YfuVA0luO68WmJhxMEoGW4MfoJqB+g47zN2gKLQ
Y/e1NiG7Lyk7V8SWA6dfJr3+7B5Ai+3SUPFohJ0gx+q5I1cSxR5ApPQvI/QR+gcxlNmBfIx+MazB
eCsApxd2SFg2Q91LkhEG3GHvxXKfGQc9/2u7csrOJ988nxFSSF9pKA2m59031TGpvN3s3zRTbEPt
qOTWSLWKqtNpqyUmlB4QRuuvjCPmoLcty4KaeJZoWBTY23e3e9niR4j65ZIoPFQadRUoJguywpTj
a6pyOZOEixDDtl4eM4C5DorJN8Y8Q7tteGa+ebCAEK61ELIwmTWiQpYggILqt/iYzpnxsl/ClAVv
WFNpnkQ+Eq7X/6iD0u8Vm2EjWX+S51Ri1sUsMam5TmyX+vQSM+fRKJ25cCa9LhwOtfy/daRiqI4T
bR1cFEE1a6Yga5h1GU1FUnTOnaEJxXn+PdNrF0E7jCbTCTnGAN3kVZtRzR0jgYzpLZxpwffecSTs
sfCj0oJ5riNn08EELaeExMZj0W5Zd7NyJ2A1NEYkTFM9i5xK3/fGqI6A/MkllhJp1WUPxY16nRj/
lVKES485LaGUQQMcwr3FKHv1WongIiyroYxomxgRrY10GKFqV71IaOvw7DOj3AtGQ1nVi6xeKrrO
To3st6GurXsV/l+8pWqaKd+JhW8kGOi+HznQudxg0gauzfJEEl4WAetxkZObACEf9QChO8Pfr0zZ
XXhIRO1ZqyTNfMdLSptByTsL6Xe7AsvSFz1Q0V2k4vSDZPEWUfMYQpgzp8fon19DvJ+PSyijHeab
S1N1QH663AKlkLDucDBgs/x/2qJk1HC+spWw/uOvp4/8j5m+kr3t88/M3FBF8RbHv2G3qybt1k/R
cG96v//6jcSMXiY6j7TWGI9PxE3UoobFJQhcANYq+DIz5DhPlltvOp3369H64086jY5tDj2khd6Z
8SC1fAyOdpDYuiZCLOFoju5oEXWCfiaKtIYPUjdBY5Y9LUsEMrMgN0QVMJWTplRrhtqio4K80bTW
5uXCud6d+dfQsf6Snwsp7nbbiVze37NgonY2tmDLMuJyW3M3pbBPsIPQr/lEFWvtNxUVGAc/lf0O
n+hd6eYVQEAdUV1rl7hR3vdA6SppeNzrdIPHfzxhnoGhJQ//oZoqO2NnIYH8a9wHU3YnD4J+N+zV
EqzWRaeTgxKcvo4jzUpz+yeOoHozRQXMpkleL8SMMfrVBgXk5ltGXXE6kVb6s2QA9PjQ8vmDFKoY
u0eGFsmyxceXHXBlDTN3GjlLPhl8NMT+3Cl+AEB8+ucNthDMAgEW29kC748poQR7vDPwP6HQ+BFv
mQyPOL1g54XalF+wLipZ8Y6vI3lp6HJNya+rZ2AfZif34WO9YJQv90N80vjfz5cF7TkXfWAZYWGn
HxvClfkipZ/iX9bc8JErP9SnvSi2EgnNEmK52h1ogsPePO36lNRAESIQwk+/wTUTbsWIxiroexH5
1OtNJK7A1ottg+5zOHzbu6/6qFYB/8nGTIfrpgP/BrrzxEUC8koCpQVzo3aJVxB7cu3Ta4OYuCNA
9SxCBfN/ROqm+KxzDSZJ4Qlvxe0KHZBxxD/Z3CMfLpkWJE2e+ockACNK96hbfwNUBKuGPqlXJhPo
gTBZ802fwUz61TeVlq3UY0hZtW8VOOKUjIc0l0C1SaPF8Jt6W9DHv2CXGRLNZioEFFwSTX9xQ+fu
lUFbISYp0i0Hx6hZSh4lKn6FeBhZJVnoik6r1L8qd5hwokxpGRGVSWzc91PgAzqwisjzW509pdQi
7Yn2lq3+pxIVwR/QHMc1vbQ2mV1h4fmpu3EoQGHM1Ix2k8kWmi1qNdRUQpc4pDFO8xJSLbec0RDX
uHWAT/GcCj3zhCrKTI+kjYVr1EEOG19o9dbxAOan4qhrP80DsBnH90zMe2JsPPGSQInHHemUg6HQ
563PYmVsdaZf9b5XoeVfbNS88k62TEP7HDtmIxt8lIwUU6l9gVb1BXZ4YJWPXM0/9gsuolgb9MZS
yJlfR3otWW8MMikZw+kBs+Dd0/Aul33JSR3Tdagj+rwKjp8q2TrMQ5ywXpe62M0mMGcUGRvI49mT
QD4TNB4ia9ORbfqG1t8zSptr8A9P4LibnluQEZM1zqOdIN4PnZ/I1TuDoyXVBfMTRqY+BogfOVc9
Hz438NFoufckwQH0Bi+Rp1OzOWWSp+o4q8OhdEz7JfSX251eODKYzu7iOnWxYU+7P7j2d4KxVJTr
JYVO0l+zRxRpyOpOE3JKTw5fBWSOqx7ab5xSwkMR843LwY8nCm2CpKroj/3ySifVKuaFYHTumqpa
pXRDNjpdjsUQ3UYZMSdyuln/IXSxal3KNbWYtWA+2MEQT4KTU3O1GkeUUa8XREMo6UjNRAcnp1LP
bT0eNeWctSLg/gBzWFtZM78lCI7VHu4k0HH23dT45sPzjM/saWZ0ZIxTU2yzStdieSVrxzmkssyV
7YbFiWsl7i1ezbhfrlvbuXPX/043V11fXSDtG4EEhRWUMpE/sl4RqbV6/pCWQrsYgwYo1YJkU5s5
btV1U+w/PNFO5rA5NSkza4cyvJdZEmBN11zi2SZA5ncgq/y9OrKjQnz4tKlU0ywSFHQ2cULIpXyw
u6EA3i0YWn6dFtxC1aiA+htJjDL5HQmSQHCp9NbyOjQaDrXYfBMly11q7VvhF8Y3/FJSoCSiDzGZ
1//XCyH/asOp6ckML+Uyfy8xofYy+HuIQCniJILJ3Joaw7U3tLOZsTkhdv4p0ppvhMhfdyG1pzDo
vq+W7T/gWPv/jKdNPbsW7Dpq8cug3Mg59CPfYK5PnurhYg2QymDfaylKERFHz6+YvM1tERGsZ0oc
HSccQqYtx31nVSgO5rHD8v6re2aAksu6jNa/J2EaJmMKY4Hk/OEly2B0QkEIJjHdeyD50hcthx3K
vwzIzQQYR3b1Kay4z3Q6VPudVg9SzhVMq3/zzMruZkomGm70Xy04g1iYjKUsGkkLbTq4h7rmsLwR
Tug51sL8NaZtzWCRHOFFVUyFo7Te2NtL8AGJCjv3pZM9KffxmD+0IhHxQiabNY7yxYXXj061JPs0
H5CjdnAFoCOVflns5doR02fdwaATYseBLMBHlC5aT2psDlQKbOU4Lf9mS6yPCeeuem/Uypn5FXpe
WMUZAKo2RcyxzCzQuZHeEeyI9jzPUcIAXfiPOASBV9/pMlaZG3fgzulhjKn46xNvwvCE/FJRFZCf
azy7c3Lhj2JJKMkNJe7vfPf3GV3w5r9kXHBVU6OCyVQSOvTTi+BqtayuY7kNV/Ri8P+r7OCd1EUq
PCMSvRB6GUnSfDlbQlIx/ctcCltcQ+b1ZAlIRueGIl8hHo8tia2zcaGu04NGRbn4UgfTuzvH71rL
QF7ojjTOUGIwuZzMd8wpH9DvSoa+yj1lp2hGbA0gAIhc62buxRykkFFFbAEp58LAsAq5aq/UpVFY
goNwlXSz2kxyNIVUhnX9SdlRak3aRdA9UFIudad+SN6tWXOS+sXS6bAOv6OTltjY/aCq4maarg+b
yFeTxJcqx/qEwVhNiLTO8UK8gJQDZEBgWUWSJLIA8ZCOWhSmeDX+yLfLkadnWcZvzszMcuMFdvXo
MSG9yeDqZ6s7PfSavZWqygENMuVpKsOFklXtrEMjvPUCVhjX3StGBl7lZiOyrmYG7MzusZH6+maE
afGdRL3veM9e0SONlhyn7wMq9ekRtxbHNecv80B9Ci5usvYFEnmeB0/2uQCEhBeiHpVd0f6LOUi7
xTYA9CNslh3OEm8vgK3+MNr+kstVCUhbbSCYpIXrkaQD741ps1+k8+pSP2nNqO5Ct1CmLcPFYj2b
njIF8fRSltLXiurmjbXO1Z9qHdPw2q2HP40XzSrx4O6sFZE3CRjqgDF/WYXgfR40vXrjLdizTyD3
mKHgAJiS/Ny7HcdS7Uhcpl/tv++jAKEQAoDKf13L1f2BWvLacppi6u7ed+HGk6+XzHQJODEBNUrn
EGntPgAXyk/aSxm8M1j/dTi7FFX1wmvbpm+SCFb4Wju2Dahktfn35DEwPhyZe5QHmJ/QOPUvY0PK
EgqyzENRwdO9KutCYnVNGBm00/JKZrjlBdQj+uiXgX/6pjo7prqUvT9ilaamI99WaKN6AQvffaNJ
aKf/X+0/6+Xdi0pLZoCt68o+sb+Uz0n1HU2Dx5ZBuwnGKaxgiGDeTsXYr71A0lWGFtLhJJ3nu0Z+
Bsl3w5w+DXy3ZhFjDYvjIjc8Vr6Rd30uGiqf2j24BN2u3ZjATHldZeSti7oh76dxwfrSopFDNANt
KTad3sKyoF99Pz1PpTkHgyz/mrRllLitdLuop8o7ET8muysVRBe4+xZxT3HojCZTdOCX8ohiIaRk
DQLZ8oGkdblaOBrZn5GVpIbcF9bFNsuYhlKNnQO86Mbkg49kUgC9z/Bj55XOgQLQ23ORn+qSM0wM
NdC42f6n4RlxmKQZmJujIKWRdLgNHse2eS6qMUThoMSsxmhSQjs140IfFRxoSXbLQnaRuppMZgcZ
l62Eskm1UidDNZYDCHgQT02bNg1tFw5jtAklCDznLPVB0xyCvmcyUgWdkZMkYbHV0v6ycGVFVqBt
4lKGUDSqpjKTgyLCpZfgeghiDiU7rKACI0ANyi9hYSN9qjEMvAK3yGxTY+2ibEW0UtiBqtNDLdVg
uWqFC4RMxV/3XF9/bC8TnNxThqx3bEzQS8U5v5JUYy9JnKtnESgA7bxOuQSWesYMAmH7+loksCvC
FPHpsZ2ywwItEgiZPvUdxkoZ1qQdg9o16bkiV2lKxTOjhjsHOOYGgo6mS+EV/baOWVupUMD5ERhI
9l8T8U+BBek0EsBDANra2nlNeGM+6dAzFRN5FoN/6/NmjHqKdSaw/Ed0a5gVriGoQEY4u0mP3TkW
rtvUyUxhIQBMSksENO5mY3OIcnE/av0O0d0zcfqDw1GWx1HmPKg8ToaMDC5v8iooM5dzsP68ev1i
XHpjnylOYgJbBvP8Rjbq5gNSq5EKo2zV7mzjyq1LBA3t7qV5ktheUrO7GDelyRBqT3isjUdGXYTZ
cWl1iMXMcUCiVM71VNJLy7Jz0Prwfvs5n8sNcX4qbU7kgJ90LkOzUBxwt3ZHG9JtS44MSC60zg7a
+RH9WJVO5rLJq/yawD6MS/j+T/pgbhfjsPC24EQsun6cACU3rcs+cshIE2AKcVhPDT6O0JbvZ/Em
rYJnLMhTHjok+AFS3r+p+Tg3oEMNQqzk2ng6k7BIXtLcMQMuQS9S4RQKudi04NnTFbIpf13/AbHj
9PmbXa+Kz9eEvaba+uG/9iP3DB/0J8Or3RaLZJwYygLRSBZ7fODnrwNxPIm6NQy0oSndtAtMS66p
rT0D4ngZ+YCsw9wpb03S7jvA0E4cyHUMyE38B2wXCnFi44qf0Tvcw1EiKZalVI8X+kBBpqFgcsjH
/1wIcSZfC+QYghGm/wK21SfyMs/HDpLCn3UtLet9KSu8bdbhD+m8Je8akMu1tWwjvDdvBvmXnzY2
ATr55t81wSDxZhXbP/EvPd7fLTtITgixLPeo18i0dSbjwFOENK++YdtGeFHLDeW0RP8nD1JxwtzN
ZWBZ8py9BmS+eaCgvlmP/5v2/YxaFYPOWaLkGdYrzFL1LcfkX35p1Br3tM8QhHu8g5RVK3M1ao9z
I+e/lJ8PwqANX8jZxudk9HxzJAUL7dw+q3rCHgBAbvZCahwmcl4nCk4B7ebGd9SAE0PZ7j9sjEm4
Wc1rTPGneLBEET1KYYUgqTb/6dCV5bCZ8qNd/3sK/n4LcqPsOQEp7xOtpiuZGCC1Hb7n87uSfA9C
uYeFcPfzqJPVAcr8KY0UFsLlunKWiWg0/JFeh1Cvf+4HAdyQEuoDnCJGNCTfkcMt9SBkrxQHrHLT
RWif1NxSPri68FQAVmvqSJ0fXzinwLTRZk/Yk3hYYW+nLUisNNJpDQbH1vCv8t2vxD2Z+ogEtoWG
4/L70T/hDBX7PqWzI4nKC8J8yQTl0aBnAPRcz9+8Br4dYcknOV5l86F4KXtSC7nmhR+fddC0c4je
B6rR52bawd00He+YUQssAICexeNc56Emxm5uanlxh4uf2e1/isS+nv5rVB4wtKZhEi+yTehvvaEs
+BPYIsYwdMXvuqsv3t0NP+WrHRyvfgkMiQh7L9umfeLuv9hjMLhg5+STN8ym4+HyciW4Vc6S6asm
BCWJVcBe63xdU35uS7O/FBLy3AHvWkJHwfSO8ADSGR3myuYYUJvUtBmEeQp+AW1E6ltnEn9+Eb5W
rsQ78mq1/ud/OaP1fN10EWqw30Xir3h9U53UwhyseJG99KVfIVhunEGxENpY5xr855kFBR01uS8o
c2Ibp+dIvMdlkLd1bbiKzsypKpaKjBk4miIRMVunTm+LJ8MFkIFd1g8aPxPHuTqMjQ3/PD4NoCSn
oEPUmOyzuX3BOS7GAx8mP2OsCxvyhwD2HbqhD9eRgb7K3NyYVYjVO1NZG5eoCDrKq/XTpF1tNokC
UmDrjai6gtQY6gmHNWoM4/OB1x9kNU8kwzmHRoDctYHgNYXu9LP37cSXrJJQjEU6MAAxSUH5Xvfh
KFg9j0k9Vmx5pDi2/AbUgi9qH+e1RHJStOJ63A/kSeD+lC3tAYl3gSBisxBPBZ/tFmTeJmSOG0Eo
I+rbeP2SmONV4XhSMcC8tLOvaELT5yqM/uE9/sHSiH1O0jGy1IsK9toeyLLR2XhzpXL+zn5oJJfx
XGpvOF8bsY4NBbbwEVoxT2ybpmBPa3kwmZE4q9cGV82lY2VYktOqCbNZ11sBjYT4Cc77Ujlam1+f
8RcVhuedmO/UR94/dhN66qwOnKFhmf1B8Bp8QZ/ytltXQKn1Gc2nHootbFTVEfjjVrcE7rNVMbC8
CkLHN4JiGXlvpTbS3o9fLNsK14q8sCoc09HXWRxe+ZikrCqu9VUq+HIxFk+9jsK3jN4kHV9cRKsb
BFPYMELUU3D87JhsgKUwmESajs3cabmWi3giKoND2OdWonhY7KZaj6ADAFVCxwLxEb5+6KWFHQQL
UMJgdeipdm99OyfHY+11fMhPPQ/OKMrLUn4pvYUmZVoi6eD4ZK8h/LtyFMo32PcAD/4YfV0Ibzz5
2KcS4aSyfkFxD9y5WG84WnsbdC7iR6ntx2vorRPP316SZO9yDW686g/UdUI+Ot7st6y50++u5KMI
K5QAl7w2+gGI2D+s8HO7Bzzd5eIshk7OrKf/bB8+4pwR5cPX3L7uDmyGReDJCjG0/bVQqYSVuyJE
LPP21hhCxoKZ3dFbhGLGsZySDoZrBm8rth06OOV8N6hfMVLnYWrvxfELPAj8CfajYJQ+KpbYJ2A5
WQHSi5ef2thJiSZjkyvdBKquT57TA70XpFKorB/BsMEFQkoBMQGRzGzjfGS1XbS0PeWMDWRjXB/a
+hhPz7+E/H8RQzF6PRVDrVpAlRHvf7+ho/zsXdBcI3a1mBVzRxS+xRZyVgJNBKQWXuSbU+Mx3BZT
AfGWM+sWfczt15Wpllxh9uay0kuJqhUo8LSsDAzkThYq/KuUMSuGQXF407BgwJDT2t0CWBBZJB5l
WhBpSNPRv1oXp6SJ7YwMxkGY2gq+EDsaYGttuhagBp68ob7FGkOnA4ZidA+Eyo5PBClwgi9Udmec
mAikDYQw4rpe0gkD+fP4bE5HxxkJemwdU8a+KVx1ep1+JUv6R+FQbFcb9t4jy9LEkSc8ziLU/hnO
i9zczcE8sUgrFz8PjCbLt99+tPZN5/xc4xfyeACHz0m06sKV+gv99/6UnBRAxT3NCYIP6dvCU4kw
nn2yF8H54rJTJWn4Jxb97iQDbIst/I/4OBvBe7iTZ/mRm7LtFCQab4BKJYcDiIMfZSAcix9bSI6L
k7Loh7/rL/7/1VVmqT6/x9k73MkE4MbEtfqkkD6R+w2O7YdPn6GR/z9Bt6k7ip+hnN2/dkAG12ZC
yVEelcYScCjNKjUrvc4VDLxza0ojEgPA9timbH73Zz4em5RWbNpMSx+rkDW35TK6WR6IjBMvkQhL
AAWQPJ7jr0vZtpnHazJ10fsq6/kkNXs7LYfWiwevlwLOiEfiTwGKlYN3Yh7yf/Psba03C+8sWDtd
GbBNpOcH/6bGkwsWOHp4kzw1Msn4xzo8/Bf+9R1yTZOYtfanwE7NUTWWkVsL+Cb1OFTbRmuFOzp4
13qpH48G1jqnGBmb2Pchg2ew7u3+580pARvFO4yXAa/Cqu2Q7Y9FwsWKmxsIFGcZwUsfuQR933W5
unn2vNY8pVMWumvOm/6qSsivt9NFHzZUDMyRrrXJtn1bCFDzpGm4fd5KUOUFC8wKWrVnaEs4RRkj
dh2KpzaQk+CydYH2ngTaAXALI1Ahq6wphsxrMOkx/nTl45moDarT0TurN19AB9KE6rkyWfiTbJ2z
FvWpy19MpIX3vWDffsuMbyjjGWls9sTdRTwk0uKpyjnqCInibcYhn0nxcGMj/skMi6Cx5GWD5yZo
p7ytyYWnnxdUjYmlfSeXU9NNnkmPemZI5TGbvTAZ7HCwjmlHHKLiB+f93NPEXceEUy+XsFkN0KAA
Go8/nYWHDcDrljBUWbrj5sDfgxqvRWXyVL9+myyu5SCIQBF//DNPhen6xYp1uO/CleKCk+vVDjr5
PZ3TMOzj1iZLtsux9iebGZ0XBElTZFKlRRGiu5H9RjWifVHd3auhcdulLqblOpzvOEHpOUcCtkMT
EwxzcNp57RG/VwzE/OfUVov191YTLJKVJX/axcpvFzxin6fHT4ZHq2X/tWSnShLefQ9fhPhigSUf
lku9D0Jz7Ylqvbl6BpZsibz0G6cNVUB77TI0TFgrC84Gb9fAen7E0J/31IHppMOwpycrO2kALpzn
YSJXHzA29IcFtqKJ4mPgYwQug9ueZUZdERyzUXdCFYz/txntUKhJk6ErO6b7L83d8A5litDiH1q+
uakTA3DFWLtDKcWg29AIAMFrKeHhF7sCRQItQ6W0x/WZRPvwX3diJ8CGOsWBBidrXQYCFmxklhcW
UUb0x6gXDRh6wxgcXTEb0uCn0/f5ntzLLZeg2n9rOOsYkM9/oF0VWfgX6vaY4SdQeYZ6EclIOuat
/I8LBxfsb1LSgfmKdftFZVpFph5blSlWQXwOZd7AeFMl6CMzadZ7xZu/nWAlK1YXQpFLLn+a+6T/
uhXyuN295nwSbyGZTnF/k+FDic0Vpbqzi88eG801tjanw3nEWVeET3kKwYagCLcQVoXL5ue+swIw
cYpiaxaorL6POnJVum3yIURUw58NezT5KlMEzHCqvQPvvjPxnjOe+skreNP1UURp+NXY3UyZt1a/
ZM/3B01fSzNTJPcVqSJMyQi/QbW/6YSmBpYDnHYHyHibraPKCVd0ducfThL+qAVw8bSvI4f4dFeW
X4UJY0uN3ER0+15xzgalMxd74i66ppD/MwFLRFoMVEKLx9SCPJ0cCLcJ9yTyzQjPtOq9mo+XriR9
MIXuIuSk8PnEudLYBWLgN2tzpbYuMOuOkLRBHbt9V+JA7F3Oe/ZhHgqG4Uaa29DBQFe9hJtaLxT9
L/pp9LJ6h4Har6OoqI+fKyHnSZGJ/8KDeE0xv43CvjJiuXHe0YgM5dOPdtrrqIAwaVkenV6kYBas
pheneMz7MaFBW99H+n/5zfsC3B3gOPLz2zDtPAxhW72IRtIcbvBQl5J+vddnUtFIUakQhv6aymHX
g7Iju16nwtC19M2YZiyIn9hygBK1k7gaqwAiIHnAD92lFr0Jq4JY1FruYHvFAAoHPmuLFnwrAS5S
qAP1jTybY1+sW7GS4Y1BOCRRPoSbZvVRASb1z0nXBweWjlK9pDvfnsSFsU83j0B2hrtc/tZGJR76
IbPHIGJ00Kzp7VzIHMRcTnLDcfGfBQ+F87I8iscOIYPKweBF4IOuRbPzwlWrLWnSffmbtXoOiuYv
E1u+oGApcOJS3RkXEriPWMCoJl3fK898BjqBRvQZWzw7+e41djCpckn/yMhx2iH1ILsSw2BJPmlH
mVaskVtV6MaLniMolLP+UABnoMBbS4Ykb4IIki53nhJRufx0vdrTw82llB9gGg48zDzi1NX1VezJ
qt7aWJyXihar7SHmomFtxi5in79mlKX9gR0WuAcHHLAbXybSHLUxYs3Kq9VIuxUthuW/lyg9/MGZ
3zyKIHnmD5xYEahMzHgecLQPDYUCuFD8pK7AaG+PApH0t7qmNswwKTIiCqPWCkMgSvhj99LZz2Vt
Hm5hjwVZ92AfMp34ZeVB5Fwx4PFb3z9127bTnJ9Afuxwag+yzGPSnipwoaiuQoUfyJRrZTm35921
sS9D66tOnpr7/fDIfxuUy2T6dxuBMig4nvfvBngbbp8XIwFS2ajuvaMOIyL4HmUfdh2H1iKLLJ2e
7GH9v+U8Gv43SKyzFKuWdvyYfNnVcR69kX1nRqFxB+NrvZ7cvMcUZb2PUP3daWO0KgekFGyxB8UI
udNVbK9mh6pyzYr2++anS98ex1AMXLZkAR0DNfi9s4zVkDQeCT13vuc6QLvQnL7IVSVJ4ubXc7hv
srrazWHUCNcURRU4R/EzhfJA6Sum3clhAjKxkVvQjBGihp85lzRY0vw3VjiozI5X6aP9VWYgelXf
Fbk6xs6duPhLHu95dHL/9/8bDHsl586k5yT5pHKD5qBteDR7Uo3JNzh4ms4H/GSJk+c0txsxdUPJ
ymIY3L0D7Cwlimr5yqCI/n3dlxz3GlnRT1MOzPoDrKUwqnrpuI/+FrMR73x39lyEjgY4tN16hwhe
khO2/KKUwrM9zbDzNBDjVxQj4ZlKHRB/aQvybk0T/iemXpTTASOvnn6+SBp5BxrxESXiXWVQcWPF
vvSqPPsppziRYBUe62A34sGiRQ+zeYTPyHlEUxM3AEyTpsL5Tv429c1FYGySs9Lbkw6Nj/I0prl0
mG0ST0COs7/jH1V0Gal1aO7hV9roAI33GDyqqgGqoXzEvUPYFlpY6ZyUXF3kuouVM7+ehtR2rj7L
LkvbSfKtgXzyceZJKJ18x50YZDPJV6BItlCyC3rbVmFPG4NIbE5AOnhRkSZfzqPf/Iqls6wVQBer
GBPMs+YWYzQeClr66f0d9t7VGFaiEyBt8P4fQNY0TVs3U+wna40Dkyf6h99anNiT4TY9je7Og6bV
mukoNShytbev0cFROMTykQtoe/WttD9LExjcCCH+hxkk5W8W1QBjJcGMyDHO/oQEATYUkZKqGBVl
o4m6ULdkH/nb0mROHnKvvgOYLP6NLN1qYNGyo/Kn/q/aiy5foZohdH7ZqydepeRlOz4xCxChbaXT
OF9wpfHRLV0kAHVi0zWaHpYKOZZ0TB5dce6U5+9jSZ/7uYRU5w15FZ4wZYWIAi7V3Os9ZD85KAkB
2cn022EiS0OBoxLp1IRmmOkjEz7FDQ9Al5XkjUd17kYoBcMo4bj17fWs/cPpMlkEQfexrPcXfky5
JnYghC+CytudLGZGJTT5kJQRqQrxfPhz7ILViCnkL4W0b8n/KSpcDhfrSErfu8hbbEGlj1IAxmSj
WuZ2whhwi8Qtvj/F9ORFJJy8GhmPTH50T4wxAmIdh7aOUyyXsqITpwkj7gBZrYNjJGe+zSgaGBUb
C3Hz7bE9IA/Y202ixu+HycwsGpEumzkvnTkJiOZUkLmPp04HpF2BlvoP/YivT6s3uruvO8hovHqh
1IWRNpicDC71tJZOfNOKxGSIPuH0annACGt9/KFSsQHeZ3Hv4stv8kOW+qiicoLugMhyO5TIlgWD
q9Cs6yTqBXC2T9pn63oO1s4DXmQ/XBzRo0HZd8A35yyJy/Rt04WRfwyij+BhYCwgVmxCmyl76M1b
ncKyf7groAk9WG+hUpKDl39oNsX2GuGESNbi4OvKM/lT96ss1NMLmevYdaQK9nDxutxjDBVEOybY
bmSBaQPU2E90QKCdYccAPXXOM1Q6dDn/L5HwsKeWKpT+tzwmZ1zfzx19TZH+PC9QYJv6T0WVGUvg
UCdMHdBcq7n5MicgTdVKvcvPlsXnQcsWomEhcQFBdGABfRjnaijObiW3Gdj7yPgxc0UBAiyVdtDX
NnG3LGD0EvO8TgZnwY+PODqBbFwlmMvwYo7s07w64K+EY8agPsNRAMnhmWTNK8c4++46zkTx7auQ
uQSAkhCxi84EfMpI0xsmDCn8xpsqtC5dWktPK9+6z/LbL5dDlsxnH/cSQzFP/jv3e4YgXsgE5/pT
q/dSqt62z0zht5f66Ify/AB/1YX9Lg+XJ7pECZXs4L0GjjiV31j2EL745lXEeRjmVmRny4Mld27c
RUe/Jfi5UkumMrN6NOdxZ4kw1cs/UQGUA4cFDxwyxWzz5b0RUVObxA3ZMw5LG83SOUFc6XcxQwii
vxgSw9mk1vqRgPJaKEWdPfplpcM9RyAq102MB3gORFLAqdsrnnqCgBA17H9ugkR2zoxLQM9BkQN7
5PROAYW6otLXGrWxxAE4mvLc79ILAjXVbGwrU7ygR1B+s6MyG1DSG/AK4QxYqs9gxSk/KmBhiGQh
r5Fehg6n48C1jKExT7IHXhNdG3Hn9K+Za7AqhR1Fk9XRQgn5xfgP+D75M6oJBx+ho7px/roYfgIy
OGVSAMj9WPJTf7DUwn/0NPdmy332kTxFRiawf+dh3g3x2N33FpMyh3YXXXXEfNwxqWPlkbv4rlo8
icAsbppjXBnaOEWV0mBeE7zSHuA8Kb7bzcLyBgi31jtJj7JqDFlnKo5OnVYaBJmlJS8Y72XnVHaP
ElLxA8rgXgXBHu8Y6qaSy2JOYLqi73r1hq0LVpKr261XWo1A3+RrjwiCHGj9b3x1JUk/0TJTJ6j5
3mF4Yp/jtOPulbudA6uNxlq4UYOjuZABneXTTZbsBlTSxnS2DCqzrt/2JanLgqOO7/K3vZG84538
6zKMV+xt8JRZqh9qR6AQL7iPuPjZKgDS0WsK0RJA92ziX2GxN/lHePYGIyeaznH+tGB1Ad+EqjW7
+4jIUIdZFFUrYhg46aX9kJqTCer+2EucE7lB3C4CkfNvyam4isY3McGst+4FUrYEFpYCCaWdZ1Cf
RGiFhEqw6/OPEoKbhNAn97HAil02W5BFP/yly6/UYIv1Ek659kokmcH5f6PLx3taT7TZBYhp378h
GBcCm89T5+i32dFcDalw60ydMDd+tolPWfYUA0oOJEfuxQ1YOa8S6TJwS6s0JG2s5SxZMBTbj8LU
JkynMP5As4KXzOCB+AiH54uyXuSt8SaRO6T4ay+Tb7ngGAJHy/CW+1TxTFkLmDKBX36XiF4ocTMC
4WnrI5NvJt0OU8xcZgTFUKp+Jnm8zPCJRvlZqTszvKC9A1kaw9TKMp5ZO30z37mwQfFCQQ8kuT8w
WGSmtUhEna8MGXpRS/9Psu6vgK2kLhili+q+94AtE4ka0Psp55llEU5ped3D8sKMYvG/E6JmcJw6
6YauSMoBYDDDl98kg3vfMzYk3DHUUUMp6j38sqGpSzB06f68lxTlkO3Xw4XqKWlKhGnrGslcfOri
k+BaOTh70eJukcAvLwFDE+DxTXIC2iVtQPdL2N9Xgfgwy8jBgn9/tUj7+u8roFli1Ao2KFpEcBnf
bBzZOraSXGizJVZzuAdEW6RAFwfs8Lp41WoyGIJrH0kaEvPq1ni1ovNkKYp7PKqe2CzP+vEOC+ww
Hl59Y2uc1pEpKO3EeSTofI6E/nCvGQrffCqYuCojAXeWMSOseYz6x/pAPOugbyUvzd59Y7sA5z2a
pV0p6DQS1UbAe94YNbkQCU9XNmoT4oecahDn04GkbKa6zuaiGTZmOaGlR3kV1g4EtrQon4tEzBLi
qIcO2GGEtWrid7Kz050fqnbfhhzeab1CRcnqpXEF6u8GEailpCj42BNw9wr5TbOtxgt3hui9RX5i
fL7KSNjRc7z91I7ccumrjIYs6SfZi5XoNNXdR55utx+AJjhlosUH8f+nnbPmubLokhxbwDUb3FXF
AXFj1XQv0OUKxLUMUXD6mKFD2+JsxbU+IqKFIcypt7tEQ1wv3eM5yV7e88etUsy4PJpsd/LNKO3T
77DjYJ+5pTPkEa03zSu4f6ohrhCjngsek9m6rVs78VgCVXxVAPw6HLEA07KhWSUQv1KmMnhVEeTk
+lGFKUxfxzboHln9/8cVQ8uD8bQdCZ+COVubV5Gi647vdT587x/rJeO4z5l3GbX5ZcW3stkUYyLv
A/YwKqNVoAC8JHFDFn+hGf5l6HhWCnMAnv+mUzMAtZMNvUOOVvXlKHOhizQwVpn2A1Kp17hW6B6W
2RzGCfVprnHq2VkmPQ8S2BMtvQ2DEubU0Wht/8KWMBpL9omxn+wZPbmGiPUciEJifQ1vPCIgj9Hi
qppyFlzR57W+be3I3gOKBB9HQySMFT4HNZ6/Ww1EoC3ka2meJXue6+wRHKLBXI+fBX4hxrc4quQn
h/N3HTpKgQl5DxD3vN52E8kNbtZQMbt5T5Dde+sE9UtbD9brlsUnmNGn24UAEi2V/PtdREuHlAeI
TUsG8dmAsKqNxP8mrZVX0x9boHQswpy3hhXh1rbZmolth/fxgNoIz0qC2MvhrNzmHQU1hEhVNXiZ
XVFrM4scT9/hdffo316UE/M1/YOIkidxb+o4AXzVnc44OHT45vjXkFc5qmBJ7IZbi6uYl9DtG0ng
XMSF2yRuuEe0I3QDisVUc/RnihVK7b4ZqAoSQvEUEKwSQJ6Tqf9FeKmF6CTjw6isuUq48t4VPjRa
g9YLOaT30dKuerwiynhy7Z3JdekSY9VUqz5nz6mmFyMAvzpjawrXEszUuhfNW2SC16dHtl7b0cfF
a9O5JJciHoGb7oykr35i3hjaH8jwDdV2YrBU0unpNcZYzHbCTkcO5hLxvYItL4flkpsbHdSzTZ9/
qXrzJLtCYt465ZzksnEDJaEcdupKOh0BPbRDmyvZa8UTMToiNI4878tlFs0EAWPSinfhbaa0RRWM
oURY13vWxdFmPG2krLn5m3BeTe9Bl0jdtR6EEmzU7832P7V1dIrisnJYFdVhz1PbNVtOBsEkt5/X
0KAVuRG0/XzQSNu3LSGTFasqy28dANuF4z4k9gBRDpldCkCto+v+gNxKKsUKPVSo0mLw4Fy4Bvd9
41JvRu8Lr6uJKNAdYxHzRynb7RLvpAJq7+BuC+NUn1BkuUKDbImETbZzwaOrS97XCZpxWZB/8yfw
8SAAV9y8D4O1s0P5ZJQ+nMlXJm2+FQwiUo4ooEaGOaPWcd2j5vMQIQpdrwBqA7h70r3zrG6uuf0m
J+Ka1vfT+NK/jxgHqMRDTVLgRwqUl7Pg53hie8aIEIdxsu2eqSu8OdXHqZ0AMiW33Wi6e4/wJuGd
AKc4D/uZlffyLzU8aVmoBL1L9j/8E5NI/kFyP8mSKuLEO6j3g8pNCDUX1yQZisjZjUpB67MqiqCN
adJ0z0ofrAl6PH8fWQFPOUN9NCoBEG6uOCCKowFPy7yOJ5Zcbv2OwJ8cCmIxLpbNCPBz5IXYPiIs
nDoDkYUZU5OWbsGLOaj5vV0upPcOi5h9V/VIJvEfBNfNR6vPjmkD+uXoF1x7FXdaRK0cqHeKXaw+
X1JFeWOKIFV09oYHUu35ogJ1GtydBSbP37pe2b0PQAjAAJEhgIdjjOw7LeGLlVTrpTr4KQ09zoa0
92ezAVfR1ozbwwdqiVB6fWVTYbDPfLUT1BJYTFeZVLAT5AbqMpzLweuzoD52x0VAFGCFdxmtH/Qa
uXCEgCWFhQuz012Tkgigw0ZEEMBoPenUOyvbpTqq+MoYhk1GDA78RZmsZkkmMnElW+0UNte2+86z
QKXtHznacBLeKCi9cnq2k6/48fOTlE3gJsuiTyBbRRMghPC7Vj24O+6Ds4Nk8bU9Wcp95sDSleSD
hydwb3l6CUaCF9eW1cJgXVjlFSrtw0Gn8yPRAALXcyXJ6ax5mLjc5WBKQ6z/EHFourFwBlE5hkVi
3N9sqLwdESw38GTE/ICHbR1DKV455QAuLRua85PRz3uZpTdPDFQBwik5sCALVGb4CxwAe7NH6Xp5
OwUrE1eqCOZSeVNvcwhm1F+FE42IRUTwvbvFOTdJsznk2U6y8apNO/eMlo+bRStdkPbsiC+mHoXL
r5ptuIyzh9a9QOjOKVJDrs8e0dXztSnwVrBurDbFPar23roXevPVlKNbIxK6Qf59/0AwTsaNTSqv
oHzUl85ipNhqmldvFlc9sNwyxaBT2BGcwaLid3/hrocYEEObMS7dGVR5k77qi9I2Ck03AaDdY+dB
h2KKyp6U+aAegHnJCSyXIGFoNyHeA6g5eSZPfMAj2QJC7ihYShA71aqxzAKBcGYpcVbxnDn/sfIO
UiIFq+g0JRgoXA1OCChju+uKFP5kXHnwqeb0Lmr5QlLWTTffTri/WFUFmWG5XGhTQZ4Z1Qm7Kear
6cW/+a3y2PG1BYn1G/Sf3smH1swbXTqIq9zmL/dIuKv/EDA2sHbkHdHgG47Cct4fnnM9Gb/imzk6
SuR0FD/+xy776Eh1ULSq4T+bqPbmULnrPGJ0DpDMdbZTy4vLdHovFdYgITdjkzLmWLWV9CyJObdA
4VYN+InXEYslJhOnoVDjBEscF3YaarNV2X14ZwSw5y0k/IFlm3vnFNxWfIPgbn5Ooj1TlM3JTgYF
FdijIeRbLe1Mp8HRwH19fVoXcUNdTIly7Jzw7hJnnBokyBjDEbzTtXT1byWnouuuh2URex9tAwVb
/ikbhnBNoY5IFjIncJjly3jPpVjt5mq+YaqyQRaW2t+I20NoDiosq/fmvlwYzAMkF6DmfNLbkTFu
EYtGUlHyVzlSq8yn47uCZONVE4/80mvoSlY7NfQOXHDeEFoZJwFDmNaiTO62D8M0gG0/X3Rbt/y2
Ob6L+bAR8/B8ehFQTRwVcAQd8rav2GCsaNret9+hX8ZPO2gsevVxDB5e0Ua3Q6J8zHZfV4s+JVtD
MpnS8siBMVP0SmePT7MFgWDSNvZpTaXnDcuPl1+hVGGL/E/4ccJJpdHZc12/VcCLY6eMh8OfLHBB
gFV1qNMBmo2h38N8EXUJAWT0+HXuZNvD0KDtxIPdyDLzA5Bo+gPep+j+Rte7KgEgIMktOpJno8mc
th/3aMpMrDBN4KXAcILv/HxLWIc0kwlgIWMQmEQw7XEyXaqd77/p6rIeee2E25roax4I7jyIWnVm
66KpVKOiaBR9LwXSvHOVgmq78p76AsT6gFFTbHhRojOg0vAhSQg4Z79AANfglVDARInoKHlCxx2g
4BhWDwXx5YXgs1begJFVhkqrJZtx0VloOkwGIPOzxu/sQz58ol2PelKhIEkoAVbkxmLCnVSp4pU4
cLOFzl+5qi7KWKZUa1drMHS3nfL5ncGA+hlx4nEYNIq1LQ2ihlc2cppXmT5uavu1Xd7TTZozNEhn
qUw2XuZakalv78Axml60+FBZpm41YLBJcHpeqUsjwTb00qDNglVWXfRGeN6aqT32ZdASxO888a/B
JXnZPQKL83UbOWWfyaPDbZ1s2AIDoYvWa+E0ZhStd/GWaRuZRtTh97l9gpsSNXDoPG/g4yuPN9Xh
UkJtgVSysV52RNxShQbYyeXYwmIzsS93L0/uWOjjVDmmcHPvVKZlrB/BugGntqFnjAjvkJMErt9m
4fIjST5w4qLu+rkvdbprgXlYVKuIAgIxLoiSCRLkrsm8FRLCZ2p8pIyr5FzviSHc5nRUKnrfSBuY
ze2+pKeeZjOnxz5Ik4VQm7I9P1sggq/QFXqqZrsJ+MOcMrzToZERdEFi6j7H36VZVkzahXxyS1Ch
VST8cOl2g36Rgt0cLxFUd1xtNiAaj2l697EbQEMymEgGaVHCB52hyfHwYgqViQxZCfJ1uhpxbdM2
mghModEAM624qdHZkiLgQhoemmExh6BjaaR3thG6Zk/Jknko4oYCg0tQg7mRxrBS3vspvFz+4RXE
1KK5Xg8HAjfKsAqc/H2t+/wbP74ueWm+6IKmcOhzTxI6LbmABHPV7E8AeFZDes95gmO4+1vUoKCo
UnMavPtCQTfnWY7flCcQoVyYwXpI+Jh0UJqtFW42RkjLmiSSIdQX3+vN8ervC+bHMN+kBp2qAw8Z
GtYJ7O2wLApqMo0U9EfUjMeOSoYEhYXeLThAdYpdxBmqCdkHt7ykaADN/U2IxzyM15d2jKD+pnYz
qn5lxAIrZh+VGlB7Cknq4e4vmK9Y5RW0nS/Zc5RWC06qM5sGS78SO7XzHLSUH2ELQeoqbJzPhmWs
N9IJm5AkMNYkjgP24nYxp0A28XuYa0ZmRFkkIN65aM1iUalVo6Y3i9oKaDNbbMyosdKQNK3Zr+LT
FbrUVmxXqAtLYTUEwPgnSl3zYafjssg3Lz/zsFSdjIXsiSMZ6GInKJIrAKvn3o4O67pbENDLH0UG
wPNbjGvah9hVu2LND1XdVC2zBvyT1zMKxlUnbzhJod+6P7H1XAgolIoSQug16a6XqND4BjiLwNVX
sa+4SIohX6qYpXFgogikQJ+h5Ph1/oq689pbN9Uuf8gZ6yF2agYISfA6Sy/hp51qggrNnvbxN9+b
+hYKrgZtf9JKEzZXE0gwey19PcFMWhggIckYHumyYfxmCKDNdarBdwFA5Dq6Emm5Qyg8XDsVXCit
SPFII690f1qz3dZnQhsfgE0YCjv3Pdhenm8azVxDRkzbsYLilW6mT3CCq8ICb6qDtP/PS+2QkC1E
StiVJJ1apygmrL7UMWN2Zy4Oa1aQ2fnoi4x1pj0gBz8AsQjSmbDi6H/W/m87ajMmYAxwdjkrTaY0
GS3Sax/OxfjpaBADMNjAMnAto2G5q9Hp2JllvvHmLq9YbKQxnJWnw1ChZIicyvCM8rJE5skYe1M0
WTXTEoV6fkW8rgnSIyXSpnewtZx5TCbjWXsu8oL6yPIE6fh0NjKUn7ufxeEoNPOg4ySnyCE1i7Fz
ZlXY2Gm0QRyJ6Z2KEQEeVKyCvh6NTQ0LpGLVWWKMEx2/lHXJiKsVncFBZ+RE7VNnGB4mlMnETSnI
8K9lRFiWfJz7p1xmlfWwQRkEqN+SczZyAKVWn1tDpdUc83hMe7d/0aJPMu5RMxs91jDVaR0jbWVw
+US7yJvSkopNjlGpodYT5+ZYwJ4GKDpbrZ3uOZM4WcN2/a+ZmESbYhSrgJ3uy/sQkHF33X4t56Jf
T7jse3y1kEPQ84PGnVM3X5ErxaBkTNiqVlv2fmL39vuk3UmPlTMoIPcX6DJSY7DMMzs/sQczBYAW
RcOYAjhu+UkxUNlOQEQqu4GFErtexyci/0p90ivGZEJIOg+Ulqkvpg4kzZ4O+ONa84qeg/v2U7S/
GEqlYAfW/Hxz4M8RwkOBRH5EsAnPDsiqKn7suSAN+nAZT1nepFvAQ7CKtMV/w8yf3+7V4e42twT9
OnRVAGR1Oz3/+VkBfZPak4lmmUeKINQ9jdcqvioH1Ik5JjrEa222lXvfVGQZARwSOGH4Cm5TBvm3
FrKziWUX+EYlRKj5C/43q03CDfaNK3IiG+gtEh/v7/rTbXWJRb4WqVtA+Loh1b16uRbqFczEcpzJ
Z372XKgk9fUbsSoUjBmbPYRTIGUq2erCwspu6UU70s77PfQDyY4PQO4QPcD/GVMy3IQBCbRG9o46
EvYoxooX3GKHJil0LwN8YWO15xDasV9MIJ4zaiwOD0gcgQHIurlCN+Dss6d+7gfH5VgtET/36jjt
QIYMWO9WRu4zCn2MFvYZ4WMHsZ5f508BKQAbHSbtjshMrfDzeezfWa47S06WZjEuxcFRiUJoVWKD
g7/80JANjs5FKRZMp3RH+iRYD7O3Aanf3hVHiKxUzWFNGRrdVyljePht0MDerh6yp66uK9T/DpoW
W/iOz4/u3VmugCqVxYPOahll1DIj8hZRBo65kSA6V0dnsCfgI4WI+YvcZdOfS/ZQfsw1puMZShIV
CTinuns9yu6g0wW5oKamZDHbp4QRcdI7UmMoew8c7vRoQLAtuofrHfft0jM1t3cDsDY6ra5GtM/1
cx7Yz+HyPgZs/cvuhxmtxN500VSpMnhQUboVJ/BDNRdDnFcgc2NlT2YxhS4IPKd2YvpeS6JNAf3A
Fm7XQE0YL/c+lXPgjabqvHD6A2Dz4X1f3JSG73ERAlZUYVIzpwNK2FooKKwxHZp36Gf4hhHNY3Ok
wqbTQtdGaG05KMdJb8d8bBAVcIv8TZhT1r1+0eVDLLztVbv21WwHGCqeZCDk6XwSvHZDBXhqgpMl
aaoI/+CCbQSyjHiya4gSoN31A3IktiZ7OmSANk28T+MvWyFuBW2JIdCRd2uORddxDJ830/SFSnke
uxM5VajuePAPiHB91nBCCVGa+qZ2rbxmVu5OmcOUom3N2Fho4PV46klxhmB5tOAN8qzXXZyD+ksK
gfhjiHrFklaTVookLkx3419kJjc9jgME43nL7Erpr4RHrPGI0KnrBGLbxK9XGJS9Y1ySvhcE/vLy
EEJFFYMSxKwWJRkLWViZlCC2ICPtHru7Fwiwy7R0obKhYXy2C5YZqHUP9J+hL4ntkk5Tnr1rk8cc
ovE2Feyxjy9AD8yAamJUuDsdvjXGdASd2mxKUGWemp0wnFV/0jt0CDRk+f9AGL6sKR1oVcfML+PP
SdsypdJnHH+RggKdpXmyv7kJCtS2qRCW0AweQuAZ7bZPUwoI86sMdnWVn3kPvBBOnBA6nupGmkb9
7TNmsrkSCcToQI0pGUtS2RLrHv4UehNAepj0nnO4LLs3yJCS0pkpfJOucssOOuJKDrhWA6EkaTJZ
L4+R0LDeEpz8sgyG5VDvddYuiErK13f56k7L38ehT+kcZMLh8t6zpcoMUOJZjea//8naIvXeFX2P
IrRThWVc06itFoS1abFIblq/99ecg1vfynCQ1Z0iHaG0AJAZsaNPM/R/BXzKSR+C0Bw86qqdky9A
veuomNGVwnR8bqKRoACCWqzdPBM3JtFBfqfH5W9MnEhQhFe5O0d2I5fnjbEcgVgKO7+BU5Xv6Ysn
U1MJ8xq3PE6r5g3PySW/QoTKZwLUmVR2QcpAalzZJJp+JAtHZkKjqVSiksTyjvbmsHuBo/n+2CZF
yXpXMTZlgfzonfCZG3NpFfXpy9d3ER9fY3dFLT2yzQOvx6VoWlM4ZI+pY3G+ZigROh62iOL6k2Uk
9eUXYrrbbxpPuOWBQQoBFN/m7ibUQaQ8Rykq5XjznGZek51oo9FbWmN7AZYXxuPsYVlD77EzBfPy
TJVYzb3mX8GAkZbLtp1xVGqTvot5lUVDaOnWU9k4yXiTnhmwM8jwRttam/lWBkSLs+Af4itk5ggh
/qGyYlmDBhGKuGqe2x1A0Rdjpul5BjZl+Y682fUFoJblYgf1WkO7CX0XYQzO0DDhWTT0SsqbBNxD
2SVtNE7IJ+9+PtOVUrNEA9K+5D2q/8UCOgMqzdV7o5WCyobqAHcoPavvb3le4gXQtjsc1+2i8ENW
8e/ldhc6a+Pb93ArdzD9y0KvVjLxRkDqzCerWu3GVSBJoTQNo1J8ZJwb/j24BNsenCb934rteOd/
B7T1OAGzyVE8bbAmH3B1Z2sU2GRAPL34xI0wR3ISfOdrEawfG/CgMyvBA+6YEXKI2PyHMdVYjCTF
t0JK8NqdyXhdnZq0mUbiEnAKk6+0/WTpJCFkgfODmE3vCaJ8qgRCx62SFXEutC0fGb6fjonOSiPS
3GlS9pR87kr3L2H+3+Pfq4juiIYaaQ/6Uzwq+KW9wQryZkx4anEi0FS5hMQgpPsJli0jM2mt22NS
ja+HLReLBi5L3UpBJXg9L8YO18Na4EU2w6x0MJmGZtnWrKh4S7kjCE+tBkANOA0oOgZ1EthTGWx0
zPCfRCVx/jMWzeg0eoJkt4sJebGkEbUcFliI2ZHcHucyfbUBoeWFK4G/8USqcJ4cMhyHF+xJ43dp
Lknh/u7wnZGn4Rap8ZA25w6lKGUWQ9lHyPVAmlCV1YobsmeHF7AkRM+UvNRiSW+NMeeY0aLNZBcj
73IfqT6KNt+mAxpj8nBxYc8aIPnzVjAwcUx6DuhCpj9rkJ697WvrJjtvOArqYobOcVdW/2qpjaOh
mC3+6T1QmzqYaeAIq7xcqA/AaIJEfG88hqL5trAT4EHJ8GXHRbkw6v8f297XWGKrRtABAor5dBnY
s9+KVXSJ+d82/9TmpENyEWVsbHK81Ory8I8Ls+U3x8VE3ECfZsVyGl5SrevoBvKu0x56A5jhGd+s
8r9+h1ySEVH/gWNRWByIG4AEvWObxGdLngVh+LYt+16AFjM4yPJIKJI6Yl+UP9vBvTR0P+/Fn84k
9yJRij5YDmbEm0PhXg4lPc+iCkvG1vPcAH5XmEmFjOd/Nxbg51lJNilYTSMHdMq0ylZHa77ZNRAR
4g25apdvbcruXEHL1OOlHHh2xsg20UsdRgx4ehW3FPbiPz/21mb4Qnc5N/88Gr7nJLO2WIiYSmUq
GaLdigEy946tG9p4MlPj0ZXf+uyfXKn/eHQhHoseYRSzGkWu0mOAzwsRsq3+qSpfuQAFSkvcGPmT
lOFY24ADs+qsd/nq9AffA18ug/XceLY0bX5XpkyW3gTlyuZRCGtLNmOo5IVo2xe4ta+zULDW3fKJ
oJictVXu0aWeUmpG6B+00ASxF780Huq9CbLlCaAVaof6IXeUIZA2wqi12sj9PZN9Ebodsc3p0/KR
p4H1mlpueo+ahC8JWMmyHLdm9PUow+WahOB7ljgodIsBtfoRMNeoXqApbjFt03XMzFGTp3UwOsVO
z++pdVx4zEaAEYTxohzWEPlSpkTohDabDB46GoD432TFAJYSvGq6z545MRJ608S5YYZgf0iDg3QQ
aDQ2hjugo3Cre9lhmqKeXZP/6sQlvWeAtPrmTTttFcEv7dEyAQeCjdoJvSttmnElaMn+Hh7abJyP
nk1iFwa4pRwjzwFJalSUYQiRtx+9FwFD2uPnVRKLvggDAujJ/93S+QMlA2vN/OGjxkSzwOrMCZd6
i4CS7LgST8g2OWctfpcqkyL4O03adYwy3wxJZVO1yN+imG2KJDQZtDDl9Q1cMtGoRGbd9Frfd+4K
KxZr8e95e/0KDzibOeJHsk84vDjjOby1f1u8AarRyn4Wir18SGz4wE/dOPFbly5GlGFEK9x8fmqu
oWf+WrLoPS0nkbxQPTaR1hpNsqEMycH93ATEtCc76fO6/klGsh/LFfagBjVXeESaVAtfeUvaVA6a
ZiWF2EzM4/yAv4BF4+hIr0jFGHTt6Ozn6GpoUFjOxL/W+Udr0e0rkyDBFxWjSsudf9YvK4kPhcVv
tEANZ/V30VFffpuy+DuNMAdoP45kskkbgBYdOtc1sV6qya4zN2ljSwdqwadxNj9ZeQuHrsfUVOzc
ZgQvGTuofVFR/h/O0EA9F5Xi/xocecX+PsW/SrZTnHgz2T3+SpUafRE3dRNm4h5jbov6fPeXCM/2
PZCWV4BrSKX+h5ael4nNRU+JoD3bAAqtZSK6kXnnCw4S7FmGKiwiNM0dtEr5c9U7f/bYjMojl7bA
xP0USltIFZzaM4rqcxxkRbn4XFB6gZ9N4guGhwCmNB9lDW4gBK4bHp6bi/+LIC4p8EUyWVpKENRg
cjErsTAaUCnUTd43Wa2mQGf7jHdwPEurLqE3MV9INDVi4BVZuljkMm67YjB3NmjsrpLKCndeywyM
rNFBVmP5ev7rCtgRg16h7hFO34xZ8e947FtpTERqKkWARGTnRP/UbYOLaUfWKNDh2hyBuz2T9d3w
5TWeqhzxfte1BynpGOLo68HZK9OCh7VIOblz1UpgtkYvwc8kSJz3Fsg+Lf1o+25cNxCZ1ICZ0NYO
Rz46G6i9mx45mWa98sqKy6MHcVKNv1QcTNiiTU1+Oj6suWktXGx/UWsr5umGw2Wdg+oErxgv3MPi
wP/1OZl31x1yyapmaePyG9EUniVu9HmUB688Rz5pcf65p0ArEICOjkL35JWI1SyPHUb1/BJqlioY
Hpl0MyJJERNJzWp1sP1l8lSe5XeTRUqA9gvaPIWfCSFxTlTnIc6qndCiPAOFPeym/3Yvl6pstwrA
EcztRUKkFtbCaC+F1MLXH+kv2tOA8nOKhjhzn8iqNi2xpPJ9a4ZYYzHH90ysiBbTgBnHMvF3zVlM
ThAmwSXQy+AKdGRgAQ34DlUXc08Oeu6cwSmyyUFWN2wl+fLul021x/rDMz1PFWXjcvnWIZsaRY0Y
tNZYzqe8w7fFn0SwPl0te9OeCMo5G/G4LaH3ScQSS3aTgXLe8gRvwaMJ/3wYvdg9TsV4XbVK3AUX
xPzrAc2gL/cuOR3/lzasVS+rItuyKERBG7ktGuTUDyoYH07L7Qv+D4VQ9IjaBHb4MwUz/DvOnzgI
fAe0FrM6GzM+KxDxnn2Ia/pCO5NOHgxOZ3Ok8HJOe1XzVYQle6rNdL5zljt6ZwfbWQ3jpJN/w28A
A8a66JdstSc7PXv0YIe47INtUKoaK3xeJOwtqjNd4j10MwC8fHDbjw1flB73iwFq7Xm8mhPSaf6s
NgAshSfrHVbb/BWdny6CMRmGfeJ8h5FztRbag2rNU3U/04nStGGbT3xNEdmjn5+cXIsErDLGmvtN
T4p6+ON58hzO2WiFXtNG1m29wFOciZHDwaDLTzbwPVReF/B4URQgWnYqFp6gKPZXvEXb9e8iz3IK
9uYt4aoOUQ6swqLeP/bnxvw7uw5HIUGcz0jeD11W/aAZkqINp6nqjclw1D/5cCmb4poo2bofIjqc
czHRLdUv4UywlYQlvQM2gGy+DAuZfmAwbUJlfLiL1GnNSCpoTw3mILaN/iOkqwTTrq6Ri8oV/KRL
bSxPmseiNmbs9d1eKBUtTSy/JKiTfeQ4P7cb0K4pHkqBsfq+/1YnnOPfle6OTkDHUTAruMubG7Hb
FLNEQDHuZivKVmqB+XDnkPlpRQIimhfGpx7+3tZY9JjcCTn0uQtEzHPBM7MyREUztXvmzXTkzq66
/7ZtUJMAl3KJPol09lu/wl9ZbHDLRzNbNMAoL1qh13Z3Sw5GpMdmJh4q9zew6mWCl9qzITJX2Ui+
BfS8WtpZ32FXfo/SvZORCFRmI9hdpjI0tEdlorrJxTl5wUs+vu6Qay7N0mm9By/U1wrxzJL1IliE
lYU9ImeR/0K8VUdGSWR5Zb95XEutOHMKglW2A+gN947uho9qj/q/I3uXBq7dN/uKZNJTMyoBhkmT
KNbF6JSoejSgLSBMGFgEkyoQbyiabODBGyV+gNcWoIuGpfMr1G7Mf9Lk9Y9GASCCgjQutZW1j7hp
/VHfqNdEY0YZbY0pIzfkqv8UTHKwuk62Xcbl4dfBLfj3gEqqfY+BVRIFO5Om7DmNAQFYNS3dsHTc
f1ywpa2SOkjYeiNlvQfdwKNd01xg6I226K+cxinhacVqTDZ6qmRwfgILHMfzyZbGZrS5OJnlbYGp
8Ne+5jV9cyrapUSChBLjDl/Mws9WfXDIePlQXKBzzaEsM5pdL6/51QstU022sNqaMYu9CZ4JLlCB
vGk3rf0FJu7HGrSa5h5xd9KoaCZnUYtSnpSbd/yoZftFyoZoM/aQW7T2OMNR5BrDiQNYkplHUmCN
wfmsP7AIxQG9ZgroPew8Pg6VNH5KqYkjJDmo9z4a/6jaegTGryfMPu/4OMPcoDigG35k8ewflCe5
N8Netud7ewF2j3cvDc1Ds8qt5Y0ns/+d6jx7oJ9cjr/AxtA4ON8ekfjkzxBV1KZ6+B5ehT1Yygfv
52MtD+g1qzx69JuZAAiz1E7pyCdEIiFXqKWnvCpGsPG97kli7MVw01zeeaA8D+/oczEMIAvRO3nw
l562oyTLharQy0yKt9msYdJ2I0XAP5CXSQ3I+qUmW+ol8plvYWb3jKBydCvxoepJIMS+sq690scj
V4HhsYJFnLtXmHRJH3BncCafRVUwVYI2R9UvHaJ1G0LAhOTeBb4YMmARsI8cBut4d2G2Zr+wvMPl
PXAhSHacdZdSpXZ8sSMFBGKolmZp+WAnQWHQAzouQZSy42ZM1yyF0V2L86rtyip8Ib3KyPq5nWqT
b1pUgzhHpIP70z2yQcJAV0YjZa72W1NCnAzn489DWRQzwNuYnwEFOvPO4Vw6lOUUqb890mnCK9B8
E53nLSJIdNd4sI64nWhI7FTYtqy35F3faB/rYghAriTTlD1ZFa+ZtFpRbZr5Kigz6OOZXPLVh9g+
hFoNu8P5lkdZb4pxbNsvYM0c57WBMOtqV3tvTDEgr0aYa77PabzFhOB6zLye6g7P1QPAT+pI2arp
oE4W1vWPG4k1xbYKVSUqwyEGrK/Me7x4CeAzelBB/YiyLSH9x2qDrrQgyX0l4C+LSkieAzff3dwi
0uGSRKktVm83GZm/8id8MCEGDArRD6MgshjnFRytKDNNc2Y+qqfboBMvT/tcvqgYpwlgktjUHEg0
vzbmEW8pApLaqTu/ASxkRd+t6IqaVOO7EdNnymkQJ5bKozli3zKVWfZ+JP5bv9dZKPBF419xj5df
oLrn1OiNPNGanYsZxxmjcJoMRe+SpYgwNa/Kd5UK+yWXIULaqeG+1YGxWZo/bpzJV+959rteODGP
NjqOcLDphG9NG9mUOXievGtFWlbd1rUWaUDtgiA8zow/Tb4q9SFF8XS8jxyztNiPMEXkM620zEKO
bpYJI4hoXpIeFWv5xQ3BFSrgFxOSLuaFIoChZc2qljKozA67C2XLfqPDORdgidcVn+BQH4X8zrwX
KXLe/qatE6leHPN9gatCVgsCBjmzE8Yp9mJYHzmH+TwopMzEReasLL8cmu4UXDrB32F1QN6jdAha
LzCgsiR8Vw96PxHvjDk1wz8GV6TCf6lk6EcNOM4/uULPi034B9hMbQGggbHeQ21585phzg/mxSCy
yEUomaEAJAbGNzveDRZKMiyTVEPmynksjnaJrZ2Xczg4gJb+KnxHNjBUcYVPbRArasYbi6SJSnLl
pPfeYzSOc7Zko/8aw1ahhAL+y7IuGVXTrS2IxliT+NEd0paze+6YlSFprOmmQ2xK9tQlBUP27Wn/
oWnHj05G0BUIH3GznDBx7MGr8vL+Elui3Q9LyRKGn00y4yxlGILDdLCSl5Vh6IWsjemU3T3SMss7
TX6FT3QGUSCgCBr3kgcQsCmTr2LbOLhTMRi9T1kt8tZw1ejEf09TeGsk3aeXBHeo/UuCx6TsEnro
5tjW+gAhlKKSqxa+jmz9g/Li9yN58AwZFVzt6pVMlItSmJ0k4VE1QcWjPGC1PkS3/RzK6MEVqXL2
sDUm0pD1DnVi6xazgRjKsyK8iYVWuAGmQd7XeXt7V6lYV2AMM0dZM0AaiR04NIFXcHSQFT66CK+g
XRrpBPNP0CFqMwuFhwgZrwWc4pJFwlVULQTX8MH2sq2w+lOY8n8k1XsZyCD0NolFqk8sulnDRNib
Dcvucne8e2DXXR4o8WU6aASD/WEmgFOgyQEIvw2RqbfeZmY1bDwMUH8O7aGsQXHCI4oofi4nhdUz
DWH18BV41Bb5cJCok4JgWihsgMLHzoiprirLNmq4DvxRk3HJhczWEeDDjc2U7uRciZHhsBI5ysDT
BFYnq8+04XaLrDMjyPirK0H7GFd4wDTAGvdDpeKCAhY5j2HJK+mAwQWWPZlOVbpp46Ia5sQZIFRB
fcwio1IotVRgGe1u2cUW/UrIqgLodZZ9QgOqbattfuM82yUWThQoBqn3uBHoY0AvC0h+UWMckfWI
FGDCn9T8kHgXNUEkmnKqCuKteKYxLE9/mgeyzQ5buqydyKFkB3aruyECovCPMHW+/D7aDQFA+xzP
KMNX/hiY3c5KLfa9JjjM/UpIqSaFQJ4/Boaajpp6ArAt/jtNxg3EYiS6p0mND2Z3Sl+ArAeyY0wM
jZvYAMYxelPjmRb6eNWOvKhuNSFToCpFQGpTiWD8Wb8KsUysJEkAA9DzkBNv9RchVBKR70sMB/El
kkBZcZCy+AwhTsaMWOI4PQrjZ+S6CT0q43lO1MYgnS2XDOu7SMg/I1gGcNYteVTSYL/Ssc5tAAhG
a/TkF01YQPd//K6MmdQD7igSTMz5E1rn5dhzOpFmTH6cAScbNtvor6pZKc0CkUCu46Gfen3Zj8nx
N8Ae8YUSAezgaCU2jwyknsHjSEv4h4hIl6+rRIVmX0fA4BmPMD+1lt5ksPd4lNZPZLOFIQO5H+w/
lNlQtjVuuObTVTKrjTPmi31i6RZoizRExdfmS2R090giqF9WQWbLvY9tcs0o4Xb67fYPyx//7P7f
iZHu3N6e+SG+nXgdsxqj18dkDUrmQZo3IjXkDpNMd9u42L7IIeUgiNCaI6FWz+XYWr7Ybsc7ADOV
wuyD5EngDSHqtl0WusAR6bykXFr0d/48so0o70zzH8SVfICp2pDU6CduVroniTpBhtRPz0nKXlDC
koupt/rx5DBpD+Y7nbRABewpCdXDgHUbHS1EiZOV3YqUan7JFrI3IKXl9EH859y/SfMuLXzrvj+E
DAA8mq7iSBwUYryYuObuY320LQMA7m2bnoypSDtjklgm5tGK11tzoGe39BP5gvjLZm3fl7lp9r2E
CeHWByuZt+TjB4/kBB4Mk+3xjeCXRxzUeDVdVzvdIi/F6D9Tc/sv0z1fK3rVVBY7tfUufnyYlmTV
lV13UkuJGKwhYN5Yr6Y/kwBrm2ZWNPlojLnYN5q9IBHowyNCbLae757gc29Sg65d1ueM/wp1DbKf
GbKZTZ8rZGo1J9BWVF+QkHgmIhP4QC/Dqp7wqh6nzJXxopK+mz4laPHN35AoevVet3JMCd1X5Lnc
RCGHAgG9R+B/OaJ3TXJW0R31ntbub+DbN+RRbljx9iZZFHnt3vGkuNEksEfzMvxM83hmxKTKC2YQ
hT28lc/YSTKvxtz5m0bzDxqXmUldxSlDrrWNUZo16AeA6lyENykxxVpTahhB9ISFIon+4afDb+j+
QSos1GRl5dFzQa43yiupb8sCvDgSNiug8NCmv+RZI9huZQN0ec1bbl8ZYb86HS8azfCnw+2b4faY
T4QexsbisoTzZrvC5p7skf1jk14cfj84arjdzR8aoO4UaxORfRci9hgb72IeXLsq1pk+7vxvA/1e
Rs3jrXsDIk66O78OdOySVrQ8zgVBo8BKtYq1HU+X56EAZYZMg4iOmULfdEGmGiV7jKs020gbgM16
QHazaLg0cz7kUdbD0Z8k2cEZsF3tg8MiiseUfBXLmOJHLRYOmV4NZZNPZVxKi5T1T9VfS3GiS5zc
S+l5krVjhEvSTl5GdwON2NEIYmEMhomvKzd8uMYWqII/DUcxvd6SMgG0s0P793YVZwhSKz7I8ZsB
5ytb3aWfPrFcC7IYimWnVPyAzhltGTyP/laMmxhLWac36TnTcVH5/QLHmPASwcAUnLryf31TYTX2
kbucoB8DbMBcUcOegUv0cRAAFA0e+9GRCgF7+NwmIiY2WVs0WO6vgnSozGFx7XC+jAHJsj9QAq9R
8TIwcTQlleS10mZ0lg0FtGy0E2TYPdkI+vO5BUSbigWQmE9pid1olZOXpzfJRW1Pu3B8m9+gfiW9
JWikXjdOlnVq+nmZnNXjAlfdV+8sn6VFN88KCE6TIEHVmqpB1tIzVEFDufagh0cd/QpEg87czcOS
Eu4+h9X8dIakWOq9kZZGAJYBZBQEWxUYfXIJTNMnpXHnoNn5yQ7MV79t3ASRobx2mtDYx1OqR/J5
3N7mtpUf3EVBwdazxrvWzPNnZ8FpiKgvFGW2G/VDRQq/o5P3mg84/+Lmd6TwCvqw2riZhfhgYytn
tLHDzVL/VEf6ykEaw5bbX1aclh6X6pTsmZJ5/kX26qf1AC/pL7r59mXg6CpcX0WnOrpWQySvBULO
iUGofGMbFAK5/k6u94P/rsxTXazu0TbslD1s3osMA92ZWiqWDDy5itsAkPwcEQXL93KwpK5+81Nm
HN4tztbr1RJJ4uDF5J9BxiVvQJQiSkqqb/8y2lf+2498BzzdnYZeGeI21DkCErbmcfVi8p+yBcYo
0wtPEfOCaIRmkSgY12KzDLgwamqB+vfZOxCCJ7WDlukRkRiPAVOj/1cpY+5FsuEsYTBuUJOdgixT
zopdQER06zMwkCawnjQVLkWeU4AmTGm+Erwp9nM6E1ViU5pr7Lq3G/rLpzvwIKYQg+/MZfk9Cb8O
nFxj/bKoghh0VYt5zg1EbyXTHdqLX6f+ZiZLz7pgUsoMjBmINDWf4Jp5JgzYFrJyFZ5STQYrI19W
3jvpJspS3d3+r0TCNRD1LTKD/K42gBk3RiYUkdJiYN/6/Uq7iVTEGmitcrW3NaBbDN9xdyRq2Ksp
WHwV/fiDcIoMNb8E2pi/r+eABF9wWHevXvaZ73V1yiQ1SGuflVz2EfxtF7pGinL+nZ6At3n9nyXu
I0S9C7rAoRW7tWWBZIz4p0nEq6Buo8/rc5QwqOodvtVqD5gN4Rh4vsNuAuuGTXjbP3MIbU0YQR8c
cf9jyHQ4AhokymAkDzUNMBc9Zk9p0oUc/e1RKm7WTXsPl3AQWpY0/mEdPMpibaLEz5XyZlVydhWc
y9v6FFLwXA2IiAErwBKS8U6xYmpuAwVG8f1NLgAJBq/GAxtXG5gY7SqQBr1BZfITHpx4HwudN65m
q4VM/gH9Bs5VwBN8feYioEbtZFZpQfrh7u8/Hh8g/AwINr/wuYta59r5/Jj9st9FZeZmx6+1rRn/
7VQXAddFapXi2ECMVl50vSPuFOkRpOHmfXIM9xsBD+aLNVHbwRj1xB7z48WZlcR6ncmq7gtiZz6x
cY4WPvdINpeTHD97LUfAYeLj3b6zI7NBvH08jyFS028BTVq++EkjJ4mdMB8kACEcplHs2+cUI76K
fUkX9W4xj2WmWr8wZ/voFvQUp5oQIWpt4QMKQcd9vFzY0VidAhApmJE4352LhOs85mFWWsf3Jclf
AyfEo1tXOjr5vrBmID9bHVjA9ZFKnT7a8ztq8xO3AnicRS5+/OnFsoQ98wFK+xm5F4RjflbOn3Rs
c2dxTCu2m3OScr+xVbYecxGiSRC/rudpdlOgH5qnkeL0RUzwwEFNdAxtz3EkzApv/qa9RiJvyVW8
MSJsvx/GOK4GJnV0aX3WUd1SrQLKsMtIBX6Bk8dnC5K8H72MmpYPOCztDalR58KPExxxOna4nsbN
9Sezmln4fkcGjSiSQG/1C6NsWgXyJtV3kFx+REIPFlT62ykqHLp8CXuJ8MY/JQKb77bpYzWxqKkU
nqUO/xfseSPlxVmQZ6XJN+Xcs2oA61sHPwRqxevha/1fM7SchTMwPeet7FvnfeaUjXzzcIwhj+lb
YtwRJD6sNwo/SWQnTk3aV5YtmdNba6EXDnQQu0P+VSsuQk3gFGuSJWfAgg29Hw+ftFJixNZ/lWzN
0jOUH7eihzuahXzsVXbzBWlH6LNIe05uYjHoHOC7dUCgTRRG3Xjtah+SZBBOaQzaBjf1+3PoDaa+
PTvnzGrD8mwVFCwAjqmxArx1ayAAbPA5hgjkbfCSRp8te35uJ/Is86A1k4Gs8uBHUjfEcVC0wIra
TzHs4IayfbNsgnipuP0DGyEnZn8gOHec/Jk2SkKceC9YRKTG0yRuqu7rT4M9a/F4s/vBl/KN23yM
je9K8nZt0n9OvghLZgcGaLwWruvgY5/rJzcQD90IjQIr66JMoRDTgb1BB3vGMsLBEVy+4aumuVLn
HgfXH9AfKQSPirRxFUWqlkC9ASw1nSizynf+W5Un0AGCI1JIRY58FgcJdJHFHLz4Y+9hjsIBvlgx
o4NR752dP4vWougJHPoQh7o9aj8GuwqF99y9o0siZt+HwImNH1C3Cki9DPolCZn+K4hEHYbm5TcI
yuQlKLwW/QUybstYt+c6qpOHSozvIHsAO4GcAfEXBqfhBNQeewG8404jOn1OslF8yYrZ7gW56FrN
KUqDu6rfUenAaSvapaetwBLDcmHXBGRC3hTSkZl79EyQAOtttqTeIpTQlhe7qF9wNazyCutP8N6D
n3SjbxKi7f1wVOfs7OH4/CbVGylL0WIe4RfNkxF2EzmXyUtCyLW7gQ5WhcMpZL7mHZafzh1Vm7qd
PzClv3iSbSEROQG3bwapsYfKqRHYBooGfdzqjhKAALovjsFZ0Pz92cyFVm8kabeGhqpjN9vHosTs
Rb5bz0k8xS+kT7e42AndAe812nPR7ogMvFC3JhE+LFs1n8ORV7FFBqJOYXJFAN3pNJcozvSDYsti
x3cuVyNEJw2myPUBpL+H7ucBgZLlsMdIMGRBRPQR5apZjxldlId6R7/7/cq3uFbabDBcrvNbpg0/
/cLmrwUvVY3BmK0ozknu2FlP+IwTz9j2U0Sv8bZYbR2E9TUt4OH9SJFPIDx2LpnWN/l4wFiOYtpZ
M2zWAg92siXQ0+rK4ZXBRS6p19vnMcnTrwsy6cDu0baakQhSNyMpUG4GomAXEMETuE7NtR6VaP9Y
O7tHP6ZVn+txnRs98GnP5KthMOGMF8/8iM2Sz8sMTWv3qWRGR1iVQiHCHOvn0SfMVe907gGkfcwM
c2PUSR4pDXqCQBbw9XdLwxHJKrmfikT2uAovg18WTj6y+r/DKTThp68EZTE82MY0bZ37aVi7Fjr1
iUgpJInIpKmhcqK4Zr6VPKQ0kbGlIn3I3JbZLwf+Te514QpJ8uoHe5gLt0kTg9mR9wqxkf/f5pJb
RxyUdEz5TnJK9Ef625S21vLXrvWokCKST6/6WuoCUlbCoW+bRmfNhaWL67/aq1GtfAj6xSj7T6aL
Ms3PR4Ynk297k64/jn+hwACYLTAlNr6Dr3lTSxLs1DwvjTwx5tjOdg6HE+O4Jp44wpwmymeJlR0u
rILt8XU89pfz0XASf0YTvBQf2HHM8nc8gVMW5XAtpZ1lYy2VJ6Mfcqnf+Rnh5UiS6dwh5LiwApJ1
Hznw9IgiF9QRJ51JuNLfd4e8tZHFN7CzN8H38Y988QLPDsz54ZIDWVG8T1/O8j/DVfOURq5WzUud
BoEnwLA+EP8PFTGN560pkxyllQdRYZNiXKBPkfMS9vfXehaV3EP1dd2twbNOBpH60Cg4y4M1Z5/9
nd2ow1TN/AdV+XYfp76/dWUBqIP0gGxJpwVClMnlsbgixJkOmwr+QXV/x8eX5R2BILw0iElviKgv
Z8DJgy3ytJvfAaZ8X4FJbYqmBBMAt5L49idAFNd19xdKTmF/BhtBsEM5asgBw/8CF92gcjZsWbgV
IIUaeM6afllh/uDU8hjkPlA/9bprqtHlcx9ois3AvqZi48w3qFdiUpyDX6xmV/Lub0fUozjNjtRN
SP2n2LNQ1ZGNAcRYY7aGc3PV6gYhiAVe9CsoI0hPLJNCu2N1YcWDZ/4AWNsDmnoYrd2yBOOwCkTe
h6F59f9ZJS+WFj4n2MOhjCASPr3qX6jxgzefx51QGhY459naNH70vQ3J5JT9VQWATmLF4xFcZkN8
krUu0SvZL8Ac57EGFWL8rgd+JoK+uObSBZE/FbYozSChcBR0G4VO+jlv8LzkhDpMNviNM+Zq5rs3
4n3XfV/V929IBcTbv4iD+TeuWRNyyXnC4kn9iT5ESmXpbnTfDW2OJDM3iTCGwogQanQNWqq1v0bQ
K59ErX9kq7I5znfNnYoKJjKi0LgxV3KCLKdBNB4TDdikMM8+jHCCAZOX2uln/sWC8md8Aakz+3Q8
AMDCw7EfEx2oD72TSGUBtQvHKceIIEyg7C6M38YxbWu9DaHhVCGMdF9H4j8FN9HMM0EXPyRVmR68
cFtwxuJ7aqVu6FwOobba8IfKabEqr+w0g6t+rnOQVKiM1STT7Xh08ibfjuanYeMUzC5xphgy3l6+
BRX1ZxxzeMNU+DY2xVFacF7GJPuxRqovZPPhnzRSFHiVyv9GyVQfnaD9mNENEVy8+roNrHGPHSPz
yI0K/namUPorIqwe72+c+tzdG6DZqipcrmt4wpHqmqBGyt+oMOtsFUj4+OLw4gPwD5Fkqqiv8KyB
Orw9ohtDIN6LD6Ohpy8qmS/GckWNw11Fm3jV93Xj0XGZmpJ5cKO3TpmjNVMltimFDxr9Wly3j60S
ONDyeDeZpXYGYQsULkgcvioF8Iyou8FSDODaHhpCfX/l2R72JGK/Aab00NKod+OpKn2PtLxVXXha
HY0/sXSnqFlUoVZblwfI6YTMGSqoWN4nNeSlU9kqhvF6koIG9MnJPPK/qLkrNpoBrHCLZgIRGLWc
c90ngAyc6Xa5nWLptZTECafjDYqKRwlYP1auilJDaixC0/dXrXTRp3lCn7fbKAJNyZaFWOWl30iL
6gAfQud+0oQTEFsCHq2QAJKBNA0jQz1nIZAAgwm9ErKFB9tlS8kGUq9DQtR9pSYPwn3npKHU3hP1
lMOx78q3Zz6VzD2XkwXPxFpPEirtPHLzy6Y9ja7yfiDz95tEYlsA4TYxSNPZBywWpMpb0ZwXgkmm
b1Jj06OV+lEC52+/SoSuKq/pMTVSUJbCU9biaW4cjxBFhcEARkob09h5oyvNbXKAz8nhOoI76ULN
FnnqdP5UQxkYi8c52iq+h3H+3swd51F+nSVRlQlMG4XybvSYBr6UYDJrQJhL3ZXT60dp7QbPyI+F
ABM1l+Nt/B1xv1n4n5At0fVocV4JKszFdb8K1a6B9/MB4yxUb3e+MDF0C7QKb5shclYqG0AQL+fQ
LSZ35G+pEiSPMci/NfFSlJwyNeSgVDlIYyDhKEeAzzGXMxtIPRaXqZBbPyunZWyit3GXDd2n/MKV
OZtfmgtlNc6B+SAiosucPwqQG4F1u0JfeCy4xCzV0fUnnQgKDdGpUBd9p4JC9Tr5trQeIiC9hwjZ
z37PTT9foVrKwDbLErFHgnQOwfiNnVLyUx3oZrgjYQkE4asShjamVP0aqY0vqE/oDicjj3pgC6iS
zXBvY5x5szmTyqUSXSzbQk1F9yUz20JtA10D1kDeGhcAbz6RODEOm9yT4gMDgApat3+ocj8XsJ29
kcWwQAWZOMM78Vlw6UsPXMtUaTvQLNOA9hEava6vOpdDp8quQ83h9xME6Eu9/8GKRIYAczw+Sipp
BYkJaVE6EmYAdd647A8EWI0PyXB8foEF9M/mlrKj9tjmA/p8ksblSbu8i6fYlOS2rSTEnDNYEfZa
mN7/LptaJPuFbNPBnUM4ZtbQTCA84JqlD0WtpXxCf9dYq+BZYN5LK0lPuKQX2lQu+b7dFuKTz1mP
VNSGdQI7v22qfcpjcarYX/HH2Ro5t7bPjKy1neb9k1V7EI9imIVlihw/40Dx3Z9Txvinq7WQVv2A
lrXP4x7mk750hkqbza25PKi0zHfhQ6kVVMikqI/ovXGqBu8SNxY38avOJGldsggMzhm48yRVTagF
zrKRMVXNxy1mErqXwXSwhW+5cD9KVtokVjAv/AztJ+zHQq4PApADvEzhZp+O+rr3hQU9eYqOg/9w
ZayF9djkPYZL4aV9nd7fMtPVOkXxj8/jES+wAe2tX4PLG9fw4eykvEXDAbEqG69mIkN8OMghsxjF
WKEQfkikN+uVXQ8iwbcZU3gZgK64AdHurVsFovK01cnPQy2QkKww38MPtFXyXtCYa8YESofxraGY
SnM4ZDctMk51xYZtaL+mpaK9VLM6PHngj5s8j3PUMTuX2zvlcl8/JyhVf9UfxRcWhuS2KF5BG14L
3Op+3xGFCDDeWFeiOVBiWnu+a4VlPXopW3mveCWHQANTUgAj5ycrODortjX6JRmmPw6PoHnj4nkU
vExlxh7MLmmE8YXuRDSngyZmGdgS1IDfOu32RbS591MsECGuCv/hdDQOLq4uYab0NLNIDNYmnrnA
0Wpvf3QYAh2f+wUcBEObZIKcfojI4ZWF/+HZAPOiYA5bHf09VgBMMt6N9RW32T1lg7kn4V1NZltB
enOTolVETztESw20/0fB7OowH/fKJbgMb8BWVdYh9+1rytyJ8YRd8ni9vJUodLwQ0M7CiwW6lz12
DLbhkdkwK82ks3ibalo9pBnUo6nR4qxRAELt6SG2OjtrfF8fM0epD9R2EcjQ+K8gufv5KANiUIET
fMYttEz1LH++PExORV8CvOkyALFut5+tKRRz2dF6Rottdc+SOOULHOYVJjk0HSsEkS9YTWgRE3tP
lopdC5ZgDM8RwDTd7v9H2eQ6slQrwX/oyu6GZu3LQDfuI/TwG5p+nNPnKSJbbIG8sfvMsmjKAUIy
A3eGpWg4C+berLN1h7LryBmvb8Bsf1pnpxNurqBPpZyTxB40Gqs2x2DCbr/YRPBDeJnr3SKgSWeZ
4UNpP2NDc8v8vA51xfISN9/9/T9zf5xEh1Sa1dFGfO1cIhw5NAc3buTK93kfQj8jvZJjK2X59Vl+
xxoMLSCKCnhdi4oPAKDLWD0yb4MYDa9lWc+qbpkLA3gu0l/MX2/eCkQNJxToNo40EI28yfzMB2Xw
s8jEs7mx/OskC0BO1SDF8Ti9ZGtzjjJz+lm4t6iLrajs7ZP+skFhz19pc/SdCqtHfw7J5CWZpeXS
TECkKAehrMYXR7x2nSUTfONMFEo2pFJCUmAHjaVU/uMw+zT5LXyxtnHfGOhZ7KLQwezkjFJxn9dd
wmTzq5bPece1xf4DqFu1BdfCDSpL2jTcXoq8UwFOZ6bSUXSX1P6mIGagyGwfOFcpr+JOv6lqkE4R
R/mVzx9JSLGm7WS3zMEtPsrnzJtw9IrlmQNMIGtER3wPul7de6VrOgbh7Zy16dqC81x+JDwLPiC0
psX8i2XiiuykHbAK1wQkv0tbP9srOLusmsfdHYOWqGwv8nVwTcHclMUpL6XNxHhEZ9oKkMTNujho
SWO6A3LtP4jQ87f+BYiU98l2xWEKq2kqseAzAYqwyI65gnpYZk0kHi64vY2FJQ+6aX4ENE6vUIPC
2/tDaEijOURQ6Wv8H67OJgAbT+pp9YFk/l1LgaA/8oddXQfgV6AGfEwyLkhfvPosXLKybpWHGLeU
gTZPp3/7bF9shIwjqF5Ae327vJo9Yogg0cHJRHXLmDPGsalZvtvfMehrKpcWYhpRyYkb/le4uRNN
NtU5wJHtv8usPhgTnfFrLAVG53qkuhOHCbMd5JFBso8C4yJsEtL5DrRxqp969TnsbmuuN5QMXwsq
+2c7qKnT8plJSc5WCwO9cuU31smTPRj3BQOYZ04iI0HUCiSR5S/Cn2IFu+PTxfxspPS1anEfdJCP
g0VsIoWnyYnKFULVlybycSQXpr6DFvvmp/KkDAEbrG952f68QZsht4TyCZ4GztRLtWRQUAS03/rP
rCXfxQSRF14Q7v6+NFpjCv1tJweryz5xRZC9h0tWXdBKKTssTToVMH/tdL0AzGFcsqq2l/O3PPMy
ONASXfUv4KuDSjgQiEc1lRqE5SVJ5rW0b6J5EKwuj92dG89Opwp/ovKQOvz8czCa3HBzO/9aL24x
ER5zyK8XuCUh2Zt5HqjV/LogJX4kbOzQi1EaIlNizcr54BktIVQ+Di75k/bfJSQ9DvmvIJ5CxFtZ
m1ii1IuIZo6yUK6D74R/Peco288Ef4ZFiSIL1HMAl7ZPCiiOZpkWP5ll4UBdUELDtr1zW0/wsUO+
RAPNlVoACOs2G/x7vFwcUGs57a3vAm9D9jHveIKZoBIiPuRg0yrIKzXUZlnvopamoBA8ffwOEqEs
JL4aSPfqLOmdVcOkj8wjCTwInYppyuJ6X48Hvja+q2fR+MlTxboG7V6KsVIVzNAszFxcDpHpaxU2
LNSW9bfYMbTZ1m3st6uHeHcVtz1fOXBOTK0zdUdvsoh2Z+OI3GeVVr0/lWUVM0Pp+8HBzV7oMd94
91QshK0Z+awLdfmA7YkXlKsWymnemUfJU8iUSE6svgr7AoKNtoRxPrMO+wvlxr2SSkNBVyaDZrX+
jwKxkwh849bVl31iLNpdSq+8nrpYHFD4lKBiD2CeQ7E2rosz5lRR/9M1py9nqqPk+ZB1ek+2McDW
tFhU9PrDfr3OnCdXEGarFLR97tTf6hnmpligD+H1dlvTGT02kmhagt67qmEtMRnlsbWTfLqNqDce
0TVZI+KVCKqsvN9w2RMXZ8Awon2vjJVVkOuDWYDZNO4FQLg/y2G8u06JhdqNRBAe+Xp6UxaHVxTB
1QddsjS1mCaeuc6OEYQDKAGKh+T9d7i88sYgUftpLZVpliFNxVnZ5j0t6UNYCVV5GrJ++YlRsIri
XGIek0yJUT62TYZ06/1Bb9ZbQTc3O3Y8CfCuIfyLdA0sbsGb9DpbiHQlcLVWOAjEW2n35VgfqzqK
xRei+eUGBktVz0Pm+aKf8uqZPbNBTEvBrJ7YFdff28Nx0wUTmi1GXZZV845V94rdqFFEp9g0/gqi
clUYtKKSuhMw53gv6n3H9mHezQlV8zrofNPxlfJVFXTE8TJiPTdyrYbzztr/hnPQwb9WGGrXv0C+
fcJQOaHgtRHnLwtmrqUketiQSZ/RM07YrSa/Q4UAjkE97jOtyfQmvTerUWMTDnAwtVWvNp/uFXui
3Qqkf2Vyzg2zL6teQRqs69EHVYyH9eU67pzyZKRgQLZH9GW+C54VZBNB1/38J3drFlFytFBGf3PK
O5qUa2j9s2K5O/2rxX+zQ0TKQ9R2oTzmZwhpOleDAb3MYi8NsqKqndxXbvDLmXbq1ZkmU57+vXcr
bm2foENmvV383QVN8wF841q2TzPu6ZHFRcO5LPoiESnWrknzJvos/AUdsHKuqhj91Jz94iClqaBf
0CdQvAxW5uw9TmqWTWu0HBG3ueVqFNHg9xd6CxODNhkJuMRn1s8SDQzDoWx/k9NwEMH7z3nDSmms
cowFQEbjoJDg0pSOYCLRNYsTugjc1Cm8Z/nGdIjYA9pkEfqraW8EZfABaLvO5adzvvES10Nn9Ux5
8cVohsoY5vGvaNjlcvP3nequ6ieU7uLZHBEBIAymK1FhBAFH6MWPPon7IyTHzSBn7zuakwqDmZ9+
YV8+rK3hJYCgyg2rDKiU35k1O3xJ7SxCB83/wvj2UyFy984BWZh16fcb6lEWMWhqUfK3s7apBCuD
32bcGCVCNOJsXWXbToGE9lyq8UbkxpFcDOl2WiCH2VwDrkY2ofNq2D6YRDGYfSTh3fZF+FCZE9HR
WWvBiwkKTygVgjvys2QMvVakCUfQYrx2I7Jq5802a59LUomhKKemnLw4x3A1nttUuu+fkXzw8ZrN
AeKG6DXtdYT4ZSuqzbhURCD1WnGdocP78lfURj6FlEQhW02/j5kcADdgvLo8DM988XjLMq6TZatt
Om2yc24jk6KWaf2Ez++M8WFrbycZLVnZIbBiHbHnQmOkbiS0r91Itk6rvKH64X5X+zmcqEjrB9eM
/6drvKz/9GlZZ4N0GEjtRefCHhLr1vkKpv9O2JD+4XFy1c3hDbMjJNOhoPMo0LL128EBZALjaUGz
4AW5Unr0HvKEqmO9d6q3Hv64BpiUS3c72NUbOTDsq5aZ+yp+hdgCjdXfVAM4krA4IdXyQj6NzRWn
3HcNRH9wugLsdgSBNM+SO7rBtZtcmKV3z5LnOzbSAM5oAuNrcoLv7SRA0mbII0gTvY+i5Kxm+bOU
U0374XvwIRlSGYfcbymt2SwUpl0a1wSjBylCa+MfSEhLPlqbc5q88gVNFZcSwoqWO3kwcW7tFq6n
q1Hdav2sKXp27Ib/a91dI1nRxwWUQKCqZ4mZ1zet2+ljX2lqg6YZJeWcN+/ybAA+5KbHRBFjI5Ha
xd4Hr2Cjn7Ex/VpF1trRBt7/sxKvq0zA6fO+44ow6ScXvZVPZnwJBPGWdh7b/rljR39aBqyKS/np
mWCggAVqDD5wbvg1VlsU3Eq7VLPtJt2WUKvZ72MoTdycOG9a4YqdPC5Xj+lk/D9PggFgY1n9bfx9
3xRhiFOZCBs8K8Q3dw1Yl/5ILwiTJCoJOn20P2Zl0WhZFkOSFQcEWTwA2nTLSKYaW1h/28apvPpQ
UVqT7td+nN+YeGzibgGZfm1sUtS2L93srd6LlJe+i3r4w5sr/6H7E++q30y0N54mmPyOAIWKrZux
H7hecE/mPV2qQIDLlqajy5QNthbdaY/VZ4PH1MKulqCq04ih6PY3Z7t4eNzZ6GFmeyNFd1H0iRp9
OuesziXYwMqinw4kmr340xVIb7biMqN6NVJrZCyhjkE+h2KeJH33mKtmtjDsWK0Q8iTDHtPlRUyC
xJ6xbwr0otIMvTFMKQ8zuuqRN+N3DbeRay3HbkE1q7cQ1nbC5/3R/sBI4A4Kp2zTmlNGzPmfN3E3
peWABoqzCFcecS+rVi20ZM8l3GGFFTcXN5o+Rbt3q3ifYX6LYpu6iF7V71pLzbRo7HXfs8rrCfBJ
ujXQlqRaz2ofB34mtAQrsIF0dNxo+04JDwAXfHvnBigKK0KpK2YIk9OEt5JMB2vXXAL1cwo+kg+z
Cs/nEM38u8tIyBgWncM1Rxy39EqV4NHPIS1OzJm4dOsGDKyapvVjk4HEX0RI2rNQfxcwqJDbNU9r
UNrvWiyTDBiGqui7Q42UBJ73YG3Cgx7bxB11FjBnN+xKOf1DoDkibsnLT3IzlVhq5MJeiLdlQGdA
UmKPjzSh9S/Mht0PAc8eud8OhValJd8nNzBjZ1LESma+GDawRmYLa1jUhADN1Ob6DyG82Dr8VsPQ
eT2PGDOSgU6lAyxJRdr8/IDsXLRF4qFvFg//kMzWr1sw2Co+lWVZ5bE6kUA5Tj8tG4peIuT0S8nl
kfx8OxhC3qpwVALRs4P9Dz6F2mjPVSLKbR89sIJvY+refbzCUC/T7qVaUB3vwf2R5dMEP4AImzTp
iez4wdn38Cz1Dw3kpZkp6PAyDI/ptmrmTf5BaPPzARWRJYqD8fJ98BsaMbjIOkQfrLdHqDxa3JyY
2z47kX5A/1EEfNpc7m1qOzsrf8muyFbeCyQEn9xwZK9mZvofdI0ilIZWlQOT7NR7JY0SMvfN975f
jBTxzznwP9MADfdUaRYbGtlkSppTF3nKI45wIn/41JNLE8Qp4glV1I3AD0kADgb4KriMV1yZtjM4
zrQ+p3YtydPW+FQ2EbJ/wUWOo8n+aP+yY7FeQgUtSkKUoOwTNqQggg/yOOUCubxOBCtAY4jlm43c
SfpNmZtueYfUeAPSxXwW8z+8rve1OgVVV5N3wAR4eUjiSEvPSWJD9uezTl0c8WPD/6dZrvQEiJvv
WFdgVUPOwUqIKIcKiz33PSFgoaooJ9oB1xJKHpTtKM8moyNgDodboiki7jLS1aI1AJa2WI7aw0pp
u+Xqs1kYiPCNu+vyzV/hTCCN+nQyQ3oATDzLXIsU6FqQ3PM79lloiB9wn/JtUgkSAGciBJw7QnkS
2/ZTlDWC97c9s6UdI/dKpjYdjo9ckkxZXEXNF/ftDwCFf4fXBDpfg+gpsT1pZstfwwjLnUJBDZi1
6LvSLQbhOUaUd++OVnSHepg6IfcvxG91/Bzsln1Dl8xO8wonviyLTvWbMVJ59TEWgk3euFIV5+pq
rt83zfkimLWrRSfrq+P/oAY783HtKriRqdEh89vB5WNmw/27475t7KUaP0ukGmT8QWJp1p7Gem6/
zqvTlFiHZ30U2jCs7WZtKJrfgs+9DkpFMmYD23vaWFQ1I9w/HwE4e0zsC4vFfJHF7YtbAl7ZUsox
vKuXoXP5Cyrp4TbkAOroJFVMUoQ78VBFydPq0DTNZlmO+f89zYNJTycWlfg/4qPox5J5KhK99wEo
cTqhj2+Z4QJKliz6fPjxBx8DEsryLaRdNB24llN8wjUrlaHGZihJrX/FNIYpY/0QqJ1Br4HneV1w
D3C1K2iYf/jNa5HS0KYM/NSiIymxF5FGFm9TM6sp5ECQIUzzdgyeQwiuTTys/09vjJt9rkeSTRcM
MavjQxaPG+joSBG2zuT2E+k5OZBo3Bl3IZicDwx7RZ0wdx7rsboImpcZQBAqLOdaBhppyK4DxI5y
idkxf8cG/VbBZjUdCxJQsTtPzUMw82jYLRtMUrAxARQ31boV3db9rhfbYStTZvg8KotB6IgVtLVu
kdoovMZhDmLV8nA2vxz2c6TkGpUiejJ84XFwk7f9YRuZKBDUzTDQ+a8NxaA3lC1ANifnkPtpwfbE
9FPnzK/1HvLKZeotGhd+SMzuyScBVS7jmpFzup7WkMY00HNSI5YSj5QB2ny7CyF37zw7ZyFsEbKc
x4F/xHuUxk/imQyJEszz/5/4Ab/vHJIGBnc7cO/lKqPNyEvvsIe6ihGj8sKP9m5tUp/QyrYendGI
pgNVa8YByuP/Du5iOq8nDEtDT+YMBhnbW38erdyHyA60G7ZXPmlZnO7p/RAU9H87X7FRq0VvW4qh
S8D/7fU7485/5RFxsOWyZmK9ZhfSnS7r/geOonoVEDDOqjp8bcJM25E/Jngx7Mk1qhuikveQ9/pP
K8ZeWBgmA1fzJV9bPGKHjbvA0o0SOlg3VXPNtZvWYhAHzvFz3kPFSeEEAXJfX999193TX82i6+Vs
rwzlFL4OTA6ciMkudK4cdv1eyW+M/B1EJQx5YxTCRHQOvRmwzU0DHI2QFGoY17q3byZUUecEuOb4
vukpE5enYZ3IblHxZ1FbCLaqyJQDriVBLcuQRbTjAPt9KEr4lc9t1xO9xit9/c3c/yc0SKT7OlSS
ewfWCoePbGaBEYh+o81KzjRkJSBc4lX9zwDnRNazXB1zghz89fVrkPN+MT7KjnPJeuCd1OoExKcP
LO4pX1clde6tEnNk8vukzAV9O2TG43xEwUtkKI2KiSrahRiN5kiUFTo/ncZiQf+wQxi331TfVHmx
HO+Lgs4mdgPao3xjBw9RxznjCpAHuzWvpn64MBym6sVQHHj6OqDB+yo6dl1SkbrY5eYz0Mgpd1hW
3VYVwFw6t+QThkiGrEOM7DZEs+ZaeiZs0azuMuFU6alycl19AH5UUnLCHBi0H+vMUJWPtG3P3ciX
iwn9Obg09Olf2SAESwKYqpZgETXrwDGpzrtOMxoHTYeSwtTC/hxgSwsFCO8fcxG27jfPYtDEUdXp
ECTFuQVgHCJelVaUOM9/9f+laBBnc1yrVPk83lLwhOABrhgS00weeyrc2kjZIkWf94iDlYbxhi6D
4IrZI4IRBECmi9u6yiCT9jMnuZg4uJVO2acFB/opcY93A8neFY8Jm62GCvZzB1qxtkN2/OReAcPi
dkp49yGavCV1EIqaqbzCICwfJZvqHWvPApiWXwt3TTc72Szy96zbcB64wcuwv2q3g2tuSvekSS+A
xWV9wrPzVzKE/6SblyEibEVdOyhRvrOx22QNIuzsSl5+WpUrzGy1MjsYc+iXEvQ8HWBlvxqsrcff
apOXmDg64dO1pz+KbSnPRNfnbqKFM3Gc8bLyYjgJzQtPH8Ccxxe0ffDEfgi1DGqnPucxlrfc87ni
+tZsE6t+Fble8CkeGJvrH+xrTeENjzrEMyXN68Y0dnRazGg80FZi/vu160MRIty4wBtxY5euZa/G
LYj6hSsfcHS1E6hn445jl8/eCZSo11AtcIvKua2O16xuuwFNdTYflBcR8bzixGCwCPwEXOw6Moiz
uleRsuoCxKtFeApp6Cw+M27vD1ELcflxYmjWVb7/oYKDuWvJMXBjn+sGvRLkUSoxWrrHkqOSyueo
3tWgVYTcgpzxpP0kWKbPztCTdETX9X/NA3fw1OkbLIBCRwWZYaDbkVS4deIOXP6FSDd2r/2cDeTl
ML4uCVJ86Qgy9Lg+fZSVdByFjZBW27jdT4/0KIeJealNrKX7fbJpDhZkDDCQFwpRqqwjTiEmtW10
M+qNHVKjrcOgzt/Xe9Fm5+8cB/VmqUuLVqYhRoewAZt3PdojAN/hVA6oM55/iAjRC5kKl0/xqkG8
g7qfZqhCO8f5mqee+Aoy87+6cC2znApTW2DTSXJzHl18YXcp1KfPCof5i9aO56+9R6fI0rZGYaGY
6WlGYIxoy+crIKS8S8XlO1a9yBXn/NNVNaNMCnHzm2z1/3VJgoTpwTLpN7NfT21w5m9W+/zYjz3I
7lYfzTclWkthH5XZUI4nUxy/eVW2++DLIbQwpRCQKLOnDyHNtSYf5sXAWZE20DCyUHTGR4D1cVbp
F3Nxu3ox4bptwa1db2NHu5tU2VIpWQUc/tzQWhM91HLF0wUWJ9VwtuAJJ6LAupEPiMKN9iCoxHKn
erFq7sg17OO4oZjdO06h11XaHWSMxEqfOjXjqQsLWZGuNilwenOGbBZUs0qFTwWy75+irTxGuXC4
1i49teAbzxU53RHku0V6m1Gw6YDT5YGHT/GxqszMoxV3+yFkTStmYx5Jtnyth22vCF4zzNlmzftl
3Sruq9SOuUoxzSj8jC8UDXy0XPLJDqkjpHdqGIzwh0oo3i9IIggISA0bJZPztARK0qP5C1pvAEv3
lJkWRTv2t9RZ/zU2PeIBOKtlEhtRq51HqytF2N5FiAAJjiQYnHnQnkGgYB/nZ89QPO/NV8E8KM8d
qqesVY0nouaDT/xnCmVQtp+YRocqd3RfRFgDcIOwdDyvwLIleG7a+JkoUlOIQBlbXx4KgcrHpz6U
K+/YTWI9WNMYKdJtkffmHGsUgSZOHcM0AnmiUu8GYGH0ERjXdAhx5ps8t/Sl9pcV8q02qR7zT52r
jjuQYDEv0/LXsL4jlFKRLUnLHNimOSYLV5IoMD7kdDIUuFlqZvimMJANkdmPQRUmOH/Bh/MAxtu3
lmyjy51/uXi/FYLFNUiEDFAJ9nvMor+4Ve688RLTEd7lTzTuuEgkIQXz7RGl81OJw0uTwIssml2e
7Y/w/f7A4P6AKmyaHsR9cIbGCuNqETELgWe16v/NmYLiMYq3rgl+Ak3HESA8Zhmzokq8Th7nPp/S
Qrz/idrca7B7Z/VK+4yaANpZXH3l2Wr7ugwPWyPlWUn89TowFyZ5LEv9YLHYAFLuudV0cVVlSkPG
A13SW/IZXpExSin16SJfsGSTVQGYJc6r1j8PB7hyYwm7FWkl6D9ShSxaINjE7PaBohRfWSNAlY4w
5jXV4oDdlXo/e3E2xInbbJN9wEoGPk3YOODPPBzqbA7GOF5gZlGSZj4fQOVdUvA7K5gjgpxyVTZ9
d9sWRtNHWaOSGLJ74PeFz1f1QGhS8bjOAG+lK6LCIJ+S9uXc/fnkKb5lwSS4DMfhX6x5lJ1XRBIq
R4Nls/iQQodBZwalJ/owmGoo8STNp3U19brd7Bpt3bW5tUNCMHaTGTjUFBoyJgTbLtDZcuSMQvjx
c7cUZIUL+FrRjRkzgM0laLl6wAkoqs1/8SsRTW7hpX9ruNpN4cJThGtBhFJJ290Y1WAjnbEOE7SI
Pl3PjtGoDcVQzYhhPk9oqYIG1tHvgrf/9CAw98BG5mVm9WSKUIzTsiqQSOpey5Bw5ADKODgJtY7W
nE9tklJ7QmwG1ZVUb2mywQPNBz1cYNTH3co+lMsBaug8AHTkhlk9PI5TpCdWD9ZUJxAB/nY1Pk2X
umFCgEb3EifNU135IYgTnms2LhaG+Osy+VfLBLsX4e3snbfGhqJ2OQFrt5GsgV0vYsD0lOvK6btn
MinslUB9fI+ENjMKvAWAjlSnwXxtG4iXwJ/S7PXhpazLorv+uORZIG0y5tMA+P50UUJjTaV2MIWX
bnoKIH30fafwpOcZc2R4TKeDh/C/J+NsOxK5scI4mfh9WK2Gby1sVM9rQtyAvpTuzSZ9H/9tllMU
5JOwB/7FdVTBj09Wy5NpI2sVOXqYkn5RxnEM2Rd7aMczG0fgiQz6Z5n5ZobjVGD3ehQ/L71FKLoP
xV/OytjV6UX94QzP1TlA8OGV8iHxkCVCrzeXuRr+AjFu4qeBK4HdjKhpvFguH5SEKZSa2mXKMuK+
9ttNf4VJs0m9m5CYyfg7ObkLh2bsbsYLpuwZw0JnFlol0yQV2LjV05iK3eW7I7EJbld3SneSrH2Z
bpHnrYxDZjHg1esVQ6hVOqiahPYlZplZYo8ZnaZtsm46V7gdQTfrcq3d6ha6K0nASKbWcFlk5B4N
+1uLAIH1xkUmP3vaAL2RwkTc0RPQqSHgB9NHPLOQJi4roIItWA2C7G859l5M/kIYCXZATrlXznsy
smx/mGKgYntipwb3kl+1IMzQc6x7dc61YbHd1LiFf37FZU4PQmIpmsfw6bGg74KFmHblKzqYUtvu
9En8pCcweQog2ruxT53ARr27nWzaYCX+VS/seikfPJzjzqwSPtxMgxUa053VsGIsu7VHDtZLJVtK
9m41UxNfDXqEETW1/Lpfz8Y4jom2Ef2qve3/cPad6htptGFDcZZeVjBP+65CyTjygrcDCANzXwja
5WvFigrLZKEUnccioO8W9CD2300aUXJM0OZQ7IunRnhh3RocbyVGagu8pRVsfVckEb0MyH4Yp7sT
g6966xT3xcp60oAiRz2cY1082OKi+wk9FpNItLC/3n5czOc77+gB0Ogufda/P9ebGRJFnotOrGaC
G7URK6fQmCm9sCEIWMitZpFBAIf8jO8iJeCuUi3/zC60UBy8TIWRCdK+h8So9mh2TLBZt/iyk479
TWG7roUhuU6CBgQ36B0O1xQnQoRVAZYwUH8Z9vud787KZ/Rc/YNNHNox7nxMf4hqIsXyOqEX6auM
h3e8zuLig2XmMDDvfuxJcU1euwTK08spUqmuq33YC02wDOcoSBZ67QulOya3t15NVbnL/YxJpyk6
2WC0Jo+7E9zNxrUO/vBe4ytvJKSTh7z49jiasiKV0yG4uHwt02rT+hSGrxvMVFOPyQEk574Kjini
R/TGTSzpzu0Gh3J+1HgePck4LI2I5oFI7N6q7n1D+ILwtk6VDJQxWpYYYb7Fs4E5O40TUNa9+AKY
VmhQ9EoNM5C0uYeRSwsJKdPFaaLWhUyKoTA8LyfYR/5bXT0tyBmlC5NLEIaJtb9jvenSHXROPqKG
4opW+j9VA3tzS47JNjBbWZtrX+QZMURsCze683AnIoLwGRvTUDeu9V2ZusjvMcBdU80/resykidV
j2YT6YAhtxsPrcrqaW41SELR6/3P3QJqKr9wor5YDQtXuW8Tpbq3znoms0agcMEtJdCHv3/9UI4r
Y04jI8vuPfAQgSBh56xAP8xhKM8eKaIUCmdCT9OKBsaFmbq0hPd0UAHcZ4b73hvHc2acJsIZzYEH
Ky8/+qbd/3RyRxFx0HF9S6f+2HXHhabh3LcC0PteWDlSeoH7E+b8CWF1cYbW9/EQsLwn2oYDtiYr
oSQRqNo37w+WsDZ93vvB8T89UM13zTHiD3IsAfcA9ODdqBnS3q46X0tpPpmxFMSvPMCwQuFNtQGW
QUL36zJi9vaJFeJe3vdogOTGz9LOyds4Huc3Pl0FChqI8qRXvdVwGhISMmeV1indRVVp3LHE7Cb4
3VPt1Ncws9ejFZWTZS9bjAyKM/yf0cW/kKAjaLyDOMpVfeZ4MGG21mloUK4BtwbPWt9Cm0dpH6Og
bzWrjbsdQXnyvlXpuHrZcmfaHlAjzaaplg20hVlygVNPKSMxmG09p5wXNlK/ychDudhBt0n3UnK5
G0Sb1sFYn7ssBNGd92NtD+wLUUcL5ZDimiNpyYsBu44M2pLMdt2eZNMdtZ+IW7qniXFco38VyXDL
R3wg6XJSr5IRp5N3I/PSFsfqVdfreFrzw3y3PX4QYKrZoEX9SlL5CCQJY9L5A3MRLEUg/7BIjb1a
FGNnmY2ZCj/jNZl53/A0wA+hrWzLO7Xrg4/TlNXLT3Um4ycFBByVanYfpxFPC109PtCKLDFCe4vM
Nz6IGaYkkoAox603XicH/5AAsjllv99tmHdwJhqkelj/ZO3jPiFBYTeQV7GdCwIpSK/fBWNA1VQF
gJNoVSm4qdbFVAsBojDEQ16TTcDhZ0Yqw/8s9jQbp1IHWK+HI/NEKNdUxCKeKXRr+v3431X6fSqP
huDA1tshC09Fapb1kPLG+4baO8dyZP+TaVcWEi4/ayG/0hiYkIC3B9GQbPX+dAPXIhgdpWQ6hFZu
l6jSHiaiRLpKqRARu4iESazctqe9mU4Ukn7wbVw1SNasWV+Hay5q2qTZBpxxMoEv4cvZW1loOxB3
AefgDtcznwyYFO2w1Fj6VvSv/MVey0NfLPxKBa4yOP4sEt5NhYVirimh34YkIEtLvTVGFlGpLuK/
YusVlADJsNWzBibQZjpTeJnCJy5Mn3csPE3xtsnJzvcvj7RZ/FxPI658eIWx1ht22bX60FdA0tZI
+IWb9rHtV9faxwnJ+xLr3Vq5e47izziARG2xjKlvUb7lNq7+0SXcylBiHQEgQFT0VZsEYbsAJYEH
2QcrUbnT8PCRDdmYy9pm1tBAZtBsI/fy8qgstQ0M2+BsRcDp7xNrD65Tuc9uiUllZzFosraqMD95
2OXZlVU3fp8GnCEwsyRdarv8yi9Pr7Mbmsp2w1+WPmqzvIYhBVLkUFTitzJwAd+w8CcYfhzMh8Xc
fa2o91fi9BtSMSNOIWmaDo0CqzoFNfLgrresdERvN9NHnnGQ1imWxwwtbgZ/d3MFVJdcG2YuCG7/
QbO+KMq+vD0Ktn0i7ElPX6He/vsT/WiE67inWhMn7M8JsZZKYpZDNDpwp54B+0Dvc6srND0148qA
DmRf2oZ4syBkWb5YhXIzDJp71giKlAxsV61epkeyk30bu++DdyE+yv7NPHtKuu04hU7W85p2EUhD
2JouP40cM+mLCvoLltJuOwy4fJPkh79uK3/ShbDFPsMwbGskFMu1d1AQzJHDs9Qgmj+AdwgElaoV
qUEe3oS2Lrq4AviWyaeKpqRqndz6Yd6xU+Kbn0MDH85/Ci1imeOw5y/O1h/4fT/C6a4V3UT9iv/H
m+Z+5K9na98gqimuQXdUmxmqEofsDA741Wo2I+VMRDbRiB7HCEKhHyqfZ5uiqyhbHdUTLlbuExln
v9qfJ369j9JINdZC67BbO5Xwy6BEj1UU2qyJ+elrlit0IXuPuImJWhxzsBmcx0BiGAim5T1p7OVy
pKpLo2AS/zf0PlbcsQ5bLL/W0OHLBHg/+zMmYQNtdknS3AKKglN196cJaQKyJLZ7157RD1xSdpSb
CMfadnHKhgxJctNfX3cLg2wFysxhHtMxG7vnOZrchGfwk3o8fQnVgasXimv6hkmMrKjcJGWE0vez
rlwKNjyhfYMp3ZKsZQFWwwIYEuQ2UqXgQT8HkqawfqZhZHhKPilcGkIgOaYyaOi1hcaOZcbphGSj
wj6ZX1f972oyE/H5WAeV0nsVKiY2qF4ustMRVEuW5/nOazO78TVikQ80ydd6kK2R1liiyUOXp1HH
10+tyesjWxP8KTpXNg3bW4tOdonGc+GyJhkNAgroO9sjyZ7j70RLBtspPiMWerSSXnm3KTE/g7O2
FMAj+KnqnhP7+YGToYll7y8UkrO8EyeyKGQjTovYPAQr23BCzERVEbhAqhZT0Pt6cWuLgZSwUm8L
taXs8kMgZo2oP52pLZhlAIZSpulanP+cGaKQ6ufS+DVjYhjZdClUJdZkhESKDMbnmaN9jsjuHsPa
D2jDc3cAbZ9cIGLyNIb53zqxh/Thlxq3a+lYeSXtYuxMFQC58KqEHVxepjV5Y1w+wg7xMKpDXim5
zPpF2AjlBGlcmiXLgblST80Dfk2nlylwt+4mTFXO272wsMIDGQwe88kRBqkwAKPJnlyEkCg+ifK2
j6qKePIM1Cra1YJZIE7EnkzT1JN47Lhw9WEZr+qDvacEAvoZkAen7E0iHi9m8hE7mOp5sc7e2Qug
tIaCyAMyzp8sqPuuWk7yXt9GVoWTA2nhvqogitiAsSMLjHytH4ZmuyqcvWcI+fzPapuaET01/zLL
/Ac4PNXfgGmhAvBpWrsDp+s+zfjQ7IGSwtJfYu3n/G8wU6QeWRprVzgWf/psp4P+T3+as/GkWz3y
0/x5bART9T6ENLi0m8dKYIc+sD5EaSAtzNoHfckAryZ5dgkc/WkhBcmUAHhjru8PEjBXz8rDdbFi
tLEdkrVPbfsd3dga7BObib8pz5nyFTHUx/HlX9rfRsdGxWwy1tmbD2s5ANsjMXx4K8LwSz02VqDu
hFptM6XLie0vkaOPp1kX48Ii2icuVe+BPthQEu9JUGZybrFNJjfXLo5UtSsIiaUeW7QZvrBRIH8B
MqgSoZdvhxQ+rU0+K1RiK4TDpzH9syFsfyE7oOqdNIyjS9qNSU2c/Q9rH/bb4b3jg/7kcrWZLpCS
wWlsdNsPAa+2FnpMzkHhm4m1ef41RJWJqF+3PdP2Vgk5fJTBgyZ0buNboAIvN5onJtSCdCxHl91u
bNOh2Uv1V43Ctxfm3lI0jsdCm0mWpgyuBYCOigRj3GhhtWTcMoejSpNEOstKATilr5E3/9T8wL1a
A622v8pqhvDjgjVq0MC4x9IImT6CJVsW4JPg05kyZtmTQhbfwSetugTcYUH4dib4cs6nV1KiCdCa
aoMdiTE4znLugUTn9pYsVJ5+0tdcx7f+3ttwUnEjUQFMEtaemzoad1InYJMNSMHb/5NWuSYaqimv
uaEKcxSys71temMn3DKMaCt7/+BXrsG4IpdwWFIbmKyZk7KKh+jwhPJRb8TJElshtFGiLl8hlOEw
s+b+hM30Z8TrGoG//CE5YA/5JqIu/MRDAd1Idsp+fid5VRjQi+klCU5XFCw91Mj29rATNImpo0Cp
PGY+cx8ez3qPLDiofUS1a4r03R+IUJ8bZpuqFsK6qpnTBlpgboTOMRn9s6ABl9z9HjAE2PkUloqE
LkIyQ7K4HCK16Eal/oiWm2GMfoIociHLfDT4XYl3HE9+Vj80UHRg7MaYOqr5gjgNdt5D5vVTA7w/
M5l/psl17NU+rK4+r4ZJuK1s1+RU3KbO4LyDyk7LlNZaG5XqWMj7RRnuyGel8IDM5VSRylzb4dcw
75lizAZ9mc4sVUBbYooEvS+ZvrzXMvNKx0CBeF4TQ+q/uULHNFs4PXHa9C/tiUhhokX0G/lzHRjc
EsOw1ha7gNp/BigFAiGJnynSNDwHMmfLOACLfW4SVXLTfLpdSUb3RuXRfeqlBzsCt+/l2SgNge3P
27MWy1aCIY9z/f8jKFnyY4WXmOkpO1M6Q/7Xd95t7uwOfogGni4IV83CY3YZoT5CBgRj0FoOADui
wAY9rNE8tZ6cK77NBLItj8AMDRkOFtzbSnRdmQdpXbKDzVZ3jogH/zzbJYPj5I4NprLk3wJN5lQT
6EyCaYZHYa9aYTHLRa11FT/7aht1HK2da1gzIgnzZt0tw7yxmkZbPSj7giPnUTq+Zei/iC/JuDgy
pu9yF/qdFma3fJ5V8CVtaZT3AngRXJMyYDtPq5fOh6OguYgNVk8TspDZp61sqh+mjtDvycAG3QPC
riejzzrkMkHXcor8f43YPVDjnTFyenZck1Unn88C8waEqZX6Q9SoFQxEDrTi5HW97aXaNHsXoQo7
OmofqK96IKYxVvmp7hEgAoA2/j4TWDgbU7ByHQseDRqAVQeeGjfwMKjWe23wrz93HIOIO3q0l/BZ
urDH0tsouIOImUZX8Povc3whfDaCXXfPernac23+HPk5g1s/Ns33SUirVdTQKk3eOiM0AKf2es4H
jbkGlo9jhvocIxK7d22ndhFHMTwc2n5rfwcDqyYCkiUfH090Xxn3gO1Z2u0m1YG/M8oT60IppyFm
52zq40K1IDUDtN9gi/aPHljfgroh1rx+2AM0RvNdJqzDf9ISA9KkWV/S8qvqx7w8J4jC6RyY4VsK
GSP+c1c9TEfl92uN5v1XEQBZl1asMBhk45pCO+QQi1pHT/edYDPjSqGGJd62WYAjw8BED10gh1xl
aUnHZ9C2yypuWYp4ZZ/nKnxL6tvZPK9LwOc1H1lUYkfQuhQ5I/BmIYFT3MMXcS0EPaiYqtMFcBlP
DclQ+O5xIaLV9Oq7xez7xVabjJum2pqT46J/rY8BFJ0y1dtFUwQZKSurLYMKbWbIr6jniVzAJkrY
cHXihtLegBnOo9cC0RPptmljlQ/4B1IDaVGzd4NoMa7q6ZaCd5AsL4QPKAF8EwMsuAJe8ru/xxp3
kXLXApb4AgSLdwcje0PoZXBdeeaTglGeKPdICD9xtaq+gflBTxdObgzIdFTLa8cs6amM55v4ozK9
FEPRQjTMr6Rt1fKN4FUG/EyYutA3OZR6RL15nGWbH1auzgv5DE4DoztEnwpU7RQ9EARs+WgcMTPW
QbSti80/OJ1M7cBX7wDtG8IFHHrq9EBL/vXnckAJMVzI4tKrBOPJxASYKyBoj9JqLiEdtxiI8JLN
Vw++QPFe9VfznBi3BENN0ufSnW8aJ/DpwypRb3UFsJCmG6BlsPZ7Kf4lBLUb/yoD7mdRO/DVzqMw
qu0DQD+/SvW2KxkEol8g2A5H06YTpQrA7gm+Hn95kqvze/UuM3TblAXNocMcf/mDgdl9zWNLBf4X
gtbjI3HiWg6EyQ4M7lBFYHw6BoF80HnscLVtJmWjyPqf/a9mtdNJ8BJAl5BMLV041MLSK3he2mgT
yXwXX+NkKniU5CKbN8QCxuyUQJPkpqpOyVBV10IAyLzSvKhDH8IAMMNHQjz2DXI5CsGNlXvnS/+x
P2Ln1oDCKk7VIIYjIY24Tj9YYzpl386yYHs75tF62lnJchwcWT4ILtyNI8L/hYuK0txuf70PNDR8
l6OnaJS6qyBiR7qi6gGtKbMdzXxf4/lpTy/sKFWCIg2N4UtwzfW9oUvS0Ul9CC+05FGceqS7O1xP
yiu3BZfePPLbZScAjLUchrXtpOWmNPGXZUTOpwnBGVE/FVTvYd4inmGpNi6AeKGicSKDU7JpD6pn
535Myi+qk9rDYHPtMwfpJP8GUzf89oHDjvKg0MgCcF4xYoZp1fI3TXYp6Th1y3uvNQnAkKg1qVc0
a/MANiZwsRi3XWd9aLKtRBysgQRuue6nMwZDQ/AUDmuz51hmdc1pxAqEqY4yMphVECccewHl3K59
GCnSTSlTE6fzlLW6YTmGeQgW7KMzaSEWKJVCHV4BLWcspEOyPpqKoRIttTuoSDpDDXn+orsnjspu
TLNW2Lv6qg5TFh8b2lzNaqEhVNPlSd7Bi8xJ+k5dAEGgqDV14lJLZvXZoovDq4Yfd6hIm0SbxWCI
FCjeYJC/vg47KNJS6zyoc2glnOrXw7ILFfBXEDcnUsu66jQIDl077sYBZGd1+2U45x52ZcVS3Wn/
MpHqL09QCjHXfZe8DDyQMqQ212car//57ffI0lX3XeUdFh7p96NRY5pN0ZPOe6KFWu7WLvIZdHvN
ozrl+G71IMIBcvZf5HYJxDX2t6PWGZOZ804Y8xgTxTAthtt4Pf+mHg2xeMHUmeWIHbKV8mUmirO/
7AXQzqe05/z6YgC8mZvpLqyM2AbNfoXpRErgzp3RqTVtzAmhV837S+qOTuv8oK9bWug5ktJ6mzJ6
CydmKhsFLjLMMqLD4jds0qS8wdaA2TppXem3veam3+ThDwhgqGnI7CtJ7pn2FAt/xMgTpoZjMjn+
MiSNJ/LsV2bTsPBTEKwmB6mWsshN5vX1gst4/uR1LA43C5EOvL9NoB1ygJThS36XagMeX7H+rraP
xWr8+gdmBvrt9ySbRZyHbM/wM+ecxtmyuueoelUBrxN8SALPNCRzV/NReeajjj/EzdyhSyAV5Op8
xopHYuUoIoeNTsHf3yoJwzM71ccIp2EAN4Lr+vji53byw2quTjfpQiPxMugcdFtuOuYcbYbUzaTn
v8HhVXEmbPLv5JEa/EA4KToIhugcIwydbSKc4DHaA03jUAPCrOsLyRDY0R9zhQ/rcZ8MMnzd70UI
idGuiZmNI1Ad0CLlxWNi43Uww4pXcARUCjX+cG7UiGKGE08I2R/MFNco0+FjDyeZjBqVru/ufRSH
4mQFUZbl2TESLUtR4o7Qg0EpE+hoibLU/cnL81Bdku69c5KFq47R8/rOBZ0pl5saYz36QgwteRAX
6qchXKrzPPs3jN2S4WhPSCWgjAts9o9KMJQxGbKhXfIg90CMWRFTifxsNDE2Y9wagVGLaB/ZripS
BJe1xWXmbTodpYca2OlckFq8sy1mGJewFiVYJnYy7mR3Uc5p3aA7+X5MvDZsc/9cLt0ZBJ+baKKh
3No/dOrscQXwyjc4gjFuP0zVbpJ8vp7eEQMrUE9YaaxDwYm1K/yaTRHZdyXTkl9k6rUm5tNhJg3l
oSdLF8lDHcmColyk4qWGUkv1244496qxf1rtM1zr3D12zqQi/UmERYUKgwjXu9KnaVMwHmGyJPrG
QnWT/whVO7XAACMjyYPvNnskHX/+JJ9L2QzlAg6EqFaDU+zhZ+9j5Oh5/Hn0mu4zvsBOnEFyUbFk
hIk5sBx8S6RVDXryUB282HDM6yA/1wEuKKAJTuzQaqN7g538NEjirTSgKaiutIQQ2ImmKSI32tzC
XNSoffoxpzD0Cz5KItsu7KpsdfS0cYTqi41KTOtaxr0ZNZ9E/FJWMWOX88D3DyzdyLqBze4q9e3D
e2fHecFTX9EcpGb9F0hjEWUKbi6Pq/zVTKAq2wMOgy+tgP42V5xL3Hp2+LYnEvT4wdXKmfX99FNC
QLR+covKD2tP2BfFcF/tav7qnY3qc8eMZCf3pYZ3+gShIu03AB01NoQgrIrMfYdTYlU1LMR+gXhH
8eT0hWA7CRCak31ch9Pw1lNOb0m/HwOMPoK8SlfPos5wYWkPwG8LTFiQSeWFG6dVJ2PnWqtEABPK
hsJhW5KM6iuD7BtLodhXdASvL5OA6JCWJInX1cfqYuwksNR41GPU9L0JbNQZ93ylTJtN2OgQ4lhc
gu3ycsJY9m2PhNwD1kUWAIA9qz8Ur1zhyZj+5RwodCJmZ2hCbdia1XccnQoX9FhkE3U9i7db/O/Y
uHV34TYaJU0u2CTzMUpF9vCXmSUlhQnVxIdYv0FGHoi62RQizxHva8GxPtnIb7sXO6PM1iZWeLWN
uzk2XsQyVrj9F4xT7IJYtd+FtsQVhMeen1n1bL/VqjQ3j0ZPylMzbraP/teASK96IRg7ijHS/bDL
0VmaZS+L1MEyPl8woraW/7wxdq6tnmU7nac8NxtX+4TAUziUeIpcjn7Gwb5mEbj1ufLIq9vYkWi2
o9W3rogs5V07GX+IwJiylYGIji7zoIq2qfe6IOs5GF7yz0VnEV60YpAz7oNmZ0Xe3yBamphDCSmp
tdOl6T3QU8vzQv44JfwSjA4K9B0XltrQfN7EEfrVXJUE3vQYXCqdFFn6JSrYdPqlvbTlFPq/n/jb
0UNqQzr1BElh3Zh/qPtPSAli9i8DsgsaHDAL95aaKgmSxFpXRLDQ9KyTQROnnSGmdFsHZ+HQwhJk
/eVIvBKe8baXIZvS92phjl2m82fAErTxHuirpZKTmQIcuO8G13D45LmorPtx9mzntXlEEpRn1QKm
KrY3m10bzyAFvlNgn3KETTEhUlq6vvTAshmlRSsNrGQ+1LqDoI6A9PM3LtIDF4SjHZa9khxeG7Wi
iCxbXzCaua7YxvyGrMPfqbphkwctvxUuNKmRD+Qj9jPWXwi24R/kpL0wtWsOv9/8ASrgART/RPoK
EqYavHq53M/ZnN3ngSTGXXaXqnp7hJSjPLDyQF+zwYrj3b35bC87uimvsDdaDf3RWjajTy2PDOy9
DiRhQZglKLEGJ/Tiz14/C9tJGfxnKPUrbx8kpHhIwqXzbC2BT+mdpTNj5Nur35uY8O3LgGTUHZLx
AnrBbf9s3V4cM9c5ag7NAuqdp9yB90rUGgLUOd28SoZM/pz7Q4KlIu0+QQBqVlXjrPlh2JSPmM1I
XxuBbJHnjqr/pNm41Rqm9katFHDSWuc5rJ/kMqpLiSi8PtVX8gjYFy2tgqiDyNZFj4PImM0Yj7AB
d67cYLNt7NGvSSf4Oq0+O5xWpjK2gUOUu8hrNjIBhGp4hGsQw493DnURkX03kYLfObwxZVE7AYki
UEqyZx44XFdkV4+/h7axJdAQ0KKlKbTukgUQD0rJzHwAIfEMMF0HH2CncJDDWyqErU8PHWDi3wgs
jp+mCXhpEo2qFY7LqPL5k6oiJlrZXL9JWFiV2EERlDs+QYs7wKq/JH/gxg9QEPYrmATxDhJX7G2i
6GpEP5MhpriYLuzlXzsfoSQ+jL+64Xf9MqaJUDAJ8oqUvtmhNYSIkkYx96yFZxV8pgrLcdWHYCVG
HEdo63TvOtC/7kaCk3Ia/c4oRNIWfJl2Sr3/OBwtjDDcSQesuvWLb2yue8ukV3EU6ZIkCSgM9FYy
c6qXUIp/f42TBoBoEunLK/hAoVv88M+TsrdRPkGFluA/ukSZOzQWelcycj46F3MvSmYSustdg3t/
MpTEko6RbKRsszJfLKRzkwue6VT7M68WuwHEoT+Pmi4xp1QebxFLgkyOFILoYifzqyewHDBfYKbV
tlG4xbVl1dYY+oGR5I0zatX6+sxrbONRiZnzy/FIpuC8+ftWppdOZALKnhHnqbsiWvpOWHUa6QSs
A9+5FwzZiA528rPwck3TidhqMExTXlyxqnSXzyem6MNAWpz7lSP/MRdaGtJ8i6w9dIjlwp9BcuFx
2TLBEsPbj42u7jtvG+k/SNo7s76r1zyv00A3wW3JQtK9N9mEkesWrTuhh2zAloY4LA3+3HjexMrV
w8/fdYP48E365bTlAYTkOE/P/YF38+6OUXHYjEY1FhRfnJ36t0G+C/rfqhf8dYXq9Eunu2dJzyAf
+Pmv0w1CgkKkhz2vOqoTFajpVxvpnXWPrLXe+lewuaN4dOA141ozUjxl9cLXhWJKrNnNIoqZeRyz
r1pvOl+bjDC2pf2wNvRR6/+NBincw0J0CbhXuVT8Msrv8oBiBP8OCeBzmkUURexCz3s9AkQRMKsF
eMP9iEI6oXdAKhIOqBMvPZXmbYgPAe6nfI8nFdaY7R8z6mdC06nRAHf37g1BgVSVl4czcqD6OAwl
wDuBAVmp89usMWXLTEAhJft7tJpI4nzYc0/bCZqKRFxy8AqLHeT200V5jvvh0wXko0VEv06Bfo2L
EPX5BIvrVrK/tD2TeUgRHtl7YQvpvD3Clai4HiVrpvxZ97Mx9OMlSpYtJPuu4c3vWP9BvRUJt1d3
q42vO5a4vwjyix1jPjjyF7UBtzrrR1c4DWV0C3ownZmEheMN03CvF2nN1WEhPDS2eCvVliwRsPcU
25RjTCn4CHOe1lzwRJw2cpT7nFvJZ3F4ONG0dtvkDlAJ5W2aubPgSVjZtFMJFXoT7lNEhGx4Wlro
shhmWODTaZ8x45thM5sLDItuOLaVUk2NLDeXvNvbj5JOhSHAgQmpY0AIa++LPO3cFs4AaEHtAlKQ
BY1sunYul9fpMOQJgGij3kX8SGxVn2xEa9+VLqoz5/TZ6YX7/oTSy6vJmuruCxBC93I0SMhMNMUC
P6rp/Olx5v/KpVtZSQmJy2GmzmM+CSZteOaciGTQPaFYlt4ELo7cVotfVrRhjaHmZS1KA9c2olya
E9ySWLk+cg0B/2Ye/rBQzM6POIvP9UyUrPNTCzVizXm3Za/oyqyMU0v91zJi8Vhcdyw93uBRM3hY
Se2BiUSB5iq/e0Ka4eMmydOZAr6TUF7KwoLm1BgnVOk21G4qRh9SONVm26Hz/GYUbPKu19bPDmX7
4LoTpLXz72meccWK/CL2/hsrR0gPgd4mXnIp6h3sunfQISfF1FhiyzLFUuy/1lXm0gqFE+3CfS27
Qy/tKZ8jNs0FvAHzlNDVl6Gv9eyl06+GVOaFJsagH9F2yBY3B252M3tbI+flGDEAOWNDUOMYStpY
OatVz0bjv16uPAesfWL/OFVI03bbREj4O89KF/u2uUywpm2evTLNmFlvUZRiwpromQmBLIpuF/76
+t0CwXWq+8poIx9pP75rYDkFI8PcKSVJJJyRUywohxjJ3sEBNFe1UYS93aw3Y/KsHaXv2QetxgSi
+sFl8pTv2igYlCXxMFyauzVFBwvh0vo9tiM1FNCnQDUuetzNHcaxDAa8ftgnAKVtuSh1d1uJFNFy
Ly+UHm4aJcEypUrbwzw5ptzW6DabLRXxLtwSr0V7gRZGAGZttOpIDacUyLvaDHBUFwexVvNuH+sW
10jtEnjJ47/Fvw+UGirrvx8HMSKQeb/NdilDUon+AbFFlnU+y4wCaCv+yee0cybfZkMqJjWL9w5W
X7xJlgwncPP6x+Dcjul5tMbZnlYjcbEzPe5CNGiLHR8drEsaS8iYjDY3iyI+orTL4VzTRP8yr7Bi
Sm47I9Mli7GveA7ESFZabOhc6QrR0btwKtmyw1CStxdRN7A+7qholEYIRlIOqUwifOWzqRgj/scO
qWTs0P3flJz/7nEsAO3go0I/zuhViOXPG4W4WcWKjQC4hRejpa0LYAnyHBy2j/qtQ8sxiPbj/j/X
KXL+tSrKY6jn7WTsc0dD/71u1udcSr6aj9OMJVfbpaRPLYkcDLTsBPLjW8kMuqYaEKbrYmTBSfVr
h4hFp/SNHif0/+zu+/S2vpSgb8l36sHcO8vzdt0Pjc5I6DDL6F1oR8HXCe0QJJKz4ZNYD6YYDT+U
ut1WpVwg9fkG0vfTHmruunGDSokZDtYzTtADjsNBW4kLUXnTqThz+mlkLvC+suGKMWmHrsS4Be5W
xT0wjUg8mFY/qsDZLx+I132ojKH/m5bK+TZiQo/BsBGWPD2DM4LhpQBggy5vnHsL6gt0Qza19rUQ
8wItGpVOEIjAd0+WVrxwBGWiXVCjcN76YXCrpQbSPBmWMpwExtC0uma05krSoh+nXrd5c4ZgJIxp
Zxxyl8vLAXi4Q+QDimdgWUc6373CCiT9cWC2Dw6jQgrfeSQJFyeLjEwrktVxhq5Ug/t7tBqsUudO
3PD3JUnVPtoO6d7gqod4FD2DsKBDDOkwmn0tJeIpg97dBg2a74ql7IGW9Mdr0DH4tvRkAo6CVw3Y
EXAd/As2sWsv+d+L9hJOqp9UbjWt2JcKEOnzqOzyqdKisyuk8CPNTZLyQXW9qpCsqkuV+AkM4JhB
zLDorsF+XTfmAnrE3KAmkM3xRr7Oexxtb6da7Qz4dHEKvGkpsQz4YyNR/oskJAr1Y7vD7Sr+k46Z
TVv+ZzojR3CTY4CFLvtH5DzLds/IcibpzoJis8l1j0OGYyrNN+KuBE2dFMrzBqrhdPM4zBWCxgt/
s83PD9OPr6GNzBo0Xce+EimUczU1oU5QJDcE/VmYFlYO+laOFTKlOq8ZS4SDF4T5DPFFE6Hxk66D
uN8iO+tBSCXIaGY8fLS/4ZMM3PRwM6Khul+o9NC4wchHkTy7aJXvtfW2QMu931PqlhX1bUTk2PbX
R/iWDACUTxY010zT4VdLVBDu3SZ6RZY1qGT38TDBRO1sSGow9BQ3dOLi2ly9Re2GizUlGIXVxt8Y
hUqsNTTZKL2O3kQwNZ0ykzTrL1QPimpkO6r5+k0McSjQHbJWb3+VXQjUnZqcVK7k3EIKIT4nGsi5
diRnN6nNNkT47+p/4pGY6FBio06g4ComgwiPPoXUFgJ0h9uataCUSOox8JMShkQNYG2govO9EEM6
yU17gk+V3VQjd0gTnd5CXSNKQdrOB/Sc86IIKLyLjFQXQSx2AUSaePYnIa61lOtFSb6s1b1x9Oa5
xXUNJEDItaaxzI1deDXB4uGe2bYeT/hOB/D1LWq65sDALRFr2MdNV/+vlXwFyf8PIpjYaL6uLTbc
0QgmNGkxgxaFHJ17pNqRyKT2cRgYxoK8CUYlEAt8zXZU37Zg7J375Kg6Rhmahq54m/nqYY1WFbBq
32vjCQ7+0ECIe7d6x7A6HUHBtlMl48FSpNS8EY8trJk37Ww5OX408RgjNZzlq28XJ+8npiSJtb+W
QwF5hlimKTyI1j20Q/F0XHNnoNComtHHp06v/AdsChv/64E7dW6m8oo2JcjuWcgEbUG9JeCUGxuj
IaPnCcDFZ9mo5DNkPPyvMSZkd/UCKKUOOVxudEudvsfoR/OR4vFVimIrIKyaMOBCwOKaamVKBmPj
hF9zZ/xPwHG9vipstpg+MA0QJeGz5pI6oSdg2Gb+7NTqMNuO9OdQBiE1FNOo652VKDMtAXA4jSYN
QiIDPiNNFuuVUtNmPPC99KqmX5uL4zIS5yktQNi5vwzGCNzYT9aWfNnLJ+LOy1+2PVFfnFCO8MYV
kqos/YPxnkD1cVaFLsnsIhqHYsxcPb8ZHoalaiNQnb6BAGKyv4EprLMAYqSYX7XZANc6qqNSEtmN
8Io+cFnSxvU52r9dye5cHqJnZhHtNhUTmSZ6xyKexVm+g+p6lVF0PSEFFKY8m4nwlmXwusTO35d0
Yx5abDZzN/rTBz9rNtYuNL+aoh+p5MYaokWm7sIcTo4aIXK24W0peD7wWhnwqwEKiCk4BCqTthMl
SXmkQmcmErOSUReRVI5CxNM5w4aVxSZqrzYWIAimLWJannfyVCVnTjArOVOraXjP1ADqgkdPbhVY
ddpiff8nvA69WHAqo8UOQ8O0AgrfQ1XRcQ2U+yhhJCOtL+n2P9FW9/mUZEOERHEHiExe8KiUoZEy
sRBAHPbC9Hy7sS+/B3patSdPOI/wj2PSh5Y0GOuiH/3EP7wEeaoD7Id4bKIu4epeWFzqm9QIszeb
uC6Xgl1bYEO+2oDcxYsVr0QrTlaFNYKwc0yUM/ayOk34kZrQ1udnbZoB3VQ/ASss7UC7ie3MSHej
MRWF86mpH3x/i3US8Mc2rHMXIcWyxLGOH7xvgOgRvIFMYd1LoOk2N7HF62vJFjK0jgrLgZE58HQY
E6T9i7dRikFqwnlM06u9hzGrDevBe+QYqyuJEl8IoWROKKoLXdNUfQPaIu4WrRJjcizCoLLku4eV
w4DIflNUaniZNxFvQpLy4AKHLT6uDw9bWLexSf+6LUN2fai+F5ROKLruHn/WqIMWj0I/pJtsZ+OK
NZYoZdPRRdGOpc2mRPqgBQ/J4QwQQ0TQ6XqqqnSAv3WxOxjCUXxvUYpz2QChtkjaeCLdPrLplyY2
7HSMd+Mrhj1ked0hMc+jw7VC53FVm2QvH5nwZtKGyYp59MMafQYveH+pTISQ4wOAHTdAZez1rsoH
m1T4spe5lMp/EPvSJsy/aqi2iry2uTmJDWhxPj3s0D57D4tt7VdyJjFp8DohVWpYh3Pe32WnfaW/
lh631qHC69ujz9qGNDBkiH1aKSydLjfvBOaspzLiv7ZGDSfENJGeiuePB69sj3Y5hmhN2AMa4Bcz
/MD4mxKyU3lfoKiWXDljn7BPQRBvWvcvgPXKlFSuw++l2k1ksl2VJopu5zUZf/GE0/KzLr9UqNGN
nBf93n3nToGBsOS55PXsyIvTvKYEr9rMaWyEcn+G5AndXx/ntpvm7HreFdFgwYA0wvmTjRaMKeFy
J/C7NX2CFSpH3L0T/sM3y9BXy1i3xzrck0v2cMUqyz/PYcowij9IvXe/0+cc9fT0ISG5heK87+4g
kCsmQoZSqcqqqwSImt3nIIQHLFPyv55L6r+ixrgYOtSKZHsYgeBmfRDDK8Y7nOTxBZidKX2FFcqy
6+tyO7hnDicitfQjNTV4GTWRDhmXvGAo3XIWcOBULUbtaAcdFIiziQGNF5LB6t2tmSWCmhrms+Ua
AlNFh4dNdza3+NJcOc59bLWIRRFwHOcNDoX9d8w83oLS6sxrdYwwgzyI7o1qjW6PvGY0Yl+8O4/Y
YAuCERsTPXllhCYi+vGob5nYqXPCD8ZHWWHwJJ28VdXBonF2oE1iLqNYGOdJpmDux1ao0MTFfY1c
EiezSEkhPyjhcUtAT6a89f1gUyElE9+WjYgLKLeSdAaQND2yAs7Y+uyn+by/q6+2e8n3QRiZne/c
m1Ti5P9bSCA3h7y5T6tmvsCRAKkifGZfx9k6tKuYA10PmzO1jLAAbvcJ+Ye0XYmZQb5yP4BjE64q
zbR0oCieEQjzBBW2a1tfPth4vJKtHUSc8Gz8cIs/TruCk71L+FkdrJZRL+sLfmNT31z2k1ANxWWQ
vrYue9nQmZ6dhIFUon5NOrUX4EbThvWmTm3R970NyU+FNDkppJvw+ye3pEvS7+mEg/8Pa3iTDpKb
960kWgB4K6/2NpCTyhF9CqLuZaDcTfPe1woq3ywq7ZD3ndGXAOJ2+MmLufE0c6HFHFnpOa79dNO8
Io8IOS3wL7d10VrNMRXpd9o4qjPoIKlJ2jyPU0RX7rIQ/1htvDtvX9zNo242PXvZcGhzwL8EVcWK
8lehjtdiFMwc1KLG9D9+QrgcFfvPLobLvq4N3SLpFya1qVUj4g2WkbmJNws8ra84NRKtwQJRhh0g
UWlYKW1LzUwcduYONtz8euH0HOBy1FubmlkmaNfX+Y5P4R2pi3RTChcfySdjW3YIFBUO9uN6HrOl
6+YP2TKpN0xcVpQsR92aNzFGEnnlhNU612bS8aXOVYLSI/koJj+ptwF6JUMj4rYSXRQL/5H3UcuP
ZYP2gEVHuS2AXpa2zdQGOFI0qBQ2MmYuw8bM3PmMt9hd5O3Yy7PMt93eytPxFPHE1K+HX4C8LV9K
QEiJzgrKnR9CBfGNHGCPTVxBlieVBk2cGpOxXyH8NpDhuXwi1gLPHh8KjW+tGyYSyywfQQ/XLx6v
G8uRUn5X5k/3tDAV0MaTKBc9EWAb5znZhbZ2/4sB8XEM7nf8lRYfAXoIoVgvZDw3RCAzrBq65RGY
aW+qoYa3V0m7EIRptZwxy1oeWNY1PCrncU1QCH8uc/minxKdNXLreoUNtGHF4jVGnbkk8PxGoQNK
Ns+ujgjsxPUy0OePxD0FtnzwTQibxFN3Mv1uczFMMl7Rj/XqJbwaWO2gw18ZnkvMcGV33MJpUu/c
BTuH3QM89OPyxk6f6kw/LfEAICX3qbnQ9h9CC4UwUCzDzlju4SyxmHtu/azpN0/ArDrSIbcmot72
hf4lj0oP1Q36JDYmaM6I8SYeuwfzocIrpeoUg/rIRtmaT+HQs5qF0UDxFlZ7fOHcIexVhdF1wORc
IZ81JnkVeNl5k8dpD5ZqjtyA316bsLSn7Oy13E0tvfuH2AWveYW+BxFyA6ZKnlk7CT05lInlu7e9
pPf6+BleYabLqbrXqfduyV0HBgArd3gGmCnIrx6e4j9nZulwKeOE/XrWbTrIthMZHKVLEGtpipXx
MSv0G4STxR4CGIpVSsS0cLkBKVzNhdNb8hM8qFbu1uSlxec7p/5I3+skNhQQN9AhsqZmQieIopYb
nWgxiMQ/G3cE6rHWJ99PVvNK2NM39GBU7MDzv6naBAiTI7Wns4pxPthpQ4IH97qTY1TpFGAhQa79
NcK6/r7z45jnkenXt/GgE/Un8wWOOI7VDZltbMH5+6OReLaw8iAJImh9I7Wmd3TpftQbltTLTP52
po9doFpka4WqHMpmznWZwTiD5QZVJrXLvBfsZtK2FPWs6QcJCJsjtuuLRtHmRpmaHVUfy5d8WZ9c
wa9wRhjNRhFGq6nGT0Vy28u6blNsVM3g0YegVeyzYYzIbmPjbQI0VrXwi7+jokKEqAxrLovWhT84
hTsKqYeVeFrymjDMCJ01wp7khe0EUdmj6EItMJBsg+z0UC2FUX9RvzAinelrcojycj74nzAHw+HZ
5BToaM2IfBtAW61D2kGAUsCu4HhQyTSMLIvL/+cJmGuPeNZDiMilChRijxmjGGp04d6d1R0xDZ6T
ESQ2jcnZ1XqHjnNydwkUcQG4QKUKQKZGNPfnAN/LRgJzENZ794dF3Aq4ue0FCGSqgixAZn4Nzisn
Gz6fnIyJWpYUrhZ9R/UDKvOYJeTBGdTW2LzvvfW7Ii9wMj1WIipXLP4ZsXzq5r3bczuA/XsZ+pU6
6z3x86jIhxYNuHUlk8qVvTd6nxP4mQM9dlYFN+I2UdTycloDm5vPCQeqTLwEHF8BFXLPpGwAF729
Lb1r1g+i+ylZVkQZoxHd3sQ6E9Itq52SMaht6UOtnY42bDZ3THcmH0jn0Q0SUUsErXcwCr2lzQLX
vTrNzZxl/BWyjlNawniCBlVe+fBl3ZRasTE+gzet3baxZSpUs/MobRMD9ZzheiAYkIKkOttzUdH1
41MQVtu3UJnmsuHraQxTdvJj4O+iVW5ztIXpoy7J0BQc4UjpLYkSwUKJarQg47wlApOsIHC4+Q3l
UJehbWc6LAUY0A1+jR3Bx0FzRR9Ibw4lFc4/7BETiXmki4HUrXTYykTRO+2703r/cAX+0vdu4MvB
Wo4CIvEjIjMJc3kv2vk3yTA9v4U8ivtFmsFdiAMM25P+LSZnshaBMV/Wfy93JN78I34K8Cb0QqIh
7untpMG5omuPuVQcFI0HAk10BVPPGhip4VkRsxpTXCfwTgPhjnUSm+/t9I4UNUw84iR/yeFm6SYr
bEVGACNDyqtSsiB2frOLWXzSjA2HCj/uTBIMv4YGPJaU+OjuV3+wJgz99haKtYA861upHC/4Z2ap
7wspe+EdgyBYmmH+u/m+JgEuGv0laSRxsGUSLV2yAVyOifPnoxnxZjprg52TtT6LoGyZ1fHptF5k
bE1iKiiNH4ZckLbj/EEkJbEFGgQ5B5WUuX/m7OPr20bGda4w/bjiuqtNr7Y3bJ2M2FOmMIWIuW7o
6TgmBlvRKoC5SI/cFbw55wQqJZLEss+LT+kOorPhMyC68d16O+GNDoQYtN8VU1UA2jZu8rZeGKzu
linJ5TchhG01J0+dCrAK3uWuZf2DXUQVD6DSVS6IFHlhWbZXWPyfb3bkUTDE4mLout9vO1ek4wNQ
OuuZAySPMNiIiKGZs2MJBzjzk2gZc1XseRAVEsfqP98vgY9aYOJYR5yHv5YX0EsqH2NaSKtrrYum
9jhHCH83wOkarSxl0TWStwIIHETBlYmwZDKdm7oFIsc9NmANSAjFo9REcvlwhfwW37Feu5CAmacL
QSRonEzpiSonRmWEHMAB2xGaU7898HVHoBFr/dE8urtp2GujIWsXYT0T6hB9M8hl8VGLldr347JJ
Urq4JqQvKLekE92s7Dz7bYnlnhOUjzRw8BlUcOygfMrP5aeICOeMpt+Rcd/k/7ST5Z0Wao+Xf0uA
CJSlNJAmt3ccb0y6cZhxMuI/1cn319x3pOrmKo+5HHg7sdVQXNCHW9nmcHcMovpZNgFgX0NAyoxF
6jMvRYESus5HscFPs4Xa3hTDXifeMFkH8dmHZ9fK3aximrYWqj94mou1J7TbflJzQzv43imIH3Cc
ZadKUncIe+bdWpxgMEWU2/6vjtG80oswMGOw/wu1H4oK5bVTiTaDzxyqRmwSxulyTNaePPj/yiXS
gXCyP4wd9udNZU6qgU/lyz0tR0A2EkLrQjw5gcLvuitGo2cQJtl7rTI0+dEnnebakcU1EpX1jAbp
HWlfNyd8Xat31PnoSXmuQTrqdATwDg6bDSxjtadbdvo+g65z1759nprmuh2yesv5DD1oUZ95ugmj
QDnaB+EmZzi0/8WBRanm8tAeK2hM+TQgXyHb2uY5tu+iqj21fYxOvwJcZUPnNOjTk2QlnccizdXR
gmv5JmYUELC8jC4soFQTOr8l98iBA3Ij0oG9jJkAVKVmbK6d3gXU4/Z8VzXTOq8g+Cm2YQ0ynglK
yZ8TeF4wKrRm0Q01i5vb/B7T/EE9M7t5MGEV3N4ITAnvmfQr9VCAZNbAmSo5f2o8/3JaKP4I7dPZ
CK+8shr0T+t6wRHB5lqiwOkVRGjDH3XlFltTJfrjOHWx6JCvxVb5bL15l7HDa5e+OfbSYgKAtcNP
1afMD3a+Ub2srUHdrIHt+ybL9v0OKYTk/lYy69fW4Wy7kv8z7CIuJBIomdi7730L8rTRtz4MFTWq
+q9+MED0c7fGEPkJtIjqDT1mzUt5jZG5SHPnETLCoDrH/8xdWbVijEXWDxfmhZ4Y9C+3ecaPqtQN
Qxwr+uq7MaEGuMDITYT5Q9MJ7fZx74Jsb40axWq75IJM4SAmKndOV0Kb2MED5fRIdKt5YkwvGEic
ex0sWcNhpM9l549+shDx5XSO7PKpy4fnfbKqiWH/oDTx4baRxRGnTbQ7A+gtzX+voZyI2vRy8DrQ
6on+Fji1ZBQeih7uc/n/7PSsAIiMA60RU7ej87oeTV6zCu17bXChHQdeKswjSBJ5p94B8U0slHzj
yLWbKnohxeYcTSbm3Mv7sRjYJhyRNvPyz6i5smfzqxlMG6KzLvlP855QZkmw+3GOOOe7hkleiftE
8mjr+SFxIxpZGe61te+PcauoyRPMf+0LnJDoYIKAKnJbgJ2zCOaWRmG+7FxrnJO+jJwpQ5YAf/Mw
Ao7KVnfEDzQXa+ibWOuoSjoEnNy6uvx9yOJuR7bsZTixanyrbXS/FGN8tv1fyTfAfZdDrtgbqD+P
nCP3gkxOJjoIht+tYwqWhzVkkbVtoj/JyGHo+N6qNWjdHHLRSwAU9j06J4Eov7IhFx711fWMQ9li
3dk91+tcCniWCYOYSr5tnUr/D/r9XiJ5nhASU7H+hIKelpxLstc73W8BKpZyccxXcmJC5SZnO5Is
LXfCJZYt8Olaj4R14gcka9R22bJNVwb+CyHp3XkxKP4fp1sfy1bPs9ijBrc4n77GhtDheuHRBvu8
EcEe7MEU69N3aOLTb+fBuyzKKD92+y8A8eAUWq1VFcf9cuuBuMAo2BhZnxtYeFdxmEl/PeFu6pOy
m9fn3/kaIkXUcDnkC5XzKgoadnahiym76pmG3PF1XoDyHmeAvNL86Rd3U1QqYWtCSs0e0RjodVx6
4rVndRGoaIihJu5HW42O2/IcfqtzVo5s7HPcIpsm6cYHJCTlIImzvmCvnFVhT4V9Pf5gu131OEiI
7r6G+sUNHzklhRjxh2yhELyqDDhKDioPVomnnLcLIAzjBaKRyKKLVt+CZDWO9DPBgKgYDMSkL7Y7
IOIUJ6y+FgxPpjCibyFFdmVUF6lXWUPIk19QxeqX5+Jb+VeL/TJLrf6ldDHmPGjBaboJVCxsWO5Q
zuiIj5Fv3pVgyZfKeO71K/7uWAkq6Gh1yI6zWYvT04MMPrfwVyz/iIPazZT2FUTQLgovWMKS8uge
jVayjBg8aQ8oVx9SqKQW7o3/U00a2QiOPByPNj5UNSeoY3ZVVNB5mpponOGLCW/CruMP6GPdC/p+
f7zd+P/Nlt7p75tJH2/T+U95vkMRS8L2pVdyhMR7LYCo/HtemPoTGubUrwmKV3DJsbsSo9ZxJT6r
uTkudgmLrT9RyMu7HzCr0W9J9DPjrVPPHBG15YKNSZnrnKTqpZeBcY9RfsF/mxnmc/viqXGkts4Q
5irP3rJ/VffHAzhLtup8QK0N165Su5dQV3R+oEG/lJQ4PKEFNDm0GADooTQA0lGKcyXnOLWjeGnl
KdUOewEcjrS1mTv+uzuy7hpDKUb8BiL0+LOdJUpwG/fd1FryZwxOkpOIaASQuW6hagoYFJJr4zw5
4rFK/HnonQR/L6mtL2uSxGv69K8NZ3tbe7V+dpggkAYceUDIi4966998uk+z+1w3bVqRBhKxcTpH
eiAwk4+aoIo62eebyStwlXlangkeYRF8xmIzhu/IOKKfJSYZ7rs5kVjP7w9lJPCQlqCWqr7tJhbn
CB3D0f8AHTem16/LT1d6CHdIdLx3h0+oidxcpXE5Yad2EowiK748BGosb/pxX7e+ZCnS5eK+jV8Y
TZXklbRbjMD3bBJF9OSII7lMfxX3CKW7cOSXPCR4iUN+gwLKO9kIr5Bf1SdZ7GHCpKZpwERrSCif
is5UR0wX6yAnqBv03Pa1KOaNa89nF2rsDGyFzc5RN/CJFYh+K0gI8IrcVg8WaDNkcQC7DFthacFN
2O+5AHbv0vFJ2bLb1Q2WICgH8JoyZ+Snswp0mh9enTnA++DKRMjcNfcSL8u6pK//6XRdyq8ZG+MS
B7+d2XU0oTFZhk3dZJCBRj0i76ELAbDxr1MiiRboQF267eAEdpdXIs8pkkHLimRkg/gX0gs5SlMg
+OjgRk0se2wtdKfOiQGrtV49dnfRhVz85t3VWpp6l7EIjXBjV3GaxRu5VVUZfl8ueoBnxPM6dJN3
W98FCVwXIXFAQkzUUa3Vr2axtH5vrTRvdMq8XIHYq4+It14L3qqzpgwbMmkX5nls+kUfeFv34hiZ
9jL2LTvrZUatqoeQPtKRJ8OsNM82g4N4n+ofxtxCJaGoTiioVX25ePoR6q7+t0awVkEB1N06JDLv
BWSJZppznUPardqtBEvoyr/y5E/Khr9WMITdCBIayzoiXWGGuq/0cHTY+vqIqMi0Sccp28sSXByk
W6jLlvs6gNgcffp59Czvt3R7RimwqIwgH0AkCjMXH9L3gktph57uiosuPjavYxWnO2ClKE9LFkfz
853NHmU6CNSLxQ0/N27uo3z/HCeTBBHkQQ62h5SAz1X9SIs7PDA94AyA2FSPkzjooa1ZesV58HGN
KIO2YdPCeWaCrOFY9Vt9k2EYCp7ewv+vCwbk+aZ8sC2UVCQBp8XeJBednR7WdquBVw8RfEzOSt4U
viNs+fIMtpVBArXYuuP5Zc7hGr6oNfBPS0kRAdn2dbTTt9qmxlZdFKPpKnKwjt+Bv3gQPLWIa5kh
r8scfx0s4MZdFXEPV6Z3RMLo7+rbnr5Lvw6ql6iyIQoi/Tb0glB25G9OxVv15GVpJpdwpyId6L2y
P+wEZPp+ERpTxKp5ehZw50s43I6kxn/dcMnKZHxAXVDh8lBXYaAoqz2ST40v+tkqrWeddfW0pXJG
jH/kRMDHzqwAMT69D2lc1O9QaVBkBayZV881SJhIu8iaLOYzx53uBqArEsXwg7O90zI3zDMLSN55
MgfI2g0u+ufu3/PyxNA0zM4qLYn5Ltrd49vhq6e85JPPeNG0w6nMYq02ZiwE9tisNz7/CQPDAzzf
hmaGmjIgFHHsCbR2Y6JqFGtWkc5h6xHRJJMdCfheqVlnpGAuzap8GSqMwrHS/+RYtMm8xbgTVII2
uq6GSy5v8bQ6cCzykHMh8eom/Pilu7I8tcJSyf115e1O9mTy5ntry9TnlkSXBVEMaALDi1PFnSoV
ZSOXHVANlP34Ob22pLTwcFhtghspaGB3/LKrte3DGKvNbkbbOhnryuOQ6tqhTmlzdwq/prQKEZf+
iSM78xQX0J+95f2YA9kuY4VFMpOHazw26Fpavkv7hNJrBXdzQxdiRirwQ7IbjzbSwnZkg1n/FROw
PHHb0h0mV+pZI6emYfiQWqSRUhOzj9FeRFe5GW/dE7mI7VdrjD8ZIpf69jc0qc+DtNdYK7r8csuq
A05wA67j9l2tKozuF4DRUqasZ1dpUZDxk5+ntdWZsDepi5E+DYvbhw9P3qoU1or0tM1+Ij9FBE0w
LG3Dukh/3w0xT39SlkVBZuj+3xr/uyB9UvKYkYlYy+fnG9JX/VD6P94Vhbw3iaJjUaXZMhzShoSo
et7w85v/KZj50pvwfNPeICUdv/31LPiwBKnH5yXrWql+iGkdDCD+KBDvrd5ycKEVV4ZThfbBrg0d
2ctAXi2dxiEgxvI0e3bXZezFAOKZMK8q91mvrXw8l0JFb1hQ674AZAd1847wvAlQqt5jzXuN2iFT
fn4bRn+jnVve5PZqnR8XBOFMrArzA3qRPRw/6JlSKPQY8qJtTc4AJ/NzZpu4ZmC6NxPSTyQYOyMn
pWSpIfRzz+4sxKXbxt1tW+UZMCQ4PxJmND4F0Q1ZHQC7YDJy80pcHM3Sek+oavsubJsFg79o3Ozz
EIOzgYzJ5lqrCiD4vvSgjBSfW1qmYk58rKf/LyCmtMFgPad+YGIwkBnOO741V2/kc0oCgoek1wbs
+WP6mVVQd7yXrogNmPaChK68N1Qw5VRVfNsp8G1DQv7djsXFwN9RE66XkQAcOUjjlvCPTJUXykl9
sVjTOy0IiYie/epyv29UR3aEw1Bin4CJNCpcunY50eDcqbFC7mr8ZAyDNuk2aHvhWzvGaO+5bZ4M
HmTHm9o+N3LNCbbPWrg8+5nP02dEwlNY/KXAUmzWTRzfjsLVTjmx1A9lmp1Pom3w4WFWS6nrSHbe
ikfZ+vW22lkdj/QWC/QA449nwCoakJE7RMy7GRg2i7AYQd+jMA7LB1Vd47mFLh1elRf6StYrtgAA
gsHp997m2Eu3w8cOvNiHS04fm95QZL87BdtbcyXiI2TgAgoT/kTxwHBFyvEE+vOmlrCBfUh0PowB
SMavUDaiXC3RUlI9xZKH/ZT3cApVW8ow8veZ+f6vTGxwa7Sxb5bhsbj9MM37Jrfk0DbeDYM6ZV+e
b0VFZyxnnmkY+GTeT9GcEFel0LJsdejnYBWVwwjrR0DpVjZRxzf6NtYQejy7o+30ji3g34dLc48L
npqAbUViDMwUoWnA88qqLPw2252S3wenLMtLqL3IvwVf7ZSyOlHZDY/+EuV8TKzSy3vDdGHtzv6k
3IbjoheHIjA+eNp83Pr+/O5/+ttc4l9OASilK09vjpOcdvRImRYrVNkUWaHtgMcoETzjLUdtmWo2
l69tcntkKIY1YofkB+INEQnUIAgna77mIQbjTaVGILGf2Y2n1entkNj+V5BcAlFbVTVCurSGl/YA
13CtC9RhmjKcUJw05nBnmIDfLsji3NamhmTWE+9jdyAlTbO/hxGSgVO5rR63UXy6OuWO7ANhSHOd
vc1Dxhn9aABoCqhFhbvt23htZwT15cS33aZ2/YxAphnGkCEEJ2dCdsCaIAcv2hau4UFfVD1mW3Cp
k84qABb2wl0Dh7sMV2iRL2oq04//tFcVdiLac13mTnKMk4/Cr03C1xpiKKIHqEYq9wxOzQXoG6T3
G99QCqGwxgezazDOTgxMxK1QoEpj6xaz7DD7SufA/md4YiWtX5gdXnUooUMJ2l5e6iOLZrbWlzo0
A2MjRMu54JPRpp5nO6XTJwZP4W3r1uA1Id92uM2xNNVf212/RRKDbPb1wJWua9LOf0O1LNSF9mUG
AN5Y8d9/hS+oJttELjt7zCXifiX1W+mH4nZNq371WD4NVLdXu78tlrARNIh/8xx1noiRClyReIfO
XFwB6lxJuzQDgiC+dMhDGGKRu5cITZR+W5xQhzCDjfZSEANuVxTd7GWucQdRjJBlIX3EgTXo6yq+
l0jlpsfRD98nR9/2mltJk79AeijSq9yWI9rJvFSHFIdvXIF+ixjS7kwnZsL3mszEkJ9Z5tkooAA/
wanYh8RmvwumI8KvlpXfWqvnXrGnGTmLFwfcAflxw5qBeWw7GG9I8rPQKE7dQSDpEARd2YXpkNvy
JCPD23mx+MV9suOnRdX+Jrc7azzpvo05PYmnUBOzqFjF8iE/chckaDnu662JYqngsI4G5JThWYWb
xrzMFzynXOolm4j3pDlkENIRLLMDNuE6M3GttDfqwMuwmzDIXo6fxO+rFu50H9tfnU8PBHJ8WTNQ
rZd825nyrf9e8SbXgTZikcsSjtULmiIgw1pBGwgZocECd1LZCDqQMrbUFiYFQwWKE5rpzIQLc/2X
woQLqLRfCaeSgfBM3BdywxPAA13jYDDpXNPUr3uSWb6BK3LgpNRNX7caXP1vevNoEhpix1xv/g92
0/swTjjuMkiZMWxfmg843mk9tTk8carjhVaKuRbPNP5S9b7/7L9zG6gR7cvUTeSi9vLHYdd6kkgC
Z9LeI2QL8xI1POU6tNB85WOogztRFa+0HN8uzZ2llUFea1vuctszlDZwSkFXjeY9ujaqsy4/f5Vi
BpipMivu2EFnauVE8UDu5ql1PA7mWFOxoloVFYnexPG5Z7YYaw4panOLPYTOegBWqb3/+82QcMbw
LX1hE6Y184boSi+/V0U8C4h8t1QKbLxzoS0/FcHqQlupY1G4PuaUj4sskFecnJBAhbHxXaxwFfSq
lHiAfMyrK62ATNzKkFPaRzR9L/WzQjuDZCwdyp9MleT8/5CnPzMjKB63JhBJ/FZxZ3o1ItNY/epJ
JMpgJCMyUVJNGdjc16ErxSPX3JU1ZJov/2MdduQgSPkEjSUatI40eUX21IT6rtsGZA1oc3o4Wt+1
8LaiPqEzCvvqbLf6D4rR7QAqg2lpCRu/ztszxA8UBBCupo3Io0ATDTF/xF8qKBVW0eTYJyl0GEs5
JIg5QAurnnuXIPs/WgNy6jkist/pcBkZg8WbifHnDbzQ4GpomG274daKPefQiE5BvQGYYBdvYCls
hRzN8I9D3SDDtvBQ+LDGK40CoBneQjFVLtdz2G6Gk/bJblgVpFKkDQUJP1p20BIKbcpUYXw0puq+
N5T1DVhB0P1/n9Rmj0KskdFkh9Kk0GgJRb5S4UlHI+lJ3zCnm5JUG8El0xDo5Fc50cMclkajoV7L
bMqMeV0fXZ/hDfZcDPP7tlXW1HtHH+qWGHl80Vm5CRJN14lWmjRDrVgxls/6s6lADd309rxz4tDY
Si0CIvBsW422sn9jEpu9a//onkvjgZC5e4ReoV7EDcdvr1nW+8Efztbzgt+dVHHXxrM+wUiRx6cv
O0W0tVcTITaOg2KoaV/EFBmve7QcqGgFq7H3RjK5Uqa9er43U5SP39dxGgqXLLboda9bz/fYBYaR
6pzBYjOv/1dA6sLmgshx+vFtyFoMhzbUoocprDl/hc2tHYeZDfDHo4AK8ZE/xJjvkbEOdWwdkGv4
5C4VKSfcQcBfyrcXDewIMcjZ8xKrBa3uQZXL1pQLIwqlv6t1M9FHkEZ0UCXvig7NhBcslkmUQRqw
S5fgmr+VuJbwOYj1KcszU5Wfq5d9tpRDwRPpvh7FtJN81X1ChwwtsNZYV8AQqT2zOlPXCRO+1XNR
dCDEvDozPv+LNjRjepUI7wi5uq2i+xgnospJ6X8gj1SoQlMZOJ0aPay6eTn2/TT28yxRREvPKIat
WbEoBpiGzHoiSXeDPI6zWX/ihHUETiPqTdh49ii6nQECQkcJp7KirsPgiBxnzgyzmFJxbVRWqDnb
UpQyjTt0M2a9vxOVfadHNtQo1wVBKpptdjI5Fo+nj7eU1wF0fz72CugXs/HXzOU4dV60bu6M4DFW
fC49LfPyFOddAj0jZtZt9u1F2/LN9Cge+DCpeCJ/BI4fgUUc0TX0RmVLUP8eXckDL3mc+cDvZg0Z
JTmfyaqBU9ryJxQloSMhX7Fb9hprzKSV34xmby2rzrFIBkvI1YRiaInobs2UVRG+69UzwJSBK5iE
q9DR4MI569KvXYkxBKQ/VBo8plA6/NakSp60PKBuizqtx7t6GfIjzhejAW5IBCJ7NvTVSumpdyj8
o7RVTzDuE4HLNx6AmzFrTAF3ha0BoYF2Y93Joxt1DltNxjbERippvcvGs5KtOhO95mhaPD+uYHWB
KLXMLeKoYvWLmuf2zEshkXZ/auEBUmhYJSQpIGyu3Gah1DWsfno+F4BZ1QJ+oqzFCnTrtT4+Tm5K
ec5aNgcIPUxsrGJ4+pE97Y68nSCP0rdkK0LL4WM82i4Qx3+IkQNFMQIOh5KvSqY3doIWORmOZ+1R
j9kf8lG7ADFGiH3QJbrOBAnFZwu0Cs87G1GLScsosfpHmRFq0cLrbmwu1lCumCSQq9mTna57/ZQf
QM1iUbdqNozeMSGz+EN4oYorcVIKeZwEApT9Tp/BrZtm0BK+qD15bnugrug9ghNloRlHTZ4fexJy
Be86eY+U/4mVsDcwIBVJN8I3bgtt5lkzIk89jBYPGvdWvgvGMf0eOd6ROhadbfyEPlEO+rp4sxOb
PGuK2LLTdP/VIfEdviBW7SEVdXRuY4Y0SV4FcS+iFVlLp5BB6iZty6s3s8BqDNp+nx/6IaWP9m8r
goqM0DqjhJCzv/6Xlq8aexOu/GQkdVlKmMVvlUKqefk6DIXAZPzvSb7nWYbOIAF15wf54hGQgQ1Y
TxkRHABRIzXRty69IVAkFBYX6AeX0F7PcB8ADrzV7hV0je8o+FGZc/qIK0PxDcRwuvtZeZXGCaW5
1J3RmhDeuxj8IldndOdFsJmoUjDurZzZv4Z6f0ymEccevbcyK4OMfM3RL7f8AJu2wxU8LujTVca2
CXvrO+dx6ixLROyTn0ujsjJeQ7RjOw7hrKAl2XiGDZARKSTW9dZVXBCOjsJO9nWHzzQyVjv5ioa9
n6OSo3OabIcbCPW/ZOP3rs6vU0ljzzg5l9v8Ko6RpjHJyHnAzee/fJbFiBth0BZXPf/1jpg5py9V
Y9DOBK2vN2m6gCCvCv3xc4DiKlO7S9W9GexgF9m+EzKuKQYjWQqEtiFEKCcFmC/e0UkTLDKCInm2
z+crM9xm+GGWbWIF5pAmHe4WDLbgYAW5oEvumbtnl11IITWoMcM8/43oojYl/vTwqcZSlt70w0Q1
3AUkp0Qx36CUUO/acl8k7qAH7/khwNgkkoxPbpP7YJBv8vHLBWX55AHPtbCPeq6K5XH7Czmf5EPb
bTHC/khOl+mpDaG7CSYzLMWRNP/cAqzj3q85jFIHd9SzUD/q45dBmsQ8bzbbUjYKAVal8gpZuXZZ
7mjUOiyv+4NhjdK5fxkVB1Ve7gtPnKqHc6h6zW0UvHwSSFKjSN6XzvQwGHmdHZAtu/aAWGsWJUgl
O8F4pJQceKNk/ASWKTmFtq2ORvK3EsYWpGElQ1pUZbDrHCYJhiKkUK7ARScN1/M3Ia+ICSKa7wKJ
Cw0SV9pCpM31Te7n86R+8YO+JVPB4THxp/EkNi5qZZDQS8v+/ajYqZLM2Y7U1GagBw9WYvU1YEsI
YXlLWSxhAf/B2c4Rmk2IiIIBgMAnHJIbBB9dlJEqw++v9amrMZKx94Bve/lUU1zqp2oCXqGdOB6E
8FtuJwIWsbrTCGoCBqpRCDsRtdLfoSfN4Th1MBLhkK0Hq4uDSWpXDY8GoK2IvETJOGtQkRYHfiUJ
c0LofKLEphVzu1266jW+NixSVWGRAbfwzOJfv/dNBbFP7DIG8NKUZs57XFKIAS/7ALMAwJ6QA2lZ
1Rle/WlHR1IlzKILTx3bVkkawP8lKxiM/w74cGgDDWM3H1PX03Y+4m5joavVKnMj9YS7dABdevtv
BLOZfW6XvaMIFSpAIhO4dJb/DSofuw/5eQ1gAvIixeyF6Fk2WiiXk/yswiAgwCUHHHdq/Z5294vV
WHPxIje/9XtBy9w50Qfy5urquKU7YnMhMuqpupC51gZzmBlvskWZ2nKljl9TGC/16WDtdSCZam2k
JnMMYMZp3ufiwCqJ6cb4kt/GysFFcfqi/0Hd2O/BJrU63iI0kGIT7kw/Vbgp14Co8Nmp7LX6t713
E5+3QQ5s8+5tr2xnTlpGr/nK1iygCJE50VreWS+IPmTkDvZc1a/JgxqMLCrbfZl4lNBMuGSWuAwD
crYhaC2FYbQnsxtV1G839R64HWd30/yA/EDpZ9yd5lnykwia1pwoOQz5LvuOIVKO7AgsHvOyQC9v
uc2DhUM1/48mDMHK6F/ZfzuNysX92Gi4FfDZtJ96sfnxemPQR95V0CucOS99ItDoA59+VCRQXcq2
TU12GTcyKSjSH/k5HcAZLhQ+usHdJ9+hcIbvbJKn/+/N38EkMVRg4zi7H7OJ8Wr/WOyD46zl/sZa
pEO+uHSQ+e8suOUNQ7TbtzojozHBhJdwASsqFIwqmaXj/Y2Yi5kPKJ85QuJGBLn69H1sqJ3HnyJO
9f5xwlZ9XEjshwnBF2kpOodrX9RP2WZ9G2Q+5AZSfvCmTXI4xabxxmXozRdMnLfIJfcUf2oIngYk
6WYiX4U6c6NCFo8Bn/ZY7YdS3kRQ7pxl1/3kgDGIj98eBfsywmioLp+KSXBYMVlgdCEhhapY4aCF
IjGwpZ6UaD17CItiVXuKkoeJ5UVSjige5p6vVv62MAEJd++hAFLFp7Bqia+jbNbZTUBmmyVoBnAK
ZU/OqVn78mqzcfw0YBRieVnIlYwMN9gPxL0TcVdLT8lbRE0LLFI3nqZSafEs0q3dJr6kI/yryUZM
UFRfrNh3JlH3fusyHIngrQ/q5yIoxs/Gbdfk7OWFL0jOsBP0NPKDNTLChD4J6UKhiUJTagqN271k
fPPFfiNgHoP4iPCtKQqIyKwInitrDdoX/xeqYueY5a1Wo5cvaSfacvnVlen68qyZsP7/bB9oVqSQ
jJPbtB+rHLEehAQxPnXAYQmAykeWvBLDVFDu5fcSz9+18H75i+LFTCjJAO2ZXIIgr7U0SOKmMams
l2zjiJOgbx+bX7VJgIbazJNqSu1FPe4qG+XeA/erAphksvvifnswFJgJE4Vic/rYjCTnnS5xbhMM
ZsNFy/gSRXWztXzz5vsfhp66h3rtRo90mruy/eqTIWCL6HzC7r1/wDvGEwavtSQEQLuLn8TRkdCg
a2G1SEVhSnf+Rb1Uh2XI4iJspjB/DbmoYYFU3aE5rMhxqXLNdZ6rwGQ3Msk3c7WiqgKnrZyRcotX
qOW0tkFPr55zb66NWtOvpFOzv1Pp95uHhMD3Qd69uuF0Nf9jS6ADaMKEqvp9IiinglWq7cZncP+e
WwgkPQ4MvAAaI5/n2skQDnouGbkBbjfNAnZgdHbLP2C4lg43acI6W/JQK+Dh53q9UKlP1y2AkF1b
NvlnVf66K05FEWaY5SZ1gWJChaUzQVH39BiiGmCFbBLjNzl8+XsJukK/zcTNuy/cWvNRexrTosLf
6zOYUbYBFPBn9h9j+tKUT8BL42MfmLLlEYNTqCwrW4jtqDzLzamv8akgG3Fu9Q6mBWE0uMNZhDcp
ADpbvB48yVN4izDXir2fVtD2H6lf1LR5uTHMQbH7DUyC+NNo/UPQMfjzX3NDDvnDvcT2wbx19eDc
IQUM+ubhdMGHq98ev6PLi1aHlUI7efeqsqEzvffc02jlplN6mC+lXJLqTJ4ZEc0w/g/zt1g726bD
Vguj4NyjIB+vIfxf1RZkJn/kcglATkT+2SvApUvdujt0tPm3z5Gn3VwO2r4W3DJvB/0yIuM5UmYB
RNBSiOOlZTIFoWfI4FwR97PxenVBudrKSKb/WubvJoC+GUcunJSrbGoRi7h1uBm31HeVwUvjn1j+
ZELLtehXUTSroMGBduXn2pwX1iA2dXofJNEzzDcXZ+8D8pFfntms9Z/Y2hglo0jDN2OD/R9bJrT5
DIDMF618WhXReVcWj0KQAYwg23LSMOL/XtJyBM/l0J5gnX1roQPY+kYkZCrEkp64x+cHF2DEWEGG
efr6FXOGo3ohyTARm2WNvlNX5yejvpE1HaX+k/OLa9TDAJCbREE5BDvkBLzFGi7QvuPu/aFQYLB0
dAlJF3m9NMN0eK3Vhph6ySOybnsF/w5lcQxljAe2NBwYBGAP5itnkyDHVdn59z9PcKWD5Yi0tve/
8VF985vN6JkXhxCE50ZhKJ/8fGPH3+ZzHeDhKEyrDOYjRGE6uNs6hJug80Jcfoo0YJGjghgwhZWf
Qzv5yLvfpi2qhUh8MGsLt99Vvp26N9RKPXO/j/RWnAGPZqqyNLNjmkVIjVSEvsoofZflN1CFCoTU
U58LQI2e/fEQDrytGhM0m0wHVs/L6WYdhb88FbzAx4P0ATNX5yrTWCWOcVB2Cw1pOtyhbmst03MT
dp0I1oT4Zq6yHPzin2bLDOnB/vVJsG5OahtKj03sA6AqylJ2J+n8yPa9y7qlSvxMz796UFrqE4ZA
qNkXmjT+RVTSZPvmXsz0HmMoYSZWE1mNtLTWJRInLmNNUgjqvlUO2H+NUP8IZSOi7K9dtaSXTmTA
gtY/ZtyqhvQtA11P+IrNDewrnWyocRHWdpzqXU57wTy+iW07qI247AnKyiGKACrC/Jk9apOmkEo6
FCthL7UZB60G7HpLS9SNjEkuvJDBkm3xV4v52CGFfr7ouldApAHipMZtp243K29ZbxWOe0DJUOQ/
hFha99kNCi4dfdtCnwzETTSZnCZAcCNHxO6QYB4Esc1e2O2ZAKkkgk8+RLvpd/RDSeLFF+fSBer/
nRr7ovTA3WBbNz0D7ObV1q1s4hEAnxnpM3zO9qWS4xaFCMML2dedWJ47zCBICSi2ues8iebQ3BfN
bZcsW6CjWSXhY7QQIYpyapLdsHSOcy1htdVGo0I+ZCEP3WfGxCC8riRbJDCspkR8mTklSV0dNCTv
AWO97npEyZYrh63tA04Jki53dN2LR6V15PqqGu+qssydLIUcFf0fWGf1ZQ0hxDOwFfxLmsJIFTVO
ivo+MJpgQNhFXsPH1XbClWjlhCGrbBF6+Z5VjGbm4beOr0whtp9wyJnYe7Loui/NCtTo24E5jYuT
frk5IwcWc4FeGH5lM8Uezs/2jeXE/ymH3k/AzyrieKHarIQvAoVLbMBALORNUBLOu1b9uJ+7Eogl
XxZltqzB6vZjYekkQYLAiaLYUotbTPa2Dut0GCri10ar/Jk2xsRceuQBssIlJ2wkePzzZ/jHhBf3
ilcVR6tbPgNtbQJUKe8snc2qyJ277/kKkF4ziYykGcsshRGj6ZkftqYFT53ORGsmZ9GOdlr3KmUS
eY08yEsXnjl6Ko5HyOkVQDo0X9c4GmZnggrE1TVVtD6vaXWAO6dxs6DM9+NXk7rrua28+jU23wHs
TtupoeZCT1ETddHlP94lCZQjfGmy5FzvCxo6i8pQFJf6YyXyKuO7DX8EQi3UlaIiz0A1NQwovibd
KHiV62XKxqr7DHdk1dYK89aM8ecTsPNIEBorm8wWQS1E90YAfNCdfKKr9twpV26VDGrfj1gHynJZ
JZQm4/J9f4Nplw3DrJX61mAOOtw/AUc3cb3HCQy4xvCiTe8/uFohkgA6bpLnuQivfiDhigEzi/bS
v4fUZw9DprLWMMnR58/RoepenIS14MbvLuQRMCMVJMaKVTMQJm4//swH7zjBmUYEH5tLL8Z20QWh
JpY0Hr7uf91IZDktkxyIBEgLpR5DD5m3xwU+3ih9kZoheSxntuM8yvpU0/EE7zudS1SdOh+Uf27H
o6zv3hkKZqHrZ9YLvozgibebRJI3Po/Ui9CN8zPlr8nXv4fSu3Z1GNQpBVfMR73mcdjft0B1e3ub
eXNBTYNLVnFXSn1C6tklw0ybRpGy4hwlzTAofjPpndOkmHbhpOSBBHgR9mKNNBkjAUe/3git+F0u
h4nAUzCUjF0CDiscr7w5JqtiLnvucu7I3ufOr9bIs9Ya5cg+1Uijika6lyGBqWL6zyX4+DAv43go
y04Blxf2XTwN/rIc+prN8udpivyfLQJ/hfLzi8rfYaw+UrZ6FTAh/5DbKt1wdoSFbgkzXyH0iOj0
0rwKvWayPGmB2fb9XKhwGezU0rkQxqyDTJu6vM8gXejmp4ISx2X8jlCTL/36ckYsqnH1hKLTFYPR
iTV4e6c31MAScM7LzSObPj0D5Mqe6SibHa5eZ6/xJbUC+/9OPzgQ9mssgf+j78IoQ4ZqoBwVf2v8
ej9t7n2QtvFOPicLbI/Gm+QVvOGxcz5ZOG3rGJxn7pVM7TNCM/i3nwNpS7IVa/OnF+tmKEEXyA7C
JW3MluXB/Lpow19VLFsoro4uXfJ45U1YLbSUfgXifPG4aviX83x5FWnW9vTRIQ/AVIWnrR5UficE
43FuugcTUOXU/npeYjoOUShlQLTFhDVm4IQdOfdb6/FtiYvB7Z6Ez/UiAzNuInvzOjaPF50NGG1H
9o5f6LHG677UqTzMg0x/xESStJ7Ke8S1pyCVcn0GoSL2Eg6o8IGYAG44v4fvCa/lVVIsGo2CTw6p
yZPBTMW1/VaHPzBhK175vI/3kzbT4/Q3cRiAgTiFUY2020OjfsjKHP1C/L6TxXWSWMqIsUX78Ow7
WZDukpM0cl0RYoI79ai1+rFwRKIFehF09GQiz699tnjiOd/TZejjti/hO6wFBsyE1HMbvZEod9+k
eRuwp1XUhKLfaYxgNagdqhCUelulZhqkV6BfiPphuMEBU+fd2XCzGc4bNcrSYQXV94xJQT3Yq4Bf
z3QNQQ3Gh9cZ9MAtbSw7xox01awqCU8yilHWSkprw+tFo7PmiIVYPfKc3H/sw9vsjh+wfw1sog68
LPBZJCfp4ltkYjtBi/ru+mYWpXpWqiWThPgGy1aPMZ/ycI0HvE5ZiOCq5SkGnY2lYcSS0LUzooMC
7EgdrFFoYosncU9bJXOXYbpaQlscdZ8DC1DxlOp5BL9297pzqhUY+Tc+7I6aF1LdFhVGyftU7ZAN
6YXNWk0IrByV1RyeZpSTse1DeEHOOKI5knWZqC04TgoEXqQEcEEkY0tRO2i5R9wVstCxr6fFrVKY
DSX5q94N/6kb515YOGfW6h3NRJnsNEYXJpA8+pvhN/NaRtvCPtjrnJyAlZoEQOst/ZqTcURT69RW
yiyLW0/IcB+p1+3bbjymkfF94aOt9WTdZJDmu67Fr2bAxMwtPewVKQk1Fq4YCTe4Kh8idw3L/ius
6vfqIoOFAnq3vngsUQhr9oeawyary4UuvXWiiFYTeU0JH4xDb3d9G9dUdEB4iodfnS5lSsVu2wea
WUAmZJkexHcNA6f/MhKxVCoSMo1czCMeLl3Lz3Jz8umC8JrQ/sA09pyh5uRBcVm6vbhrPRdNmgpt
prZjhkeHDYmfQ4UOoXGepZ2HyfgFjPSxFy1A1yZpBHgzTy7OwxqA4MtrhQkB3lHXan1lmL73VlwG
H40+lRgB1VYhl4xInsIBMqZYbloroHotEMxgVeojTe3p74gvdZgJNpEWja0j6/xiruR3U1NlLXc4
vcjXSiMJ4flFeFBvtA9UeaKU72KA/x3Z/OPBNJQ8/eY+L0PhLy0mnryqO8skwpMyDAOq8qh6dEQC
xcqr1Xq2HSm+g/Ft6myTNxTTUOmQdHULV2nMdLB1ZDGrS+nLGoFAJOV7yL30t6+KZJTFPqJmCxFx
cHN4QYnM4Yt3BEbw9FpUrZdyrzFoXzuZmKNys24+xGd3/HNxpOTpePV/7YD52NUCzBqu3hVZLMPM
4MFNHJ5kziQ26XhqRhBUpv8OVaOatCSMh552qTBjGqEu+4neEdnVabZyJRnaHXt8R6ziSDNnURxz
EtsMl583aLm1RFXzuBOlz5f9oMsW15e9x2WK08YLgxa2cJchj4ykldeuvo4m47eb0vS0V6TeUL+j
w4FKcJ43vtP2WoLxfyGzozHUuPW4RA+ytOHbCtbp1m0aY+xpBn98OpzTLz/LWmidNhs7mXfbXPNq
/ZaIUiEN79qpEkr9blezA6MR0XwTKJgTZMmCHv45uyB9lYJ+BAly4tBePETqtjiS4zhlRfhxAIyD
wIquzNcAMv+U6v1dFUzcx2tfJ+ZFWOvjyDTYH+Glrqb4UVrmuxcuGDEBRaNPXO4eaqYno10ogsOM
2bCmpad05i6vfCmVo4Mv33UPdDNWBckNSCUIBMzRAwWjWFUglI2d/p7chK3RFbwyV+XS8d54/xQh
xPLXAUl0ITRBd7rhnmQT0fTHHHt83FCto/KZRX3WOWXFh6Y2Z6Y247mZ6ye9ONT1w6915IhXk9eG
VZOIs/WJLyz3fqNK7ZuwKuUF7FQdXL5eFPfTVM4f+x1X5QeEmlPr9ReB0dTsrlc5kdhHBVvbGahj
iaf53SgmU/u0cQ3FKjCF2Rg1JDXQbjI1muuSybhg7OBaL38w4irmMqNs6EB286590tcuCwqRvGAT
WJ9UadROXG2X7LCnagm2MBWGLXSLQLns6CD+VZXoL1dgkaFOKDvgLbrrJKoUDQTHMVz8V1lkbsR3
BNRYuIBtCbGTnDguJr9W0Fsx3ua/4Pa14vWTHccmRX8tSaaGaoZXbU/bAISjkv2n8jEmkOxa0I4c
XQgS2h5mfnTaFDpdFPeH7A32h5HG503ulisdgwwQw9Fsy20atc2NIMhStOP090Dj+xMC+qkxftMS
yRQ3ZfbdhwZFrAmx7kUY7ma1C8wA3FRfOklHsgqLEAY3/sXIV+3eesFdJjkpEilrAQ9sDaDhejkx
/+geoX3z+loTM7TCnAkj0o9Tzl9QLDqVxRC2TWZ6QSK/X6teX9csVD2kyERdoB7Xly3F0Ydszjgg
yguRxY9GyQCxiATPRuO8KplFR+KgsvTS9KMmnjlj9+YI/RCmcy+QP2AQRjkWcV8YqIux84DhV9jV
k6yasaEpcA2/vVJeE0DQpxTcSeEefwZwOTsifKi2xxqv1Rcj9JlzOrHH6SDjatlaTs/aPr7RAryN
u+zd68h9UB4ia4VlNPSor165e8wSwtbbozbE1cEAriwmtj11itj6Jyh86EZAIR0nGHcyJFLlO7uW
bOQhvWshZptWmoHJFya4vGafX95Pr0jbBbasGkNU0OsHd8M2EuunGrrmTsRe/lvnFckmwWHMFdMF
DTkiGvjxnXmdIbV6zl8ewPP3DoIFrcMwV9kG0BHaZwLSX1z+RjFxWM5EsUkfdhpplkFtZuRYzh8Z
zHGceknzofAxi8YEk6rb5qbwU3fd6PAu69oq6Sj47/ExcuzzABrgzOLOUgaFM0n0DUDygz29vE59
+9HAl7IeHEmhW0bCY1R0WBfO8hp49eeFf0neoYSdo/uTFwA5WipyurTS87vqSV/4DArmKd5531nq
D0dvgm4IyFiAzsPhkYM5JpmbK3dNZHes/pchEY/eHpkbWlM1VOJXvbxaBMkRXTv8GiApeXTjFNmD
/2JHfjukhQlDzSG4NGuc8snmgNCblEuLerCNrXXhPFMCNgHayOPqjxCAFTXesAWCQgrf2AwJk5C4
KUNoSZF6MMYyg2d4ABt8RV7pIEjIGIVxx+kRBjJgU/wGYFOZPB3FgWZoR4Q43ulBi8ijAQukO1qC
Rju6FGjNMKVegoQYd5VLUl+VRKA1RsiTbUcr/UaTg+ErN6N/arK1F9TspjdiXIY8sh2kGh1Wd0ZD
Tw4IFvxp3Z9dI3pt1eYSVHZcwZN2e89ZOnRVXI/qsaLeaVWeU0ydUEy/ALgKhhllH8Bk+DG3x1o7
NCEMQtb9XWUOqk6usYaDh8cE+gu6+ITZlzonRKJDSmJk+4kEd4TL3JvbOggwpcSlB6K9MSYIkPQL
BMrk1Q+VR/Wi9HVVyatUueD+2pWl2g4UiAxEsUhKKHwlb/5YhQEg+WEjEZhiVM7eYIxIXZ6pf2J1
p9gd+HNTGxv4Jsl8yFh3j4h5PR1XzUOFEtVb+1OjsQJ5tk83C/pCiFNKDI0tqOaxJP1x6sFslZsd
YTY93PXiqsBsn+hmydIYqXD7VN0ljB1QFFpfT+kot4YHv+pmYohS+M3Z3ovuEVZnT1ShmZOoAbJ+
/afDhKOHr6uK/07iyY2j/DdR0dLbI1qb2bzk/vsV6+lR5T7/hAE9WH6Ghs8318kOlyu6MGDAFD+J
zxg1A9nnjJYw+xeWKpwvO4LYi8STQolfo9qc7ILJklZG+ewqCmkV97DcrPMJGlnFqEKjJUCgCZdW
sqzH2CvO+CcgcmaJhWBQCAxeL47QZJRaY+sdzYYT8+qoHQQL7MWgrPXNMmfbPMy+MiX1/v2DFmR6
3zxY8EuyByoiV9HcMiP/YNFuw/Uzadp2iQaAURkVnC7l4T4oJddBuvCLANBpcMI2biQxu3dP/ns7
pi7VEY9hvF3zQ0Wd1SuVXjTATm9BA+oGMDhkxBn6yoncs7Eq32xSeRJF1Fey2ir+9OJCqSbtuqxu
+8WAX3QB3uX3Xqs3brwiOpOGOrZcvwp8Vr/+YVLo+Uwl/AMszH+rrfgPL20+/YVo1jDKFEzanVdO
JaGOYnYeMoHhtV7xqUBL9JN3bpUvh0O69WItRfErDrHK7CbKc6l37Tz20e4R/BtzJhsKxcj1k9CO
m2a5q+Tu/Gjd7p6AgkRWsC4PP19TK/H9EBW3UkgmWB0G7c7Cx526RAgLIQ6sAILSIBU8Bw2sVBfD
FHNIKxcQEVT3BQ8Hu728NvXd1U0QoQm1jqBbG0yPajQ0QWxXO4WOUHhK18Y8Q2TFgWNFUj7swnOM
VHukBU62B35ztUKZAXSmfPQFkGVR+ia0f88JgOH7D6YcOYC4QL+sJqmnYG39P3jYW+BKKyUjy6dA
McOi7YiNVPNVjRmpgPUWZFb940F6tNSmwxJ72S6vnJTQRK9RERwXI5eqk8XYNYQCr9vo2YyWLKTX
FD/YiJUpdDsLxkQai74kMUV0rVIoSNsOQlJT7jehdMIU6+I0W9tUoUTG4+g8xmZulZrLDPpK9zsH
wdhvAZf17NEzCRF3rSV6wrSKH8NWvU3tvnYg4LgfCmcpGBIrvJvFwPtfS5JxZHnNXfD53c65Pc5L
m8PECdPBSmPkjn5+NVfOu1kG3oIr57wtbbKA7EP2FMOj7H/BNRQNQPmd7UUsBCJD0bki7QbrbKlS
hdvU1JGL/hgyX4iCj5m/0w2HZ3Z9w3FJsfgj7v7oJoyUwaB+Ib5h1M2alTCEfBop7x+B4Ljm+N7M
obIqRgMYRm+7QICvnZXMPAeJlZKaIrqmJBvTRRJ8VuR+1uKXgkqcPDItAfIXWOkqh6Li4xUnZk/S
85xGOEJWGUXkkBic5kfwrfo55CKjaqwR/jCxixXXhOT3KsDBCI1vA7dxKgrcnvTkF6+AwzM/2/4u
PqGd1hxcAYmlwPVPVgVBeiJP5O/j1Txdk7xi7RCSAzI/hwnbTQL3a2EuizE5f/ice+3RXrQHquIl
8SsgIfWOSBNzdi2UY5meEdhUXcPhEdOF4ruAe4FR3mRXPwm1XDjmTCCRioYHD+KxGbZ983RMo6Ll
o8fSp5nZs5k+Lcu2e2ZLwspYR4HtaGZ6RN+wjotFnMS01RHyns4kFlCaqSPYGiTSi4VLHAxbP3Wx
HOCp1h3P9Jd37xbfmq6bNd+yMJD65LLsFjsM2U5dJcRlvp6pSyHmu1pmLb6Nlzjj8zPw2KUP96oC
KteyZZX78VcKSq77AfOcP6HzR8rqU0BN61AYf8+bQO4P/1aeQ33v0QSwUX6R9KiOKDnI6yE3wdGv
kQLyQqs6EtLAmy+7bPlpNe04yBAhDx3GLMWSY/9O4tIkx9DLQBlQ89KcxiuPaNqeVoYQRZLnfuCs
2FucM0IQLfnN5Hr4UyeY180iWYEibNThm2YOcTOlgXzszGjoeXkMR6fjtZpIm7CYXN9PYrtVvtBO
KCyBj2svHyUDVxKah7Bv7lU7/8Q0CRdQZbrUTbO6Iu2GVemefsAwQsW9N+CiEz6zAbWO4FbQMlEM
ldKIhLAkYYEqzzp6kKKae/xmpWzl9AQlUpWwu7TIFc6/7XhfSmXcggHWfROSZzf+mp4FiKXXwZH/
C8hwvP5ManKvWwrOM6RAwoHMsj6MlBI53E2Lrr6/5i6NceP7XMEm9vPHAAvzrv+iSNJ2i11Sr4nC
lTAPbLgWgIcefBVz2ZmyA7x9fwsGGRGMlArk6kgDgPJ3JCTy0S0suxP6NZnsBfyrvFWHhZVQjEAs
2G3edS4p7qVQ2VYhhva9lkF912OWbRAp2J6pOf/UtoBFI2Un9uIzhX3E1Y6EKSth5Udyqmg6N9QX
yw0bdm6FyvCRdW0T4gpIGcxINpZwCKzm5/XNq2DIKZLs7pJz8JiasUyQTKLPe22X2e9q8iHal1S9
fjyx5+a6l4gZPMHpZpHA02UzcNUOisi7IPlBnZ+VwRChBanvw1lkQcKv6C/Pkd26ib4S6kqvXArp
Pbax1df5ZkhOWDKHfTRssrdwAGCpbA/ihWFKv0JB+cSBYgntgYVORDP4n7xK2/N3fVq59dAs+Dzp
KSZMxsgBGoWocozkA79jOZd/Z67OYAWFyIDzQZIKNAVda/x/p29ye/2tUHWzDXNc2WIYfX+7SDWW
A8ZOr0ndbn7Zf/P2xp9l0pweFCIXcPaZTrt9dMtvUm1Bo2jDcl+H2CrnONWSYAs/EQA7WMMawKYm
xK8t+l5SBBTRSnmo/zvl+4YiIWnyxFmlfxIeogHWTzNJRTgOS5v5w0B/HJm3dguOFZ2UDNndINry
9PXwKxieoIsJyXqdRZLdsQlZT7VSzqFxqls6X2gtE8sU5hXtDThSksYIkdSl8yqsW70E8j3w1/Kg
0uCYFj6+5hYwo4ribEehkaW29Tguew6wiO/rxQ7o4HsO1FCxGDWWcF7+4zCJHxk0CGGqpiBP8UO0
wlHLAWZKQtLuP10HUTRiyzOpcXYG1d0ZIG/S88AXhK7CCVEXXydiMJPbxeFvF3u22TMyDTAfDtAg
LtYwWeD0TK24x2QbjEDcOdEunMeQgkOKeYogme2wGdgACF8loULXZyS2Uc7lL6gGpe6tJ2AuPYJ2
sFy1vcTIcfhvaghQzr3vpHFC6m2frTPmA1xWmk17lXcRZqfGHLDMqyRrHdc7qUnw7l1MbR4bH8r1
1lzze9jsEvhXC9kKTFic4Le4J2kouTrQb/wiUi0HIRgCOuSjHHWXFHQc1VZTBFbJbjRi33SJsjfK
4IneL9PDQkupkXLZAzD1NVMi1MdMCvBzGYyz2Amc9s9vOpk2dFciriM9+Nxu0p0AzumXxZO8j75P
dLZraCEu/a10E6Y8yiDTlaocCmHXvcJbQ7d13qq207dayoXVVri5FKjZmHRZfYzFsCwp/8KD62Wd
zg4ESnu2RkHFX6GLId1x+PrLozRLn2OlSvAttmvVVSKpXEDD1twBvWjuVRqW+Kkt//a4hLJiMrmX
RDPOvL9Ej8BipSBiL3MmwGROiPCwX2MxQ7DgQCoLg/VjSrlKdraWOd054+gFTYBGuBtBDBJbsn0+
kMAeYset8aHi8GeDPbD1CSxxFK0uCgd23CdkF65lCqj9E12Wz/byhNSntfXvUqv6KQ5BfBMwEsjw
AaKbND0LHFHWxweSYyp7+sYZM9YYoDBEbg8n5QfMeaAZm4rY4MemNaaOGlIgofMvx6C/7Knznzgc
3VH2vtYHLJ0ZPB6Ury8c0SBv3pW/Slq1RF5jBSiLDY0qePC1NyVHLClLEgiZB4N+1ut/mgYq97KU
WMglYAEq2/GNLhsqCFBw4XZAcIB/T60VeoW0Ai34JVYdyk8sNM+FVXAQQbeXR7+uuVTGFNBb1c4M
QFmxHoCm7zHRmKJi8qxlQNOyQ8NaoMBIMe4INreUAYlnqCye21rdZAmxB28JEE9p8BiTuL+JWD6x
9MSYLmwfekKw7sp2SzOqi3zkkwQVrXpLXjqaP4e1dcQv7ziJ09vD02uIvCkGhinjLAnVGg5N7LKR
Dt1CcjgUQ7tIGdlBoK8mTqwaa7eHBQ4Upbmr/UclqUWUoZtsVcCi8NAvvhhwciA+ODUHv2vPQzYa
N4i23IGAjpZHo9Q+J5EKjiB82IxU+a+Km/2CshmnCeIhqWHdkFgpoQHphgzym8LWIGWF/puhKGyV
T54PoIzQsKQkErCaB1mKSbD/fCV9Cd5UmOvAN5VrdlSE2DtjXJnqsI5GnmYUx8p9iFTS/TevFIzv
bl6B/XVONF3SFvGMntiCufyc6S2UWsren0ERAYhuE7x3SgcSch9DbeLjr6cAlOZRey+K3hIvQWVj
6hJUT4pXZDP6ssMs7aRxMSMt8PhQZ1tduKAfHUki1GC+l9Mh6cS6emDKjkHbJVX3kB8GNno7FUCV
NbP52aBwDsATNHGlHSQFcnUh8yjUCmMJdaT8v2GzMFMk15Q4FIj4b8HQHkfYmlyPrLpAtZnrJWLp
8JljhsAujQ6OgyzmRh5+Yv4xkbTwamqlmYuwbAVuV7sfW2rKb/whcY9bdRpSdQSgoV/XRVD+YVNz
ZCJjafp3VtTMoTBhzWXyB4hxtFWWXJJUy49EGA1DoSYlgnVtTxegvJ9qHbeP/YnfOVGbjJPoGU98
s/N6KQFptj0Hju0TdVwdF3kP+rhNFpbd6lW1TwlxqEEQ8NtoX08PUhkxHIrGUqVlQa/FjhEqcOdR
Rwv9pc9RC+POoncvP3D1nJuEqrFGbCoOrIyJ4Mpeng1YrcacUqFd2rvaTTH80hQG0fDm/GIdo3Jn
0UW3yDvtNIZRgARD7UEZ/fCivurYUPLxBXrOai3YfU7dRH0D1nOPmnFRCq/IWbTUfwyxdl/H3i+h
tK2dCfM/QnWz3wTCAeVWMBmIXCMCmmKpuS4qsEplq1ty56Ikp7m6qC9l4W0TEkD8h4QNomwqdehE
iSK74dBMxsIeWa1QIuRzRW642+OMp5OdFqDLu+gaiFPYq9hujFy8QRf0emBqcrs7DcjxKOrIvt0N
4HHlBsqHPFP3HAhDVzz/28Msm1X4suhMse7RD7G1fbU+H0s5mKBQxSYy5uxmG/wAbMTm0cYpe3Wq
B+N8PYnEWtDyQWe5dqInk7kJb+w2192sUWa7Tkzi6WOatuzgklF29GfJcjf2FAsPSZqATYTnkxwy
qXQ9t+7guutpfz3Cw0p98evAt9FTb71IZpaVGLVNxqdfuw0JRtJXgUkvaFrE59QHK4MQCiP0PiFi
FqNzzXLOUFiXOlgLJfy2zgQdHoqSO37twEdIoEkWGL6+QPF48Lb8yl6qfOfVjWbcT9mbXXvBTJGe
eXJT2HQAOW+OMszQ0++Vegh6n1M5i3awm4q6vfk4HIiftaGepzxDjAwwmFkKtkNxqT7r9J3DH0SX
NiPZPyv759uwsetBk5l7rFJdrOGeZgMf+kIzs7XC+66jNnwnJA2wmcOjwvUXgUfLFdQCr56Pl/5M
MXTIet5l3jZUZ362RdPFxf2fYc3XW2mVdKTMdmq/BeVivGKfEjAjprJaBN4FNl8IWZx90GuRCUL5
AlPFTzs7OIHLn6PRAaN6t1x8dgxIcya6zYsAQxzieqUVMdJU7i+KKIuindO3H+0h3wNBn2gOIrkm
P57buCiCAwDJKOW9COPgx8fCt4eQybZldtZ7kz8JlDDU7cSvuD4RVIzfA1ZzTGXw8Ev7IitHxhKs
phY7Uvk+6h2lt6AT2VKa2UNuX1GaEdwbHgsIDC4ONZUSIjgEgYbXJ82AAcoDkGy8NYr3o9aIjY3c
ZNkoStQaNSFiluC6ru/yhSqkYwwhCcf9rvO4mqm8VN4JNthZHP4JvvBMoq0GwG45MXUnzOl406pg
JAojv/xwnF3K9dfQcBhWPtqfBr7SBFM+MpI8EAG6O8zD7SKETPbexFe5G6hptR0IPEdcO80vgFUg
ZgnrwrnvwHZGhp4gEehCQfyo7B30Rg/R47o5ynAkSXa/Us2EdoSE5LMZz5ybZR541L2smogEJPHD
mjhmkPKSE5xYnEKa+nRrf1FQg/77UNHBdfxgo/mXQQkp5VSEPammvSsQeoWznrUvjEZGWGVZgfDY
fwTI2IEBDCPFMUjW3eAfbmVM42/kDAlBPh0b00hXQI8EQ5sF/G8M9PxjnYbYrYri0iMbYwaZQAbT
QooXl2+SFVpitifvecoLgnDiG3d1Q3dCNfzI/sBqtn35ahaO0aPxBcak7FyNbu7tn3mnYxD+R9PM
QMGREYeW1decfO/mQUNuALKBG5dOgg1LugEmGUgkTD6CjiK3MAwuN37Vod2kTJYPjDdRgBE2Q26A
p7G/5PTBVDYx6sOKZb14zxSjYWrWlhfPuskQ/TC9mTHBGXfcsxq/X6xLJVrwHL21eTs/qjJvip6k
xSzHOW/oAuxa6z2+cvcxMVjL/0Avr3feZPfQYTci5FEgu2Vv9bgMSxwqxC01NRVVTPZGxMIQpdDI
9NnxeVyBFuJY+8XKaF+pHqVSIwpvoAvhb3kh805gGUn5+TruW6wQbirJjk676G4SR/tcV6TrLvaJ
XG0MaFvUjFJlbIhYnFJD9Kc01l445+sCGfJUlDj1dZxrEBXIVPAMVP3qzY2oGG6TmIS8xdxKMSA/
Efht0dePc2IW+uPj8/owDLclalNBeAEF7cazXcZnEnVw347myaUU7toNMJo7Wptfx9pfzQagptql
gvrCB7HPxevn6LAkHl8vUELqbFiIYx/kkoBaE0w2ZeEehEoZgmj9xaxPijlSP3I142dEZsdWMeEC
NXMIJceLvIGRlYWr/fZUjQ0kZJVjMb7yfTGjHMsLJmePbWbx15PC80Z8tB0pu8iE4hI4sIVFhOLM
3eHvUSC0ksiWe83zGncPxbPR13ZRtZO9yIvOifgwrPKcnrKakxBC8jd0ofuKfktlYZ0LNEn/Gkaz
C/B7Lz/IR4Tsmc/YGNIFsUr+TkNTI/JQhz2zMwfaW4ogDSXDWIQZC8BG410eAWjMByTMO0SJrO4K
B5ZDB4+sFeZpWxFnPmXXmL15p2igmcswTXzCvNCLU6j71mC2X1yq2JVNOYhp6R83pvqEQpblasKl
YxBBo6dmL3UIE/4zuVQPZlnKfVrGfAUkL1QIJ+bzanToXFfHiotY0fSZDX6YhxQJ4bBLP9kQN1+d
qJOL4TpFQzdCnuInKGpGEbAavEpfW4ZLMAqDZGdkTksvbbfWpPjq3DVinmIqZPP6fKaNk1vs1ZIY
FN5168ZBF0dlSPSCZsNf1Ka+1D8DUwocAmnNGnZUcirNzMItuepDzxXkHmccIPjWGdLCNVdXV9ub
KrCxCIihATd3HLcu23oaJPf+Jt4VilvmpY1licwy+Rzw+rJPPyI35B1FPl3Jaj0ns1Ms5BwNwhMW
i1PyhBEUsGbmXvNktID+K5lhv+kn+K4Im4HJJW5FFRxugqHjZwL4UsM3zRE4eFLv4x5uJ4OjkBLb
D6QJf8XXbgNKd2ugg8rB+AALrWXFLKxnuP0ZLu6eyrg4jGM8AupbYfJHtOrEZWy44JSY7N5GZIu4
hZ6mi2rvlK4icPY2+FMXMlTB9gfDalCGXCp5gcQitHN5rMvLfpuAyoh55DJrosCCDZCbCrLdMqj6
ILYz8UmIDQ5l0HZjIbOAGc/3NGM6cV+3iCfnrQyaSdyBCe9K2GQJXoTagVvGhfBpBBF1HCFP85P3
OsbFNqR0kkR5x+uPkpiSBreF/3fE1hP2bFUHDlYBs3pPUqn84mUQ2gXAGe4G4dsor9XFvScICtOt
xtmPuk6yMPhjMwDkZRVkv7AF1VZdAdUBAZmwx6E+xMNdfSdG6RvnGpW1G/FafRMUe+ErDBiXIfmw
3EPKM27M5aftNYcXC6cnmNSJJUZTcSjZGdLEs4eJPwKI4+AzFrbZW9PPI2aeW5NzYPk8s7Vi26E+
ZUjOZYRoe6MaJJlK/7dunnl+EBAXnGVTaO2EZPTcrbHwqKE/PUnQSh9cqpvHqce930KcsBy29HQe
Ts9vGPjtiMyIk/uusDu7fOiQ+q/RVJkJYJHghHuB4DLoparc/xiQ2f/0ILqLnx9AfMuJbt6g9rRs
g4bPbHby76+HolDvM3BladtbRM+UurOCU5aBIWOFH0kwTvP/wyiumgLDcfdvNcYslDFiJY2v5y8F
ezIJnlruQZlM5J3r2No6Px9esI8eZNFwxjb8ZTHxXQgJaOrJKVJXL75mFqBI6H47pbYopOYykCCH
Xye/hKrEGEntIZkgGv7SOfyJAk+8beaH8jAFa0HmXY3TPF9xEI2O9hsEAKlcKZ/0ZDZlmXH0xQQp
5MjniyRNBROQiKaHMugydECMR0AWzaXOyqiunlkAq6cXoVCW/KJDa4vSuWagiqiFk+zm9/C/meIS
9YhQsE1qq7nYyA+bJrOQRIkNRqNZQgOhQ5FkOHXu+gnk2q+uu4fKQB9O6DuB2ZlXaomxckYShM7r
EBfX7VL4qRqkMm0ZiBu+FtD5cJ2zf9JOBNzJWoehX18YRQuzFQN5CoczrLTq6ITr4XS4SKhW3QA0
jH8VxTMQ11dGeSg20TlCuGgtFJ+gF3wxoC6tBaPyUajKf2QUrcTR5ACzDFblNGuZzqnfjI18bg7P
uzZj+npjEuQ/ACfXY3MkfWZplt5/eId0UjRO5pG+fro6/2PrkSZ3AWHDYyOm/R3tWxtJcrjei8p2
ZttuXxA+4pJaUm8AScDDFtNNNlOtRnW6wpqeAd8xZmX3oeUeBodx4p+osnVDsenAW65L59gHDF5C
f6uZIcln19VE7LP6FKYfCn+Qmo/TfDMCGRiu8P5p9Vt5MelMFUDditMFgeVtETz35HBKDhVTWSOf
8R8fdBwRIRjtL+hpO/6Fj8LMjEhtoyF35v5d/zy5uZNY7ak5vOjupEPuqZR6e99MnM0i6+JP64/l
ZX5nI7OVP0d6AfIF6YAoSI2kb1VmaZkIrA+Vfm8a/605uqUjORLp9QC1mThdbH7KUXIUSpFMh3S9
QjSupUGXpHuDhxNbR0LvqqQi6fgMP6DLxnCksHnWDZpsAVcQ5Lcsb3Hxl9qUkRv6o7ra1IpI/3Mc
dPLnw9DBwctzfYvGRECY9MOxCktoHoc3UkjMU03q0Dfhr6/gceqLqZHfUoQ9dEMg2yVX9cdXaX0I
2OwpvnPc/YVQu7ejz8BNWvBO4qy9BcxsGhwr3E2WJZFKMBfdnR/swWa7jAlTdcGOVmuYgq3uavux
01HNMaRUmSC1cXILAFdm1SjlE3IZSnpvsnzyB8j/Q7UcmFDlmiF5u0Qls2nAzieDWezfiH4bjXj7
UY7ig3qp7eJmw+rJgM5pyiCp9Nq4fzoLdMK6y71srd38HxOHJs9K0wWcFT0hq1YrpVXkSFrrY+qS
8BOU6z3PzeQDsQJu/gb++2f28N8hPSYkpoEywq9T50dTMnStYJ3K67sHbFfYPXRHur9Q56lo4WiH
PBiNQyYNwCj3l+WiAGUXUBdXx1D+d21yeBYQ9Z8ajdVcMzAos6OWAvWqAVo0g8walSlQ92fAyibD
uwNwsrkJc1+D5TII0uIEoIA4QC1plePUlT9emsDiTA502/2MBrB3ni5ZSKFdHMFvjAZLr8B5O7JN
AbzNxnU1UAnjfN78OLWi5eW3txG2ZvU5E9ToR4/lkJIgt4UXH1Dv0lh7aT50qwf9BA9UZln7snUF
npNhJBfK3XMEfMhPHaGLp/XCYGITPsdkR0NDlpLWM1jomA6dkoaNPhLrzK9M44yOVDVyZHtLgDxy
dh+BBrBsHJN15Dh/+hf2ucbZQ7hmMlmzSWfy7ZXbDNierVjUneuIARll7++HEJM56VoYKH8loF/3
ajkjqFXACRZPDc0IDjawxyPMedoTL8TFifz5aWe4Waq7F6E2mMXRcEVZVWw5X2IDzOnxNi5R0VsU
67o/Mow3lhfru2+qZQRKmep7RicvIPLReQvgq2VYP6gZH2Avespkqf39lHshN2plmKQ3apSNqbGK
n5EkQFwmR/elA81kDlSRBsnB6BI8aShaF2I6DVQey5TUOf91TMFPuSk0dJ84zB1Iw8aynHrTfhdC
SLaCwZ60Rp0w4nmaPYrlf7LffYjbLsqrEOPVFFvfIaUKTcqczFOLq4jrUXow9iTm3rnXwu3LS+i7
nqmMCNCL/k+vM/dcMnfWheoFb5aSd7EW7/UWPADfvUKYPM68J42As0aXAeNnCIhZP/PpdRnoo5Bx
RsLCNzOTzWdUx3JI210fucfKvysNRbO+jcFp0RdCA7v1+Gy5KXsgyvZnp1jmJF7v+bskSFqCiVIW
wozvieS/r8CjwE5bmgoBbjB2s6zQ2sECl4Dpt3RB2QY9ydGgAfJOPq0656NE2MqPsmfa9UbvBnsu
tjPhylVsYfBLAYcSpBBUlB35SB01UNooogbvZbr1yJ7LZlr7OpmsPeUu6QDTkq3+U4AndFPXIrvh
j5+YnkUcKzq2oU12CjlfRd9pzzmey7NkkpeVZaamv4gGqxTQNLQR9mRLPTQPAhV37QPEW/ZCFtQr
3Lx8aKjvfRh/0uq2C40eMO8ofK7l0Zmf1BWC+tYHa9n7zraB3PjRGNmH/i9h2bNVmiBP218Qe08A
E/4X+RoLtsaWMIAeIU7djYywaXQ1uARis+n6rguQQhcvJm/tujnlwt4kr7cz2uV6ne9dQ2FDtDH+
JwRvLe7w/w/0jOWbUMzxVocPFtG8Zvf9aMwL20UL9qB84bIjNdlxEFj2woJf3p3iNtJ9D5capyBD
6DHOjSPFwRHlbcnIR1pT+B+/pgS26I+NMfpBd/srG+qjn9Q97ptcyCME1C6xG4zMIX7unOwP38MR
xozWTqK8HMBj7iDOw73baoYQOVndZGW83A5aC0+5AllhsAENmc/kWKQmQUXeR8NB+OuKEIFLEU6t
1MZDa0Vs747P2Ylys6KzTmljqBLeCsgz9B4QrtcfLNmLylwkJoOCGKbBl+CxBbF1RJORDTWv16wy
C+Q7NfmICqxlIT1WCl87eEl7kvEfc6zu6CeP1GBx91EnfaEW7Q06buZPN/uHV9iKmjLvdtO3kv07
AgCNZa3UfM8IsVcuMTt7WxiApaAdKHDcpEvChml9ds2BGUTZu/enAng0WNOos2dcb1r3bko83jQ2
ZDmGUo3zkLnF0sNuhaS1COYg6y4rOW0s+FTd5Wvep+BJYQ8G4vpoMKv8V5HwkkSkski7xMK/71Mb
wF82zDf8yOVS8KZArShFr4atwnMFwbESxmp10XNGs8RhqzA2c5hrQ/VK1CCAC04GNj6alPw1zmVV
DLfmUNkewpCIiKoKhjfZtLv1OekdUJOJPSdyCe1MJhUUMNqrDJX5HPwAcCWt+N4Oa6WLgF/qbm+6
0xW57fSB0hHHkHvb+cjxpIRLsisp1PJbVieG5D5MbtbRVUfl7sVHF50Tzyz3z3Ow796zcgPfp3SA
9h6VhURRYO0Ab+8FRRIdKb87ZVmv7WO0hHsa9tdrgGYw2JN4oBc+KL8khTci5jH2nM4OllEfHsXX
F6bSSqeiHNrnRb1xaA4u1aW5imWa/DLpRrmxiBSRmJKrnZv5lh42nFbe1QLcuUvoPSZBluqmzUWB
SePMXeo3/wV8BeMITev6t6lbrOlv+P0XjNnI3RK2TCvr33y5YWUfGkYFSuweqFP+t1ICbMlIYM5I
FYPMiQtJIBY3SV3KDetR2vC5xFUvdfDCztG3XBvMkGeQ2taFSxAX8UnsWOT9ge+ihLP2wfkb95RG
92M/LCFUKh1YWKBWuSbP7JnSXIVWbDRDYhJDh+KjlwzsbIhPnf4Whq97wRkqd2IF9/OnYyUcfewI
UHfZBEpXSpNOAmo3q7FroBmKz62UO+PTnrB14oKhGcrWy/8bYRArrhn7YBjIBHI6vYMeT3JHCvem
cLPqFip9mNifKodxsyD67k/rbjFJXt3jBHCxJ1GmafYWaMFiz3P63YxtiSd5TPWrfdKJNOMJHBQ2
AHiZ27V20BcBPyhuZfGE8QvU6lzltDL6NNxd3qXrFqIsnioeODGkyvFUEjYXTPgjdkoF3VY0/0+N
pb357pHF3UGtdtTlM9dwUxX9K+Iql33hmNV2sc1yC0kxja+IKQGyKBRBSItyIKXCdqS5tcHbz1Gk
7qhsOI5fQwLpM1IR4r69dQTVkFRXkzbX/eRHmhzEYPsXe9B8cGd1BM8QzbZxdzupsyIoKieno6kp
TQqo2TUfs6nydWbzNqZXSEabFT5BB2DrCWo7CRxis+7B4v4arFKPPkYBBo4oPRV/rh5bXCaXae+3
BEh1YAU9ypPgY2wv3C5nWxO64trC1gMezR92+f0BF5YmyXOqcqcMKNBb4vxL05I6DWecaVwtT0sp
V3138eEN5Fs/A+qlWvmt2NLRWgr3VzoTevtnqtyPO4TnyIcB0lHfYQtHhM/D48Rn0iQIQkKGCG3q
TREqdRcTif+evjVGuE+TPBWyJYjGpyUeITHhywyyI0LIzjwQVVzWKgXH961o1tLuev2R8YxsQLtl
oNgJJ2I3yPNrYxetWwNDIyQfPQ8HEVzUFqWIljX2caBdo8atL4eGeLvVgEHtfOFkLnANWlDtOwDa
f//umn/H6iORsQJPxjjeHGsnVh43DtSJi21ZRUIzGEqhAR+yngBvy2ttVDEsgu9qHn5ZRvQ5VM/x
6v5Q/YHJdjBfL5NQT9P5fM4AZKqrAIgTp+uirO+SAZXdH5+fMiYfQGXXpVhoPn2iCloYqOmuRxKF
XusKNBgXkwgiAxgsSRXx94k+zbNtNC2dFxVAytk7hVLNZv/E9cZVPd/ZqjYuKfh/TsQzOPteYCSk
GRy7m3NtRZFmI2qrANnuMIMZua76gVLQJFW44PyAyjnTaOChggQZLIIQaO9hRQs/HuNxJqhito8e
7Zlico1EZAAM3MXCk0z1h2RoPJ1qvMnKzbT9DO5/3PznEki6Oa84YZ/iPMCi7+bwYcB5dtF6B/Ix
Mp9k7lWqUvwQvgbN/KXa8YxYHXO1g8js6gWn1Gdcl6uxMQZPGKmuoq+l6FB5qfNJibVQFTWFS0G1
awMFSFyIVG0OKxNkckeSrtj+ojdwlNKwhC/KH0a3HWKW4K1+PZF7cYiekTWXUE4K8qE1ydBmMRzb
0O9B5fj7ViszVc+e+U+3C74uJYBBNwWDGf8idAJYTpEnC1vFGgxSaJwLwhnzP/fOUtPJHtHENiUC
/bNkNUnoDE+Ef2f0KSycTBL1s+SZNw87/xRZn3RJ/ljeJaw9SZnnVl6fE7aUmUgC3Oo1M2qqz3ct
zYkA+756p7LZsxWwaj8fJVAUR4EP3ggQHOpDflsOEO17cONnyHxkNYWfjAy1nQUjouBRbv4CZR1E
JCAAMo5RzbG/WxEkm9e9gaDl/N5WXXCaVIC+xWfnfVcJwSYrXcctvZNzRKC58mKFryPUjL9pNUA5
39ZqHMPl79n050xllYDpL3aIYpmh7okN14Fq+ItcACoEpSwxTUlw6F5y2i7rm5aDoI+RW3DaW3MA
oyF/NCE2KAZWeLpJzQrwsFpe8m9g1Uh08ds3Dzv7peXfrQ4GzHzpFjdwMh71GHGwn1VhHhYy8KmN
fh5O0MkH4I82MLhvTE3JEQegq4q/5I4+IbwsT1ETQHr5ugz1x9gaowjXYfLjR9WaMpXNa2C5aKNK
y8NsXFfqli89MHS3WOfsHv/+JBB2bvkmjpBxQ7cLlJ7y6d5rUcoIvPnXgIadwCfdU1ImiutpyTr2
vapOKHcz9jwJslSy08GSi+CNgTxC6Gh0lexw3YW8T5OVx+7w2SwYKJLo3+N0jrAauG6LCFLqdRF/
Tm/+EBWu0Q1oIhk85e1dgwsQMISinUQhGt4ocrroWP3cCUTg8NmLaRPE8YCgnVN+HKOBPfnsGJeU
sNMoLOp6Vykc1VSTHlG2VsrAUMHk1gpwFbQv5yINGI1MQh2ZV6xHktLyNx9SzcY8eYArpKTgcl8m
WAy8tivrbrIpCaFJYhmV/ZjhjXvVC42Rk5Y05Q7SUcR9apkff+/pf0nCtMLOv677o8md6fUtmRt3
JKvVbHEDNvqAieHNIl6/zJFncbjZ2UdcZaF4puizCKni4BdyMbNijhdvluHgNjZVpm1zga8NH1cA
DKqo9lF6HgSU1WnCXZIcjji6p8cUKPwUycDP0b0wNjoZFF0EPJ8TXrBEoQs32/B1bsT90ZouysaC
nnDH5706mo42ceZ9vQN+5zyPCCfZ2k4o48gwwuCzyhWjiFmL5qwt8LmguttiBsK0zR0uVOOe5ysP
D42HyCdByzpePkSJTVuy5jBjZb34vddrIR0jhNSPIGbUYdti91mzSvKZbQVSGv1uz0Wy1VB+kWjN
LNPQHNImtfCZ7Cahtic9CBzI8+wifbkibxQtiYrcVKejyeU7cGDxsihhI640T6gLT8GuVAgSwtOj
v5cgWi8IVDcml9nCXTVM4lTr4U5UmlKY0VxmvpGDRge+pSSvQnj6pzwyzjLFV+DP+ejH6ee9+8Hz
3lM9o+izHI2/JXEl7kVesinvM79L2g93fSRLkHTHpIPhNjqlLduhwpDu3yh+vlLyJ55E6iurxShq
6gB2TY65lYHygIsTe0UqYsrHH73AeUIeaIQt4A60ucq81u3bDN+YyEMh3By4RfsQzqEueuaIpi6E
tnHN2uuK06tCoDYUhvm8eANxyVQmOzVWkI2toHvHxz+zoMRRsZ3qbNVxmHw/K9+RD79a5IMiX3FW
9dxB+unPTRXa+x4dOqR9i52U4abWf58ilYJV3UrJSwPGNIE30dLp1W0fWdT9EL/KrS6uOJk7J9YM
67Pc2Lh3GGCV5uUxiz6gVM+ovsi04UQurY5r2keNbWEZL1MC87LanT+rpPhz55XtsR3aDqt8Ytgt
3lXjEEmunidk4Tz+7AdbUDE0YsT5XNLCrWpGWKq0re5dh1g82hUlVLDpf91FQ1RsUVjbvVZDBCov
l6Bro9IgWfrdXoKHC+co7iTv+F9EsyT1IMjffmDQdroLt/WCBJLQ+S7fc/PhfVFsScg04Ke/rMm1
B6/ENSc51pne9SkJXktrN21CU5Jo/i3XsSK+NRQ9J4HlRNIAARlTwyXsuFaFs4CGr3l6MnmgULVZ
oqJCEqCbJjhFrisbSXky3sme2tmLFhTKX3hHrM+6Q7UHAIdlMF041G+IfnCsZGli+2eViTcFeXWL
6XlkEOsh21jlpnDIbL70RUbzMnHSiCPRd+7p3c6tDdZ3pLPzJZT8HD6dhAZ7NxsdWBmDjtQ3U+gO
q1+XJq3sHYKHhY3ZyvnLHBM83NNzL65gDaHxQYvwBa5hq2GLtANiUbMH9r1dcvAAfRZ1MDHXNNpk
XM7Ld1O3a7YPFHbiDqEcZVSHKOb8fPIb/wj6MBH5hQ9kBnt2vtirwP5Ba6+E5/uDAhLJDxcnwfLv
Ltsjq1oM4Ee9NPt2gnpOlZT1heNOLzIveHlseXqhl0rbST4Pw4lTUNvzBKT4TFXRfSaxUbcP3162
wj6r+6JjJ8nbE+ai7a9Z1kHa+BILupO+LlMq5KrhH968XjqK+wA8ZvOZB6A9pCK04LRQflZjzK2g
aO/toGWkzcW0ItnC8AOUiPh7/pi63c/sjJPCbTcw3XLmzHAaaQ9Q6ekydaEs8ufPE9yKlhrofZmP
4sELElGo6F7LFNujs+4x2XF9VPRYg422ER/zgpzepW3aAiSRD30JdKeMvCaH1BasIdIivOKR7w0L
yreoio1T/GppZKHMcF54P+h2+zSVyhDw1rkcwWvD/QyuvBtQNY8bBsbPUBQSKPRk960Gd7BkJOdV
GVGT1UqL996NxVGbfzIuQTk36gJImjeBgn6F/vhtddkhwlzbfTV0erupkYm5YQhego2I30aYlWLe
Loies46PSKSjQMHRoFBCUayXDdFwAbFEtOmoETwnOqFd1t7vylJbs9eIYL9PoH8uSWswxyVHbg4C
j8wby6ybBn27Fq+fRaIzD2PSDOhpiFqq5vmQ05SUZEhB2e/8Q72kf/+wgiz+v1MyHzLorsYSnEf9
DmXja5BY0lqINu6bIEUGfhJQFseNzhGURAjmv/IE0g2hMVzamx+yM3Ro0ZJfbEy7aI+UIEQg0zXa
Ie/MvqI/BEnakUunOPn9T6ddknV2r8/S2P256HepLyCTCoaLrBC9R/jun65PINZEAL9jjgwZuKb3
lKnCgxt1hkK5o3fwielPX2AFEK9ojr/SlwvgebVBt6ieYMYSgTtptzeaNCdNGBsSXUmdXBIdC4+D
OhTTkHC0G7VrYjxmtxNAA1WNsxzAeqPeDRWRvl6DCHVk4dtoXtVKQZFhbYAEYN9f42gYeaq4aGAW
dmJNj+Pfs9fufrAvC1ki5EMRn3ICJ4Dq8ZGF6hKpd+x2ZBG7HZCD+fcVeo/vh7ApJW6Uq5qUbZlt
gJ4YQ+k1ed7m3QcbGImd7TzWVHMl4NEJuqN35qy9UoBCs8MdPLxyN4uMLUvEoDCSql5VbljYUvMw
eZzhyRjzBFxOrZryx813VzMFCTgwoD05/cjefjArFRXVn3tN27DPhHwA5W9XnvnBDln/A3aNWAva
9X7dgmRI/cI0gceIv8pjRioyao7XQoMi0W7yCk5EVy7e7fP/MxyULV29jU0PRVGV3fPKd5ccbyvU
4aNC+62v5Tq+/yG+ixkJM+KAMTTU08OdmxzGYEp42tniQPBAQ+8hyYzMN5cSLicPw1NUeStBV/R9
CgEziweQitLFRz9TTfNx1i7ZV9ELL61T11HsCFo8wjRyV3u+Brmi2wyugYM4PT00aaWuhrjaYR9i
E9j5V3w9Jf9Nltl1frhtX6C/kcY0gjm307qtd4d462tAibf6k876uLQGMZP29VpYultq3pgqgLw9
XAF2uz6iqaputMcK6xzIUgl6+0K3JULzUMSQyF15u5Pow12CPbHszijARf3XXeRK+cPfV8KdyDsB
URn2Lhx0cJyJUMx4AO1strvjC6Q682uVX0xHKEReias1/SjCPphPGosVVD7kmkK+nbG6ZErYOyPD
NRfoPKS8ZZ1J2CQF8bYI1oS8pRrnhJtUP3/FpoAkG2TJ3y5VgmTEtBKScEJbrt+K+7p3OZ5O20f4
Kb/GPiXq5BjTo+AXZBFISEsNz+EJMhylR+CZhWuGyBUPPPIpT9v3elJhEdErR5jRI7jzh3bztMj5
TXS+HDkWARPYyH+3zUTFO1g3g2Owz/ohr9kwGKA/MiMij1dCbkQbKpxMiVF8d6QQciHj80SSDq9W
Udnctl7Gu4tEJ2z1DFh/ULVP+QxAfzANHvKMMgSXETH0znf/1R97XDAeKIgxVBkPdo6WZXp4r8Jp
DnpUVrRa4Gk/GPspEdptiF9wRsmDyD/9oMrSv26Ymf24Q4f+3G/c/0L8cBbFoVGw8XBrohaGzDqh
DQS6qmQkgwM1vnnFl5mhuyes0EzzUjrs6ZLjQCXVBwtaShj+PCSMLW24BXLSsXQmt1COSTstywIB
YmmEUSz7lSH8D8SlUkHoCU9jSZNHzewAcsYx9hvfskL9JTFqpXAnJWaUwGDMfR6HvBLu7nIlh4OE
REelAFrkU9Tf71o8olY7Jx1hd9OdCIQyrk+3A5bADtcX3F63ZXK+IHOTYVcYcoZPC6zLze15tSGz
wcDSgoT/6AhNS3WDw9/J2kETb4kxmkS7/VqZrUhgLxV5vqcCSXg4v7vnKUWddejlP+nsqJweVrKM
G/Ozn+GemblE8NZOcI4IrTn2O2dUNdWEtZ3/Fis1EfzunvoTalC/8aln/Kz0Y7NERfxyUdwvzhfh
07otDU5nil6TTgodQAcYIhxLucQH+b0sPmKLeJAPvyZHhlvwWRNwGoCq7S0V1LdKU647PpLQfdfO
Zr9iUwEo8w0VYquFWojLPsNKP33wjpnmCcYnSuVMlkmKw43xcNGDR3HwuaPTObylaMjLkGzdN7dP
v+qSD8xTSlnnDokxkR/h1xI7OYY0B+bdL3iwqftqBP3jfiHvCvyRelYRNguGLZ5A/B9Lftf+5HPH
8rhvg7J5Bh19O13Jy7MD8RXbfE+m6V1MjQJJyhXlaELGltcg8DwvX19P/KV9XfYxQcA8SuIiAgI6
lOFf+irP0lz8XLMO27l9zUjnDdICytM+hc1p8PfV+pY+yl1RMd5RpiBzQNK/83DW48KFekjCvPrr
vvi1c72XQG0EAEdWH1xC2OShF4kaeyYMnaKzDyDw4LFADbHzCMiBsrUCiJ2qPsOZoX4rD9aur22D
RB5bVJV32oLh6jHKfJK6gfWmeGCfJtmxAhLgsPL+pjxBD0o4mA266mz3bLPCBJbOfbXy+2LCmdPh
GJrCcrcM15wNenqEaHXpiJoR3bNNIbcI3rqs96pW5VEWD+pQmJkdOHGckEFAfx9GvBXYqxcaaD0v
ZQxvkAj+xiEXr3MSg9h3TEbwBSj6ntZQqscdCUIsunbC5yWMBx0upnpXFvGGF/zmCofpwVoTA6IO
iXhXbHaFrDVd1+QBN2fYw5LaS20iTXFtKNg1yxMiinJ/FaOoDK5z5CS3JdbQewUDUKmgKcMRtCEd
+UfM1kIKQKBzxO1p0nLWlcKAhPDYqeDZTF6/wPLWmFfEnIk5UgFNywENF2ZxKyIQsyg2aHNnQjc4
001cRV8BZ3xDheCi6reiZyYY+Whl3s0vfeGNmJvRZ4foyVMYHhofObc39iFuR/4kPPIcd3JXXS+j
xyMrdX3+y1KEOB3ToLyi7SsHSndn/OTladImjJNavH8QsLXrZvBy3H1yLGozIdPUxhCJovACc0s3
vvW9SVi9pxLNp/ub5LdLzZJ9CNKShzPHj2lF9wJ6Tuq3dvxXjyD4sWapju40VHa/IKf7/UYxwx4w
MxcCCCmUagX3+T5XcDq4R8zkVJ9iFkJ9IyrIedY7WHiz8FRU5rodPu6eNhmLuc/q3ydwFdTf5R8O
ICCJRk+LlAlVKt3efKm64ck4a5tbln/wXc+sg1o98rXYdkQf+UqT1o01B5NtF8QRKWhY+4ha+1oo
oUjKovXHgeJkDIJNgGE2SuVlO46Lb5oPf38lKPE+t9e4XnhMuGyC1WtXCIc9UlCEvmHrtL6jr2OG
pCzRUNUJd5uM8K+ztKPe5wu9PrmPo+dVbiVQe1V/1tQKGlp8cxYut49djZQKdWjp3wpKrIDrYDMr
HVVxTD/aO+o8ckBxcde/LlymeUQOYxG2zqA9RVzkg7565fi9B30sQXbOow4E3RvTUgJ3JV+DRqsC
NgDbUeY1+6Kr7q2uw2ahuo/YBJN7Tkcuxec9ffw2LF0BICBdI43S/pik3i4VEg8QLLo1FLdMvaO7
2iBAjgYvR6uX8eSH+2sVJY4NAVg0QY04MKi4sNemkupFabvXk3o86nDv6OoyvUWJdm2NU3dzMNvS
qjBG7WmUG6MnhHpo+7b3k/wEYw37Bj1N0g5C2P/ocKPIQBRVKunL75GATrua5dQJShRboNxEIPf6
DUWsvYb6pQLRJ6Poktu/NHE8vD+IbPQWxz6EihDqDuBHvPhuVCJHU/CvaYR2OtPqUOLQSmqpP4P6
92SY+IfbNvEwcaxhh3AlXU88SAkTH0zIQV6Dlozg9luyNsFrPG4FiJeJ5sLjUdiGkZ9/EG/lH6/I
iVDC7J+kGsCS1zVH6mQywkAMgFzYuoyboLwJ3RpRPiqKmuV+nvRvwRciFCtZ0TOBJPg3RJf9CEGA
mRkM3Gp6NGFP44687m+cQQduzDBg3XF83WKdqWwRYKPEP5c/hgW+n3usfmeCDZra2rHkpu/9wMTW
u6Ic0hpEvj9YWfwycuLWqlaaiMVmhQQ/OetLj/Bv/+ZU7NlLrTZHO89UDITkiZvGLjHmb9ABsG5P
cHG5DxYmbEk3wjNG6m7kcqchuZAnTXq3RWC+5kDlr8MeSgLUTmhjCRYRp7Wr/eGQVgo24LweMae5
lYZKPtGoT2Is4t1z/o76Ar6HOpQ+BOynjqOqJY8mYxXtJfJW2c6u28U1L1lwQRVtR6owzmeARW1F
j88q2Vc5qXyUPuCyjkLdG0Ez1rSLzt1WqayROVPKb+BYKQhl+TM9LvqxBJm9wT3/dOCvyE9kKhx1
gajhUwB/DM/k5a/YYcss9SVnnx9AzdMAMuzK4D2PkjkVaOVw7VvmAioZP33g4yi7ilsOu0ARQO8k
0I/2inILr+DdsyYcwd5B12hi1rBvehY5AK9kBenX3Rl5j3cRyxumymrbnqhA43cBZD9Iksjw7yVR
pbagAB+9v7Fnt+qc4N4zAbE/jd1m+TEsC7PIOsd9iEiguJeqsXhEwR830qW7QtUYZXDKVb2CUEqT
8bhT3QKAY0UEdinVVM1BciNFnXwWKdv+A0nZ5RvdWTKnncJ2mbpZFO4TK62mekOBqVZZEhzb0M8a
UifIcGwSewOSRSKN549MH6cn0cybVrXO8GQCbAgOefAXjkpqngEHsY8PjCLrKnizfxawUBAf6ERg
pGhdtPOVAvDKJQF+SUX8rx1QYiFY94MGyfXKVjZ2Px5SadI7v+D5SobmG9r1URerOAR6/jM9u3lN
H0xSZe+aT/Xupcigm2ed2NzIcwnofAOuND13e2acaEFQAenH8tBQ9LS0fdHE41kTcFXWAI9zRjPi
ecIVjAYCWW4xZbF8qsPjzjxVJ/oHH7p96z2NwXenUOIx6fzL0Bp1c2vO1NmyIqh/gUSUWtf9N3ne
7mI9hCCPL8J/a3VqkWlS98XSs7qwoWLl/9tbjC+ch2l3pNeYCjhTuZDk9PKFupovGtuyBloPr+63
HYNu+mVsqFHk2hP18TCD7oq+yvLivOwUllY1H1X9wb8cl+zD8Ur8QncZoZ3PVUFdWZdsKvMyrOs4
IaHTklQ9hWYhb8mKOQNMSgKT7k6IqRjCdJZtJtOV42N3ER1eh8Uk/AsvBnBqcpkkRQQ9DesOt8hC
rmi8SO/7y0B8CTMfq9HD08HUlhEp3sHu+qnvU3TX30904vOhrsfof+JzLh8rCvKleeIFLxTYxdAv
YnmVI2GOqz7dn5J/ndDROhflYQEmMdDLGLo4VJY3l6Beeuk/kYIlnETsIdiqrMiyaenekfJqRX8q
gaAuLKnCvL3yO9vFsbxTuZQGsQ3BYrCB0fJke9CoODZneNoAWr2Hv8VPGh1fzTQH1ubffTlCLYDp
0Sp+Y/je/31f58Bc1OmfB/PePmyUJnFubtnvVweGRwtGhddk5prHW6LsQOFO11FCsdNWn5ppzgPU
HZsif7SRf/mbgXfXjyQvndgcSa4mWevldUi/ELQTygJ0vhbLezFltqUV/AEcJIo0ufdwjvHhRUi9
nAy+68uJKlzpTj+zAUElHFJYV2fjki7IvBAINdRVMCgosceEBiHFOFClBaYLXeezRmKacPV7aKtg
mKQep2haNCh+TuLhDZcfn9XXqN8a5Yf7WrYl3ZZJD2CHELiWGgW7gXO7d/uJy8Q2/UBOaVS7cY5K
27A/JFD4iWCbsxKMRPJEDTZfVOIlAF7EAJtKj1e5Yx4W7Berf0vGfrWfdYXxUixk1ZK33DXtyYbZ
mMOlaWyCMmLqKtKVN8wq+bBpXGoiMy65HerwbNirvzMlarJ5cYpEbFbGCbbH9TfsCLXj4ILnm4NB
XOYfS8VMILManp37Z+O6HWsIuQWoKmEP94KhLl47BOpoYtRXlqQUKY2zJkLZ1RrkmP4ueMvpgoTb
O8pjAAXzJieCCeafNe1wIrFFLLwpYKTPBbwuam7HnxBn5XWM6ctcb7Yjcky22MAG1lZMtO3bZd3i
LxdRC/XPZmzqi+bqFK5i/Syrk2Hb6zMQHANHEXuXgf3v+pRonNfDFMr3L/TmSNiEPtCHOi8OE5CD
XIRsIapaZ6xBRjd/bO8YDBXx6TOeSYmNFvd1wzWAO8W25u+SYjJ+C1hykmyY/NR0y25y6RWpKb09
1OHEIMZ9Om9JIx6yHlao7ZitDEXbKrBFhTAjcpvcewlYoXGe/P+ODX77dSMDbduyG23ZZ5KRhyUd
S+Kv751khl8VP0ZzP6if94yrwOLjbhdtTiCpa3E6n1zE1wrHmrCneIvWpOJOUc90wE/ROVnQ2evM
evAEwl5Kv8P4gGE8thDLvISBaq2AFwNeedq9HER+ztpFth9OHPEfeTmJBJkqSvaPxOb4pXGnrOk9
lHnBcG/OL9H8DN933ItL966J7cWJuYjNi5KIppGC7zmr5MEY6qsD9YOnOJZptQNHQj79fqpAtxPw
kvjkWuoFBTKfmeZ+mLoYYQBbsHKC25/AF91JnFUamJvxEeTDxBEh77WWljDR5zPGEYw+JtP7qRQN
3njOSX6WEOhW9fk0j2QswDNB7dUpQJB6+MKBhjNxb2ApI9swoPFLPA7IkgJW75vHafgmyQ3XOPOy
EHj0dK25Mwnwu8+XLD+4k3pBUVlzDg9CXfJWm4W2XDMzwx3B9+A3Tj93/s+na1cxF3bcGddlJ8dm
GKb/yqahwGtL5vkRfePXSp9vYXazaf+7uTJ/HM2A7pnylboHoG2x9SKg799mLUWZzBf2rpEvlUmk
0+F1WeJYLzYaaMe1tg3yAosoKzhwDu0QyUoE7uKSLMAZQz8r7KFA1b3qFgX7BFG/H/+dwKmJO5Jj
1U6hP12+lRzd2UC1aDx3e52F0YPj8LdVfhbnURICmjbQ/JAErJi3S2kny3Y+6faBs9kOeSjumoSO
rnhwXJv6+H3n5ZPvbqYwpzpea9gSR2F5Id9TuLDqEVj4ydcHv7TxhJaEMBLKeuTfyQ5aUvThESCb
Y9IgSrPKzy2yaGq6hVTiCCF8JcX6qQ1xyycJYQrngc6XGJADzvBeFkSGpDle9dqWyVYHV4QHfX4A
wBuSjmGI+53Q+CYaXZ+mb2QRPbSgcXNYa4sbHFmxNzhbWjr+9iheeECeEdkZKzasNLxWgpqbMBCc
VAhrCSKzG+6Sm6s8G87XqXlloUeUGRCYZDHmUYKOitjbgj6i5jGvbg8kXnmcp4Rvnt4ZKWaVIU1m
jaFMlKParQTeU2AwSlzkT2m4Ku6deG3eDQ5aA43i0yLfFBho7ffdyh9dnq4v/i7YeKjD6nBYt5wZ
E2jJ3Vp9eZxsxk+61vuZFeg9gtBr4kX0Aj88Y1KCTq1E0wSu9M81RyFQUeyGxLJb301sqDRwiTUc
YFZheBSG0TUVdt6eJpIaTjewxmCcbsWPWXEOMdTF9KN2Y6tEUZLNKMmdF6f8Ctyeg6hJmFc1sWLk
g8Vc2wh8fDofatBUikYbS2dhHkpLm0bN35PieDEDrD1L4HY//Eah37pQrvOpPiMhbSk7BNhkOaWF
LD+6m51uWPjofru71BHHOhuG/aZegebznB6WF61O7423ao/QLzIaBpTSNecJJv01PmyDVckMDT0K
IugtJIcxAh8ff3ZA+I5gb1R86M7JFNTv+rJ5L/168hbUjobWqjKPZZ1ZaDGsnbEHndhJS9P3G0q4
5eUVRg+VILcHWAsHNfFXGX9FUlsXJguV3dqs6mVSx2fNxJeza5s9cppsXwjgrRFrwEGTsJPFvzhm
Du/GAR/ar4w+W9ji58f/EovcYSpmINp/adPmxoNVWiWRezX0OyvASpRIPxMXVxCG6Vl1nJ2INc43
X/V7EyyP9k6JKco9jOxaSiTGnBEN8lc1j1QGKYrp5sQpDY/W1wwQqQR1pcWWPtu5IAwxhgNCj+gN
o+phBAWu3M7spcKYGkfE2NWSgbiMuot1kzIpawNiwqoICyQm1kMHOmhXorU2vyeDmU+C740P+QMs
95Ssy+jb/CdmFr1VGH2Xm84EbhtZzj2mEOgDtahlGu1w9MkVFOkbiCEEIsvOdIMV1AdKcsWG2mJ5
8mgEL//XBBahi/q/XyiYpI0/KpjjGbUDP6FVhyzBh1P5UODjprQVRtnbgZulH+adssApBLr/i09D
SkvsOd4MfCErjFGGmtlj3FnA/5aJA83vEb0D0FVMMAexuNik0Qxu0cvLeddJYES7xW86Pcn74Saq
xljSP8BhaFVatikoO2ioDqbR+1JsTczloQ04Yf8+wNVnwpauF9sirYMaN6JkY0CtI+hHhKay3zD0
U5Ifquw5EXbQ8Gc+AylLwn4kyFJ9lV6E6cLMYb0fkP8EeO07jjv7R8IVDTf2SaqatqfNtMayx9aL
xXCD5hrKbHiSsrpnggRNSJNvOEboxzvxxazIqzeALCZhu6nLdpG5a71kmlOELgmiKiXGAqGtpo9a
O+Lxp6GWhomZleYyrebEWZqrfuxxBqoqQLLN8PPhHRQ/F+X7hWfTZsscKaFaNAIis1FCvZ5yAVuC
JRIqNNglDOX7q0NK8VWyZHB/PxAI/YZjR0H+0HFmNnrVGu4SzXuikzoivTnnHF/p/D19h70DreBh
9R8Qx0uSfxKFSe5H4STsqWtH4gI5KdtASvRfUOIVcm+s1yssNrz7TkMlvqu3tJNbEKw/KWGNYapD
gduTbhWisXzSst6Y96Ni5lHkfVQUCuqi5VylXK1FIEa6ibTIFzEXGARdVhCUBV58+0Dh9xrI8oXz
gUmNPQL5kbu8C+2g8VaT3UHSfFpI6YgUecK8/EwhqYhI31HZ6nocoDlA3ZBv0VvQRmV41foqe0w0
1apuMJKRl6m1m5ummr1sB/jJ5DEHEV78vqPl9aboo4ge9sk1U8lK+WaE9ZWfsdL8AzOcZVDTT5eo
AAekvRztcjRiY4IpPu3t36AwTKEZLiBDZtLcz7WFaZs4MOqb7kknf03p4cMwFdFXZhdISdLsrJ5r
unHg2OZvASHhNtHgCXkVxVdmVYC4o7ldLEOfrH2ULBwnu8wztQlEihHhhgM+3Lf3js5cvs18a44N
i3QPkeZofhjDyImaV9/mrqvhVfnddlbLK1UORh6ddlJMm1JXRCDKLuKhS27v+7OclQDh7gIV/+QP
Ko9nChsK1qLfWf5A3dfewWSPHiFmDNJibzhpkIYA56EVjr38D3xVXhc30tPjVMKKYvkK4HcdQFqE
4keftd+iuqrnwIOUsZJu12SOKCiiTcgFt8DpS462EcIlC+4Vbj1iWQ5sk4NgGMfVsoqn1b/syxFu
W0ONzyI2NgN4BAqOacfIxowe+yS7p27wm3KciWN0uBvc2qoS0k0+4fwB8Sc6HyoVi116oSuHOLiJ
8/3TNEUE01IhUHMwa1ZY7KzjwDpYfpB7WNbLG886W5DUUPd3dfqK/fsBRxq/txbATLlEslXm3knL
VU1FrkLzrPcR8RulavaiOJCC3zsNgPVcpsGmC/mHEe0Lk/pwUJpEEwDTQ1jNqtnc6zYZJW6YPUNC
HlIIx3tzI3TwS7I53awhKZx0u/R06vg77VUfVITqk+m9nnfhFvCMsvjqcX+DaXI+U3cb0scjHkph
jW2k8w2TvGJKduhwnzrWBPeOWwX3Suk+OlUOvZFp2ti+FmnXTbwL3arlFeE4YCKCTg3UOUg7M087
P8a+BDzlLISdtZOEwk5N5Z5YedvcRDbB8EK0J3sV4LEE/74JTW2WNSptYSqtVrT33D4c67TdpNFI
9I27WyS2ZVOwmezbPIsElNj2YL7x7GIIpIVn38BN+q2g5JZtUaX/U1OGGITIT06v9ZBCOn6tnFCm
aUvN2NrgGmqhHnx98EC9EtTLT7DzCmu0RQuYqKCFLhktIZ8Nj5NOP1Ufz0B1ZPbyGyI+QOtslOxz
pGwwOGE4NDMW3Cdg+gAa1MMjVNIDSO9PT/qrQqMiM/YH1+46732ovWwSv8Mb7j/cegFYPfNdosg2
WNWk/w/mjKn4gY4kDiYpfi+IC7zShqrwuh/1VhcY6LV9+YrQqi4FR/BGoGbQyNX41N7LfwF55ksH
6uUXtloDGOqM7yHO0Mjs8N+2nbcrdNZIYa09dB0GxZGQycmG31jp+Eq1F74xfMfFefQgDB5i2YLJ
FfvEAO1Z1ltumGSP02cQ+QgrS72cmEKTOBH2XCrjFn9PwzFkJb1EiyQ5X4+R1keC4w2+PPzcBlhY
q4LYq9HuvxXBbvp/KuJbSglrefjSPJ/4u8bcdaKD9WG4Xw4fZSrMGbhag0fS37OYreTbfMlLwd//
G9TJv71BMNaNz9Rhc+BXebZladFrkKIgS5gRvIOcp/yImUKMQIVdUsjKOjDhSe/XT6DXOK732Mb0
N7D+YJatI5eDC2nnbTf6jHIQ704w28bqIgtiKVhK9BvM5AEG3gRDhVPIqK7hVS3x2TnY23q8fVn2
MLz8HGCclboYXeoPVgguWXaIq7dvtFMiP154w4rIH0WjcAPhEZTSaoUDMdWVJUxGKcwhyWKuWMbN
51386SrX4F6t1lz005dwKgTRLb+/m7ws3Jout1/IBhBYUBHFyoKVEfZ3r4AyEewnmn8b47cVPo03
Rl328ILRqV/qS9fAMVOog5eC7NDKreg9UPIUbSJenDzWxCVmhgGuo0jw+LUfyv14pAasTpNduCWn
LLFJHwQ5mg6z0BJsOWvp2ZLjT571xS818xekmXKG2WUTHv34Usf37lv0sCoCtumdfDyKD8+7MrNq
sTc6kmLrTRjt4/WV6Mw1iGDGUwpvevd+D10BMXa1CrDGlBAKABedXSujyT1b66Sx8E6y2IJHK5YK
nG7IpIqFHgI5G+VJqCmJ3KI07G4QBt86K6DDTs7PeoIR95CbnhD67bNaUJuG7vdtBIDlW7NiGK1d
Qw59lAoCw9ptfgnry0VGfWMRNjW4hUlMFqgzQfY6rbh7t1jBHJZvrElwWMPa7BintpGlw8r+Pulr
JG/xttSkIelDd3JJ0tzL/slieP9lEx7WnXxndpH+0dhUSS8AoEzB2F9UVpHSSxJafNgmimzKo5Y+
vTrUpvgH+VvTWD6+7DBE2L9yqOcj0yo87gEDTMc6MAeI2A13PBk9L6O8kVf43IW7syLRMS+elbwj
BzBHPiERjrCWZtuxBSrrCXhu5AGerREUwPD+eOizb0oGRvjVKWQzx9WL/Cpm4dgizS2jZD+p9Ru1
+WMgXDOsOMA2Ssz0pe4fkBwqapQiuac7P8hoWGi7WaAAdNO6mK88J35Xa48lfIj867z/VZjlNsIe
sBZMozQ30/j3eOztufA/E44e7AXDVcZWRwa0IMxO913fn9avD09DoBCUrztmVBfzQ9gcfTDfNSkf
2ajsyV9kxo4JDnaGBnUVcBdGZ3C6jvZt9KkNLTV+KWESF66lOb1xcuRly1uai9ZviO+lWH/85UYM
RbwpPpYs0q7PVZOU0lJJo3dD7MY5aoAFyll3toYHDJ0hBIn5Ey4bPb8DRuiE8UFIaBQFxBqGjSRU
xpyE2QbmNHJ0cpAC5eQFBey74JKkYXbpUNZlQFM+xiORhzSoTRcQXTcvmEmc6VNsigmDL6qWTzk3
wpKBghM6U72glkkYS3KwZj4FZRWWfhIcN1j4/2+ACqTGbZxZ5tTyA6FE/G0RHIUPbP6LGqYeimXk
+1wyNeCtYjkOsopQO52sLlZGN81aXpSR/Otl3XMkpoWjUunHkSR1xfwpruhAMRMYlbsRGBtcrjmS
NoX/8dgMha4K3vvzzFjaWv0SjPtywbVhLJBIWF/pGeOi3mHPauuNJbjQ5WDw/F41xPFmMMVYJ997
zovQIwMtvHTK/G8qMF+FlGdmXZ/ExJKfE1VI2CeYk3uS6Zy7XbH5PpD1y3BT2XTipwnHAzTSqVjH
77eIB/nqHpTs6JcvuIjZfKv9Mi3jZIU8sq8ajtKMGzocLrm83z8TPNYwBw2Aq+BME0h2J6iEqddp
jA4wtaQbZCQNIVkTsKtc+gGPlxnRkhqGncy9r8bTPrFbphftXk5k3V2/o+vDKTnG/C7NFAsgmwDR
MexdLFd3U36/Pz8vcW2yFdzsxIFfjCoJOfhClCiXCeLXZ1NqOoOzFR+fKXbGw9RDyYG6bw9uMIcF
QyHooRmVxA1y0OxseWG3fAol1B7mJN9d6YqNUvYw1jwLAMU6Eu5t5CNSmtBvhvFpQeDG3+Tut6KL
c+m3m+xGIgF/xDzEjp5b1yITEwrl3cMnnlfJTf/4qaV/hvoJtC8seO13JeN3LKS4k4KeaMatOfip
p25LlJ1sLZYxQeQG89azKwOjYOMmlIkKM82MO0LwIzRAmnecaAvi1pARZwOcffW/oIFsKBtqnPBz
oCK5gkoxtb0LE7vSVp9XxuyKsS9OK99816kBRpdx8Mvyj6e8kuzw5jWGTS+PnZ3VjAzhz7c1nJNW
YyIAtIlbZ/9GDKkUimf9xSuUXV1N+xbWfoPMdU5S5fxzCx4LA7aGekA9hyLKocJC6p6/ondVlj85
bih+ljkts5eoxjmjLSIkJPmV7GjrAEK1VTF9M67/A8X42Oauu3sZAHtLEvBXjPmyF/d8JD5uXSjt
WPH64kyj7mXGo2apYEWYLB4l8bWgW6Iwa7FLqPTW/ptJ7BrMZskvDx4QmJGXAdXqp5ljCap3uOSy
wimzLI1Gdb6ay/ZNc5Spl+H5vUDocHrbGMGF+qLUfuuR8R/jeT6/KOZrG6NNMtHfPqunGfVhkQPr
FW4DkUKakuNACM21IoKAxFPgRuuhaN23paU7UJ1Qqt0UchT1x4mfQovdca/nFfO3zAg+UthK5uvY
6WzmBvXP/tGCS0uiwLZbog55DndTeRHg+43fANuFlXmfvrxyP1bRIX7Obx80d6uM2ik9RM2wY/gH
AbuXJnPQ7kQGP+T3L5qXRj2wU6yV5Qm3PIeVKpU6gxubM/84mL6YlhVszyT0n6MGEcPP2VqGpyQX
qaKbmVcRF33V57kXyRVQD+F7G820mo8HKnFkTrD5srywlOs3T6Iir7L0qWYpm+15nwdIRNAhUXVt
rJZP9RjZslx6+eryVYTzVrrktFNllwR/aJUMhvAEJEdU+gOIpPccl6xxIGq+A34mzDIfQyHEzTW6
eF9Ngokwv03eGBP9K6wt3R7FezcJqylxzCt1LO8nBRQO9W3j6amDDCWOH/JTwniv7GjppMCq5hoY
Fe8fdlfzJXv4XWfXNKHVpZ7tO/8OPg9DobXXrDGstTn7ZS/5Q0wCqF2w2ejI13Q8+ithxHnPxRDh
4r7I35L0i6BNe9qbRRC248Op9cJQENQMhsTI6fAt41i5c0xYKbMiIMAojB3mWm2P99vSLyzs0RBx
iexGK9mQWT5G4EiplBc+AX4oGbtWCDc+oQekw+BL1Jwtdp1RDWx51He50DQRpkltHBwL1KVGz+QA
S4mi098UsviSP/3U0cm8zjVz6XUo7YfWg16c3/zO9M5EilOPkqy/AaueB4sIQKenDz6vTMIzKmyI
VtNRfXvgNn7YNvWOqsxCAveuO4dYHv4ZPT5VLK88/3iXFZVgSjytb44heGU3TyGZSdPkPVCY1GzQ
tUI5Omk+n22xt1+bs4xYwYXTW6UOXv8XYpqeMqvamnzUusLTQgGH2/Geby4cLHBsysIjNnYEalzA
u0TcbsgsMqFmhoixPTagA76knU+CqewOUnv/sD51IsAW960QvtNmsALOEOQGW4Kwq0GF/bphut9T
+H3yN5kbc8Bp7hz13gkfwh366++Jid/UGoGYjEkdmr+3/4eppsB+ust2lntO4geCU0DtoNxWAzst
rIbBi4l6YrNBb0Sofny2PTQghCcpnI0e+eX5sZrOhspHuof8pUsL3nVIEl9C5PjLH+jiG6Jgflzw
JVNGZZjyD4EOgKTCjPKS1TnxyGF85dPLgnbwyoHIkXt+m6Bz2ok9ryrP8i31/5TuvBsbOKMZYj+E
3qr1NIF8hMhskzp1NhviWd0eeaQmFnR0U0bToHPLMYEhw+ZMWbA2RVzb7wPBnNVr5zk7TVfNtOFx
dxX9tb8P0VfiN7gJPbv47Fh2S/pU48LYCl+ElJY2pgFdz9xNCRAn3pCujd4avhemdb1toLby5aGA
u5YcrMmpm7/Gxlcg7VVbNSBj9Ry38ZppIiwKjMCCwsB0RajuNW5unw/k4IYFetaWQYBfdWEUv/e/
uw8pXfvlFchFWMgQGSGIvQ7hHeQ/yu/Mwij4SLKrmldekrn5Hxa0UovdLzSI2r9tDvBa+dOaH+tK
Slf+O3fHRTR+UwfjIBxRHjC8/0EdS7Z7GLoDNjwvRTLGFnbkMMmWFnBJ6iRbvzC73MRwlj96MnR2
67ftuop1IAXicsM+EK350vqzbwLU6LKl/wgXQgVUKJIOnWyo0CbS2HMOa6xtV/Pf75VDEdflQ52r
a5N+TKtHXw3FX2/hSi/eRqnp1DS6uqV29GrbsnN2E0GXwVcKENAJYfjYDNJ06uvhZtdzC5FgrzOj
/JdD8ZBdvdwz8DiZhlf9HrSBZs9h/cOR/2XALI+84m4SDd6VBPElQGxpcGQpwmMHktx3UWx3jpZP
l6bV5NiLIzKlr9HHLpDHXX6vVUijasQUF+srSfSaaR2DesZOgB/XAqVKnEwrcrpynkkrcdxtATTx
LzvPiFDQO4X2CH7Ua2X8qiBjpTMIIDxt21KRx2uldG0HDis2+AWifYYma3jf0L2vIdz9VuTAD5Z+
TU94t/4webG3qUjquTT8++YXutDpKA3jnrJ475ojQYmk+eYb7sMI7o8j9BZyvJcdrkGjiJPun3gF
yHmObjdCcc4WwNOYMogFJWIbTLlJPAvM3PdFlV6P/Vqr2mMcpyJ41eh7G1R5jxZeEGaEZc46k5wS
71R3Eqi1P6cWsiteTl7i71t9dehR46h3bAyMOMdSwBXAZdJXYSiZiPJCNMEKlV07BpDL2kp3thzI
HpRIHrDYOz8TOK2lPnfLEtJLw1CKRCzi40720zqK0g06E4pGtA7+MIhxgCV1T175ClbolQbw0WYl
iI3gP9zWCEn4sTdMvm4XxdIYq0OSfWaaIOZ7JBqLVInspvpo97iEXs/VxLjIERZAQDitXV8CocCc
Wo/7n/VpdG9y3clUjbJoHAuhI9v6EXwY8Ph2LP0kAK9jXFoXEL8ggYrm7UM7auZSg8RyOvtwBFSX
qb/Kc3NXrJoeEkw5t2Vp3ASd4jf8m8tP8Pw8k9HE7ln1T+Ia/ltu5PwAZXZDSTFSX4y5qlN91/Vu
zjk28jlPc3NbRi7872mmFL5jQy2oZvmUWBx/5hmTTqb1JIlPDySPRDwy+wMJq3Hyg9yrXvCjUV/U
9wykXqMvZg/BNNgJ6+Mdq8IpybefIxNRjOBF6McSOPKn4Mz8xjIAvYcd98LE+Rwi4Nb0V6YYOJYG
xHuQ0f1v6D2w/KIv5mZVzQOgTYkxZUX6+8CuxSL/321l0ouvgCMM+p/g6F/71UktswD/ULEAGvps
aVHxWCEsb4BWY7HbER9D1n6+2+5j2Xcs0hae6RrqUHaaHmJYaeds2okqpeH16QqNwImDDYe+Gt93
lS3eN7itCYZaB1w5Rz3ovpfRd/G0mEGJnRuxbybMNNmYOqu+kr8HGAy9wWmq76w/dN51U0q2Stv+
KT1JHZBftF+15d9PihKkVuNMghdf8TazLdd/VZITVEKcmGVrVDW5fgmP3yv9vdZZSdlTjShkPX/o
tE9UX0i7id3/IWCozAYFVqiIkO40mlXOfNus2jZ2wWREs5NJANxVTzaKKuJfe9ax6rAbqaf+kdqU
ta+Vi34cfHGN6DIKJLq3SO2hIR1lB5CczoETY/pp7xGmRfJHC0OQF27+SANaghvM/1dh9YPGnpgh
UkJlX0WZ2FD88R3bRsWuPHkngmk8MdpM4SCsgYGwFJE+FpKwN3CeQeNPFMi/2rkJtnv72DptlABr
v+L6GUb6U6iwkHji++qcZHVVKnsyjK0CqMCBjaNzXX2FlUX5IWtcLE6z9QoU4TbeVawEgLO2UYEZ
VhnJwjXkoJfVtql3VG+R0GByH3jMEuIhaDfcQDbwiX9YGvQtweWWqHFe0iGAUWB6Ua0g4SVKRL5+
C+rD02XnC+r5bavYy094fJOldB7NA59DnffDVIa+QVqQH2usMzO8Lnvj0aPZJQltSVBfvVdcuzhS
xHgFbiORefiLQOeOcujctCmwO+wJWG8aPBYFhQEgQGrMpttN8CzNtc11BSh9XQ61eVjUl0nYYP0x
WBFJjKGCyvHVroCnFNefAaq04sv6LDOWdXe5R7A0ZDs/BFIH0jj7y8NBw2ZFe9Qna8Eu1SccCRTe
tecCoJvXtXie+mB7jeGQLFpWSIsAxs3uCdKVdBXtqGDR3QlRWhlaLgoa90YJfpn4FVsX0lEcgoJ4
LFdM0219tlp+6qT8MReuTVwITJ7OWiC+f836cVnq3JvHoxvZgSMmVhqZLTgtyP5fk3660Pf2HvIK
nlgomWMQcPMQl4ZgjKYBYAXI6b0d/fodwRXG85MmCzQJ80+pOlBJ3o+KJyM4gN+x0ho3agIDY3nR
OeSb/SDd5xaxsUPwt44QWvHOl20CUCWQk6wyewDzsXf8kcnBkB4PxgUhbKmEf6ryx3tP39QabOIU
lJSpvrz3EpfsTOuVArK/ll0lJUL5RUiTM3uKmNtB2k4hf32WwFH+JW+M7FhIerJxTTIV3fDIj+iI
koY61Q3OeQ+/eCK6YugHi8QSCFgBSEeUZRzHYiewLLJo2sy/KbUTVFkyCxf/gzGiVBZhOW3fCy0R
oIaHHx+65VviBDIW2BwWITJWMseaVTl4wSB+UwDmHU67U6N/h9t+JBb1tyV419NeEzBGUkys8MCU
vCslfTtEV8B9ltvZKIx5CSib7fLkLRHZhJAGf9XBtvT5rU7Tm3gicVEFsb3nXVHsoxBauTM+9VIC
KMd/+wjMx5SJksdQjf6Y57uHZvcRJhZDVGX0adKPkuxxkhQ6EKIN7h9Xl5OXwa+iDJfOk4vcW4HJ
q6ZLhKh18ykczJBWHYb9aoR2rDSTB+GB/nlvM3iMmmdFErXIa3ywa+JDkDvSG4Idyxbke0tSwSbc
EnwYPeFLwqANt9sN0Hq/4YmZDp5gw6dCc+6nbbscWjGDAzLWDInHD24RgqGhyJZAdaKWiL30D9Dz
eFh3c4EMh/p3AUeRTO2aXoxvMFpWLg4raqy+02B7/DZ0srhdm3BGxMplP2Bx5ID6VtYy22tyHSXZ
pt/4V9CvK4vfvW+obgZgF8aa0lQQraQhzXgX3uzmGdg559OAa38W+yvhVBy5IHrYg9ZhZ7M18s0H
dqEIbxXc/9kCM5TVSP2RijfXm2Ktr7nEiANB5uJEpn30XYIeBAiViDBJht4XMkKvib/EfL3gv45r
xR794yYrFO3A+O0GGd2xY634e67ysVPYeMoIvUcrfTjSXMexI+neFGltusyJ05kE3XSknj6FQRYW
Hhvg5xUcvsbtpLnfYRMobUZu8N+bH2EPYZUJbpNV5befJkKi7JduZLui1GFdrz1LC3oo03p/YWyj
hCYwazMn+R3E6XiaX0hQ/0WtKeGQ3O6adYYqMsUSDVs26jn0sVB6xPyZS19+UWopFBCEP9AA3vtL
OixY3DeqRVR+lEWILwiiGLeRzQdpteh+D9MLMnEkgIlc319Pv6BQ2gQ7kNW58IQbnIJal7EgT5C2
f23LFlSJ9z7vymJJ0eqdV8kh+fLibjIFD2GiBm/jP1jCIdfgIVeKZg4kT/P9va+ym52SQdkwoV/e
Z4yoZsZneDeN2UZg08oP2JLtoCTAYQOOUz8A2KKt9CO4+saV6rcDm86Vde8QfT8kw/Hu+2cBF0y4
tcoLYmLfYGNe4j5ZbDpWPaXR6IDwxmoG0q2jgHsDoXfVbDRT07F+1uLM4A5ydp3N4um7FfKcGJMj
jX24D+xeIP7dHyl8Cwli8R9THBuz1aDw3rmGi9Q+9Z8Txow7OYNgYCYlEh+SbtDvcSSU/Sd1we9F
3Jql/rC0fZTTroN3pYzlr+WAr+aDZM9bskf+MjqR7mpHY7mBNXZWLYN04i1RIsPTUqV/8C7eMEe9
uEup9I2gqK2mOzvcjT6Z68ZG3BgQ2+OOGkE4VNAtBAN5TmSkh8SxxCOumgyvJoZ2HY804Nr368K4
+4RmF5PAbu2x8LpyIcDnAY5z+HgTGBHGjr4I4CEeQsx+i1EkBBajKOi3zHjMqcT4EGzF+qB2Ei2A
EAES9xuIxVNdmT1ZqoGkSGJkRiUU+1PYZZVdIq3Ca0Rj+x0ivODdl3w8kOqysVITsJE42Zq/LCeh
x+ZopbEGLefDFR+paQwPlNsWR6MvdMOQxwvJfJsm+cjlEOk9VMG9mWRY4XyCsKuK4Xx9NgDMMpTr
C8muUtUza6pUF0Pf49V3P3ERiCj51m0wn/q6mEhnE98MWkHgSDXreRhXeJF6GWceycUHMJ0JDMgN
r592aSlkm5xsKV5deeaHtJMtXoQo14e/JORL6yLBVa2sYb5V4J7bMLuAMntnzV+VfhAar/yJ8Lf8
kZHqg6bykK5szVu4KPBRdutknNLCiIy+wG22ZJyoZyJiz+CxkSjXBpVAhz9cKS6IvmrBtGzhRn90
Pq0xcbweicRjw582OJnFOs3DfGkfBNbxBjls2Ir4i3sPdxecC1gV1V+NdP/yRuG/TkhZb0WvvXok
OATFoRud/6rByCHtsAdqriqubazps8j4RPhkuGxNq4Rt8qOWSG5cXJStoJ4RpCcToLU5qNjegWGK
/b5T/S1FWxll9ZrF82WnWz09U8jkgvoJ+zuIYHn9ojpZalpAy90tjkyLaPc0XZWKY1pkgNf1cuXY
Av4rV5dAdSkZNNdLw8cGt/zcXVU9nui8uDSF8Se3NAdt/8glcuAlJ7FoIqS4a2ufwJkBtbO7kati
xHGDwyuCHriQdvXm40TMs/1o3xTa2bOB51kJ/6chynDLsuB3j7+dF1IW3DRabdhO9OImeFgDXuKP
aFyukj13pJsIwnCHNcMsKZip2P3WJcaGKlPYYfI2OVH/O98z4KAZhjJMkqultAhcv1iAC8GHGj1O
jgW8mwPk+NhTJiE1KcHgK+PIcKSRlN8iy4VkhI1zah2GLV1ozhF0Luw0W8GCk+JdMzBfPCIabcWc
awmixj8cEbJQBeGzAcTm9XgmjUCdh3WqTZz2M2JclnhZEL21KgEIlRbh20H9e3HZYRScoOUNGunF
5j/v6U8beQE87qZLG5l+09PIn5ZbD57ZjAgVosWcAGWz2RdTsjLIpC/fDYAZ5WjKnCsfdVKutTjh
mnzmN5vC0SgFoqQnnmPKUSSWOPbtl9oHay8Bf2IfmUCAyyECg32VBa3OQQFwwWi0Gh8fx0s8wSUY
eNnhQ7VvIBxc6gybWxNks4DdOlwYNZoE/4w4Oh9HtIJDySKxN6LYgpy1BdpFpY+oueEQEPhBs1Kg
zzgnFfZHWupZYZDNZAEAhfxiPBltzrsdSwSqfDAPPluwjTCP76YaBBzJnNrMSI1oXp3JT7CxrcjH
TgIY7ChiXSVsWlvKMBhcAHPItMM/XHqVsO4G1TFTHyAch+g9qLDyQulurWKik6fGoxt9JwIH7876
0koEHRujeMx5pywTDsOS12QHBGhewZZTZrNu60yKQqZmdMCSI4yamzEpdVSfo0Du2mOD+AUYZ1/0
j/vSp83Wb//oHYIKWHPGMErLETJr9GGyDYugfpBm9OnrAwGoyPBeiVolKPZPs5pLD+vzKGj6O5RH
e6QA1uSps5CnNLfB1cU12XG5iewNrhziKgqkpItbSkYcPNcXItlZpEb4Ei4aN8umnWF54chX08HN
bOLgkphiBTonNE1ijWXQSnljxtux2EKSjU2sCSnyre7zRrPV7jErhwe18HXbr1vFS4YGxHzsLQrG
Ny6d50ODLSyER5YnTnZXKofsqgpGQL7w6eFxpgvtZfJPAjUUg7ESfhM1Mo0qTuDuC7GTKXNy/WiY
JQsNyZGfn30c7iXMbeIpxS8GrrVmGccd4ZLXw5T+ilkbCWNWRIzPHUoH7niMY1r1yUXFU2vaTNfu
ELHm8Xa81zupfmtVBm2W731zqpCuelRrwlN0YuWakqBHyhPtctmR28PB7UE26JVq/UfDsC0k3E0G
7VpFzKbe9zJCozPEIRL3EZPzrwRNufHbGQ+ttLcUnDd1xHp4dbtp9k6A1/aeBOa2x5FXjU2GPsDF
yXW4iVOPY1nQPAbd6J+MvORiLRE+D6w3F0ha7x/L96sf/ICCeX0XXiJP2JOL5whCbYS/NI/s0A0s
nCtrplRi39e0Hf7nfrVhJleui+UUm4Mqa3mM5nqd61XWhCR3F5xixR64OlJJoKjdIRJg9IoDd2mI
DLMs7rNMQrHCA+qOEReUkjWM5xoZ9P8UerQ0pcreiLNiTO2Bk0cvc9PINPt8oEEg4EfmKHCjnrZI
87zU0gd9IxIT1U41g06ndy14XlaRwqlwZDA1YJ2SdwV8Q7/a9X4qzyiCoJAmYFnQ8qBJT+w6J+uw
oS2+U5BIpK8VVHNR+vNeD4/ISWPAeAigzhtBsanacwK6ydTB1xzfcxt6vveLgyo7zrFZjhueUHsO
2H6Ee5LCbUDMhfBIE2rxX8x60x/VYUrx4p8Xkq9M6VJBjWtupFNTo8pnAbz0K7RuIV9p5G0lILUh
zaDnzS9irSdW1sTyXJDvERdgeHoB0JZ8dVDFd3iamScX4yrd1mZ47ZslSHjuaU1X0wr8F0T1reZI
/QbgZe95rRkor45UuCvMmQ5KtI5HSgYd7BboGs45ZhnhUpBo9kjHa71qJ3fgYG7I+r3iiJLyZyon
7VvebkCjjGOqfJXD8s6RcraQzmVUydbaSLDInp8nlovZTPjaXRpb7c883nBiEeDfH10kAGAeHEzd
jjZ6qajWlDz+fh7AUcBThBaI0Mpn5M7ZpkJ9DIab6J3W5Vv0tVAgbUjImqMLh4gGZ9nAc6EGYShz
521KMv1ZtX3wCvJwOMJb2mR8f5RKQ988Z3eAqnfUfvxGZzHZffqi0xw7+wbyGyKCsuq6n+1fzE+u
faQbvAehzobbHGVa2/UGOBajUWA1iJsfioKYzWofS0I13B07MaEi97/HupBz0hDRDCSl5p5lAqEF
DDRbjcwunDS6keT2vsWknLrU4XDHxRV/5aA03E6X8+WFCVh9Eb5kFKd6ENfMjl009YFrnXKiM+4+
5Fzz/2wk3rYPXig5q8/biM7TLRs6/XGUxRUKnv7evZNXr7PwXfwk5njAszdYz4mYwTsfFzD48zOI
F0Di38ehzbqG+JC8cwuwRJwXv2SDUHZSuGpfvd9HxdEeCkBTBCT2+8pdzTjtiM/RaSda0AZ9nvEG
Sl5RoKNwOVNC847afLMSo4AOz2gk/IN53GbuNXWZHpUP/Dawz5vGxggkifZTsMU7ZecBuCSPhaLI
dJznuq91MX+PyPxEc+S91PfMDKfCRckq417rD0Mo00vJy493M884faUw8WVeZR/z2qvZf++2Lb4G
C+idjKDBG4Fp8UfhiMeMX0VLa9u4S5zH2qtNKCR0IfFnBjls1wpja4b4OTDkUU3TEBGQsHpxLWp+
L9kmM+inPPmnWAFk2nRLZUmj6VrHLqoJnOTwl2A0HCxHMKG9e/3wbsA9a9ZGS6pb5gfP4g7zwip5
CtG1W3qt7Y8OavoFLXhxLaI57yQ87ZTzFLp/z2Ub8G8EVgXVUw3wt1koYe4l2+nZgMVPl4Vwj6wW
tfvF9c/TLCWDSGC4xanxbLrSXjQa4bYk3nS5G32E8i1SCxhGjLTve05eL9s978rPqd6RbP+AeSuE
6GWWe9NbxzZolLZ0kAU2cSmJEHL/nBxGz2dyftJjelnwnKr69nJKus8iJL8/tVb2Fso0XOuJn4lc
YCPremorgIm+sqzgKz3CRVWqqtOxFceC6p6WMIIWL+6buV2O8DnMTJOCjiddsv0EpcJjVAeN4WpD
JtpgTNRFhdAOfrhYdNRZxch8703T9+k+njjsmjnGYkepeS4lk2mflmpRgK65S5DTIxJRjhytd6n7
Ft7iuWJRJs5UIeRMlqhWxPg6oXCV+4rfns4C2U6EpVPjpXUvTGhqG992EGnt7Ha6hdtKVwEw3JvP
THycDk92P2TigzDGDq3/NItAFChX381ijUQLMhBGFOIcV964Qy+V5NsPiW8cVabAi4tMHCgrbpQz
ZnngKZ7DvK5HTTWz0qgUx6HuEaDJJXc2Rk9GRHWP2IY5rNN/orYYMddVKN3PklqGAQXSt3hFoTne
Lr22RWcHUwQc8YMbPKxQslw8N8WiegYwUJwAmFy9Wt10uA9npRlcmxH5yct0wPLmwhkX/secGPpn
KwwKwXmaZdwn2DDEnPWSTXJfOU/zl2K59nHyyT259+BQRJbQJ5IC8Ce3vQjnuid4+GNlJcmMX5Yt
FM+d+wsMyIHGeV/ThY9cDFvWXob0aIkmkTEvZ+vfY9NrFj97GTQbQC8Gdr22konAkg8EmotZ/S3a
h8zQ32XgqU9U3BG+Zeji28xDzMGAd5O00wT09+ZQgSQgLUvddl7g43ZQ+AWAHACKk+ouzF6yFjs7
JZ+MJC/etXukR5YTRb9GtBp3SY95K3GEO2WIuKocj05aM4H8PnFcuMmflvUwALL/wl7iKT/txOME
XjNTF4JvKomT4RXURD8OI1tn5IOTuMy2nm3p7uBrGhoUU6BBSdbrv+YJb6wg00ubo3toX8mjhmpY
rmtT9t/2NaIwmEVZ+18I8kU3l30rIwmjE7+nrwmY5pVuV01q5bpIvKPyEposFiDlClsymNwH/VDf
+TGFc57xtSjmYdYCkIGX4V1+woYe/wGmPsEH5AMhDk/lct95z9Akn2aeMXEi1unL/xoJxJhRbHv2
h7TM3B4qmYixjyloXaQD9YHCSjBRLD5FY0wLVpQ/Qw+VNeC3lSVqlGuasG1d4ZH1jwCo2kTFkIWE
grDlQ5kaas5j5HxavDNOlHp3Ns9fz6mtzOE+GDz+3A1Q8wSdcgYV7TP2YaVI7puCNXz25ZMqj5Yz
Zq+gsh9y6IXKOgr/c3zMNuSaNILFkvN/c/pN/1a4W7hha2X3EGfgIr9xxFicgd29u5VAs2x/TAuT
WozEIfpx9kvR1wJkcffXs5L/ZvhAb+fJCRNOtgz3lLs1NIw2C2BTmZEP843Vfnr2NDla0/Ie9a41
8Kw9eTfbYFyRMPAx4GVnZKvo7283L5Qe7spZhW4u2u49Ge3v+u9ACQkk+32Oum8Je8RBM+kRDqBf
AtNCoH3xQxvq+4cZ8o+VSubVCiNdgbmmvlXbsJj1o8yZAbSYAK0Y5zklqsNDRMEPdG5bN+8LbXK3
DNZpHxY372HuvXidOIbwxRelpV72zbVwQFsLMnn6iqglanLeoCq3+4qwdoatWJmXl47jbGNBUUne
XUAnypa4CPDk47RgzHvsk5DLIvGr35Yc4yzl63QUEKFItOTL4oQC04bZkz5AMSIHsnwhbonTkyu+
Zr1Ujy7UQSz97O+GVTL2LEtgN8K2OzdLCcFwgErgjm6zYVWFQDPz4DBO0XNubVKKrn8wqDX17x13
gAp+P/XYkh8jaQ5Pmvfbq+KJzNc2yHN5owpu7TK9xLYxSqe3UQX1Oyh7cBKXnSBf/0RgF4cdeWpC
8AXqakHFAofhQA3zF9kreAirJZ1q/Qn2uI5sa5F73/kSLrSyqWBGWByvlAFrkaTn+FVEkhNZ4yf7
M09Se5JBOPEo7mRWykyc8DoyTwKHgGWslFUbtGLZPbGF5p/shayofg4FQIon2F3hsfIqjUeS+W2c
Un4VjkFr3Qj8nVdJkDNgzsEACqx9gIF8mubxIoOpazdfI9Jzvnedtmf6aCbdB8QDHFw1xApuS0hy
sb9MpdyKy2GSfP/in+ozTZ44M81X/12WO8tMGWfh1zy72B9CsEjSuaFgPV63aZ7aAfi/UxrEZC0B
5DmhkXddww3CL+XIEjHwbo+wpd/4yd1ilnazlH6oovOz2BnSxx/DrWF+OyjZlcc3FkdV6zgZHcOl
56BlUXVFQDeJTEUV05Pxkb/SqHYIsSGF+sQDkia5yB2NgjZs80wZ1NS42EkCGysq9F2/6110lccS
5PMkloAM4n8l0xMP+Y6KvyFKCuoo3mN4upBwbw/ufTO415k+N3rbBOh+w2vOip9T33BiCqtMrgvF
iuMHFoce1QOh0eWVkhawyhBiCzmLJAoKxqu6QU44rbYfFL9agL6X00ivTFiW3+JCrD6y0iWv3BwQ
4HEl5VJUsyQkYUZgeXYkzBHxCLN0ki+fxaxK4ZPUJBuRWMQZaRTjG5B94MTCMx9JqcafRkMbn5SP
C8VsCUinIqytWBI0aTTrnfIwno9hvke7kg3/ki1iVRQYTDzZ5YofWub8oDDWi4LElKBzuprr544Y
x/9B2sDDj+GgV/zKTgYPFJx0XWVTabB/FCJl192W9a8+MKSHsi4hGotLgw+uZPJnlx6Qbyj0G9iI
L1+VjqvKhv91FK37AsL8wy37Cbz09a03QO3ALv493SgQxShBY2pDT6maY7OiTO+RZmBVCccMGPdF
freTNdJZYL1dVUWjGihfeQHxKFl8OTJCi2rFCfgkfkTA70VaRBimV2eT5+Bq9ITnHi0PNl/0/hLK
aFG5mDCQw2PzUyQfJmHbXXbNa09065Zh9K5arO/FzPmXj5PJ7Uu5Ruia0YbuuWVMhesS5n2w8dyf
qItpO7JAsZ6mxiCbUUHJSzphOLRI/shwsR1eXwZQ4ODaYLdVTh5JVF8qyAt0Obi2bhL+y24hkJQt
sE/3E5WG0hX4xV6iS9mKE1pLhVYTnBJiW0v4T8tanZqNwbO748iNWfxDQieliC66dSx2zGCp7KQA
5uUELSNM+PmRmLHBK90ymhB1QDs7L/mcFsJ1VNL+niJ8oeAg1T75sYrDCBqkTik7gEWhQuYQXRp2
eKMNSZ0qaHABEtHCyfUUZ8cWwVqYavYkp6tQiyYQoz6546bJIklRE0zLd5ZbrT6gUM0v8FRmGNvI
GMwOkGLzbU9p+xbWurM8Sp4he12ahChrXrtwyVz+/f3Sou5dHBEPAbZPhC+i6af5LPDOENW6xzlb
IOOfTi9fJ/y+ESR/V+A/RP6VLLpO+/zqck0JYF7wt5sqrv5wNSdXBPaQOHSBVuJYdc8P5s4yStjE
k7dKUZ4CpNXu/10kW4D/8Qhxofg8J6o/MVeU72RBLl1wr9l6YPRKEcL+cvYIqU5tkyX48P/aWlLM
WAB/NVyfcSQKrwCoDSYwrjdr9kIXHC6ilMt/IC6zAIWkGK9h2xO3tnTD35gW4s0ahU5wPpf0+vLR
tBm2v3f1vqD9/hFB3tgIPb/eztURh1SphozUqrO/WRUl1aDX3PFspBi+WhJeXxw+5TWoioTDLM51
JTRqUlnGcoI2xltJsRPzk4VM0zIPkX9wj43MbErkuL32DPzu5ox5q8F4LcK1xYeFGtT63PjTappi
ypjrnIKZzjdur5/n8FiljoE1JgLvMpRoLVvo1OGCBrdnxOzdGuWue5+XzkrpwwBn0QqpLrHiRTEx
QU1K1/UUXz1WdsIQxELaUc7fUbcT5sDHrk7ZopycJichLDUVbA/oRlCiXmbh51Nag1pz5acZRNc3
buzmEbVGU3N0vPfFRIL4XC3jbyQoxs5JTJ5P6IdibeYWas1lBky4vr08ckE676wwMPR6rF3CEyjS
qwkZ6Qi7RGtEVRHwf19XJK18jwYeO7E2A+OC9iG+3qOt3gLHZmmeY0OeWlNv0wKYS8KGd13Prpds
RnxfpfeLJaFHqdmErIBoY8VxYvGeNSNzCUV+tXzDl2RMP1wQXa4mnL8OU6rjNlq8JYTKZU3YcdaT
0DhmNVADvG9JFsHLxNmcpWb+0KOnRsXJuK1SGZ24sha2LRdluk8fZ/RGXNL3DOZa+isk6PK/h1BL
ybnb0zVcXMi/1gluvT4MMB1M2zPZhh57FnNthIpyzK6tZAR1aEmOVOZ1zk9FO/YaDRTUhKl6FAi0
ZBFH3Diw4Rs5gdAoCb5mUSHgeG5chwKxubNjmRS3cvi01XwbZ9xgb8bo8s87fyx9R/eFtUeMn6+u
fboqfQcx9qdrx+VqA9RlodFeHHxXVHxyzb0tWLZNZTVyoNqm/wtYamR7qUt6A07jcaXV63XJz6Wl
OerlW8U0X9kdPVw5alonJciHHrggbecWcy0nuXvuajZhkftr9HchBSMeYbj5rugbm1pgZ4WVeP6v
SLkZEom/Qkk991000An3RfufTBhUZNoLEWgWzxqNnZCUp2W1JUiNqENa7TyEoDD64po3+7XCf01l
xbavspHoUhP4znop10Uk08F/AsG1MfDLSw2tpL8brxib3uyU/lucV2fdD8DgTvlJcaMYcfe138Sg
zxrumRbmw3ZUpTvFmjfEKbqCAZFBRPqNv96YfO9uYGIMmS4g29BusB/p/ZHOUYRKe+RqzTSlmS2z
41w6W9bRVFNDbgFkAHS5JCUWWejZOq+7R735GvrMQavKIfPWHxX+B3ExLHicrK5LoQ2piFoT18Gf
sCyF+T4f76/BPW0dcp+EPdFupoUfOaNnoOrUzeL/M30zhlR4JWuZumRgnYI4+qmUZTtMhIISlz7g
tmeC+7r/cyuLwbfzLn2375SFdvDaX1ToTWgwakjoScZiqL76RWG57rslAa7iuNbJCdFjrXVbqGcy
F2HgEXsttPfeYUTAYOqzyOm3/MJxcU3F6XJ0uwQaS6Lnr+FubEM0Kv3E36cubdw2kttV8ONkyA5q
pXJ+amjKdGv3XT4Gp/XWsi+xx8lf9nrD//TBNuAbfW9poS+CNkbQkwp8zsKB0Lq1k5qpmdP9ErTu
JKmaG2RaPYf+3Z0lm4Oc4QuT/iVF8Oz/tE0Yrb8iKJNcsAgFkCpb7TzUco0578sh0f90B5xAKYAV
H1HjY29cYhvGD/AHl4gAFTw5p2P1YMHiw7QEMm78TdIi8mmUerkIhEYfvkxfzXXVX1EPxqbfujfw
EkRLf6XUVnf8PLhkvIwn+o8n1b3wFDvupMojwo+GC7vFysJ3biyCrzM/K8sT8z65z/Ikm3M0UH98
nF3GYScTjiVzx9YTeblQ7QtkMczWCN3DXgmhlw55446/Bl6QRYyqjLddgapa6kDIL3ZTQ6hdyt0i
2cLZk5+FkeTj93o7VLDJKtwrkFBn5xRU6hjSW4EFIzDVkTPLp8m0rD/yoQo+Kfkf6iAzNvFlRMwb
bf3XVYQ1myvZE66fnyev/3/YK+xNb5Bk3r6rjeiIB8ReJ+JEnjz5ahLGqIgC18tqLd3p8Bgud6R4
CwbvzjNYB9GcgGVGSipE9D/qoYM+GNIQdk0sSVqauVkOTRuuo1a8rKF7zYOwxY6lV3g17qU+D0Jq
9rpSMn7ETR8SPIdoTyk/mZU2ft5S16ZeZp1LdilFyBiE0k2M21Fq2kLuoCVF0NAkLdwvtAdDfNzE
s+70KmNdIKflK7K+wbiV6hCabRbsI28GnKIE8RTzkrJeKLLZOWg3eV378jbIdZMSJaTZN0CQyWF/
mKX2YEuC+S/flfeEdoOjTNXpiP70Qf3vvJ9CRelBG4Zb1jLTLW7UHDbw/BbqjDaczEXdWY5l5lZ/
WpXEQh4JxQGEKvJ/sa4snJq3Djw2yjfZ0KQ4au+SOBvgkcc7W0/vUU04X4ZT1A5EpPGmdjhtRbUZ
md4+kTD7xLUSciPDlud6P9uivGzXi8pBQJWcmgjPBIiWddbh7olg469D6+2d8a4Ih0sUJpu59/gp
bFha5WWzDNyxqWkY4xZpna9ShN44UJ83J4hkyKrMNMI7OsfcFbvFl55pqU1MlLp0Sqt2exROhoVp
XP8JLD2y2zjP/129codHDfhleMglzt243NOYM8PNI32FjURWTOMPP027+Wi+9fbY+xzmNf8LDDUy
Gjtw/YPZBf0b7SYBk/wDfHitupmbZZ7pzWORbaqNfm4sl3oMTLjmaX/F999oFvpP/NQwGN+loATg
LCuv7M+RQtVvzmytxndogPfgHraqLuB1C+cdfOoTv20CxQ0/qaa/hUq9Q640U9T/Jj/rJV8YdNRd
tCX3hfzaoLVR3Nfoxz96j2YIo4TEm6fEeYyEJZGur7hKLFQSAeodUUJAaCi0GKPESCOZKQNnrlEc
8OPP4Kb4X6Nbk2XInhL+IDgnLc00q7/XnWNUu7+lLmR0CCsbdvLxeQg/v+9xfocQwa4LU3v3PkAA
SISOYDRE422ogaRoh+1srPKtNYoU3lvm68MlDl0ONITJBR1Fm2n/vxcPLBXr225Gil/0Jyz3ZrAO
+C5qA7pVNyJOVW7nznmz0Q/KvHC5CB7B+rkuXfXLI1s+upebYZXVqcCW29San4+YGLSZf2ltcRLe
JsWeEOkot4EWGcFviOxY8pii861G1rgeRWclf1QbJq/Q2GHbmtGqcco1dRzk13+zNxz2QVb98J4Y
UmHr2mnJlAssX+4vAUiroCypm82rUp/ZtDQy/IO78NPmIiL9EfqIu4zIZuDp7Y7ARbLV5lfQmsfm
wJ4qTcXhwvwR6rpZM0hSZDwpzz02/vFXVbGpiq7L13eTXX1JudqJI/seQan9piJ81KZFyfjIthCP
1+kLB92AYwRa+oA3OgW9N+nfEr7dt+aerWKk1kRPGXsns1THuDAEm0A/eTfee3RrHZJTBsRrVtQI
wTeqgW/cIMIiktXMKlPzCGkW1kquIeZidlOdAuLkZd4KXf4G3N4zYEVa1IDu/12yC6FBq45a/6rk
+AP5hACrtBAbH2FWxM/A0hJQxneV6i0RTnwQXM5nQK+rcuYZG0mtQnjj1jtkw7z7njbIB4mG8yKx
sJ45yZYpEPaH131AzmWYDCe2rMqGmmlrtR52IV0qHTJVM0k7A7jPyCy4E+XPtSjgxxaMEta2V0tE
JsT5fdHygxGjYrnTF7O66xqs3izcfNoPKCU09ax9StMLnQPxByerelhQpmM14PzqF62ufgV7DwB5
c7BwJ4L8nFQGU37ITOoX2n6q6nEKSgmbqsqeyeQWRCS+fCIrqGojfRB6CSaMiXFnwLY2BGZFZDeB
Qs4oMhhwusb1Y+wdHewux6gN/+RTeV+ENDnqwAF1xj88G20PMrg8aZ+X/exbSofYWNAmDHFnQj6b
/hbDggLSho1JPQ5XKCpyhyS1z30+ia3TGx/HmZaP8l5Z97KWBBArsjyBRH8evjSV0OFl0+IkwIL1
/EaSK7TRcGGlYB4dBUbBio0Oo0DD0dlR+4K8BZrtxAWEpt+haI3aXQkLtTUeOcokGq9iVPTR7YA8
lzUiBeqGwCQcubVWEjTkWisH6gbz0U58zDSCGL/0kWDKfbai0p81O7coixOSbYAAvR3qFaHwasOo
K5ig2QaBxpcC3qN82iLMQSk7EoXxq1rQ5FZaj8JSU0DexPLIseaDIDCoNN+SrxrIxzhXqbgfacJJ
z0JTg8VzLKxzHwTGWxsc3tnqJJ/VDBOHf3VmhwUW/UVgvTKrVw5DXiO6JAbZBG3FU1gxM/z7XY3Y
Xan0xe9QuMkmz2asTMklJ9aBkFSSS6MUgRdQfU/OdlgaefKrZG47zDcMpcUCZY5x1Xou6ymyeVGh
ejbh1t6R3Y4q2RjRKkbO0GSqGHM8uTNocsUBrEDXodVziG1Gtn4ZvVZW5nlSR1n8NlbiCV6hg3oX
ZN/Byl9KXC7dlnOyaj4yf+5ZyRtcKB1Ty4DRUNT4oJtq85rsez6NOgl/MdBxAsRsMuVRANwnJCwj
rDlZoNKtpIUDj1J8EmFcxRDxHt0NgsHa35cDOTK6BNMw/ujskeQ6/DX/VE3uzPopMSyqc3oBJ6fc
a6d+jOMi0xPvtqJ4hKyrb192QvicHJEJ9AC0Taq6/x05C5tyeGw/DiNJv6G4iqegcgjJg1wjMHnd
wcQKVSLIeyNcVxTL1Pw/tBtFwd08BVTBnsL85E3jFYH4XYcZlLPPigJx1dmKS+oPqMrWrmSulsQY
fgntCpIs4to/gnGrq0Ma+jd3G5yknoeA5FINizjN6t8otyjmFlGYE3DdEEiq/0g/ggYHipzwTvXR
4RDWtn5BTTrrLWJFzZxwcq/iX7z1DhzT621NGPJR1vvFW6aZ1a5IYZ38m/eW3ZZrOtKkvDNJ0u5A
hnldTW6B7rBks6vADwg5bQ7DSnlfr7zLRwoXEraPMFMt2TOI631WYTQ4Cf4Ow6t0puseDQEWZPpv
u6IP0gmV34TF8jdbopWMLQbKHXakt0wHx46vROWHXX52hQHlQAuMdvz3xp7ApnBCcD6V8b1ZCuHj
BiBh67irhEa7CvKXKdBgAnZ+uEpwwqdNxrwJKSzFCpx7rndoq+ifvCeT/d6EMvorDIWld1TSINFM
gqGmjhsotiO8CSCxGaWfXhM3bv4N5Lzu/pNZSEtgPW3L9fYGR11kApdPAp1IxJ/GcNFuNrw628M0
sb0heBfUhEPF1wqI4/egttF5A79aE60NNfThWEr8aM+w8P1aw0ReG/70part2nayM6t/m30r3jiW
Q0ognAzkk7Ir/Eeau7rqcik2GlqXYgRqLbkBeKB17KzAskW5xbgnV9NFFHsn54IR/5VppUOWe5Ke
6qiyiolcdrXnn1CPEuQnxMYEc4zJfSYXXLnwE4QWY4qTdMZ4EAYkuRXWf2vrcgsnzmA+Kp2l18uf
usYtDhDO1D3YbHRDu3LJpTcMkaKQpi8nAZsEmm1mgF5wCRANAPZ08pIdDZcFH0JnpDAEu+on9Agp
uhoxGuNuV1Jn2N5R+toNObDgvYUJl+hceEAIu2SqMYmiQlf2j8bY3IMApB1zmzkQgmz84d3umwA6
LQsetZJHnEWplpy4XZxrjqdfiS+uDKehRqDJN0w8tSAKqx7HzLYoHpjl3E4BEfdY7dSOr+C8XFjL
rO2YLpMjN/yZf8408eTSMPf8r8En5myU2zUGO5Vf8kA91HpMB1HrSWS4ivlIagRZUamxyP6mlYij
FqnoLjUAyCdw2LFsF9y3ffHt3ZWroTFNhYCR5QKR0A0iYX7KwPjJ4NdoPccXyds0n77Ayd+dHZDR
mjz70cp7qoCqlbPoGD1VfHji9WD2wCuIhs7iixgMyJz/BcwTZuyAL3JMZjJcgcgsj+kNdQQGvLOd
sJqYLInSoXaGkcDsDK3k9jMmfm0nDR5iuzZFClu/hxumI8TKq7DotdT7MpL6oE0NG7UvRv6W+Gl2
xOpmBx7yBYe/Y8/PwISfiLdMEN0H6BGYK6EQEsuXEEovU5SzwhXVEvHLyfHF4ETZvW/3q2hK27vG
zUjIaHMfMxcEF2ZbnOVBAI5QpiJnANNHqKjkhRhVIi0zMS1z02nI9tUB3Iab2YJpdU3HUcnLaY3g
6AuXuMPGuFJYG+Tu8fYqAOhyyywy4TT/NetWLdjs9uaiaYc08aa6OzBYX/i9tjYR49ylluEeGDD/
/fq2VItiLnh/kpZciLCbWz9dTgkRm1NMhUsitqg3ABQjhPTQ28sAOTs/yYtEwk8c5IdTd+Ofz757
GIeddn4BZ83BudUkdBK2oKV0zJG/PQP8Rt5j9T/gs0hFcj7Cje8kQMIAtQB1T0oBwbf8OqgjpVRm
DECfirOer946B5g7zETDXA78589ZElRQztSTO9DZ7VN2x09KU+1G3G56ZRuSVY0dnYwN9yvI+h4H
1noDkfhiYD3Kunmu6eAFK30OHDgt0fYWK7GkUy0uL6HfYJ6E/PZ12qbF+CVaYW4iE0j8uZLmJNOD
vK8wzx/d4i00xR3V00ygNZtzDjYKcUNpU+UMRL0hw7FF3Q1Q8d0NOwzL+WobxxRH07jaa+WMnhvr
LosnCM1lmdhhIUV/BKH2qm/4v/r8WHph6LyuUu0HYKxFA4ACwFNVdegUyQiOIql3ATzD7fyJEY1W
FKeUSkmx/hP6TV3enqckoNRAPhefnqfZ2O9cKa2cmNUsKPkRppN4Z76zM7uRfycZ+PTHmJq3LqmZ
Ep21bRw0mvjzCqNcmend3LzHswBcfUOMWlOuYwMpalaSnWyFht9Ga5zcxy76dMf1WJIrYlUDAyoN
poHJp0WCPouxoKw4huwW1axD2xjg/uln577Fz7EixRPQaO2Z2OY9IyP+2dzOJteEfNkfwHVI6eWQ
SKj42eMzFFBLpe2cjF0MliaeA8c0TydtddHqPn/7BtyVOZP8Vh3lU3D/1QJN0hLbSLyseh3cOTkf
k5MVFC+jC3Ck6m4FfqFVEye/CY8KEvH9QdICkJfZr0XlwcRqN2YF8BE0DYXttK0dhTkze7jdNP4c
B2FBDiUK6tryEWz6xgAbhFVmjtOPA9j15b3LC2eXjBAeANUi5AmhLS/lHsDp81pxSWigj+8NUZHX
gZihJCzBULNKglAOVNHxxsJngToYHRc9p6B9yhIhc3ovScymZstKnEXhGYaNZkx8IaOawgj+Iwqu
zQcJhwdeuNdxYZVcqYSJV0nQEpq4E6VzgrQBDmMglQS6LYLCozMhkfMFKNT229AFFZE/4AFSHEid
6PEj6wBENWqgp4XzDgkHhHKtdPKtQhnqdRH7kUu1QG5iRdaHEqeOWfVsiaqyt+m9ZO7j8EQ+zaf/
QDVOlnLTI9in7jV7mu9uQQouIbHHaAgu37qERj3iyC7MzCgEa1wzklVXxMNJ+AKeZYuwH35qEW+i
DVlB7DjdlhWbbGchRgedsOuPs6Kobpc/1gfK7GtYFw6R97rO7fkmI71U1Mp1UISIV/VchZqFX8KA
dosvCpkmnhHKph3QhLG2rZugclsbmB+V6sKK00EOcM/7zpkayH+CKKlvYjv/mo7a5XMBnuTPAAzc
xYdqk5Ju2EGD9s4uXETaVED6wptFIgxSpWPeyFH0SzaH7PoLW+OSLnZhc0pPAfIG96Du0PZDdFBG
sTHAnB0UWtLKmkEM98sOpHeSVCuvmANO2FuzJ5uFLMA/zyLuubkeuK+NJmYzRQomNs5ZlWduqlbM
FKvvvMFWMr5m3qwy9elcQ0j6kfLmRGnPZ2pT1VwhQpxgZ1vRtJrHqL78hL83W7X0moeh4D4aRC4I
Y+s1QvyPLZfjsvyDTSxcqknAOhly9TxNAd6m5rqtz4w0HORyltTO4Gw07AMtYSbGNnspn51wma5+
hNsWMSbXRrcfUB7Xane1p6bsdcbm3kXQXrikM+JMuwKxUOUjVPjRZS8Ghv9JfkccCSp/bI79XeB4
6WaFHrb2pz8AwI/UBc+c5ZYwSvroYYycwaeCb2V62NcfburKUrbNu7YJ4J0/4TGgG6H3poUMngnB
evR1MfpzK75zBOdmw8cVS1Qfyh+FPCRUZ7FR6dInvuPycQ3qmrDAs1Z+ii3sTAfpheGKVoJ/xWw0
6xh8WKuKxf1FSpzlMRpprnSLWI2xDCf0Q+DlTyoVQplak/Zv3hc+OoiorTON7Xp4p/jGEseYfF/U
DtQhJaDzsXjIgaeIw0tYxExZ8ND/WhNeXXeH6HeM5O9NR48W1sF4O+JQQ5EoY/EJKqC8usF9ZMOX
koiGyV2ok8OWQAGMsU5EdBIViUMPYwNcRaGPLIpZQ6kS1JzzQOU81a48gEfpRGRbGgGu3GaLl2b6
1/GqNOMtn0/YOhp4DlFEn0l8DXo4FNdWztew5yWNidHReDGvNcy3QgdYEXnG0HRyQUVSJ41sGGRH
VGEVHyDvalZHhEoT3aJadBT0RXLmRuiri6ZaX7QW/k1QnwvphqUi6aSWYHKZo063cFwls2kegcAZ
c3G3sv+3GNV/5sNfpP3dxTxV6/n3MDaclX6137XoMHT6zjqT0ygGHvjL5VawkMJYYONwMm6DKE/9
C2cnZZLCyEc3rk1XjOuW8+EJza2PECfHu1kosvBOSWfKkmNXilA6lSvYh6TWOckyt560bN/GVKBA
gbblJD+6Pqe3s9SuKgvmzY2YqgcQgOsxclUmO8IJRIn2O3OYj1bjOwEd/0VDR0BEzkB7u7h2JwxY
OSRHTvneTYz3pPVvK0x2Rzf0CPvmjCPC+aRVxZjJYRs/XnGRvcRVekBqZF7ZKqHlbQybXcg5Il78
gCnZBJYPjjxIREYANzux5EL05l8tt0kzOBh4fSgMf34rc2qvknUI3SzG346WGDlk1YeMFjUrWITC
eaC77JJUVKJ1/yYkfbkW2KOpJ91ujClFh3cJEqzxFssLQTWehQZHHVdU6GGFiUkPAM6TWAv+Ldra
sou3lqPz8TPCjBJhqSwV8XkZyal722dxQHivO5/aJKnaZHPACm0IynHv99otcpoQMpggP3srtHBn
JTFSlgfJw4Prsq3K10I8wUHcFNO2BMtvO5liCQl1UrpC0K+xKD4j9Z9GmMTxJxAIVeqAki0RkbbU
v9XcXxW60+lNGCCQxCqnSltr1PyqNhZ5b9YVJnylA0SiEuAJTQdh9pJtVrmAGUJeBOkS5WdF9KF8
AOY3pKfz3daTtOB47SkuRXOq4zlXtYuPcCOAm4iMPYcnhRqCu0CBleXm6ztgPcFKAAe2oQylMrjW
brJp8hp2P85j2bNvzl6oymhGP0Mhxj1sMpy5XlbNFOmYR8SHLiQkMNJ/ONw3q7HasmeprWGGqmOK
Ac+lXNgBcN0FjfEhnGI8acDfC3XX9w6gXIh5K1yE/L1GZy47ZWHcTPd62oppbLIgj9dFZe8j0Oso
yMiFwM+cx6yJZOf4/pD4LlSIrU4vDI36AZM0L0zrEGYGQzXXg3oLI2bttbsCmuf5+5PPXRmpKI9n
wzwhOS7DpQRKk194lz0laJ6ab52YPwCUvlTC6ZLua27p9vTfR1JYe9/l2m2NK7b57bcfddiZ2i3g
ISpins6HRbdNIh8zJhONrxRkEdAL8JzFhwYWLipETw9j1SCqc8UMHw9v2mECf9Akt7k6c+K2Ucwo
cGxSZ+D3VxL/Bmds29gD52ZivI/LFvgFD0K+0GKlmXcvMN59YEm1GGQlAzd+p7HLR8kbjzrqlYhr
HINwonjE0NZ0oLtDd/Eh/D4N/mxK5ppEVUdK6kYkUbwWyUAa8Dp9ESZrtoRK8facBYtSVFgNnCZm
RA5/Gk+b/uut7jnhMKLrpZ8CXnQm7Y6VUt2EtcQ4kmb0CF2NiRPO25Ao56Pt6TKhZB2fkva7zqKU
4osU7j5nzK3aJIVOxmeY8NpagmKL2ULEweAg96dL8Gt3DK4YgCT1adjUfRyfWAbSOEn8JypU//hR
DwVrzUhe6ye8KzSpZJzNRehPiYbUMNbvpTG827j2pJ3zBiCEruPZ2kqI72RHz1yax97K5t7uIpqG
K7+8k4CSN9yJ+UxcZ036u6ex4Y0YI+T+WTGC3oBNO9v0ri0VARy6thDXaFo30spBeRPJcJDMUnKR
7DPdjfxq53o8Q6korfcINJw4ceZzeFGOP0ObpeGoAb/ZndPGta4nk6Czi4+6o3nTILvnedjdrst/
DlRWXn+wHLA09tpjjTulYptjFtLGQckLaukrtMy4m4ALPG2uMHnt4haYxBL6UDvNANATPFysF7lJ
MfVVrq1GiEuD97ORgRlzT04JixBzZ/GIoJ+t3GVN9AoZh9Ckh6QnpdVwAxJIO+umQnuzVlmv/mlj
QABk96iH9hLvHcrW8hw7AdBqRO8KZZNI7MuXzyirOacXhf0V3mgx9SJjhEYE67rLc8Iz+KB9EcxR
2sW3jwLMEKPVi6B/qWNOull28XHBS/s47kMVRaH80ouu3GGDPBwwnWp+JdaRn+ifhTXyuQsJBdP8
DxRiabneDrLGRgbkZUswyZ9C5Ya+/ND+/2DQEnRC1wXXoKSkR/TVxfgTq57cPcoEvK7KE+Ri7VE9
HjReHY+mA5w3tMjGpLqNtw31bmoBonW34MqmSPkZOblprPzzlSrMozR9pbrkGCRNLIwFvRIORhE+
2jFSqeLsOqbjFPyMfssmNRHMKKYX6uCPlpzhQDYZWfbKep31HPREe3v3rJ2GnosDQqABDH1FY5r1
YPLNdX3uaK5aC04NMf1sFSSwlwRkrkKIznbgAfQZ2QjqeQ5SdnU2E/MC0sQyUEeO+/Py9mJZW7ep
0FofaJ19cVlq80NU1N029I3Y5w9IOxWhD438N4wz/SRwH7DOv29YW742974Ptt1ik3CQhx5SN8NC
1T4HiV3H8l81faxGFKoye7susTdkstD+/hbzu/xoCAcQ0c4BzCAcRlECjShDGLib+b0Hdotku3p3
PJdjN/RJmk9Bl5H12dPtnyDRmH/ERfWMCePZF8hPWaBYM3QWSvKvqtmLqcyfRlo/1BsZrQ9WO2KK
eDL04YB8/F0GAnX6YyEPuyLdjCdpK6PnNDz4N8+GLx6ZeX2YQY/EcMKUVjOcRkKq+5cEbR4dyYfD
NSH13Q2c3SpGe6Un8AEtYkaogDAFnft7NFMAvDsrsE+P5B2UNfnKXJFnMjCCz+gkdIAkIBhe/IAF
zJ9lwgoSRz4hBCaDQjt4XUPqQPsCleKMLLfTWYBfAUSo9+9uvtliqKMnMWV5lq9gW0szzEJVLCeG
Zcu8u90c8YraJ6ZH4CuXlJItJhXVEwc/5RI7hlLgO2mruc79NMzSd0zSRxIUP7T32X6/hX0/ccPW
466FOMDZakhsREiFRj5IBQ3Ge1KjjDXODYwfyFosXN5MTjIKrkiOwG3eRYZ4cN+L8CuOX6VR4xXM
rvXyNHt9tnoA/f7PqzibAuTnM2cuZbl/ucWJM1MXPI92vIJiprpSnAZOAgGkEpNBIhTu0erYAEW6
jzcET8i6/Vcy7FXGY2tIRzSWpeOEy0hEv5LP6vrVDao5ramvAJdOoHJByYg725rgzaSIWJx8Zbej
R+8TRQUXLGWblL8evnZZnX/tIFuI+myT2NWLYCzrjc38HxTZRy8yZfpaj31E3WtDM8cS1/7d9unv
9pHXGOlZvsbMarwdGWFhjn3t+a8nywmq+z5yHLEPefyx7Ok0Mv2gV0inPq6PbFXNzr3TMgq4fo+r
+TB5JuzBOwOC3o1Y4W8AUL8+pbB34sKgfNqQyirRjdHdeHpqxQbO1KU4z1jwMEPMA5sgkahw1FH3
JrWMNpgBYNmoqQl9qVJcdQdVsD5k/46Z7MA2UAK4IfGEcT1F10kDUJ2YwTO4jbLysVcbdlt91YWh
uixhMpwTylca1lDq5xIDnsDy5OZdMn4eif5DkTjGSJUIvg4YmZj0X+H4m34VLr3Qnt9YoJZf7AgD
wxd+Sxt7N8j3WLGSL7LvHAaQX4p7gcgxj4DS4z/VCCI5XN3ri88152mQFFpp3UHJMLuoQ8mUPHWX
xiZgWibval0nUKBp2hKOn4VDrTWvRyEjPRyfeDD/h1wo3w7060jX6vePiFvB08jXVnweJRTya5EO
7maJrmqK8kt39XSXjx8EYVQYlGLnnDRwaIOmE4I8YmaNmWKIy5WW+dYYXc0Lq2K/2SikelncOWdm
Q8yfakVpA25e71r3BO3Boe5fW7Cqp3M6UbwL/ZV9//yNbcPGage2IXmu9j9N/Y/C7kqztmS3KC36
DfVt+4wUcMBzqZI42t3bgnoZcO914DdsDvtqGCZDWXdzejwymz46ZQhQi1PP0m6WYpHEe6v7cb8y
X9KC22+2+PsjyU+n8glrHqkGUSMlDWcvvo/x6UC7aBamop/InF9+6tnGO15iw9dX2+ak3s+FTwWI
7EwgAXs5wwjVg+98M6Zoh114ATk2kD8Ikq5mAQCw8EDdhU3fHwuLTuSMeF3U6tRXGqpGkAlbjBn2
FBMSsHEImZw2VWPFUJSqokxwVzYRQNfunrc9sKuhs0tbCEa+cn8eJE4nXH2r0Af7KIIhdDyLGGFt
N/ZsGDVOvMDO6tM4q0n7FrRdtFK7aftUs+knC79yU00okRmvJODhn2GZeXVhcTAPt0GaeCUH3XjT
/Bop9qLYMAii3T/FkPB4HozQ70OmNk03V8CzyeFVgNuEFikn9kKCOabaRxJrwrmwouN8pSihd+7z
X/Sy+jJQDY3nyU7bR6x2h0L3OzJRJ4eh03+1CCYNvbBa5Fy06sRvSTNu3r3Pnutu4ZgIBb745ht3
C+A92njQ7UjyQI6wPlWL3sBYUQUYbjqScG9XwBxIIDayDFt6HmZXakPIWbwKktRc6tKSFvLSBfus
8pGuQVuNvBGk9jlQADpA3nUY+UEgD19RK4gxPkOaM2WCthgN6z1xiQ5u3l2TlrHjXBTIrzfbPXER
S+pB1WqM6cSrRytr+FFpILTtMy5bK7HKVhUU62+b1/nIn+lULnYBrCtn4JPL7rxOaokB8Ra9D7pU
gxpwe1A8QzCWFW4Uw3Jwz1UVJmVWAxBg/tLzhrTnpY8LvRzNl1ub5QuysuMYB3avjkOuPr7Yun5Y
7hHiQYo3JUrjm3ZbKk2eD7f6JZUtpdxQcTR92wbLJpxf9vwVUr5UxtruIifQCQy9VhDf24nLuSTw
a3l6qQLQyPHJ2GIbtsWnTuGfFDGqgbBSb9Fc5raIY+aZxoBocMd/W8pyruAdIQTJol1NxYfSC+k6
czVMIf9ImQEdxwbPddgxpLeLQysDiHU6vksQ+j2WE4XKAgd58sokWgolgqUxdBACEnXIhAKO7tYg
hyRlJgNVENhk4EQnnRjGrZz8N2Dt/+ajTim6yuZZBLgRNXrYqxW5TrioBKS2rea8uCvbQCYq97vK
WiY+nqwxXasUkyxlC7wHjIIYAR0UzIkLoSjzmBsTREEW0ccOsjBhVQrNCyvJV4Xls/UVfWcWa7/r
U8DJPaSUFlpzXppcP9TK7tl0pFJPg8BVSNV3Z89IsLA6Vcqrat5G7MV8BPPunhGnCoJBGRSkxmGj
P5kjvIOypwaWd+OI/mE17sUsLjBybmEHBw2twQA26wBXz46QfkchKt2lfvJk6I35G+r6DNdxMuGq
bja/bHaGEbG+H1DxW3RVfSvMzfnJ5RUQ1RiCdMeNWTT3o37koBapltdj3sid1DHUs8lKFVUmIrEh
lPN52bKHhRa0lkObRkkI1eWc1WRIxPgN5JAKlUHj4QgzTT+dG2wuj64X3RtBnc2z9DU2aP0WkRgQ
Xi9ZUdmwOj9xDAkQ/3CrfcRxiHeoiXPxNj/sUwgHmT4fbF5fm0udD3IYsObhBF32GWbhE31hd0yI
v5QAp9TFVvfI1z6xhUnBW+6itNIjd2O/PK+4ZOBcxy0MryrPSF+KAGS9YiEFPtNrD31ITuZ79Uqg
noN+j5r7xuzw3+OlEPIc7/OCwznY816kZg6RKMuCYvfVxzs6uOYcmKHud3hsXPbdvnrmHjNp23Ty
FrgOLN1LmRaxGZo0oZ62IcfPgEdrrrgu+T/CpJb7pRwFZKnPifkCqyAGehyNrt2/czLZHGUgspSR
RYrADOKw5Sf/YwrQqIN5N44HqFFjAPPgcK4gNJiGDk+RBlavOw10agOguQHS6hU4gET1FDWAZxET
A+psYPMWytx9NN0gXNhJJiZyVofoWQ73evwSnLcx131vMFcWVt8Kzbu/kQ/4kP6w2JOWUu7Dd1eT
pksC7l0tYCS5MJPHR8+UCNmibOPlXby5xRvHA3r9lijF5ziCDcmuVZETU8UxkO0OwhlcgOfGSpoO
Xhk4Puq9PlvynI9CNTatZ8q0nIHkzg2x6pYBAXM74vdKhcAlGhDc5VIo7Uihb/rUkICZE832Gbh4
pHpWLtYFMmEdzvxxRQ2FpMt8XA403H6PV5Ta3W/CHZnRBYu69n4qqrtfaaSShXPg/fA40urNCgIh
b/RRZhsn/1eh29j9Rzw36NtpSgp/kV0Fip2eFQLPFJeq+a7PCahl8BTUwYAN6ZuFt4nG5+yaw1os
m3jYdkI35tbKHX6VCv9L6Yr4w6rTAKILOz/INO/d/tfQ0A9KS3mOD2o+dmQGhkVjGsyPC6bbdWHf
XUSyyVcQzYpr7D5UcAALbXV9PJKGFz0VguI/G1C0Xndmtw1RJQzqqelisIlIpZ9Wm7F/qTxjAGmF
MVFe2UQKpELTSs8W6cgvcSKfaqScNB/xFHVGfxqieVK4UkMP3Ohp8w8o2EqH6j8x49jXudlfPdec
vgYiaaekrnNgfolZhHd3OJ05/GmsBZffJ5pZgWWYB3pr+zsy0Nc5+vmSXTMfwaxo0CPSTJFAjddx
bTZ1uULNtx1WimQSMuSt38oKdtEJCGgTWCdC2LqzVU8E1x6gI6WRmJfqqcVxix0Z96L1GP8NRosn
HDZXqfQpXpwtrMP2S91Yetvk2Ssd5A+etwoMq+lZrxTpUwPkKX5PRDbCZAw1eKqiJ5Omjt/AUgI3
12UNQDYDTiZd3AdqBdphiOaGD3RLcNzwPSQYWOwU0YjdUH8NE2fupqrYX7oH49lFgtQUDO3sLMGv
gEZcPATHNbBqWF7av3KTMIu5UmIwScqWlBE0chPVofd5FH5d/08liBdrkP5REMXhoPoQvl18MN47
1QHpjIHnn0dnVIhZ7cbESOHCXqJGK8CVe29aslpTXAIn4gRbGls5HqfRhiwUjOoRJ5G8BazQeD7v
e368grjaQV4VUixYK8wWdUQC6ZhDkvqoEcM458q4musJpY0t3CO9I1dRfRCNJUF8aGY5UZI31cNl
0p7VWN+FIdsSu9PvL1Y/7UUvkdKvQaS4uRWb/EU09RX8dnT6GLtVryD8jbISvl87bwWV8fDpyP5M
lwUgC2hDsIhjS7+i/93MrE1cRflpHpR1K1ayLRBW+8Jdh/sfscjlFiKpBQNvCEk8krqu7Jv6f6tS
nzqk21JVBm3Fq6LoI2VIqHHSHUHOVvLpyl3TYOL34guefDR66T1noTXOrjSme6DxqNjXyPMcBCso
mQvG+fdZiz0WfsGmv2DNmC4AIu7V3QXj3B13EDdCvsSFTZP5KHVPiApw5CEIHxQITRYRONx8SQf/
i1oc7rL6ldUlvWEw71zzwKwCRtYDd2gZP+DPAqEzxO2JmAFynF2vdsXzCZODCKvOrXEQZMvTTmj6
rXJvMa8Vpnnwf27eVGw3LqQMIlqUYlaxJrQiY/Xhkuu4YOS2JzVSMgxx+SJnulwZf7IhclDviErT
5JTYpRpQcgiLaLntJNYonDglAMMTexvfFknOWfctkNGAc/phDEMctfP3LyZ7vZFFFYZzsbNgCju5
C+sNAy7/C9b9JftlfAga3M1MymyGpeTusFoBUEbtKzIjXaBVY/6gFBjZ9qnKEJxPf3qR2WY0YIWh
PPYLpBeaAiybzGoEvDxGvVwUQ6H0IRlX9kHbsXlTKnKdlZzqwaV+w+9fglzCr3jqTBkbaltg9CMe
CjrRsE2noE1uwZ4JCsMoTiSDsTrfxLNiB1fg43dDIlv/QI1hbOjYV+CCKDX4mEObBOVjptKoHMFK
Hv208lyhCqda9SD9Og4xVbPC26lh8Q9KF6aal9NXfgsn3o1a4DQsmSGOux/EGZDZNWX5gBRwXgV1
KcLB2pveFea9GINruo3qzNIR4oW64qzQOlLqBdBuOcoUToH+z/3Es7z0D3h99ZHfidm1VQB+0K4O
MwT5JwQFF2J8EX5wjDEPkYoW6dA649CS5aYfIeHISv1FzHwMp4GdCD5LhfagUCsMc3Gr3k2jzqf9
CERlDQwQzSUdKaAYaxTLgBjPGCvPceU+Hqpa8G0jmrlfJts/H3z/P+CTQgFRtp2G+7O/c142qqj1
XigSx3zNo3LJkf9u6sP/ZFwAI51t8FNmyitiR8Wu3AuKvzskjT0qx48+muK/hU8Q/qptO71MOpr7
DnS+fwrOHKuapiWUIWcZVG7OlqAN5ypxwFyKlx0xN569E7CwaeUO6Zp+oNaarGIfkUQgAbTKa1n3
CTQHEH1D6TQaTfCQtVh82Nkkg33F4SOsefLQGrZ4BeDMExqSMTwiebtC6ncOAr24hpPKFCv0FdZj
MikZpnBhH0o6voQA6fnhAnwHrAN/t1bhEEKT9wWdBm6sc5L0UlAHlXNXl1FqCV3cYAIS9xnqu0wO
/h2SaWg/E3AnepAYQz8gIdvrQhuLOpcakhk+nr0MzNZG5CpNYlHO4aEwiGA9Htl4pS6sMdra19Bc
tIz41nS5IzE4P4VOmIBb4IKKarRPWOmt3xE61A8+QPbx2pk9tkjEJ47VR04OCQQatsdIA3+Aa4Bt
PF/zlHL4+pYGAgzQQomjkhERZ8kCkdeWCOGpHnr6StmHmjM2cuIxaOMmQhKiWJe0/GawP08XEYlS
NmuTroBJ0dAOMWBgBGtLRKPeY9XvcWYAqpipnX6MOB+U800Uc2OEhFeOlHWhbt/HDlTGDNDauzsJ
gCJE8F+t3ZqHwGWayEUdIHZeVc1Mdw4cuyktKUcG4nUSMgucSY3CwyFQzOAy+56lEKeslDQg/j5W
mZGe+Hre+PcsMiGwccDLteHZ6vPvb44znrvY9YS7oqBnP2qbHFqsZIuKLDe3nW78G7fced7lOVZQ
3HsdycKZulTfmVkFUTLo88B4iJJvs4YMviGDzOWBCRomrrbU6cFfFhbUB4MwkDtOXLaevuoJE/Go
+aTBnwmYIHueIU0oSU4gWj/AG46o/ZfI/5nOhqL/C+4Qvm5SWv2w3MstTcjwKaOJShD2MDOP78el
7VoyhS9Adv9p/Kdl9s56lQzSp8WvIONqx/BtrpLeQDp50WvlAYzv6gM4N8DG9TP6ekWyiu24nltr
M5cLWh8ATLJGWL/ucIBk4Cs/bxDRl0HP4CwrVX0mNr2Vo10yIbVhYewxKPZiISpgfhSqo9Hf9i4D
Wo9W0JPua5Hfr7GK7WedTZTXh2I4ZoN80PqpfMyX78VuqngIFOgt47JnYkU/PA9nqLmC7IZWJC0n
2AeM4nXYIMEL4imdXxnugKPT1NL1nwuoWuFvfvBdfmfqy9spnWoaxp6i51lbPD8OqxhVrZRa9rvz
I/zp0WcNbJUpP4CRRB6fCfQnQ7ltvRRguSsttBccIabmt9Riy3OOlrfSRWMQkHwSPqLNGDxeTA6q
nrUcp6q8pIXGdFNXQy5kp20FfHq1Z+0Tzm8mmdGuX2OOMEPtmKClrHqCI0N+SYRT34cCQkA9OYEK
orX3PUCLkzUigGVl+HRN0fHAhj1JzHBfrnhudwqhqA50d9ADm4qygrNCb7u3jwwCe8D/rB+0Y4E6
HdqS9xZ7o/QKbYbM78NdB7LD13lerZqjDuUKt0GG5JJx1KiBxwE4H3eaFqHByK2s6+LmwhSTzGHG
Lcrie16w0/TgMVMn3x0zpi8UNEFwhektU8/fI6Gt9KA1R6aDvh1jmhdz0OV1h9S694J53BRDCyOf
0NQtJX0ofviwbgKljfQrXxX34OuDciX9+Ol5NukswrFOcOZbYiF6vamRT3F9QozzgJtS69Hx/8L/
TchqRYQsPLtSMbFsM9Pl8i1ZiWqyF9clJa6t2mMy2qz7+ZcRPgeYruNL8M92/bHinUfrGPHulsIh
8oM5JIO2bMSAdVwVDO/GcaFTSPcIYpwjbCqK7m1eox0k0vO+8Gye2CxSvPkDVTxIODpnNpwuyrCi
rfNhbjTj3NQI3Vf2lBfTlsyKlEv1sTRpWe0Z4fILJFtw9MXLN2C5FlgvZw62TChNa4rj84syur1T
LlGmqMFb7cB3bBtjjtGar2+Zo9SoQBo2DUYB7lOCbQq32c9byETFSIdjinyfBy+DMWGdSSRNpmD3
1xhBCmOYxj2SFHP8y/eI8e6Xkwb+90tcTbkQpQPTAs91LIuVQ3EBFFTSUVUNs+iCTDEZfL3yQXYB
HQ2R2G9V/JYqArKoeghZz/K6w3xwo8NUULf440EpYql2cuMPp1vRnm1fYfXGxN3t86I+Dg34eiqI
JrH9pHUGKR3KDiiRdCTacGomU4bxx1JztnTHtHLSxOS52EEdAgeEFMk0pjkhmHymyuVMXLxsACzk
SPNhyrmOsNtSyHEi/wd7b4fQ5nqNMGDNBpaTvu+mkpiov+nbJxVT0bdOmOCQjflZF/e54foZFjaM
EcVt6mFQFUc2JIsC3KdV6LwDklbWnKMYq3sczyFXEpeShpz5PJJ3oi+pj3n5W/rtM8WfeXsdjjl4
Rr+FV51iZZhSBOee0/4J9JOd+ubfO+xQGw8w6kf/yXHq+0kTKp4jwjGjVCr0twrznr28zxtqcsEA
HL2gj7jWkEBLEsIFvFwgiKbzLIwsLofaXBhaXsIr9JDVjigoupycH4dHvp+NiZhJdvKEhaqWmZ/w
lBNVuuSw2tYuuUD0TcSBsbVvycDg4V9UqXByCXOcUEXJo2oTzbR1ZmcFDro6gzbv1nTwaXfuUg1Z
fBXPEO7OT0D3Q3dcLSRtHAa3N5vVJStMM/32aL1tNoghTyLivafkqbMqfFQaMM6oXbNPpL0FnhP0
YBlMNncfzW/GPFurp8S9G22C2qSkuMuws/7nlRtjEK5NsFBqbZwkuF8ATg8fZrO197GS+kYhumvz
gqn52v4XGt7hwvMGox5aOmgmRVShcLNSBagr8nlAj63+5DRcRx7M+UG5YMfE46jeuq3brs0OFJaz
8VjCw7vSE0cAWDTYcQHwWz/ERlOt5awz7mESK4rBiiIbtOHj259S2NBSgXLb0yvoeCnyvd/Dj7JL
fg8SYWvb7hTllrhadXIi7JeW9H4i49+BIhYZL43XA+mWnFFAGPe+T5BZQjG79chGDNuL9kAkqbdv
i7RTj/EvPBuWC4GVnJu1It0EjiF5sfzM1TpDjyzD9A4VZ3hPkOjILB+cVpH/tap5hbDdK43DhI73
aFao68Msf4f64x88Wif03Pm9yL3GSqvUaQMvtaU48K7NCy7Z3bsvDdHImDAdpVQz8RNCtyyZlJyn
fHBQBjIvH/QqM7g1dTWtZhhczqhb7S47EQq3UuGHRgS/aheBC3qs0U3onyptDsryMRDbrTGe2n/V
iiqCKDcN9OFiQwCjYYUKodrh9TU00YSva4Fx4qcoiBUQ0H9GvkAaqqO31C/7+Jv0epMTUZpBmUh0
Dmo1faV/k60i7OQ41UX+fhoAFPGMaZVpLAgdr1lCbPO4DchxES7MvdL/RIX7A8nppqt492Lbe8E8
fDg6pIV/m4bxv4OMtQPrLZ6QZYERVFNZswM4yWjF1rrfQ1UDIwDUES8jaw7IYsS5GQRol6LVzkK6
RFozjj4MxGx5e5G81LxTFmh6gJf/eMxeFSabN404bzFSh6G3tdMkLXHcZwD8ZK3nRqvKK6vKO3vg
7+9p3eezYgU6wvpuX4MTdpATtTlmt8xiZaBKSwYTnsEXT9P+zopV3kOCXdOwo45ChXXRheuSl4no
iuy+CMhjz2TwMiwJqa4Gc7EhvtdBeilckr9vpKVlUavJgmTEqafMzf+0pbQ0Fw6DDi/pr1ApQeFa
UKl+us/hlJ1dM+5t65ij6cTRljgkym++0MVnZqW5X9VmuJTkUz/pYpyOAHILk8Eg7g3W5K704DLE
NlEBtn3K/9riwCB8ynA8tWXzA77MXj0ZZaHUDb4NKBJzJFHKdcvwjVHXWRKLyVcXn4uz2TOl38/Z
D7PHivOv4+L6IEeVy7Z1h1PT/w1pp+T+SZb7dqHS+iU+slWl/xBw2z8hJQnoVFKelWTp5pISaATj
qR4kp8Vtk1j8dd1CR3N8xdqDaSb7jxC46BHfc5Pe+lgzKhpoYZLBatmEQgGLQra2+blNkkSZGAgD
Hl+6YUCQhvFGyR4BOMoF2cam/JFaYN8JPzQ5vW8GGUO09dpCl3RBPqgk1B3UfDtJP8B/zpU1pQHa
dXDYNQw2zxQweacihaIqx3YBB7yuvI/a/KT9JNYZ4QVyTzIFHfRMOf1mav8riQNdYN4ZeiHVF0DZ
TyC+pfYmIBAXH8BEP4MJVZLaiwECx6j4cBzOzI095HUb9GtgpPORJ9hmfC7gvsyFb3whf1e+fnSC
qpu5VH8kFY6domsV3NXwfCfBUEtPOObEe6fVmPg0RN79pFDIMUEiN8qqxk3S79w7Me3fn0g0zOen
cup1UfNL7CsA6tJBlNhroRiK8kklZ9Udtay7zLN8/ySAOXGsmDWYPqXnViZbjJrcswmAJRZ8gNsN
HqRDXycYeqhrEAx1nFpxSS2aPeY+3fhDJLgyIOLmpY8DKEiXjon56unjvVewxKyO9lmAl+WDciEn
LE6jdyaSPha9tl1f97VrKaL0JNJL0JBnZQltklgDdVPGz7GbN6BPULj0iCBx3xEOB/zOSr+iwsi6
QUrznBjNWiK+HvZybmYll9f45vEd1mB3Ae8DFkVRIAeGRafAxUv+KIHdLu8TxjaHYe1vdJ91mkq4
1RV6e5/O2UHFaHLSuoFyobRG66byfE16DlHuIF3i1FHIGvkmGkwEEpj08fIydp4l7MhivevjxrFg
lrPygkLRe7V/S/TE2TsPg1SWbV5kLpigCoY6joHIr43KE55aNqdcLW7XEvYsbO6TOwdsBWWDsyjQ
7/k6zfIL2HnG01cW5TqPKRV/uJgPsgSqISFK3eaJ88wNDY/wVhfgSYwBqrChlS/bq/BF1yQbBys/
pBWIGzazY+q6MsBxvgOqloKF3iIGNNqPbJr+EwH+OcBWEQBeSMf8RicJJLI7kbPeyDGrDlEI1blj
Ek5yXGZAe4jOU74sbSyVQogbooAep3cV7SEGJ2DpmhAbsNGv78UVio7h/yPAp55LljG+XY46y9NU
6dfRm2KIBa/ped1XnSN+l6ACohSZv+0eiobTELfNakxtCO1IPmMr0nlGr6CuvVt3JYLUy/trxinG
9UUMRcm3uGbFOqw7Ah6sFBY6Kcek171SSG3a/Cdz+gu8GcWyhC7K8P938w9Ct6UDLiRWJiUUCm2T
0xDbXmuzp+xZB4tjS1igU8WfObt8K76GY2B1EKkF3xz5XrKOk+4Q4OjWJ97rPSTRJo949tC903Oi
nNXDBCFeTbL5UmowtVh6ychJvmFpRKk5+o9vAo14Me9R7quRqpQqAX3/zF76GbFApO4MT9wqnFd7
/ziZkZ9484Pr8m7s4CLUQIDuFVDEIm4mOMUVYRPv/LHbls5VwdnHHgG7X1/Y50AYs4o8w6yuvOID
uqdPPve+GYRH8y3D2bzxgN+fxAG0+vXo6O+S2kfMnHIojMISkagRoNMMnYTJkT5Zp94yD7WVDreX
zE5rxdQabQSO7tOYN1NEIor+u5kqdElESZn4Cm5MfEH4SqJA+hhrudOxllh9klo2Mkb3UKbedgBN
C9zgdJOk45L4/P4J0NZP9S4urLtd1Ujw9LxHdeHCyyWd7spPwIWu/aJQLOjSDVaqNwWwkgjmHfsb
Erk3udHOjd3QDATnxSR6dGnEjPSFYvLTxLrojpB3dnMSp6dNrNRj7X4EQYEDiVvkw67OH9x3ysL1
xk6UvkJ6RJmP/JHGix5SUHUT5M95uAZ9NlhdqUTi1ZsQMwT7B9CXyScGOrNo2jjkcqRnm3v4hr0a
VTN+chWqAGcpdBbzMkj2VKcqrK9vDvcIf8j6leKYWr9mCZ+w4nn+MH72r3lGhJUrES81Vkac4A2H
IwaBTw4pRoB4+gYbGEiBKFbbrDgkdlWz337P6pheWJNxsVYFNs/RK/aI03uRPPaHDCaGZE0w9JSM
0d/Wcy4L3Tca8T0IzfSMEQLXv2KmIaB/hVi2fGuJ/x9T+58lw+zCpNMy3tPvQ0Vm5tc5QiiDDiKe
3osIedE5jmTjBisEAuUnwLWzvgdZjAuiFq34dKIQSuy38j6cpSP6Sw9VSBktSk/Kc3/7JZNpXNSo
uAbo6HQsaG6zi4q2isrjV1zRwuISW4DIGiuXZaAlyQrN13gh41SAO/HX8JEHhJ/8WXREdzwhPKZ+
pfPMMYhtTnHnp/b8EcYLEzUHbZHxfs5SL/BerKFGXb96fZfHeimOvrR99E4bKvVgWaX1zNsB5RuK
O3x8s3XPXLaCbb0CSs1VKbc0Fp4oj8oMBdhDL58Zf20mW0IffZvJjTBfxhxnDajGLjMH9AENM44P
PFQ5dsAs/dNLEsQYuXW8+Q2pwbnTlSb2YESzxPl61X1NyruiX9Car03DR9l0HSRcoFNhbLGTTM84
P9FpWtAR0NkYJWZh2rkEAEIF/GGXX2eE4VqhCtPv66caRe94npxWp9LmNQU/19wYofpKzXZoQ18v
Lin3K6P4B8YJDCvGuBtApnz+/aQ3GAl/wzFtVVeqiJu12/goE8QhKUKEBR5tJLmCQ26UhiUE13ZY
qULPv9sWoQHD5zG4CtkoLUylmvgKB1lnIgLXG3Sc+iV1qW+Wt8Sh28TwoJ5XYFytvn5aW1iIAHoy
IufIlinWnkZzncJihyH/1pvuSkaKBeGfa7yP35likl7x3kV+e6Do0+z86QqVJTXNSRP3eFXdcgfZ
ri/495bS5ZlZEZC2ev6EE/8tFObR++QscwIU640FrXLUAanN5Vh9OhdyZNoHNu+4Q6N21AHOuDWl
tvJLNa0vQDB/WHKxc3SoMoXfg/leH4UR8m3CnmHQ4laMq5fW7mRcBXEBnCdT7DqKKYD5BuwlyHxv
i6y44iD70Y7fEfZL+CsJI3AG2w+Qh7XWKeOjyDVdqiMp0Cax6RX04Q8yBX8PmVPOmy6sRXS33giI
zRNW5qjQ57fxFoPd6RiXWeoiY3BzB6MDe2+IzAIETu0GGiVI6pyNC89NByXpeIPRZWUZy5BC+7YO
0lTVgtClEzjMUKVBsr9JpIKkBFFiuRssQqOo2ZxvUTvrfHZHHqaX+2BOYXDffKMcKbUMfy8mgcVA
gJx1oLj5E2Eke9hUVPypYXyTVwaEoi0p5nP3vSMwHuIno00Ubk607aUKG7ok37ByAwKCSeqcv08Y
Yt9g4KeKfLBZe2CvKXtE0k7INaoFXnuKNqpRJgC1OyWwcLyqlvXqxTXvumOLn7sa/MDSEs2sFKg+
4oPJjD9/eZigU/GWcncrlgtNhWim6PWRC4mze1F8ySlWmITTVas25uzrI3tmb7IQeDTtQl/WTTu9
iFicea9qwpPytALIX3LQGYu9sK0hP9duSsi3Wj3qTPaqoqb3QwuPryD5AnYZQ7ST0K/Ma4xHTGji
pMezMfHnRyLon2LjgNiAAKN0tvh+KEdG04qMHxLXj7uKsQPMmNrTQW3GemkZE7tcltePocsnfgQv
gdZlXlITKp9rCPB574Fi3Yt7XqeKaY53rZEW0sVyUqwji4MZVgdWfeobVWAa4MPyHVs1OAuPcAFP
rf+96xTunqd1k/dR7Y37/dyktB7IoxVN9RqKbYq7nAbzlZbaX/AAmD/kFDepiTHi5qTet0dRjXK2
SpR/Lzag/id7I2oJ9eCvMKVTagoZPvoaWTRlZsCnuzueyPNRyeXOl4wEKlSBW5wCUA84yLQzDEdV
F4WRqnttdyC0NuyOTpx9rWkbAMPmghb1i3ls30johhtTTx7dz0Jb8eGqGhC227Fwpqfsqo16VpCO
tIjy+spJtDvrNDNnx0JHQ6BPqr4sr4SxAjVoGb5heEqmbUU//CAGqxuAo4MOKdJE8gik+vMlkLZ/
SNLL/20BBk0YSlRU80yh396Nq1B4IFGTUa92jx7V0NtHO0VKMFSitBifCPA4CWlIlSGT5UGGr6OQ
XGL+FAT9JVeIJdnLRRjThpYLVXDVGSl6kAAsGc331wcwuAZjtQ1F4VNZJNMllD5McyNc7ojHkdTY
gF3Sbrz74GKgoEiRk3l3v1c5GAFO8UDwRs+yeKbUry8WaM71XlFlPsu7WhUbGvSCj0v8ioJIwWBt
yP4fcdi8rFwC2rUY8FIA5zyNoQswlH5iOl0HZmdTiTXFsUNZbVnekb8WXl3cEpRemr0MfuO9Uhyx
KQPnn5gxClro/KGFhvxU7vl70e/b7Ri1YdTQ9k5s4DJ54aZxIJNP5mdE2kZ/NSxwixULsxJz7alQ
Ewj2VndFwLbGHiQgQ+VvFNlRHNVS68Ev/9hil8ESLXT2OlBh/s6k4Ib/H7utAX59CJ4U1BurQOrb
LU7+WxHpWI0kmTERtodCwjkvLQa8067wx02YFSDOZkfJ99ZtZ7jSWLcU07N502LF86xKhn4jjdk+
UvAaNuJBPxWVRPgIcmjcJZHobX930Eu/8InIaKuDMf2++q4NNIfBmUfyzGrTrsjLQEYwlxCSPhkw
TccpgGyleKqRluRdSeRZnC6IHxrIh3nJjhOqU0KF/ejphrx/NgY9fSa8cXjuuFGzpnsSA3hjHWEb
RLqGw9eWXn6rGBb/HayOQWWB2kYf3v61+eclU6ycuJITUc9TyHopLkO68wwQ2eypd9NOO8s//5j1
8UyiZqdVlmkH5KLS+AcraTPtAEjyrbMAOkEqhJlAEFyhGa9DNo9gCaaf9dm9KV7DRr5k1xAE4HVZ
hRNKPtK24FpPOYtALmmZyd20dNSzMlrLqjn9S6UNB4fZ48mp8YXTFASpg/Lb5xxAwYAQeB247Jzo
GBifM3B5GfldkQqgabS5qiFloy7c+mLvJuaGNqjkpHhlBpZxQLx81QcTWHdrTs7m5rtWC4spfs32
x3pLj6Z9LwB8YfETCHzMrXkoxoFMUTC9H/o3F4S95pqwgtagw8TIM2MnKFqVDcJS3G4Erv4416d/
i0bo2JBX4cm8iuv3vGg+ACDqq8suA1d44DAH3IGK6vywXBKL16JDapqUUcuN/yzO1tiqaJyn2UND
oVqcyZLveS/Ynro3f2uv06uMKOOfpjucz7h1aOkk720QcnN7Ya9xC6Z1rCOkTqRJ78T0XRryKY1F
ZPR9EL3HX5LX4sgngTk846c0I956GH48r/VCzhOwy9WmyBP/ArjKXQXS8HSGOvsT+sZHa/Yg7I1I
0/aktEla372aXqkyle6AUso45GjV2SocJlygtjXGfxrgQU8nf4PQhnZKxkRN/IMkNU5LEmkF92TX
D8bbuZdKGOpJx1NBFrxcV3aQM6g3ea/xGIETmCXFNcKZ7ASJVY1T/S4QLGFDLa8vQbP3+cmhWhIX
aoQye6V8R7ocxpiWKsMznel65S3Bd0C7unpQvPV2d+o+azOcE9UjRrcJJPFCLc77izhOlzknihW/
Jx46l54mXj7Btt2hCQVRFwLyKLHEftlW24l2GGLaDXhcsiDreot8zOr58aH+JetVf9qqn7sk20yG
dbxsWXX63+8XthmciH8eG16pQbL5Kp1u0PjDVbdhIMF4wITaZo1n79Y+kJmwOgLRj61PpyqCpzeG
ireOuX80i4rMJXT4U1uKJu8SUHEmww8tZKMDtKfxRSFktwXozsAU85pLJP7rfdtOnbkJ79bhW4au
1b3GoC4+2Ph0AOv+zI3YjxRQhg/bNY4HjytCMW9w99QQSd4V3PGQZ65FPHyRMZyC66OD+sgvE8ht
qvMTMzSZ5WA1FEpsGwYfywuKo1Ba6d3XTuXQmzaQQG4aNnfjsVDFe6TaB+UuoYVRCOweL9Zk0ibp
UQaPeyMeV8/+tQvxYU0ZipPKUjycDJbNzp4cqAx7sU7ZZC8q0i8Q2wo0zAWRBw2aWwupUAoNY6w/
2DHYpSux3EhabL8dz48vludvaaDcvSEzzPQxbH4RN0CLSus2Oit4n9oBr8Zkl9fmLv4AVZArhnh9
epVkVhEkktr/1ehjDGV7M28CNRVdkKTakLqaZDOwSLvZQX7QkDucryZN81wEvK5Y6gH5aQ8NFOo8
bMNTAsK0BC7bAemGEkM+VCutdm8sFf5ncyNJWsHfEB7EYVX2vsdOrm+GSnQmfckyxKUjUnNztWvw
SdDYz1VmsY7zMacSBOHAB3nMnO9IIaDKeOxOKf7+WjnuGQFGP/M5UwXSNacRRXelLxa9yiAnOmjO
IDeMmL5rc/4r1x4kBTadFBH1ioDqzDIDdg8Dws1qS+4ixdDnkceUtKRfn0HwR4UTgEHREqN85MoH
XW/+gdPvaMtcxLYzAFMXv9v31A/2yifKvDTmrFh2NxTVO+0jWiwtLGicLoODdu07G3JJxg4XIOpN
UU7HtTA85tTa+pIi5Tfb470i7X1d3Wk2Bjw2m5luuPaD7HZ7daQaAjiMbrYleLRDEZkb4nFCvCGa
NcMTFH0umiPjqkOZ8TAtBli52gd8iXcMZYJlEJ6cmk6hMnza/3CARmB+nszVn5RHSNHX7iZFIsvB
Z/HoFGfY4IZyC8t8PgC0EutniXVO8rG5ENzrM9e+MrVY2RXs6NRkWOWbUcsFlFQiQQSOGulxZa5Y
CTMVLJb/Xkp+o/RzvoSLeYz11Hd1CIGiWWdy5Tr+S2y9QxAjFhRKZv4l9RFM2rysAn6px59riEVm
tThymRCj/fRDcnEeD0WTHvs5r7lCQ/P1oOM9rnWMp6zo5ua7/oScJVYPm3LoC+XGW1AHFwrUK7JV
b3E6PvZO3SCZKoI8Kpxrmfhggcmcp8+F19srFSxO26SwcHhXE85FObwjA89tdg7+NUzo/E5ESxnc
Dc+/0a563MJWvihSGoSXVVCVyRhkBtn3st9NiybNuw6s1ATseEFqxYDvb9u35c0eIloRRL8AApmj
4+Wjp3DzWaDc7CQuM0q+IxywhmrKsqDhXfZ+e0Opp+WuvcjOeLZRAUjhM5+JiAvre/26hZ80qVxL
U/anvZfh1ad2kOvJUp0n1D/kJEEQq9kVg+DpO1jqVsKbOS3XkpQzMx9UaQCYONkYwFf26TyN9hI6
JJp/IwwYgmXdtDrMxBwa3shhSn3a9NQsWxejxRh2O89itIVxvtaMmk9ziObq4Ucmtuxy/yNY7oLD
/Wmaf3wM/+O8RG2hEFp7KCkr2m7YAz0yxXT3bCdUx8NbZLCEvm/cVuaF18oBhBsKN9jGI5oLCokb
HA9d3KlU8UzSFa6k8t1x0PxXPvqZqZO/JXTRaiy/cAxVjHMcdDX4HXi3vEVvn1CPIYXIgwYkZHYC
UfYV29hqxP4iMsuuKq+0zoWlH574Ln+xzi6epxW3JVB9SK4Fivrl38fEyiXcjNczC1+YpqdpVOQ0
2AjHvVwpFQV2pAiHLwB9oQuKPdBBPahrkPBwh314dANzSQd5G4JFkPfdN4mmBwJwak7qI/PXZl3R
478pS+G76IFyUXB3u8WS4GQ/88SFPMTz/EGfnyvKmCVptVNC26nwZHIdfUM8+R45FIdq6ylBqWeq
yCn0RNo6uRz1XgHPkEnf/3/LwlIkcQt3hIirRKd9HFpo3sRQsLDAZcfp5g9TZ1LzHbqtNwG9lWbg
gPX2dLVT1GDG+5iI/BHOvkXDgCBGXKh9uDOb5Tk0MxsZc4XFdgmyKWyygAPT7BkbDH4kt6rQ/Jow
fAwdCQUn3q1jqrufwVpduEU9hDASli2sAT+MbgR87hewtwF7NBpK7+GFCUeMo33/lJdFre8gYjqb
XcnyC60VmZloc6InoGecTyy59AW2gpBtm5cSMvhKrOyYvP0RbH86tsObfrNALnMTLCIZU9Nxp0Tn
35eiKmoSQ7vlCs4NIp+7YinbLKM8kPVEJz7cxplxSoB5Cn2fr+sQPb3nIcTqWYrzH+hrPCKb7hs/
f6oqAshDu+grCIXG3sIFD+piYkhJjOBZSh6+bJTuUJzgmRVsD7RRWhuJnEy1aLu4mzXb1mzJFcmE
r8NZUsa1M4yolO2OkmTBJlhicnhvGdz5cGrcH4dtWSUqOf1GcQbDVR7ADjSCkj/yG9JU7tGMVUkx
RyjpcP+luhI1AdmugrZ/YxnI92DqXiecn8Mg/W4ajDPw7lK6QDGT/vHdhDwUOmdpvM1mNLb0sDR1
PGYJQyzY2rAYwQ3zIQfjtTaTrQKni9p5G43pFaRl47fgtONk2x0bphaKgXugUdCh2/Aif2ohWITn
oOqPozSRqUufY4HmC7rYEAXOuM2tEnB4XxW/MOHP8ceiWWPmRPrak74xtzQOa1CJWyULm3NcSxjP
I3+6yFd7V0rUqF2sECPkcE8ZLo9O0sQZ7fTQSKXCuHB3CB1dJ2LCmuBtuq1Dc18YyUgvnxcc4dDB
h1oiJhOSgjTDbjmb+00rgM2wN1Kw0Z01EX2Yzv5lw1ofVvX0E/q+WAbt4Ekhhz8BwsmVxpFb5pbz
IbqcW46bOvGTN27KLNEKIDUopN4P+S2WRGzSkkOo++40AKgBOM2l7catGh5IDbPhnOVchovYSfjl
hTEErUL5hhhKBr/zWeTNHCOXN4DNndreEjqf7BFaDXgzdJn1BTyB5RwfQvVe8Di924rp2teAqDd8
TjwuLmw5JKQXa8cZVCK+DpZ4v1NPb0QUsHbY6fmmaiO3yMDOThs1lekZQv1YXquIOliqT6gXNhoA
RjzaUrAQWhdbHtUNSJtaRJOOc49o0ITntE2jWhHCN1roCDlNe0236j7TWlhfUym2b8kc1Vd0SNUj
Ff+8FaopTfJlsrLAoArvx9hU8j/5WwY3LZrxk7cYHeYuTU+3V2ldzuftBR7dGCS9deoF6yp2zvmw
N/hQIGVRkXSCqFG0bIOO0TmamwBt86U4/DSRPRfWYJje1fi78IWk+ahSF7YuuGQ4e4pUXg4MtxwS
RCFMkOQ4K/RBGI5WeN7eEJS1gzHBB4zjoVZeaMD+GgBIJ7E2GW3k5iDqO0gKm+VYRNMSCGdIWWd+
NzK+1DTCuiSiIRGlNWB3ZwwOSv1m5BrLl7vdecR/wplbbGcI23ZndvRqZMY/bngZDRNtxIogO/yR
4qgMJyXL/ElsOBOMuGtKzACtZ9v1iCJaa2qtccozfpTMf53RYkbGMxxuqiPq/ptVmuRG0Qy7U5gV
98sksvMvD0PeUfybZZ97aPSWW9ZIyYW6S6T0IHlZnpxu6DRcAC844g9aSvrroJnUqG0nmr06S980
kF/iG2PTdcsav9Nt/3lflDD4QvLFEb93J4xSt6t0D4Gu+Lk26q+uXWjIWjR8vYKEkff9j7V2a5Qq
pPCTc+4FRCOGIdaxTAdaR2vTbQf1MNuVrihlBkwPIAaXmlJyLoMwWzHylgHKWsfNeSI+PbWgVijm
l64VxDYrV/PrzAGLCisrNvuOjRwtkdh/wdY1F19BZDUA9gQUj3twPFfTHYyQQ/ZEYvDzbiyWQIFf
b/iFIM1PFXyHG//woJDwQPzMEUUWWP2ngcuR5eb42vYOqUR6/eRAZU6k1xN82HBCidZipYFUDX6C
NWe0m/QLcNZLbLyER77WqsbMWkCatum65BocWAWSF4GrQV3c7Unc2tviFwvHaa7avYxI09BA07jP
d9TL1yzUuvfJsBoCiPysBB2RQ1cB6WnAzpEtHDR5ujV1Vm6QDRztr2ZPV0ytX5ml7yQImY2y4miI
h7848qULoqwfx4rKsPO2JO3yH9/SyePKzvn+hIll7jiEAwSovRRhb0KJgHnG3uP7XIzSV8G1QXAV
UzpK//fQQ7dJZrNQY9g49fWFQmSoxoN3ptv+Mc2e2kZTnAG7doeTtvhmIwysM4tfWV4eoULGm1dL
31YRKD1DzEZqhZfGtDW7D/vd0b7yB2vib9c07nOVdPHs7+sWXVosJO68zKvSrIlokmTcb2JEijDp
Dk/R3wnktZ6Dqi2TITatSxhk3h4JqcYnEelxtKQ7QDwpecCsBpd0SK88K7m67WFkiFv1cL1MtHY2
Ktt+BgY9I/elwFefdluJcE8hrFj5O50v1hLQUtmSS4B8dCiKrRgC9vHvVvOOVnWRG8ukm4odeAKD
QTZM6sXC6Q3r/uj7ODHayaitdnnL9TSNsn2HNczoeN2+u8L8YGbxpuNAyb+NeNaqY2jVubs03G1S
lElKf4pWnS9qsdZGFzHqpAN3HMpfAcxgmHOW3nT74k6Wbw6wPq3cXKUSpNKE/7riEQNVfvSKvnRd
Cn+uUDiT4RaMYIVcnxvSU1k2+L7JDQoDT1qjkR16fkF8qxdQhsrJdmddlttZm7FO5X390V10kp5e
h+1mbh4CLJmexCz4ShOqDxwOSor8HR/EvAJFbn36yClUk4VrXh8PnXfSIrwJ2StjMQ1u4l/E9PJp
0cJQhPvFkTIjTevTcFzxSfvkZ/djfNdcgsMTuAI5d2wRuMzXm1ItHsiWCt84PppcQYDlXon4+gjO
cmF1cR0SK7mVnprpP48MpfsHt9nGe7ai5Gl/f9ackoNdgAAcbOl6PsmIK0lafRCu4sLh4gvNTMoy
LQusT/otm04DxuIMU0BWQKD3pduBbbiGyN1RUV7gvlXontyJHKWl09U0lx1KnrruiI2WVi9iKYLH
BC2W+1HIlnTFsDebR6xMiK3++uRy2huTuLaA/GR0o4I1jZnt4J/QR1PLaH09G6E0TEXVPmpY1CH/
u75iCvlW5wIyUlGX6tQgYMcXaDmjHy1H6f9BTUoD/kMz6Kqu9eZ+DLTpLgKHte5rZ5uaTXzxAEFo
fhMa8J7eB4xYhZiNcNeGqjuz9khSA0tw3vEG5LXAAqC6/vgrAcmH0eYpxZNZpHyKb8idGFeBfj6K
aYNwFUb6oolzr12v3xOw2klMwP9Tzgw2H0hdKkaGyVD8YvK4QnTnUd2BPI1i9rycJveEf7RIk04k
cXR5UNW8OeLerEJKa4EVrsVoK042k9u5yXk1YfuUKmnT/S8rznfEo6IwRW/rplkRKgxR8p8EhKTp
se3pHcD3RP+G5AxVdxaj2inAXhwBNg2hMvTxLNqsMSTX9400Q1TOepCauacqE/pQGJPVuoUcO23G
TB4PsJ3hTU8G8bVpWLlTAJMcaiE1PYfESvbPMj+gHSQ/4ZoA2lpcKIM966+XwCFcvP39oMZL3WW3
8dSHgb3ogZ0u/axlEza28Jl2yNhWfZK4GFnFcjwhTv4CuZIjPlDft98bLPek7omA2hRzlqH0o3qT
eGlVrqv0imgVXYN8urR+jO6DR+SXJlkF+ipym9/LxaA5PFAHIS+So4z8LyEFHYDybJr3ukdbfSqM
UohH2V5mqB5Sm2yOh0MUvBxKsS1wUsda97mN8iGIQYBkpjNnv3qfmI61/ItJuXzdKvqSZBMH4TjW
HOQ8oo021QWJfNi+auQOxC+bm7iRLNpmR/DjcdcR2NDVYZ0hqLewuh21tz+RcXa3/6xS+J7WVAwO
HW1snUz9coJcQpUdArd1ohHvfpC9iUSjF/8tuj9CLMV8eD3o4qtpSTrpCwPavUsUgKu0dMIcPYSz
UcUQEfjhaHbtZW0TJYOPE0KaZlTpLHL9UfST3NOXuHjZBy/Otv3XtrjUslM7nfuTavbKHmEuBXFj
HUsVERxIM0mqeChPTN0WRDWzP6hjUnIeyVv7Qzzxs1GueScAw5xZ2VHba7Kz8im5DUaSMYhewIfl
foTJC2JND+TNc0wOTWgeqBSHvzIsY8O5rq6vb4bqb18qtxwiRXTi9cXocsOmcyhQx8IiFydtlodT
1bNmbaUXMnhN+GpE6ANkf/CMG5KbH2Z+JPkffClE+UOdJMU4kQk4kvRQNES7ebOyDQR2yAtlhxW1
DX1Ki7kGyeBCmsaKvvpEUACPMFHydafHewvG6UJVqloFCnLZxQ89tkA2fxt0NPOD6mRp0f2ZI9qe
xa9VYVEMMmxzQh+Y0Z4BVl+26xHVD7rwi/694a1tuQ0NJ0kriVsWooQGzpplIW8ZC3PRt/GQDTpC
7xAoD3SYrCl6L6Xn9i+ke6uVKMInQ2xBXRQ0CgcM4vLF/KGDdpgxIkFzGhK157vwv9JlgtEEPSK7
io9QDblwoNw3+wroszQNSpT/HOZ5fXOEAWNTtD5I7WblupnMN367suOdsu1Wo3HFAbQ71OMiIglx
gzpY4u6e1PfKYqsYiN2xWdLZ7HqSTspNwDqsAUhNmHom9O/Ugp0HRSZuXPUlB0YKtSZbTaq/sowf
NPlUNMeIXw9c0XauqQU3dCN9upl/ODVq1JDxFpXyEzhxHzn0LGbXMMmsqZkTppaX0Kcilzj59ooW
InyGxyIRCOsAMnB7QrhhYGumBjvSBYkAoC3/qxbtnQibuAFZMSe8ZiCWlcvIi/7WqVW8py8zCAzr
MO7iezl+IishZR5gXjp8av5ICIdsMflwJRKy40or8qDyP1z5r+9zvBDCB7yzAL6F5zkoSKcZcqUN
ZI8cR4XOSHx1kVfxsSx5LAXJiBnbAOS7z39ndGKjQnFupYiPXXRVPqMco0RT9KACFHjBLUAsgTxJ
Y0K5gdquN0VpXalVvGmGl3yV1alP0JuPBTnNVUA2wPDhceOn1o6RG0lT7xv/HsVisrT2T299QAUc
jqOuQ5q8S0nMiCXz+KeXJpjhlR19ZLwzJJSr5daN9FSMcEenj4/nthgiYGzIRrelyISQ7YAye6e2
bQVMQShFQ3X2iIPs5SCczlQL3+bQ+X6RTEfGQFYb46LaGrnYbW8QPdwiUsPflAB4skFL3/w3Chvd
AeERfq5veozlTl5hVym5wXn1wBIi3lpm29mHuOQotYk+80qohJc4qcPLEDj9sd7RMar/PIln44fF
YFXr4m2dpJwXMlCsuwrKuVjFOdxA00WUV3yOdmCU51EsVSMCMXerGZNtmTlbEZrTWCxXmFcsWt+k
ZcuVeFvvlCH8y7Ez7ZqUFuo3L8YB27EQpRu26dmui2m6vBynIj2ya8b+odT+SGs4YNckKJjc3uXJ
NRsy4mxvlVQ/AdVnz4OJfAL+s4+0fytKFPd48UffnBuOtrhtaZNC3+7ZgqHyqBSQPPp79D+N8BJe
a/Z5ia5LY37s6RI5VTylvsVmGkBdRFLT1nUEr2Z5/IOubvuXw2NMV1tlWyhH/Xq0BWwiOJZ4Srws
ADiybMKnqKWGBLDSlzcm8ZGg1ZmehUzpIv5gC8mRD0oCBsNTEnbLYLeX5xDvAVdVYtZ7bDyCPg87
+EvczdZSrnTT7kz2uwiuWYSknsS6FNITMlKonorr5CwoHXMzBFFF8z3+BELjl+lb2TXL4/RXneeH
xacMnDsgvSb9vNjeh1b4y07xaTZef/6zumpU9SqkAVquAw4lBHI8PsqAZv+0oV+6iUPMCMbCvg5M
VmWwRIWqYZsg0hhEH2FAf6cGLjjtEp+wIhpjvfYH2XiM4HJYovQBSgQLw6691l9OW6rCHspDWAEU
aLAT6Xoa0EFWmIn0KWJu0CxL8MmLga6O0jeGOinYH5KXf68b2XOanvtKqOmmf1g/EQGaZVxmfDDf
dr24VhpSKnnbC3qBjBzF0gvKXeYq7TtRMF/jOcPCrmUZioDmeixYaZc8xdh1++Hpz321YLEnHpJ4
2X/Ai8yDQQesyMSPl8y6zUM+KP3OwXFcHfxejYTijcDX6rgDMnG/48+J966p60l7Fj6VNHOoqH9F
euzSOo45sEM4QDIoAppUWs0RagHtlUvBNu9ZVAUCpkJFAd2+7wd9i1W5EFzbdaGfse3of+uZ/qnX
iL1nJHlellxOtrDXkM+7nAQx5rY+fa0KLncbt4F6c8RDPfNHMSS0CJTuORwXUNiOAJ4guf9v0zdm
ysJUqIiPkDoK3IVWaDYxsTvhlTr7Zyzh4kyy5m1IuCYpQJg68PYAWJs64sodOnBqcIBIXwuciulP
gse/aBGGYOJu2BdrUgktEq+smOBSzYLhAakomLM0vHl7M0FK38ZdgNPpL/vpFGQ/uRL6fW3nw37X
yCc8Is8XXx23ulhEA3YiA9446aZzXzsgEz/m4mQqKO/uLsQgVKqh8q4EgRNwngzVDSrF5pmWSgCo
tqIlqCZMAs1J1FcAZ7ZPno3z7sxe1bOVk8ZtzrdzFs7BxLWvhfDAg9nfJoYf54guRs68yMijuvJ5
UpZSk8BzxYEXxNCil8MuHAcGCpzwDZufNr9kefaBXtR4jVK02+PQ3Rq68XhUQXp0lee+JpCnNxgg
5kdOp9e1kI7odeuq4+nd3JJaak9SxL4rovCjMwRXaXfk5ZuIPDYTk+mWKkHZ9D8JZyCtYMLnoztp
2wVZpRDos0dw9YEX39meaCpsyAIsJhi45NlKIDliE21bJaDzFCVXbCExuyoh1oSBLpEztLITWMp7
EZRK0w6pSOES/fnUkcKuxw9Y1ynO9vvC/B/452d5JlxYSg4bW28P+oLpsOctPRVbO2nQMdjtxY2R
JOgShpvZ0v9acSXdUib/XsMNpPDmADjYXGhIOilaYlQoVoF/RAz3SzdsLBWTSCtSRe4l1FPp2Qt7
jGve+MC6/QlugKfALtn4+xEY+UVXs12Lt0Iqa4dpIrUgunGdaDmtzPIN1Sf+fFDgXFRDDYYgSL0q
Ea0wta841XToGJSHltZC3SJccqdOXBcjeZOS3hCqkvte+J2bY226nD9Brmnglu62BfVfZynLYOn0
3e4P2y5sGTB3S8taCsD3TlEvKAiyIPjH5FRFr03BBZ6d/XMW0cbS5Vh+i4GH/Jl4zJYhQ8TN1/VT
l13PPH+mNaublA6lXJHFVFpVWG/4NrSXHYFUZVeTpYKu68cG3DhQkSjmBuOtpWwARjPCi1AaBP3O
ZMSsSJ2/8qY4qEljt9oLoCNi/OKWXcXrsEITJFjqZ5wYSQe+j+ae8x8scUqPwhGcaJiSyCL3DTSH
A9mXZtZ8P9WSER8y8/XGVgaWWGfLIPj70KiW8trz/RsUvIMOFUGedyGX6wtZzHBpb6rsjmgVdIU8
zWid7rsnLLFwi6VDFBdxf92hW+V9fZhQ1uBf/TtQsJ2oX5LTUVUWTPEU9+pK0jrV3Xxzv+CcFYyV
hAtZTMl1m/DTh2XeLBw/xNFYg9Ea7GgdhaWzWiYYwXJzdR/igVwqUGaG5x4J4xbpNq4KBcxK2JSv
75qpJSKO7gkzTE54QBWuvdsRGxtb9XGMFRXljtrIZtnHDeW4QYzNOL/zCwS9z90WkRMkpS+Mq0QM
tUz9kN+1g/raC5XyLzLIYP/qaS4twJynFV77NM3Di85v9HvoPGbFG8pwh3HZG5Ohb+3FwqebGrep
2TUbzarJK/Ig+gj7DWdSzLspFtQArFR8AV7k4kW4YFM/7pMTqFTJcuTvflpllZwabxQuYr2xO1rV
ioycsjwoJMhvIPJj/eb3JNXvIKTbEqu4Hr8naC9KrJ12rcRG1kRQnrUPJ5vX/Y/LhziMZGFPrnoC
w4VnpXwt0R90E74pE1QymtVEdHfPaCu8kgwUZ+/zlL4gYL4NolWvNO5o93Bjg97MXFtv/1ZpH1np
7hiFaXl9EbO0u3EXU8cvfc0NfHTBSSFwHJ+8TQVqJ18TLupi/PcnZgDRSsmahUOyRCL13GCyisq5
TdUtndnbkgvj2LKjCjK+9PSQAeN4Fl6rJEznoBt6weRiy2nkrFO6Fvo7P++zsxKWHUygXD9ZuNhW
UIEvXhb/eMAabDPAWzVxG7Q1swOxCMv3PiZm8zZq32hphxNojG1ulOvis9ZXB5NWuXXdiQKkFtdY
90e43j7/gVUV1s6TKaXLb7HtLBpRd+EUwiECBOvaQ2QFQQPCgDnz/KZ4vCTIPNyXjwLUZar9B6FD
vTMcePhzjCT5u0FmS+XfxC9gN4hS7gH4A3Xn6Bz1BFi0AfpKsRBgZsMaDiPfMMAAC4KVCED9YoG8
tRUYB8U9954crm4Qg+t5C8fRa8cOyMollGsECp9g2r68WAAFL4fsmjc4xGYOT+F056NXFJAcP0sj
MYCq9ePPJ5DDjfky5/m1KHG72gnd0YklOP49OBMj4QVdwIoUxwAIalKvhI2lMUYZcUBL68/G0nCI
cMITwrrPile7265IH0jKZEPUTz5LMHbTp5Z/FJ1OPCo2sABR1itsELqVbyclznfSWRJt1MXMekNp
9rN3P1Cno/s4hYq3zoUgDZ1jfQv9V903bzzyhRDsYD+SCJz2Jp/+zsiFenHgM+QV9ojCfUM9xGVO
gJKTg5Vbj51wEAmdTuurRfTPeOMwiXtyDL8RCIiTxbLQSoSSSiquR5jFqCWkTO0Gsn4k5s0GAr62
vL5HEv5Y1bF/xSd1duAizqDyRE82MlCC1+SMFbKddYT2k2zhKqy3H5dC/8URt89J0cPwJ4PTqvYG
mz+jNE74oUhsF2a09I8DYTvdLhsPJ80P2clUzkmYicLcbTUX440GPxSGopEVCCGKRvO16y82IMG7
lE2I8cnqhrlVUSjLP+mAvxNRh8dzYCtNd9XjRkaSMIVOve0pVjmUz6kJl1pt+q9E99Zk27I+vAbF
ikKqMDzRuF/+U5lUZ3gRSD/0tT7nDRGqfXcAJwP9dyjuqpvzTfb4iZAPXwUwPPLccyYMmeWnNZ1C
U8Yxx4YkIS9O/7camLj/X3ULqxw3BvW9QhwlXXHDa/dKAiMX6dbq+VMshW2mSH95pzUsIB6q4zHc
RPkJ1LG0pNbA2prq0wZ0hHVIgwBzEpXCuwtIT1iQkaHSfOOKHSdAA/mBWcNTNtUKVJ30ukZ/vMen
8cSJ+mDttUhmq4l8n8Y15qFCrgU5hFK73zezEhDviZ3h3I5CwkAN7uUzkqx/AiUxnd71GaI20AI6
Cw5NS1Be01JjtOgjSMKBjq4ncXcaEUpalIvMii5egAUqCylIoR+Cb+mTstDZy5v++QERIFuhJhqR
2zhDrb4Kf8JHwJVDO7PnmvPcX7of3MvKX9/U4bS7vRIwDtfQ3xjf3KztzHGdV6huz0pw0+sUiCe2
1BghgfcypFRZKarVnnUG6PvKFBVIneK51Qr1RTNu6Bp/Il/RxjEFkT9XZJy4AdruBMMPc35UL+g9
MIKfsW3Khm4La3YtOclbgXRYaCEJOSW3w4mYPmBsgKrtHmH0QQOXKRFvv4qsAgInKzsuwBRR7RAE
TbZ+nJScnbLkyGT0I2nhw5hwXKGL2obBfEB+7SHKTafuOq9+ENiS3lV0RMsGWRDAM8LMO7hS8Y/c
RFCGwMwhpPUqv5Xsj+y2y8hnaBDj1kItcqf5V6ulx1Oyyj/QfurN/jMYeKq4hf8vUpzy+jKNizn/
UH9PfHltbcFm4JgN+hzdfdib3Yy8xlNbbLfSt+aI0qI+UEBPsAHGFvGgPQdGGn0zLEHcgO1cgQqv
ORJenQkF6SzMyLod2lKnMTxLBlnn165n0ttfQCVGtP5AkINd9PVr+tREno/DTKkkXwbQRgzJrBFE
Ba7DKPTrw4rWUH6z7iy5kguX/jxMliP8XYeGgtWb9cKhiCEKEotdwhM23881n3ZteUY6wfsiCgtD
tearUb8ckHn8I5IwEGeh9XDtVSCRe6j3J3iIMulQu6JXijR2t8R7zgTQGdrizM4d0lLvBZaNCPTa
oN1DCua6pcxoFJ/OlmE2cgGkuym9aHD50BQTGXzQc5NUqYT15e62JG3Rik02TQdZN+P7/rzHjUKq
vdM3BBefyOx2v+eHBs6oNFJViUtipibXezukNyB8sejfNL09IfOz6AaMvK0G9K6PT0aXcjNKeWo+
t7KbnODsMS0TRWJVjNyxrayZpLB/B4J5PnJRY/XwqzF8LCOFGrVcDArZmTtYugI6mkHO0qTPVQEq
VQwhRky2CQBBi5w95tHQioKwNt+YMuF2jse1CA2JoV7a0nApkJU7IlMTU9rvCwtz5XDcDb47q8CK
STnsg28ySFYcVsThb1o6LexZyJHvc0b7AzJLAYj2DSZV1Pe38dRauPKTIYH3SmLEUhLnKgf7GtFM
a0WPlUQggw1VCTwPgqpM81Be5jCzONHvxAFx9fSeO/Kg3Mas2+bs6h61LIpjkue9rd8xzloQ2QAd
ridJz4wO6t8K1JeDBCjeuPXJvJj4gr7CME3yJIkUMhvBbmgNZ8pAxtW6RV3rPGZ8YJHRFbJX6KEM
pLjnRdEDykh4hW2zl7/VbWnC0Syjx1xU7kFnyC9A39/z/5LoCfgslVPDdoGZRaI/a4feB4rRI/sr
4FZIbHj1pVzIH/7q1xIg3b4lhtJcRxUDHrQvFkA2Lu7w74kT7iByBWkr23/fZxZ/lnVJ4FEZUX5K
vpRmMH8hkCDWrzk6QLMTkkA/r6LMPasqX4ve8SzQDjIO1WW5UOyX0wEVNv1Q7pK8mkPMzrZlqq/q
nrdn+LQD9lWilPTMZOlRSsDWJd6PjDnsCyBPZF1xPZK9pl3cDluhOd7sSnnBuZ2S/eNf4BrVyPzb
w2kLN0LXaq/VNVjiIYCSQ56WD+uaeVKO0CcwWWrI3j4GICaoOvm9RiO5z9Hm2BUv0gMBVeoVmFpD
a84+NbFS63HtL7sON4/42k8i90sdLXkthpgzbIYRfQLT1s7BpLJKkhua1ezLB565sUAz22AzjNPr
0APfPN+0MPyenyD1ADpzj6Y+3M8jI6tl3oH6dvZFQXLHKoAKO1e7B4y+cLiqfoBxHOAzVN6Y0SH5
n8D18grRId0LIPtHHPfIQIFOI/rYvEZZGGzrse1OQzq6mdgxue5+VIzw7EEVc7tpoJD4PUPE+swL
uTOGXNuOu4s6jIu5k07ZGxJ17oyYKhdItgFEINU7I8E1wQbHlQQ1R9jjHUgSAN1na5YInue/OjQ4
OtUnDUChFv4QSjPbCCL4WK9VfjDzqSHUGxcH5yVGGA9KgaZCIqjuKIOv7QLN9bzIcSKBC/NyhGZk
YKSu3BsB+dFyP4m103ippWSkStuzzoWJ6fCfhRvDg3EYXueAftWp+lKgojXVkndYfLnzxW6eztoR
QhZNgRKTZg/S+YiZsT+/p0uv1m3M8tfuEUA2/z+8qFUladZg2dZ57nUK4W6hYiTEATtLc2rOojCz
ev0JIXfd9XsMAdiZqKRHSPKVPvFcOysXV7VrcVw7QAgbBMQjzzOogMI/qiJMByMJYWd7NeHHgn1D
dC0PyYhwY2vYExKulqoxZQMDtJb4ocSEmztX8W9hk/Ed+IRRQDNpgQxTpoPbSmszgzGvwb8jdiQk
cnXhEySmEbhksympBuiPPUDbj/Ca0z3CMCwb0coArjkIcYL7WzQ4x/8s6OOrvtqHW4qMkEJ89nIu
qlUHL5JueN2EfRNXHxqIZkc19yBHa2ggXtzrDX07gVJ1K3GK+slChx+BBxKB2MZH0AQ3Jlyyu/bO
kVmZ1qGP4Uta9vkCm3dl5z5/hMX2w38DUe+7321grnjD3dgbhxzEe61OPGU/Nb9nkiSLhZmOWCvX
KboKXSc9jSkcZljvKWHXzJsM4J1SDRCf5GZYuezBNq9ZDEhZXWRTq4tJf2hcj1fkcsRp9n8I7p+c
Fq03TnGT3ZXnAJxhVf7FXpWxRXJUZnedSeGvHRPOvLEOvm5XGClTa+m5pfcDA9mLkH+p/+44e18Q
nL2VQC10evj60VXu0wno/B5doZJ+I96zizKevUza3z9dSHD1YlkeNEKhQe48L9+ouZt45MJSEUW9
prm8A/TFW1WVanghRua8Rmafu/XP874qNeO1f1r4ACuZW8HRhMzjHCKqOWIhypeHjEoCtekEG1Gu
Seq54EZMNPL6lVQzpkaOnXW2HuB2DkTk1I7QBWEMCIjgRsBt7p04DLu1jfX+tN1MBge9jD2R7rQj
ew3vbu3XG91p6zWEvG4NGL2bCByDnXJnq0Y4IpRcGh27OpY0YLtH7nV1IpNh+PLf1C6DJARQvfVy
EoN+YLP+GU2UHt9C1x1jYh/caLi23v2qJFKdHbkz5MNi5PTGjA7DBmq+k4U5XD8f1ML4pIW3ndhD
qAeOs37jPI914fpeP4puvFFPUqVzM8nJ77brRjtK7nCUHDy144tvGN1mPxeRbMHXCctFh8LKuROj
Oz1U+6iMQwhgQ9StH4fJVdC5Pszg/jDTRo01YTPxV6BTYOlf6NWP9JBdphG7h3kZIn8t3DArGaB3
dHSGeHTedftvidJJrXfpaf8Bn2AKsdfmPJsDb+HtY3DId4lXhw9PaCyNuv1iaGd2wFZ73qpuiSWq
tTBGmGq3xrZTLlHg5Ue0FHUG4z8b1oIJqhlTYVmFSHb/8N0v5kQggnY1h1gCpLITXdWDkFErSQwO
+dtN7FUiMcxhWCtnqbWcIJESzaVvyL1d49MEENbJTOAYC7Y3zXkLUO7CTbskvmNn5OGJZO/GKv5B
Lcyc5StlYg+MFBQ5IY/dRAs+zxMzX0bHXFo4ZMLnJZJLvn6p94ZncEcapKxbJrZMiMk9JebeFhPA
n/0sICwQ+C9UCWC8UxTFqKkzmaf08vBgsTvhqW/qnjTVKIXmk2/+/o21vOeAWIv/94v39FmU6Si/
UYL4/cxUFsNfwtl1llO2x/QerTnoRK8+LlmB0HRc4KJMApRyAHKqS2fpl7DesP5fO8ozU6l0anfL
/dYd3cwEp5Kvy9oNqg79lrDbkll9nLjDby63SZvQyAnQjkB9ibXOnw8P94CVh2/W0z1DD67YeqZS
aAAOfQL0Rf6OCXiz01+Tk8X76N9i+H/oL//TZIXYE4ksXyHJDltUzHVpmjzVKWJyd0/TTKrt21eK
tNLFiBtwxro/W4trYp9quapgDXy10EvJxXkxDob7kCDUyzmPrwWAi1nIlngANuy+1R+OBtA2EBku
10Gs3hu8HT/HpHmnAYS0ZuO7l5ZGhnwqqUULOQaZYV2677HS1Z0vACtcachndergnhY8BlTwm/yq
/cmZommXdlxB586lf0NjICs+t3BSq0SIuC/Wy1ZpvGFPxoJRGtL1RKo0WUwdWtfgXNd14lNhOLS3
P5v5WpiQImK9dTT7o2de8T2FN+6sH0kJf0E3yXmvS7NFydspKiIfVw1cOy9k86JetEAiuXDm62/U
UbTlRbMxm/nLjj99J1rUiuxrq1UIeByDkOqZC8ih6Eb7gW4o3Hg52IHOHCi/6lOc/52Bn5nNXkiU
gGitabfU9x9pUFn8uhXZnkilUSrR7zNoXz13i8IRru4qJ10ypoBXkv58TyTMjzLpqKHWmJXniy1S
em/POGboHtFjmJ633nIkVWB0qHG1EHdiobqzkQNHEC3hFmri2bA6NuUKJrMsxkWuKl0v/FzVvVT6
+sBscSMAVF22OVNaPMZPWPdbBypplGT7cZWQ35mro8WdbbCqsmJHS5IbsGC+fE+NdJtan2DJW3EG
uVfeCCFW/S1IblE+fDjzj66qB4+BCag5VWOEBdFVNwIBiz/yMvAczAFMzcpS/grNCXtk0G4XWhOP
f/9JiBbheRxyJ47XOTTjvO9T1ZmkoHljQ9ZmSRtSncEUPZCKLGL6ukGdz0SR43ytrliHJN4jeZOz
o52Ajww2H/D9wkZmUKTLzry0lwCVpN9r3nir5br5Q+dS0/IpCzuuCV5JPemrKOrS7/ZFL+mwbK5B
d8Vr2RLGhgu+J49uVbhR/jYhu7pZgt1YL1TwbwjzO7cH0u8VW2fvCremNxF5vytutwdVUKKHBr8B
AgDijUnMsVBgM52oUqvgLoRKPlY2CpaZZCur1NTwZAmE3VP9pBj8lUhj93cYITvdZwzxx3FavFGv
JaTo+4usVs7IzW48iyJvNj+r/fv6EY3wiE6cPkA/juDp7nGYxPqlaTpkQIEcxDSSSftJjxs9kQXI
qSSoNqA241hAe6fw2iHcgkaJtx1NJ0jEpT/I9AyhdcF7pS5hG/GpvOa2BimzAYrCefiaumOww6k4
6/nhXTQZSY7DEnbTCW2zPJYRLzR63mEJjUJOS1VFMRfavAqBupyxToTE/GgaX3gY6Ms4JHREzTAz
akyJazoi7eVJrFNt1cF+D/fY+72PW2uAJ4Crz7guyphKbLDKKQbHWPcblEcQAPUcz2d/1FKovjaL
lQu4Ci0E+B/3Gt5w5bxFiRhNaJBK9R4RTKgu83AdQTZAXCCltHgbQLMewtI1mfaE6u5VUXmc3QUT
uEAZEC86iYAFEe6KZawYvN6/cDzM870bTTQlFASGBt5ehj7KmSJBtP8FRuKQvfJ4XXctsjvvK9WE
NGOMGPGlvGWf3KUMV3RXLtpghgy+k5YSQN6negWdW4XOKx/qysNEoOGDdisFZ9JpNdtmsb4ZuJrc
Hm3LsA5lVgY3DqKKWWReZvpj2+S7KdiWHXusM4fKaWEO+0l6ALk1wji7Y/3vt7P/Codi29Iyukn4
fJLWWvXdbNOWX4FeIK7zKQ8ZCDIZk08ykZz+aNByFC2sGdpVpVSizRHK3qgw9J4dHmZo0RwAIm4K
0ssLz5yR2rqnAtFCffAJxXqGk9UfSMLy09LNwYeffk9m/NT+crsz/Oh0zmlKEAhWCBwuZdlUXtym
k4R2V+DiGy19dpRQMRgnz4ZBIi15CaGbgGOAlzmuBPgss1fmvjkDMFq1/1Mku75YJNW1wkBsg2JB
ez6mjBNXytGp5QqXRP6zGg7rSHV3q7NK3gfDPvniyqblEj5I4nCIaJC7j51HaX5cnpoP7h7lpqT2
DPy9Ws0h+pzXWXd2c/01hNT0/aBw48aXMXGVFdOP1yGjgn852jHmaeJhtnp1ZhoKD2nJTUDofD2C
WfYcIbuAY8TH8Ie1YtKIiMuPUBaX7cKSMFFrCfA0eQgebxiRREio7pcl6CHM+hk3h+KGEOd2ZNBY
NDRjEGeAD2xN3G8IoIRBYqkY08IuilT2JFnpeyAR0MDOEjCDPPG5O+Z+ezKbJQKVTFE8+YVpkR7d
Y9wGg/A6ciMRILwuRVqze1Uj3CRIiGsBFXcI9WrL/0WzfDXKWPRz0393fBa3AId7qBJDHRE22qqQ
vExhR4+S0k6iFXYviLLp9jX2FXjjYuWeSIi8yHZ85/3VxVXWStZDkQbjuvVaor5jkayjRbgd8pn5
wNMy2e2dTnFJrnLc9PpPJrAYrCZQv2sh0fk5DzgWROyL6muCUHSnPJEWOOXapOIoiHnPWpHxJbKI
dw4f6TB1+1p4q6cRTyLNNe4oAFhE6h104CH8trePzSsLz50UlermICsNaMHb16oPsTMLhsefoxJI
YoqX0I9uUt3QsoZp94CqNWqCjzoQwkmbNlawy5QQDEvHntTM0sAsd1wUHbyc9c2jkByMoSk+Tnd3
Rn56l3NcifR+VaP0dNPFpAflZVP1jZ+AB1tO05ExgJtAlzM3+ygyCviwZHD7RHHQ2qNi/QqZHSeR
/sx7R0ARQRf6uEGXlIqmqgta333XXMoCcWG+OK76CFQSFY3uS1w0MbxbsF7LL2vSnCur/N3zPJ9C
0lpgofafO/nf+GK3+JJ5bhiBScf7XCrnU2DPR4ObGQAAn0o7YVaJTgdBGcMixKctc73HZKAUs6+C
9RgZZRv4d1CPOV88f4KMCcMejNlSC//ssl7TYk5S24PoQ/FshPpUd+aTtHbgETF4nkHm9hj+cYud
8XkEtEa3ghwIuXCfQWQNcmbUmxxdTlgiwhciACn0nwFcFRxywz2snMEzh/WAQZXQ/RwegxL991ME
+k+6vfA/9mhHzrV++wWFoH4MxlbJjcRSSObKaz5M+pabrQYABMDNcyQ04FtbQCL+jntvSJXFQDnV
TanZ4983VJQZIk/UTtOpJJ9aNHqvy5vTTAt1OYLca8JZn0D7XBO91mxHlNS21yqSbCiciisv+9FM
G9+To4lulAz8CeVLhtLAGjUCXsC7dGuXCVNJvCjWFN9bOikxsy3kPolJz8Dze0GT5inbPflEJfBJ
6Iv5xS3WXOm+omOhZOq7s6xWdY0xudaiFUkXt0Mrm0PvQGc6AJ6bR0BMw2cplzsWSYY1PnPAsmas
79Iez4doXvRF5vLGOGJXdV/XNr+03JtdN7HYXGbH9bIK5R/koT+QqHva62tq5lX3vrQq/PVQpOaA
eLXfad6HluC+YNoKs2kXwvdqEIyeAzni0xh55NBV0MkvcMCqKHJZXbrdDEYtjM8bsknDiOHYyj7+
hDBd+KvBgtfmTtmxevoSUjfMYA/7OpG8HQbVyju0bahIFNdVhrV2cFehcD/427qkZguX7OTFApiB
cUSeG5cNURSxynwtb9pb8H2l2LthghPuxAyTykOQu1FqLqXu5vAMrdGyQ90nWklzsGNQe5QQbRWS
xCmn8ef7FiR0Emq59YsR6YC0sWnOfeKHWPJdEt9Mpt1kYUiltt41sNsHeyKZ5nIOWXjck5uu/V1D
YCj4FtsfPOIxbo1L3YW8DTYqOC+vAfkfqRs+Gsr8Hc4HJoIkZRHaHo68KCIutRA0pwQov3vc/33C
bNJhxGao7VXsJJAAUu0YUP4LcnR8jYLiL0Ex5DiGbkE3fDuH818j2l7sR9s1YryoT4XBkzTUbp6d
LQFkFICUISpKpTBDKPhcwtk+CgKlJI2fLywucJs1ZHsUSXjcbjc6no50VlIBBxu48BxC8GFfG3Ct
atHTEbBHcEl4c8TVuQk2wvlNaOSaQDIlhk+EfEWcjqZ94eSoWRBRlvH7/o1sXh1oymdO4S8rxVEV
o5lEoW5lqw6hKWdc5OGQnBEoZFyvRw0XtS8JpjUvemfblD9J8tLuxbii+FS68LFsBq+zCuq9Xe8R
EMvsLetF0YiuR1jXR57soOrVdsB9vMM4rkY9qO2137uc6z1lj4iw/h+KtqZLeUtSbVH94OnutbXN
jtZrhm0dEXGwrObBdnuULKqgRw1577nBNqlpeQeL71ZOdFdWE2Wauy5oaS3zKwhKHBYBK1Di3VoJ
Fl03P+bqEeUe6a99bJRnhCEM98T8eGuH0HdROPPYamRT5SWhQezhXuH/WKOGCmZnPvgomezbbJo5
28VaAeTOPXSJns5hGj+yBMHXVJLrVFc0lWdlSwjA1iepml9JLKqJntiEBOWfj+QsPXl/Wr83S1In
mhqkz568kQBmsESQP1p6zsAOa3hDT5WXl6YUMS+TRoDnxdKh5UzQ75YB79C3Nj9tcNcjGgQVXEtc
ztxhW0D45BK4eysOxP8pk435H4uAaOyK3zUrFMDkas3HS/KnFoLWEh6ObuHgueWSaBiKY7mlyvKP
KUPGa048VY7X7Ov8mK2c6/MNTi3gMclQH5VH8YjZ9lrBcmqXWAmGTpf1vVoad/VTpsBBqWTKGjZd
+M6MtDuV7liQkp3OdXxdFcs6Jt+hrVivsMDC4EeSmD+5qf0oVqpsia8rYl11/8co5/op7C6e6XUe
ILg4rQLohHaKtZXZrAZA9182pNdQ4/R+4kwzZQVtbODKr4VmLBBQFqqfTgzjnPMSOcqoG/5+ohzw
PSM6CPuqiP9sXdvncin+spuuKsjJ87FJYYb1SKG2MlKvdikXFJUYN+r4uX1TFuTreVWAYCirDHth
y2he5D+X4d7hR69h+cjX48tiN0rRcisDSBuJdnwvNTdtYBE/wtEV4yDFjPml30ZUv/Oo74RW1Syl
JT6XAP6je3Csl4zoEYfilIUe3PFXDLZ5/uM+2YRXaRY2wL6C9UV6N2sU1QzigQ+xDDh1V3NpXtKO
V3nDa2Ud3FJhMMKWZfwmf7AlWPaxnWlSbbJYnHT8MQehydLsNKi2b3F+rFj/FcAArOFvWf/benRC
drFZIFPP3VQXbFLUmtqEdJRV0igolB7aaLol6/0jrcizgcbGpuUIencDvJzNibBUaezbR4SoHBTo
uexcsStq3OJ9VT0/q4z3AgKuhH0kXlWKPt5rPwHOy/BRKLvm3RkspttlXlYr+mAtXyUK2XQnAGoH
BBs95tTdLyqGfxklFyzRpQ60vZeCvu5Dyh2YuZCW++ngqM8hshpBN8ZtfT4BlrVuC16AhdQEj123
w0rlmpBuWO11g3r7cEj/YjgGvWessnPKPHV5u9N5+n6ffIBuBbx+YJRXfe62azMfuVk07mP0pYA5
52REQAwLxw8dnPzrjTwNXXrlkSG6Tyf5BgrWT9nTr4VjgsNsA/fkhdwpFfkALdCffMiqacac5uR9
3bhtz+KMni4S+V9skpT5inzZF9dB/Lq5OQKWjPOPiW8PqcP/bY3T10Fu7oLsDLQMkz4PRu21hj7c
ulwb4q63Ioh7c+hz+XNCCytq9IgRW0qQwVdPkQMvH4+q87oEbpjn6vFU/2+HNwPfnwUJh82kVUUr
52jKQYMXRFJ3wrSaOV6G2E+97DqoOHtJfwmrS8VhrbVqL5h3IIEVnQadaK+36ZwC7cWD093GuUAR
yXafkrr4DEPwqR9kfyXiotgeAfRcqlbfCRRq10+4fTmqVbgVLFL4uMvzhECQlSeLXi3L2RpLewAb
rM9t90P90Oa1XWjZs6dUhzpsRmIy9V4vBmFbxcw9EOxgCQ7woj6ACF09WSqcXXEh6IgGbx0DP/2n
7ev7tvFEj7sk2qowHW72JJpsf2oY6pNAoYB8pXIHLcUZQzMBbhdQkhaR7seBuj9Odp/ynMvmMxuM
ZVH1NtOpR6JCAC6pkTJWwyVF5TP7hn69ebz4WS+hVu9x7L8JS/aMJ0nHa5hxjdPtqglVqj4ELeTa
ysQIEv81TYQ9PdMzkweFdSZMh9EtkvbuTGVwis35QjaGFodtnLvlziNHcIkXUC+oqiBbaqdpfd8l
HjVPOhSM73PEse3roTDTTVzlALjdCFLvcv4YA0TbAJjiuWLM/bQyqtLbbsE95UXOJkAvtU/56yMQ
xCTKW/GNapYauRz3O12qNsW0I/eY/Fi04cWdp1piN1Jj5Ht4NQoMO5pSiGCEUXjWbal43SYeCKMj
pXNZjBFzEv3yNB4vt6NfXSo/eD8Lxctjpvf4TRy0/Khx9Lotn7T4pVbM77A9gtbqASRMqeEbyLr0
7uYbYSlTA6hETM2vqWpz9frLI08ZqxOpes+pdi6aKEgRxEwqJrxVM8F5FBRGtgyO3kNkZmNFUzED
DL5FAcYqtRbTcOiCjabS0obbI4VINQSsMRVbFGBPzxKirWnR8ahMvPLtS2V8ENku05D1SgHQ4gfG
yoHyPwhEforLNk0GnzY9IUFsCKzVwnVnMilFb1Ebb7v9sj7ZuEFViiDk0Iv+8nnAYyofHi2u1f7l
ZreNdSCP/sA2OSLF70k8DjSO4sQmtEskq4dXlvNeKDsXaI9n1RiIlf6rLxb1QO1IjhRJy0qL8MjM
M76bS5Cx56hQ9N/kPMC3Q5w2RgeawQWDcslFCY+dQ2imGNmbXGdzUsY/5EuIKkATCQGzLW/fb1KK
N+Qi0hLtxD1v/Kr7/Shf/drYRXZA6qWjP6Ym2CrHIWXBA3BRVejk1Vv99fy3wxl+rKk84KKbPT1s
+2TZW+nx3qNe73WA9+1DPnecHwtymvPXX+yfpesalTAOqUPk21Shn2kgpvViizMwaShc52XJ09Jj
+grUXA88oi5tQ8ZGWdbf+YR9EUujBZagclcoYv00umElmDWJSBJ2fhNOdwWWyDyI+Dc+g26GUZ2Y
b/m7HquiJNRgDl4tA4kVfDH/oT4Yn4/xx4CY737iBq4OTOfL61TAKHWidFlKOcsXpBX98mneqs2d
WRMtb8m82h+d9eU6fKIqTjbdSDBjd2dGMWqH8Jl/QE/Qwo0LUyMvcQE2N1Pm4p4Tdm5ZJqdpX0qy
e7u3zvW/zdEW/Yrz6mGEgAQS0erpNhHbolilsyGhtxtf8Pus8ziCrk/OUT4hACu2JAMzUAUsjt6w
PCq0HkOePoyqocSwgRHXsztZ1wuhrbUk4E8L5Fce6qf4L+fNjijKK2jwXPnes+xleWbbeDT8BOGe
bafJAO1BH3Bfxlmgov3hMGJt5bubdTsSdFVjDnPwIiV3BYleKv9whheYqPaiBRUH6PySkn12uUNX
ZETfqeZ8zDLtw811tNoCIRE+zONHG/tNWWFFwYAMlSx2TzDh6DTqwnuWjHP49E2mTj0dMgS78axr
zsAc1Zh28ajWqXmyZkwrQZzW1b3bJsjYz6A6FOvciQo06AkBvVw3NlSMFh4lgtLfFgIM0qli22Ww
PYJd0HDsA8ApVGpv86TM6GV3dfKKN5GWU1xQ7Z4cvF1gyxNLVb3Zb5COtemRGpJVW5hmdipjHLvt
uO4t+xdJ6UnNxNAu2NLc9dopSwxkF58c2Uru/UwO4GU4XDXcukdP1q223C/lDQqOa9ED/R1+AYAu
sn+4FZdPGBJkU6QKh24OEMrNQelrZvY69YRAZreJdA2ZfyQQPtx3VcUzq/T6wa3+paWtDqMQ2oZy
bfMCGHUbeKyh/e36wcc7YzUrvDQBuJDDduFoIQY09qrxEG1B7NNsacU7Q3cBwUDnSvsj1izGwrTb
PoSaVGjC8iZbq17LFaZxxMOIuynFAPsXRya4M1okIu6aJ0226M+b4/K8V4ueuNrbx40bj+7xPVaQ
bqerdYNBHVtJVA/yAhFLP+JiWT/Gk4l+PKz2wqaXlbYAuzaWRrMbVxM8lScB2cigWtDze6j99dkZ
2NeBNXpTe5sAwYrib4iGfy9+K1vbV9C/GnRZopOOtYo+EZ00isCO98YhV5b3hkIP74SLm06crhhY
tEcDPCfvOlthVHmZLDE2LvJsrQ4fwZr8bEOkTX04XW+nkd9AL9zIkcJ79IK9gb+m6uFBzNL+gQzU
Gj0QGwa19DArdfEKgjqyXbCEEbvCjrvjFJNqWB4lG9pzief45mfQWiBHTv13la+RiuzIdTE8zHq6
X+cJ7Wb9LY6u7zA1WPwDjwiVTv0cUjwO3lIvO2jqxOOI4YssfIJmVPknwAFqo6ZiXnYdxc0QpicK
8d7PUTOqI1BCiwRVNK7SyCKdjy7/rPth5+zL4xWC0WmaKnqVALsWWWO7OLSiafA21I4vJnxFASdx
OMi8v4gSja9xp7JfJv1j7mdw3m1fOVfS4o7tmkc6pXu5z1qBwdF5rATe3C/zA1peie20e2cvnVzI
CRtOnAVabCvgPR+o4UGW6PWZ2QgEgDe2LtgErJrUi3B/UX+7o2s/aIwRGxSs73CiV7dOAeTUcxND
pJ7f23wWTqU8kmBrqSAfISjzeH5zX4kRNX/wRWYWjT5N04+LCmKTSmlQs25fJ/989/OliPcfEDO1
qFlF8tiRBtbrEObP5O17klPU6g0Xdkz72M1yQxh9fLBIx+tJC3uqXwBl8GwxGXzIEKM7CjWElsDK
kbJmypvX9oUxlJN8TcWpWG1Q19uV1Y4kO6Rfc/h5Ug5yvI5zAM+/tlrZAp3otQrc1daMre+KRcIl
CYlZHew60kZZDzumvlngrahHSP7mFxSrnaHxkHY1AHXTvu5gsU9CkZn8JAfnJGc87OSQ5OSNE2sP
d9cYi1EHkshXw8h/eFgj1IN/pE8+CWhdfB134iNjikeHRN64Q0V/hem42G9XFdEsqU/xHX9JJfj2
/04yDbtxzt61d2+riWWmXdFHfT9Vkux90B0P5IiLBSzf5InhPhTxA9iSXwYbrtsSueLh4PCxScH7
h3BR0jvw81xgAq34d6v3WpYJFxqL8z9wglaFlEPOViZ4Y7QwK4nLjAsHzLMhOiWOeBu+5LfwLPcS
f9U8/PYW7TdNIDA1xc1sRPpArV/Wg5PkIWrMdp1X+laQIdXF/YK0agZ12b5WXFtCkNFkNPHBImoC
i403ThUtcZ9YBreUaYB7KUwhhEReNU9r3FHr5FWe1NPjcNn5i7s7TTRv36p/EMD/b001xeZ3Czkx
5h8zeWAk/+Q+Z+KkC7MtG/JBu0nDNWenQhOuj74B5R/YTqdYtjgzh54mOOMdvLCOZOn4B++tYjbG
IvJYmkXYgGcgMGZKYP0r/dnzDlmcR68+YLr/yErXxQFiQVCnujW+CFoQ2ACvg2NI/yRBgkoIWMvW
YOc2+KETK1aOANMFQE/eCYTdDiDycmC3qd7UxSNpruRTcY/I9+o2INKadzzKv16FbkAqrpkjPHoQ
hFi5n1zpcwwqx3GQMsM8qZ+Pl1cKLoP1K/ODfqlwBjYIBDGgqmZERZq8YBoEqsTy/qD3VzGvCRi3
lq5fjPox+OiEuaFrpTAubPnSozQQjSBiYfywEkH9uYIwbtcCsuXimcsO/2zQic+O+7tCvAYdTDHs
w+HlyHn1Y2Ky6MpiV87bD9Z1NJpVNgWuUwKsTTKwLU43iZcH3VxTcDlFsdTVSUHA49XuUdhG0dfy
qv0T45DbvWCRaXk6euE7G1G/zENjCfPmf+LlKlD8/4CCbPWUXsKN00Uepok3RTUcF0SK9YjI7MjV
u3Hb95lRnB+3yRxYvXmw8W6DcJ+gLztJHmpqxVc7PGTi/knCDcneMGL/nRqHlUaU0DlHdJ3wNeHt
He9//sbtwFw3NLGPRJ3P0BkGW3hLdmN1DaUlacKsMNc2qNXhVrtvlVi9QTNiG6TKU/Jecq0mzHF3
Xyx06ezylpGDhCT6YN1IByceRdbu7T8Zg2KTe+YEVj+5RLHyPL+IsZ39NWor1DtKDTRHE+65xxRn
uWHqGfYHXmQ4MPGPy/wVMiSadjMqNPI+z/GPBouSZ4oB0KunQPEk3K3pRyF4dfH9C9r4NNhuBU2G
e21U1a6htXlHfUnSpMzi11RWgUofw7OmcJH59TnV98Jq7IEnCFge8OqG5WDc3cs+5BBskKflNK62
PhjLDg048pY4sBGBSlagcmvRtW8AiDkmaBiEyLjqevYwQR2U6EELeY923tUdCfzUWZmGyjteLmXl
zn0jd50GPA8JyEsEWnu1IO36ayKhLr3HXK2wPlg6SkjBw38e2ME26FuZcUslTe3CIBOn3uqPzXAo
n/hLceHthV+u4WwpCBosCNShEFvdqyKAy0sN9m1hK3Eic61DQjxk+G+ETMo8Yl0xB5wmvg+1Vgbd
9y+mia2Z4xn3erTVq9ZmSyT7P2Dlu36DyCYGccd5Z8lVuy8X3w+Bc1fjJ0rWpVwdqlcRaYKCokOv
Crqo6EAa2BSgArJG4fi8FzsztFzZohu8vKKd+qKr52jqHuW4eFw1DL4YsXQdZ8DLkGMfUAxA/ewz
2x+NywiH+HZ574P4A+j7fwyFCvGT3jYrHUKGX9D4D7qV1faOFGDmYc9UJS0D3A3YDpDErvYzuav0
8edVf0kFXT8WXvRSGr9Frq4tUtQmDPWtL7X3FUBaPFkopNUX++j3IJecXkuQ6GqMIZEtJEtpAdqH
VILQZfNNJ7sPlxkRYSiBzPS5ErWoqy6k1Drv9En9YPh2EiqFdKn7XVab5Nz2g1xVTELNcvcbgYPy
Y88Z8z/rr4ZO/92pw4k6hX4lhATALGa3BBuSV6FmCUpAjlFC45umz8q6f+w3x28/6+hfdJEI77uL
MAQHhlF1gF0ifnPZesBVhS/+/jRzcR/NhnlwwBjlbFEsMYVjvBnS7V8DIp8wisPmKqzjtVuEXRlK
4sjezWdY+dRD9khDFDAkZ3wBGlXgzTjUfG4/EO+RYExVIMRXZ3zHZMkUIhohOFXcIATGQS9ZslxP
yM3nH4ywYFJPl8hid8maF7Qi0fBafmz+JgRHmn8XpTWEa4zBJu9foHrDJb29JRl+9I3eLhCEt1WX
yOxNNK4BU7oZsMbTdR0J7jFVxkBwXmZIADb2G0e7GpR74mdVXHhLBcRKx6wT9m/lguGMH263mie4
/QYuOIgK2Q6ymZHyfWOmL4k3B62u30/AMv05HzoD3/x69X7EvteJo/KqrD75jNy/Kc2GFTZZt8ll
YfC814Gc2fnDv87f2J5c2CRvE3skctmNnkvxed0X9mtOZdS5OQis+qYBqD/8VIo49QNjSE8sUbOw
x/RDxZ46g1srD7RWfgq+nLxxhtWJE+W655XOjffx/MdR/5LRvwwRjZ6E+iv1u0gMZcteW6IvF6OH
OcjMRJADykaCBtrsteBexlWU3z4VXO3G/t9RuUN7Cej0uYcI1n7vfA8AcDXv4g2Quj4km4NVYBKl
L38EHSVe9bgF1uxvElxdP+hXrOtdP5DRrdkCJctQX/zXnV+mKAMgYrszSVbDbsnF0u1xNPHMSmqq
0ydQc7dkMswA8foVo1xkhh+TDxcfY6QLXYFUeyAlfuCSdEuSe3cUhNI5tVCeDxcFE7efmxTrXJPF
oiFJPKyCiwxM6D49BMQb89PYtiXJOtv7UqTYSYZNWdV6tSYJUw8FbzEtMwIuWtAHjcAW2KWrRq3B
q35Ngt7flcw1LC8BjEvW5qTpmOrytZxrXrFmHqqUCUYgMBDLsKiHJ+7wR+3kWSqSpoiRr9K1gRRB
crjx7XooTWqZCBpX6Mz3sTZAMkfHvWs+MO59LGUvWdWluKXkT8vjmMBWZKEuW97dlP3kFH0M+Yqo
1IGBnrWctbY2IM98pLxWz1H6/Sj4vDuaU0WgIpDXLvs/JuUVVApq+niYgm9oGKqRaLgHl1lA9VtH
y6FfQDhZ1Rpad15TNZjvtjJsLgHJSI6thAmKEplGBnZZjBK8Tuc3tYDbYOGmsM2MT+ejXn4WApZZ
McE1Uy/eqTO+SszChEoM83+bHWRep5iVrMUyUWq1KZGZ+EmIfzcqZyzqtEFdletAYP69LpitqKU4
lSNoPE1cJNJ1KfUsbzjLyODyG7Yu3OkgQsXsu6uAfjmXJ8nqbMcc7AywE+BfSetVlqDXD5UMJ3h/
eZQF2j250PRGQv7g+882T4RnbKUrxdI8SIJZ6GleUStysaRrCMhBm3eDHBosgT6CjasKzmU4RNvE
6YKLXwANNPuIGG6STDAKaE2doNn41K00e4yUT3THx1zBRLWyg4ZtTV9Pqa+7i/FcD+qQBQ2HZCLV
UQQrhSIaacpK4GZ5UQ0nNhjF+vWovqqLXygx6iZQzLZtuFwVEfqpH8/nsDWyJIqudPjCkk+ZFG/9
CLpgo7To901Ka0pFc9WhyPX0wZxlgkLtNgUCh70FRhyldYXvXML2X1VUE+v0Q2SuPb6u3M+VX/87
bVfQlXzfRcjhwvcZ0unEOH5J93dDMVxR4VCL9/cYnF2nP8vQbC1GlIYy00SW9YvtJq0mh1Hmuflp
GtK4VW/aC7gXLhYb31rejoUPJkSsA9GQT5ZJmGdCswnaqBl2eu+2T9fxXicDGvOvT+ejrJOU8G7F
Gx5MJsZznI497i3lRO7XGSD+hakmO14ZDPCrhVX7qm96sXISaHSMcWgjzwQ3oDBK802x4unMdTvw
uINXtE78rykFQVrTzV/0cv/pmSmRf17oeg3ms/g+bwkaHQIj8gjHE2dcS62KzTOh/bTyc8MU+xBK
jkVk2dXZkYSbCNeesBEprb67uGbBTTtoP0TFPHoxhepbmks+DPe0e6Cy9dBId/lwEZCjDPUWUahj
f8tFxXMZlnHacfVLoyUhN77oW5Kcqif1DxvgttiugcHnt1x+2OfaN+zJR1xlgcK0JXfK6sXuPDXH
+qnRvCjIfsXP9o8k2/gIIrcECjyeWrG1McLe9WTZvsZfpqvS2AvS5Kc/vky8UOXsvwdkZGr9+UJu
a82tDN03nH0DZQkFDhNA+4K6/Ce2DVbbipX2JvdX8IXVg1jqRFV6i/tYdxnSTFVhUvPZxLRQTxgX
aVHBLfRLIIPvrKF/MSAw3kRrfMd7vC0OD0sJiggc/LObWsHONmobZOSVXGSPVy8GsbtsQ6JE8+B9
zkg3QxZYlJrca0KKbzqIQG7iDDPhRPdNfbCt8sWi+j7h1tP/We9MwPgEjJw95JuE2i5q5XVmHzr0
uLRiF3m0SM5fUp6mYAXHduLcGnyx9Vn+jINCNmeYlJdoIH5jO7BLWt0V+qkJB6VNPygH/DL301si
89Sg6XE3Ey4m8Tc0ZfGli2sOLO8Yz9ScGeIShJPs8aYRQY246fewH25AsucHxU+QwDAoGOEy4Soa
p80/GWLK/SQTtmoJzpWlb81luI+UzJ3+IsIboNuIIzUSQxeBXVrXgNuEpnFbX6GyAwcXE0eKeTvn
Pyv13mbuYlC32PAbFoilZyxoDO8Q3FJdPhJ+ey8PE3uI1zyHqieXjrEhxmcmKj36p5YDF7dzZelx
9iCOJ2Jq15uUX0JZ0lqZVVkrOQx1tEWlJfLQB+YkeniPZy6c8xfxqCptu0y5G0yOTD4uEcGJdEa5
+eIOWacKn03dI5Yq/9OokhHq9dMFwAd6trKUlOa1VQgPYhVm+KprD2I8719DVtpsDvCOiZBHjXn8
+u3+JMzMzXN6TnIEygh2mOgI6IRnC+NvWbkfCXtLq4DNnSwPXBW+SOILdPMDJakQMo7oGOr4roR5
gf2Mm3JQqfyZGuygYFfYvNBcLOiMnGBldrYQ36ec7peWRjdffBSInEw1HClR/QQJzMZP7cKSRjWJ
+LoQoylcTlaLyZXqLrpwP66YMLnHDGXp9DSjpsTO51VoXiNH87Wa9TsQlBiubU9CyAzYOznYdaUt
OKxcvqWalT2D3KjLXHItInTArxMXKJOHxZ+QpMOI/BLcz3ijMu8Ay7POgDwlI+jJNWNBvFoLbSXa
EWalY+6+qaWJCr6T8MOUo55/ylzHFAyvL2w00pa69CxwIg/qsma8cd3NZrx+5iCkYKD86fBpJfrU
RhEhOZQ2lf/nThKGa9BfJvEUiIRoRVm87THChKAt4O2iClKTBRj+iVnQDN1Yq6pEOE28dXzldbQL
0+jnnAhWXF8w76TbdN+unBX+wLAvHZuWbAXT6QKRYOVcxQ3IuRevUpvGF+9Lz2AI0Kq01kuzeR6q
siFyqvPXOXPlM4yuyTInpooO6txWn7vxl0oXOSflFLjtHvbCT0cP7FSQfSTYqNeSM6+hHSf3wJCf
nPRdiyBLcOTieQ4DwweBhXwk4Nt/OSy//MGpZDbil6P3lITjiD3qzyvPCumDGFbRaX1jRxKYQ4gI
8+jlCEaxvCfHFIbV0+IWFpuT12WFeDA7RwEBJKCuYp8reN24j19otPk3MAkWuTQflSJ3NpGKupvn
C1aL2UAxhEwj0QTiCs4Zk3XIn0SkQ0IsrUq/FKA73IPZRx/nhwqp4igS08nDHDra/W3B1HkLHzs2
y5P4TZmOWfWJp5OgmiXAFbuRDkI/MvTWS3CesOg5HH9zY2DgtwIcPyh2bzZ6iDaCPkFm/eejo5sQ
fTKUV9/Rcw31jX+irZLUEc63/azNAfXYed3/COHX+LYkJltZ1CQiphpjpvp/7d/L1Y8NS7992a7d
iupTcWrEl7hZqMTwUVh1/6neMxphO9up9mr5waW5PNYaNMd/nZ1HPKg96nzE/wc6IYzrJNvRVxI1
GpYoD1Ge8Y85sjcPbOmWJoNRDxIRzWyxfFSuj8w1Yo2Lz6lLfq9nI0ZuLmh8eLg4Qwwb2r0FNWCK
Hi1/t9JjxamhXm2QORdI5vPzg3NBNvJFya7cXtpQpdD90RfxVubisAzfCQCvEl6OJLjHC7mu0fKz
QR/6zMOFMVtktUz7HDQeGCStVm1BWYyWZ+1zUb6OxZAK3h0CrWhnOhRARmUBS7X3dlo+YOHxy3X5
IjSV6gidNmGv7gnPThiyGHuo/elbO1/S69bUn2peLC0hqqIaJZPE3k+2/76NYWNLfMNCf7aH5IW4
v7bWSrhV6t9ktxAOWOBMmoXemzU5SXoZi5hEBDRR6jW8oVJe1ioyGBDyHX12N10eMd40PW9rVNDs
btGAJLdjjW9PcrjY18P4O2LJvTySi4H/FnQlpqLIOqWJzJ0BAjHTp1sMX+p5sEsUqR905y8+ZQ39
HoACAtqLwnJ0Zy0zTz+Oc2ocf2dV3hLKWoWqvuGSPQM3EohOvTzNcmuQfc/qhPb5EfOpgDMif/gq
l1UxWW9mfx1VQmbnaXRjyy8qCU+DdEOsVcGzEtFFi1ZsvmHhvCcRWGwO2nlwshws4Sic0FVi61gs
n2s2gWttFtct4Gud5xndKj65fX0vBgqp+d8zidnYaxp65lEN7aFyy60KQQiKCeoCK71L9wnPeuNk
qr3lS4f32G68YBfIMmf+3ZKlz9IFnJiLveUe3xTTA2eAKe++efxpcmbWdOFCi6bXEfe+CrWuax8I
HpnXXTmcMv7BWaI0S4icSTGdOqv+ZV761jl4F1+GZY28+NcbKOJxX5vdiZMOBmOFRq4dFy0VZXvJ
u6OJ5e0Ku/NNMIaUS+4K4/yvbIfVc8iMT52FrmmX8xqMQTK015LCreRsRhx9DXBxhI3oMjxW8lUa
EwCapX9mYbvcDdm2Fr6tP+NclYWDGS7SMHPbhyDngkRf4ZvjA8avqOsuR1X2AAehGHMkcxcBRLpM
GyYYZKtYTMdIQ6QAhdUeYLqHEfe3A79v1WbQT3Dlfielwg9nB701RbRfn8EiwEauD0D4ICPC44Or
th6VOoyNIr8qLiJxCy5HVmE3qbr0miQZ4/XV39TDUSBJUn5D4+00VR27x0uS2N4loz1h6s0ShQYU
NsVD5R+Jsvo6xPnQl5HnIP0yUfw8osu2AgVT+9R6kBv9v5FRL3n4Ok5qfh2Owop2glsm8Ic+I+u0
4tKLhLUn/JPsTrkEWSCoi1CsXCqF3yRHYJlKwMFudgdMSN0O72FYgt7989h97JvD54MEKiQ7UJ7v
YwMpXUBlD9Sf+oA8kin64yOE+Bs23yDinwdoklIO8kOColsTXROLdSgcGnFafX8Ex2V/vBsKBBw5
VuiRY0wvbJY7Ni5T/vax9wcZ+zveym3OCfHoGcCWXI+2UHKDne1IItjRUqGACAhDtRjjfhM8dVLc
6/7LqZIvTPpnAAhBvzTuzNevsBAtuzfnBnqQ6/QMNoc6hKFwKb2JjpqHUEEX8EvTCOU+sVWjFNDN
qzUvsvhFnI3LBD28OgXjd0CmIzk9u7RQTi4+plXvJISB8a9NjMMb02p7AgGibBJCXlHOe2DUnrhV
eOMM+9qu64MZqE9izDBBmC3iBR285lVZW3iDccwBpbdY5YIuBcGpPHe+YU2XarFDgqu9DBQxCaqM
NVLXf2r5oEkO4+vlwTTNxL+MqRf/OE1Wth1WwLdeqzUZsvwRXWtCLfVRk5KoZs8aNENwKr5WrhTm
eGCQ/gbz+qAgiUA4DcBjjF7af0+B0R5TAExZ9QMaskeBvo1vqjl7tjw6wWOoB+l8X6GfEA9pkWfp
Ip00T+2raQCIfXZTyzLYn0h4IROGqZsVFrwxIhmU1VL8AgVosDdfzPydLTBgYw+rWWDYC2BJJsjK
moOmPanMfiipvQNH/eiNF8tUxiGRRiZiUeWgfH696OFQbt0Gq4L0dNqhLajo1YyXNWs5GImWXbC+
kil3L8zBTZDuVoKC+QZVBT0Swo/U+yvR5QEwOTZaoVz5vkAmK+aKtQzMIL7jwufZuK0hDWFr0/I9
HTVJPW3Cn0+a9aOSqP0Vmqdrgad399z92haJmmtH/M2f2C27exTrI9JxLaJV0AiVCtYDM4k3xkpu
V3YOk1HvTWbJj/3iR7N44sNHWnjUUNZeRGdcV8mf6vT+p0uqLci2PdimwFIYYx6qnKmtdb4zNrWq
Vqu1BcG2n1wdfIBQZs1HHpBp2UPCL410i9R8vZ0722yGpMb8z2MuKf6cOiCPVlPmTRJpYlQ54Afu
fLbVQU+ohn2AYG+yZw+wm4L2o5bh35tc0H4HNUFskIW5qBVYVJ9oLRVR7lFXc9PlIWV5ORtTcTG4
1M8rHXrxQO7ecJrDh2/eYYCDXatJAFQ6a6IjTRiWQzk8ZPauMohezV/S2KRbpt9TsdvAZQJAuSOg
MVrLFc250/kCuDpqi6APxtXyT84wmsFvaBHLD5MsyFdRjxi0imvGfVsrb0gHouPFqqvf1LtaegxG
+HemV5zWZpLppjXQfheCtO5Xb+xOVxCMIwyEIuBnY3uNpmfovtSMgAfvnMyDc7pES8laYKS87T/u
IGVpRxV3n9mw22wcst3RHJeBFFVHk3fMgH7rjevjnSOF/W1cPlmmdz1RrVsk62uvqciA/gH+9Np2
1BLUAModfjbOygxh0ZrJIH97ElExfH1mKhnOv7de3ngeNgEllho3eMTvgZQf6rpXGyAoxcm3js7w
9fzksNOLEVjoz1uFNbTQJLWKOkuWtnMzyIHQaJXsbHn4Qx3hKnZcrXh2hgX51tTXbA+emhzdlzpl
9XsCI38igKlC4RsY41wus/j+G8FUJgTdods0mcx2nmNtXPnWgyg/g1RTcIsMTGsOgVSh/pXwbn1j
3bjgjq0XjDxgwMbmnz35IfdgOaqEWg0bl8/BulA5aUezzyeOGaWfez2dkigabV8V9lOjL2cZ25DT
GE7B083Jnf8b4RZE0bfwxlPI/Dhx9ur/cS0o3RR0tMgHVO7jPAvsMFm8MJwiYRe9CEoLe1G89AvC
VBlI/HxX7xNlxAioDJjFN834k2KT6Qs32A4p37LyZxtBRFNRAT4kLhJPGM0qTlRR2/9GQMgiLYea
T2nxqwqQTLWDwgFj7OCWIe0VDM5qznbCTlXUAms6jjV+DmEGE0W/mlsY3IskTHrKOld7OvM1feyE
RLtCgnsk2XkUT12pNDoKqR81rCD6zsQtfiEQRzXpUvygtLK3gxBFAu9vlsbcTiH/krXF7pTeb6He
SWSpzJAwLv0BCmDCZAhkNxf6n1ydG6V7iZRHmET/EY7Fzi/NYGe5S+xCzFrrAx1TO3laqqK5uBOG
wa6xYMBHTqxocwg41TRT7NHUb2G5+cfA3mIlm8U5ietXQaLbtBreCOt9SG4awm6tKCtlJsgwgUUO
LY5EXsw2YOVKZ0E8zOqasR9QkU8X7RaniZdCr+1RM3om/zQdOehjq10vhb4AcgFfMeDoJNpiVgqw
Piykksys9REXx+xfVkNMjd4yBEgGx4vHgynZqbZ9tjTIQufd1HfJc4OqV5OcZHqKhNYRKBha2sdI
HA2IJCZ+9cIXJAl4HaIFQhzW1Vp86NB7IyU9mtMBccm1p3d52abwgNsSG6mbshOdoh+Tn497I9IB
mgw6oqyYNUfOtv4kFc7g+4qIrKL89wqaW4dhV/oIbNUcNbDhoYIbniIGnToam2LJ631jVzZ1e27j
j7VKj3h0MvcfyCbv3W86NBXBRLbviZLAx+6JdSANFiF03P+ujcePT4TIVk8Qkq9YQLdqu/5QrGcL
ciSmG/US11ix/dQdxZqvXtn3lBdrOFbTQOvVifgTfBCIv+p3kolIJ1GHbZxrS+15kDelAmrEIBIn
yCubDcX09jmxklL0ug4HEFbP3MMPz6blq/ANN5nhRMXCH0XqV/O8/iFbpH1Q0KrKynP/4wL+a4XY
Y+ZqhEq2zaw2nDzlsg+JCm4gJuo/H+3Iej1VmIxPFTNYs2LI+0BYAsjFIeroglCgCQLr8rmMGxc1
Kxl/EcmOExfwgL8qxAKeVBdk9n6DSXpHgs/g8tnvK0gK7iJ5dK9rt51EmkxPAqtaJU1sxVSjy2kN
9Np4WMcwlscyc9t83nHS0iE52YmJZDYbqInipQjNFkUeNzirxeteybW2ZIhcApGf0ErYCegJP4cX
8h6EE0jHEDxtj1y5tonkMhsleFeKOsvGobH4eRECrG3SfUkP76rO7d60gTDSJk/wwvhRDS6Gk8GF
rEnZACb/M49b1bAZUa0dREIYG/MyiwoCR1fx9dSBI+gwIpzuKlJflRYw+JrR5wEkCzQoc8Zp8FIs
oQNAKUhnT0i93/dPgg9tykbJr/xeCPIhQBuj8FDXiCSE+f1jssMNs8UF2EThBJO8ONHPov4te5xw
o3Gen/gmj5WCYMl2j3Zfl/aVaUe1rMv8LvlIo4bCdHeL/uhySeFY+UQ4q+uSU/IX1IXhmeeGdxq4
saA/DC4NhxMGJcwIrAEk2+nIyt9ZwoIvU375GqaCJdwjv67NXr23CnrTHx1iQOmjRICIaenj82l1
pzuJBo0toBYBIjNqUGT9ZaMCZUhdNxzLTLpBFF88jw+GG3uXj5/vBVyyneZzTjCQAEZXPbxH1F4D
/weOz1bl/Fo4VJRFjEii2eNuyl6bUsBawhE9ub3N5eKprbZQcdKzJiMVsURgQaUlM1tvTx6jftzc
DuSRTQSIE74MYvPJr4jwjhb/FHrHZk9TQ0sBTBiHwa3Z5HHKiCxYAdzJ5DvknSD3NXzMlDck5SXC
/Ljx81UZahOJs7YmaHVDTcbzM2Tc5iTMO6YeqrdFRUwgyRQYPoFUz94eLSm9/HMKArRlge+yypv6
v9cH/a9Xc/04N/L6Mfg4r2+6dIGaIyQvc0NH5DnyEa3Td7ZXoNEICWW82aWtEs6qeZb/x1zonyj1
cDThD7P4mlgc2/J1CPsTWQSjzqtjWCxbsDB+8cEAhG5KHBvSi5QFOvQflE2BZcR5RCU3dWJklRMO
+m0mB4yjFFP3WYhpk/ROxaXSU+16NhLEyQ1JupRCaGFjkUZcok+oRS2u95+UZEgwv1TJS0Nj37jp
JejutZ8l78YpEnWQLvGwJh7XdSR4nTEAVyxB1o7pzAkLrzlhkCSZ6EObUVA30EC9vMGb4xJ6LK46
8k963qL5SptwXXxWAIaboo6Ium+r269DoV4TkjhoXLIA8jtIfIgyZPRRYvblMNFe/AXDLRIshPE/
AHEw/rLgPak3deNHE4Xv2CF0PD/795Q79cLxiMuCU14Lt9GTACY7yZbxCGlu+KUQOlgZJlgf+Sih
60EzHG/8Z3O7ZpJxcepnzD5ujq9PJOVQEPk7XNRGFScVjWa5qUB9Fg7f9VELQ1TVP+QQSm4pYVDc
vOejfxvXPh8sSktiGczFP9j3uOEMwu6AySxBS0VaqNvSHwAl1BEGS8lsvc7PFfylET/F8fvF7tkQ
vQQ5cCRemMzdzhDBnzhwuhdMMTL9krn/8uTQeovVZyNo0+giSYJC2zf+hJTrtZjaOpRfL9K24xvP
Ee78fC/cTiMdrlWwSEqtc7TafbJjsYXffqeALpJdW/py217Emdodgcg6R+kl8m+v6XLS8d83/lql
j6v+BPCtqiLugcZIfegoLwWQLaXEnDGnz+EgC3CMLjwXvGWW57wUnj/uWy0s+/sofjoeTEwRRs4E
WFUxdYagyAlMps3Y6TMyyMXGGuCwcPb6W0j+158opd0KhIuUagSkcKeBJS3pv0woWUSb9JfATtiE
xvfANUExiySi/cSLSb8ESA1f14ZRjwaKNYOtpJKx8zYzYDXPTQxzMBgrC5/wOqPiEPF/OG35SR8v
34wWHl39XZ06eSNaR+02tdEMGtE0fAqknhPeuZK3wIUQbPRzgDdSS3XwSqMg13dlzBL63EvFBUFh
Sy40Q23ocYL5pi3qFfyOwHAHAZ8yL/mOBLfz/pPk9UxGTdgcXlg4gkFT9CaZSn3Kxjd5MixtlG3T
UyW7PhFJWhP+l5jUSbd5qJY9VT88h9JHLOy6KmaPwd9oLIOiS7SBdx42kIAQC0AJZMK6ANEZ2lHA
5xnAx8THN+IUmecvkU3+/wp6q+jVBEJvrC6FSdAj2g4yG/xqlsZZFob9Py3hehMFC2dikCxSDQWh
gPRT8uY0d2+W5U0HFAZNwUHIOTSYh5Mksj1v6skE7dW4C2F+qf/u34MtjwLYeZsRIk0wRnXNwT60
crxwAcJcahbzX4FLLHvPVcvzFH6yI8LCK1qgigyPPohPKjDen0EZXrM8PJdIRqxcxVUUGImisnzR
qM6a6VTV1qqzsav3lg+RjJoQ3PeFjrdNUrnbKBfwehtKdZVoIgkLEF7AowBegw9PYelpIJKqD/Nh
MuFmNSzl+KOXAs58FtmHwooppjjmfJtKeOhojDKpYws9Ni0/sN3fr9hbRIfF+L30aAcJWHxv70Ed
4X/EfIT4M762um5g/dQ1gt+Kqxrapzk2F8/GvtC+0m3aNlf18CLUUbq8mpNnilpwNcvj5DjRjWv2
hCU0SHz0Dd/V4udXO5NbIycQnIwICPmHnkNor26Kri0TbyTLRVcX2Mu+jo0OCJfpWQA6Or/tFPaJ
XAxRcOq4qNzXQ1c1k2T9o+yn1R5DpSgQANR3Yl+sTdLCKspa5t5kRbLleYFBLL918qV2kPCQ1h2N
MtBKRf2EB3XKPKs+ZsxUdWzN7pLPyOrLXJrezLTP4dwWDGpKSxkrCJvG1sVbB5+mZ3ZLrRcLI+0y
hrkdRGsnY+nbsL1n3cTwtzGP2HmaWeMsgBUSWTGhc9HBYocRKvqNj0siscbN8kn/eGbWrmrMj7Ec
xfZCGCxpd+yHpcDPytT7HhlxzNIq2AN3//saCchh25yznDZYFG2W/DJTmhGAsxbZ5ralRBOk6s3t
HD55EAHrrOn1YdotZTb9ArdSbJsNivYybA+Fcmci+Mfu35E8TXegTDr7URYe+Y/Hhy606TSTEd/o
X/9Z9UZAJAmkOBAjtGT4VLV508gu/QNTXiCHTNhs1wQQpnitolsvKDgoPCICRuiAhMPq2Ime5Efk
rdVhw3OvnbW2viP+pH+rHUBcEWGFnbq++S5E/r6JPXjHpyYnRvOZmrAF8iXSQDKN+l+axm9SlPvL
agTHY/iIbtLBVpBMlFVWvbLV6b4oEkWNqCYaTElQt5FkvhltI6gPdjWzc6RdLPvn04K+kAC9l3qL
p2jTKpJzTsKIaSAf2vd+edP+MC/Rn65lrX2rserCJKmfIX9mm4r/BIfHOVbNBxXBSoP1EnUp/qG9
uRk+vLX/bRwi2gPwl719xGl7hcv7IZ4wEMErvhz8qU646SZDEpkpZhGrmfELTs6T6EmxI0kLoBRu
Z2aJbQByDzVnQRvantSxBU/y4VvuU+e2SRczndUyhD40BjhrsSBO7/ghGY8Ik24ArFwwFK2ZwulC
CdOLbbWG8kcZVlUPCuLpm4g1HP9E3+MpedHkn15gNy8DQBXMFyKTO+NIJfyWngNb4BsNVsaoCUdb
0+8W5RrG5U60PNzePFYsSbvPCNY7dSZWkkietHeaEthT5uBVa+jLxmit0luMGA9QX4jv+RUWn4ic
TKPcHqWJelH+RSCNvXf5uh78gIcXq3GbCeHiutH9CVPg7I/353bD15SP3rubXQ6bo8Ol3ot3lltd
eQQ/aGQUsM4kv76ofFR4Q/eUjGPi2gjYfWwTcCEr6Glb7WXCSYm6ZMdeCY5A/dZbcEUBT8dt3zti
rHVzbJDO8TpnkHXhK1F4j7s8VFMSYUY6uDir/UtQaPXsFdMgi5JH52E20qUhRY1+LYjF8Ec0S8YS
ewAjzycQtz69QYQoAS0mdYV0yS7el+MuUz/cdBIZDDvzYIu77+KfVKh3zvSuVdMXYJgG8yYeMYJx
hdogKkILYR1pd37ulzigf3shsC+gc4y7icZZLzpbTo3/jRGWHkVr05/PvjVOKY6JceY/4H9MazLw
KffLp2ok9Wwl1b5A3ae68ky9Dw1ckdZSUEXD4gSE26oLBYr4EdGZ+PpUbNFAOJ+2SXD5CKUG2TJm
hjE64C7437vR9m7DhBKxx56i4OE3P/vKlfCLjfWXu8SdYpyJQPxGMGdCKF1Xa5EojF8N4Rfv3EXE
27v6hkQDGMHHs7bQpYnj5QevB89V/veXMw+Ydp4iw7i+LhEv5+dZLA2+nBmkY6dqbTZAI6rHRvpP
Vke5qazIm4N1/h597OGukwr6fkFBNd6VEPeN05ByCMYzn1t7QG/96SE4cU5un9B1Ga7p/WakujXl
T6oBFkbJH00b+2GRLIJaT5v/DWc4kzbktFB+UIWAS7neWmM53ScNISqeZi/SQ8CCnuPwTqfM6dLQ
IHXeDRdPs1BY4scwH769BXDyVKCz0uCwRv40x82Q1yLZOzF4hrX9xJeOySeHNiI3x+EOL0GyBYJI
Mf5jkLPd0GOiwQmGN7J/IeWHngwPOqeUEU89k/Vpo5Y9s9qtFHKWmze7U0CszQI2pD/ZMZ334+Bn
oQUQShDqQo3J/KlWVrkm2zlq78kfkDuB+y7aPrHtZ+vJzySOG3ZY6zLE2q228cEpJM2cknSdFo6x
EP3QwCJMIQyOulPWGBhmC3k9xnMLh29baDEHBE/FyJAr6rd/FxUA7SI7kIFw8MtcMPaBo0/dGdkc
jctmBNmIoOyM2vFFZqvm/obIw0n7ipz7YAU/mxLSemSJMG8F6dunfeS9ePZ/aWoOZTLjVh8x8586
8XNF5Y4D1di88oQ8wntH1M4BncPfT2ls2xqWLlpxqDHjYUMIlenAqFXwK9Pn0Oc6uMr2TEZgxDdw
szkcyW7ZaQFuUE34F+LpykE4NlXD8uvk3YTi6keT+gS/V7pDNmBGAh4ESSZQvuu3ddj68A5Cf7jq
K/+HusqOjDHhG+G09BfeqndxD4+IraKUb2EulQXJnTf5KzZokDcYydpDIFQ69ACvb9IfkztuTydP
8+PJRLph6OozUufc09RTKAmsfZqnbjKohYH6m7e363eqkOGReqjI04YOSa74bS/NPbmkTCaBjXER
KmC4+RHDfm/h2WC22COokR+0qKA3S61a1bg5m2NpL3SQEymEUtvePd+3UzwjlsORBa3tFPz9C1d0
sEWTOvUB80Dl7+q8EeNXx/u3ZleqJDxok3/uinm84Qp20VDe/eezWUW1VFYIri85HflNDBMQJyZv
aLuIY6jtUaaMrHrxxCz8C19pVBMfmV1GZ/g3rpdQMrfeiO+YKw7Bb6X02H0pu/zVe3QvRYofHqZH
mGJEU78ABCQwcsRSD8PqilT5iT2bCzUevNd+At+ch578PtOeYP7XD0gYd5xJBpa9u+pPEpj2tWgL
kGaEm97yPAqRGpHhqtjGFKpoiRIO7FBMVEvO4qDlgjR3buyfv+LVfDmsKg+iQBIm6Cl4HbjvOz/w
MgnULA2/FhfRF9+1qL+juKRzv2g5YSzUaQ+xnD5sz/bm/0BzaXdMclKD2wAjIRQ5Q9B1nW918Yiv
T+61nv9P9fwLFJiY8K0cYxYPF/vNpUUXOYUwxFniKSd+ihhMNoIy79RYSpDmjoHCrsBkS6IbUsVS
TIGrP82lAWPAZSpqDIti8YSXIvRU1WGfOUFcPg5xt36CqYoPxePQCYDeOuciyD/3/0XJSfV9w6/0
Ms4zkHLsel8DHFze/T3CLBMnfFEs4KmIFnP7V47RliX9ta/19zxpv3pZaPeS4y5KibGdHy5gx5IY
KWrgQIaBRVJjj3yGwTMBHnFpD+2vclkwIyAy5urSEcnh1IfO6n7Rh/TS5p5sVGRpm7k4ckbY0YuE
leuvpSQyRSBgIMKOIHcl/XswLBy+thJCZCOyUFBAQkc+B7qhxJxwG6vbPvcgMr2ljGcQ07muyQ3z
s/4MjaWy+I6p+6CnTXg1QIimz2/rLwOG8MeZJss8qy/Ca3IBaDjshnxCK+pw/Ey3Adz9t2Rftk49
dzcEJqWDKpkM4gNxek2FZdi/LubBHF9U16FCYTdXsBjsQgE0CYlOL76BCqw1NQs7Fm/Xo7RG4MU5
dUK91ipWmdxE1Y/h4H9a5uGkpL+FiFeFoBnjfLPcPuSagnnTfIiJtrDwE47SstMKN3KSvAawDwm7
FqNsfKEVXthC+424iwbaGzt4lykbblGufKGLiZqBEKvOY3QB58egGfqX+p7VEi6k2c63c2j02/NI
NmXZIFNsFqPEj/3WbRokYFc/615p7wMIU7G+3AZ8pzSUWrpC7JlSTdHfeExttMNYhsnj5A1W+f7U
5TqgCfLPt8Xo5hCrVBTRi6SzHEHCy2nsTdkXRY+5SEY3iS+tcBwtZEbipeupMpnrqhFKgyPO6TC7
DFTgRqGcKLz9zkxmkB0DUeEGDWkzGez5c4XWXKSqJa8dkOFpq9zOZ9zQQ5ugWllXvl8zxANMFyWg
Csr1qw+YHgfrevSQ9C3H+jMves9j+JIzR16qAITJWavfl12yRyfIBHuQRiPJXSnh+wm1eFfR5aBU
c6qEpR22w2pxKpbkXn9yYuWeIW99OLb9oQ3nq/ztJlmWrEZSEsPgLc7ucI0uOBK7yWMXfeWDBnoQ
8NeF4asoPGXdFOI0Yvma4p6IL52UaVCKWQkykQSCQ57ZDm9iR0VVAXcF3EanYz/RBqlMUgpFP0v2
D6Ae+ivoT35z5VNUC1emIJ2Xi9Coz9WlYJf1vnwnPNllvpc1kaC7rLWinRrDROP46MEn4g4h9w9i
AxEsfWyIjSULivlBRbczMlcSKIG7lS1EXcnGJ3sh3HNnKM1cVPcDaRXfMk7wgo/EiY+2y80wqnWS
5E68sL/yRjTVTNDlU60gmXwyjP4cXb42Wgl9nJWxXPk21mxTjyCidQR8/vucpzkXMZ1wAAGBAtfZ
YBE6scYI1BR9sa3TlLNpO7i7q4tBuxdb8DddayZ38RlIVVZ3zVDTdESRAu8gJAm4cBaruhJwBJnA
OccYEwlCoTEVYARhc/vxgPNLkt0Br0QN6Fe3Sc+SPKYryHcRipAqDJSsMoS+g2zSBRHWsK8BLDdi
6AVJiejmgSsQoy/ccI3VvvWihgo9MdyW4LyxwL+8gRcItJW5ink+NV8D56gLUvqmSKtO6Rg8UjKL
RjPu/P4AEcyKO8hWwll6sNJzfDiT8ehJGPTGQI9HboiMhDkksSCzHrrYRke2UMbSApdIdPxll1/3
Crw0VtTAdq863xTijkpQjqJzwCym9kcizU6r1NISlW/xxhMM98RnpuHTM6zNaJ1YDFSMMfo04taB
kJ1Scs//9+b+KNQijLUNKqFXepuviSXvfpu2OxRaec+j9mvBcel5LUyQChOWEzezCUPlp1gu+Sgd
hhTtDcPVcqyTmYMl8sW7aRE0YZohCBwqXhWpMYsAN1GMyoaXw8Vopo+JSXXCN9VGMHUw19/EiLfX
+xVct7UOHIGi7ocZRTdwckHfziejv3hmvmCzSdW+YmMO8BXgdZjiW+EM6V96iwFHvTC58JbjPQxQ
7yk1vTyRkJyb6oHhE0qTQ25KxsDnETWBFQFhZ7cJ6kkl9usIcgj5c+7/htaGWyCqV0acL0XgTUcg
G+ACOfrWhl7K+1hhTd7gUoBGpFSFHDLapMmuB6ixAP8lCCq9tyNC/rU1cuQycVVztf8vclfJwMI6
LJAfuRgghtrDNcmOUL+P678nBZxtBw9eI1D9xkPTUP0BFfaqOnnlriJ/JCx3dMCB3qlpiJzPKKh5
sUguqUu1MZ4yvVoYd0xcch6h2gDGlIN6JPDyFIyyaMl42qyagOa6ZURfDAXooruoTUmJPCppgyoD
XatsTTyZN4e5NxhuRLjH8vJa3Fx1P8n1XwMir4rj+mSLUGxhUabojA8SW2hcZK7+r676QsMHyOuS
WJ8W1Yt67smJE3qXbdbyz4VJ1NC0zEA9ndYugg83rv58LVhcS3DSk/uvFE7q9xQBtys8LqN8cNSd
Gc9HjMdHNOi8X4Ua+IIhG/GiQ556aGdcf+hTsisHfASV7kCjp1YeCv6a5eCagS35PW48W5iZUd6t
s4pMn9f3w6d8ZSxdMoXNDXHeOgMEh+avqeuJIHBqA0b11q4D+pSUkOC5dQvS5zuOVvukKKNXuvOE
lyVCxt2VQYaz/S+0arlyWhewTOcHEohbTYg9M6Zf54l3SiFbzV04o15ikd692GZqNDeC6lMqNhN2
F2Fa8ixnmMxA1zvfWSroW5lEQWf3WgcLQQfEexxiHa1NJ9rLxSL64ozmPyAJAZmnnHXv+RrpivRr
HAOA18w93ZskZkLH3Wzfqr51qZCa3zpYnQ0FMvpEnstfTxreMCLJB1DKiup0OAntxJvhCX/tSZ9Q
sQ2e+d0rpO+GFBV49vRpMgkjD6F5iAUeuvTAWaqZsPjZrE9Co3bQ49H4b9bIYqQjeatrOjvmiqpm
SZKuzG0mzj/lrLQsM4LRFFNSnRBvLwyH/AzgWBRPEJ5dzcxGHZy5/F2V1tOTsHvBpHHWBENfDh5y
aHclxOy0Mmifz7taab/qO5x9S0jJcE093sqZLmwwKbBcutjrhSXQyOOCdcXNxab5tefST8NZGhcf
vKl/2z2pkGf4qjrgvZxZiJdRfAd/HvsSepfNqnn+swcjwCONopZ5DpkO5jeJlE/rZXGSbe/v2Bil
W7GMMStOAaW6B5v5IXo5FIaIbkyxjR8kPLOVoWRqVlNtZToRztrysbjH8pOrRq5SdigAEwb4jLfJ
cQgGxzNJ+B7URue0Zd9rlhg1EcC9oyHDjZYlKki2v7f6O47jFYIjpSDQuIr0c0R7/qtDs6eUsY3F
M8s9QDf7ZNZycps4MLGd9iVDqVhPVSWhB8anvP4H2jVl74XwCpL5NSBVGe5eDluIJgT/wjPk1fet
GVrxgSQPmLwJW54/c5HyWQjJF6UJ4snQ5kiyS6/TnZcEYgW052gPDWouqH41NypRURtzgrYa4369
bACdLNmzajW4O53ydE6fWl1uRPDscF/eSkqtaf2J/B5c+WX7iLQsdyIKPgOCi6HUfyr+Xfb7uO8g
vr5rip4XV8NPf//+Q9dFBvFv/sXbIbI6gfQBZpmlTvqhURCehmGWG0PEiRZdOE0LOyNTd+B+TZCj
Lsarr/XeKMmmNy+BPCF654qA0Lr1EeDpsPIrwGuLGraJplVWTn5mQfGeWYZHJF4cuhbciRBiRjNx
R7xQ/NjdlsT4q0Bz/VtrJpA4EFOblqMeRN5a9E38i/iD66R9Av4PRwjCkNgO19OIq3h4seC0MkgQ
jrBXumIKhBkk0rvW5/TKlLc1m+N9GbouXAIsP3Pu5spy9Ahl4YRj0dzUh9j4cRWYYt5crndSIGF8
TSiHp/7d2hnziP4n2e20mRM6dhoAigKfFkD+VobSDibBkv4EFfCl7GbQZHjkoOU82mObmjzuBfl7
dn50e/m+kDq03yDCBXTAVQljGZjnZ2juu4j5HChEYKM92DBueeAjfeB7CM1VmAfQMerXvWEtAJ3H
q6Cq89eCCTbCJzzHUOS36AdS2lMKi7ZDzDRdoZEa3yZ16MFFn5hzi3TSL/8/7X1kWQAM8v2Qy3qt
/7rAXf9gKvXowNvVwxI74psmzBFhpGVjgDYP9YHGWAx4bMpXEU4gIoUJDL5pUvxn7uFSLhgNFlwJ
sV+bzB5eppnWDeOC1hAJE/2ZT7iD2oJ8P8jtUMbtMBEy+/TLa0PvwDTNmTJu2rFSu5D5Z5LAl3P4
irFAJht+Bzkn8Bl+qP0FFnNaxue36090kjXkmo1l/tmhU9+cKWxOlBJApP7NTw9tTUKNvEztCsWU
//6EECuq3auPftOWdVoZZJ1svRSH25m+MGLndqc7FA65bP+f1Nw1jSMVSGCrXbdjnGywvPK8DGuG
/OYrSNZA++li7x/HIdlCk/1DfkbS6zB+76PQBLfvnKCF+QuBrm7vMFe24IN6x7tY8h7cDRP2Be/v
tqriI2VmvcNE+oaov4xM7/igDyCsdB1RoQSLc/oR1BlpUFdyHvvzBI2DS5O2v64f/Mnyog+456u3
sBDSsgRQPt4hGVFdti7HmAgNwvrogW8GV0BlpkMD2Xyf99PeGzpIHpN7686e7C1hh8VnovstIQ79
6DAFRf7LXyI+oPTCiaWasvlT9WX28S3C5+ovD/a7ElewA9cQClf3ea9+2Sor1Q1BSznihxOilIGZ
hYhEhHnz3mi3OtHF/ZGy0gYhaKKa4gRDF/lndtwaHxvVM2FCMpigJfoG2NBzDgKGx31CEdVZzKwU
wD/5da3hxIP5Tm8vN4Wzjwau96oTtbCjSX0EFEJhfo1sVVvj2ykTsZGvEFfArI/QpFhzSLkCdn5R
NIinvR5w7XPym6t1xRNCAw/NU5z4Jm+LEDHALcmEBTT5ZU5Oml0cYMrjn/yei8GcyAm2b/hl6AMx
HcyNCFNwgDMunoATm2HQMACxAY7jEegS0JbuWyjMHGflI0BLmNzlVWb+9qNc8EHtvAPE9voGUW1n
nIM/iOgdcnEPd98rZ2Po4hb/8t3QPa5wAR7t7I2Lv8a+xD/1GkJVB55aQMrSUL6hfUtBAYFWjO2M
y+d/TaV/IxcjizKM2Rp+mpx0f8ZWfAD4+H3VCbHAcvBED3d3jr2hOpwXTyfAZo48VNBeyxByAwbB
yGd2yvG9A2U7q7gutUXCrWhIvi6xddB6s4bL+ZH3Fzl3ZqnOatd7aKcXOaB9T3aFlgebY35xk5XB
yYqzUiFdKrrJmuo456WAEbR7Je4Xs7u1p+zceQA2TSHAzg/xEptI+7xzEbTsFGiYsDoe7so9gz8b
pPbqezVDuub2Eswu8LOSOturxGgqfoNZ7/x3czt9UNS47xLyN23x7Ji7+n1v/+ijOnI4+Zc5rCmT
RW42CPL9uU92YI7LvM473S0iIJBiuXtKQcNucf1VCYFGeU1sz7Dq7eKXp5CvfVVPHb7a0InT4XB9
Uw0kvL7zmoQajHGafPC/Y1xJesL73uRuRJbpqssJ6bDdlmaNLduikvlKIkNKGp7O8TY4uq6L45g3
0y73J1f5tc87gMcO9p1xunJWoxz0Hv6+UnjVdx2wKhet/IQ3unzXJF7/qsCmHydVktKnvhcg2Um9
A8uZCkQoj+7C+FiBjxh7Z4vNmlYRKAmyUI/EodfWGHo7GkrL6RTfqYhQQTKChLNDE4vO6q7xCfKB
Yplf1K18EDLjJ5007G/wGVUIkjBcuBTU3k2A0iYspUNCMSEe9Oazd6cFoobTLm+a3rzakb/yYPG7
5fCMxoHPmpLXldUrG08SIuqD56rvmHtFcvSfJT6ddXQZvr6oekbIdBdazG4igm1NxAQwHVufjjOi
K2OQJYXqlmJSs81XzU95XcobGUoGdrBfNCEk6en6869TT4RkYOix7DjPtzNt/QkAV6G5/VRaz2Dn
PHJ+znCeYcPcA2r8qmW7DvkckkUN6EEByWREUYSd009mbe5djf29ocyLqWKpWXNtscDwsT24NLI3
m8E+uTiU+eUpv0Y8s6k+LYqMPmKg3sDpolzWFELzqToL85qny2vsQflr1k1hb8QXCnHLFJmOoArA
sjHnAIM0BGUYsfFO07Lj5uD0YD+9tFMcwis7Z6dlFRXInF3PLwcC0SscaN8ebzeXRoOHuFtjkkMt
yBdEOKdfvuGohsXpnek4zC+AkTWljekZN3Zvrp1262SINEsNcjp8oy+OdM5FrHYMqHBVxp2KldNL
sC3MYT555TQb39y9Cq//1dddbs3l8VBozOxugjS3E7yXiqJfALqpBYhAxFMD+yF7OwjautKp5zr2
LKgD1FpM1IA3eCQ0fi2dyln6DQ9EAKrH3MEWnLjvm7320oxcj5abTH1N98dvshEJIxNuloIvXfRm
k+JVP/RFgCTq+QybZe6E/7k0M+eU8TQ6FF8WcE/G4zWD60Vv/AzXX/FWC2Kfsbjd0CC+Ka/pYYRM
4eKLwEUq43myNwi2kswu2+lERp+xSWb3OqjJyJarrTUp2S/AGmokemc2W2sdT+i9eChvAvn/maow
k3lTt/YapduaIrP2wq66twQHv4itD/Iz0/Nt4+cCOAxuSUq6UAVL6Iw6KuT1TleJFZeSvlddsCFp
WsTjtMTSYLstpYAMW9N6k41GyGTI8wIHV/wnz6nspqdjolNcn9O//qQFUtaYEdFcYSu9bA9Rxt2L
x2CvYiglxIDz0vO2geyMaUAHayU8hRN2ZygzPl7MX86mJDBU5U4Nk9fIDh4GXygP4loWsmZE71LI
kfbrArsTVqg4Qa0RxZAYVsLJiRhub03txaTjNWjCtHgYWUVCsEPvldjzJ957GFWUWiLNJTmSamS+
hscP7w9rM/AajBlmOUUH/rAOCZaL92mlKc7s33FZIz9KWij3VYMAn7hY0zKDlVbiv5aWTxlM4r1r
zLLWMz7A/FRPuKheUiSXxg0ywke2RlOYKn1mqkxvthCUCK6LIVVUHZpCDmW78xCQV3m3b7xxaMSE
eqOyJox4xS2WV0CIr15imkdGPbysfYtnrKbBhlzawm8LtZ6F7+f5KjuBtvIZUOOZJ+2UOM+Y97xd
9L9bIAn5B53ufsQeTFqBMVz4VSs4ZsRKfj5IscBuGxddZSOTfq9CrHOUEVkj14tih/xzjDBTow7M
2rQ/0x9tW8ReHo8h5VeD0vU06BLRS8f63WOYS8R1LZvGNYJ/ZSbq21uHfQU/G0Z5J8uAncS3YI9M
hOt2s9CFJ5oCteO0Bov3OxL/gsfzPhCQt4xIeDU7JA3dk3nCwwtKnPssbjhUtbAy48g8K+WPw+T5
hW1YeRLHUi80Rx2jlBlecJCR/QULwkmxbJC8+YVvM6XbJiUm+9QSlyIP4kDc5I3LiH3yJ0tyzFux
cCkh/nVyt/45+lWyLxiC/rz8ayRrC8Cb/FEuk7G9TGtNhsw2GYIfE0nGKOdmo+IS/GfW6KVneiCl
KaWMSh4xrmNHqzC8lWpjglG4DPNBSUWtrCQoM5NTrfNjNuOwSR+tPZXOGa6c2jLhVxiIqOAKh2PW
ryEQ5WNjnns7EMsXmJc/4hPGKWFNEISnhO0mFzUc4UyF79EW6Zugxe5AobWoltrQzNaQWaubyeKM
QhFjghendQidxAwk/SQ48lutT606kqBmU/A86E1gSOucHkEusYCPO+T+nHIUaS3OXfRt3MPxT3w/
TVxYikY13tbldkv1dT5TgA0Av20P1TVxpzTtnpEsY6t6nVsNViGFqk5+GtuSqiSapVRmFoH6g6fC
ViRLX3FKZGA6kfQEJ1cnTne2Y+XnEsxGb9X20LB2xt2+RAOFnXljEHUAZ8luozqXKWD94Tts2Hb5
TLdmQW0DfCBqPk0tMCQFVBd3Wzp57w67/oOgrAlbk0c975/++etpuDKF50B60jS6D1jBOY8JY+rO
jYhSrjfmfFQDUMa1VcohIGC0N6LN/rTUwcpED37oilNHHTylJU/7raWtj0Ch4vp4s2D4TfZiHRng
ElIOu/CI9fq5L6K8oHSGL/XxIn+SiNR1IwIAXqrvlvzMJ4z9Z0qj15dvhErwpErhPBLhQ8E7u/5N
jbFNdtqju9Sl/vasME74bKRHC6uRAB5bWCstNIaN08o05rHfuUVvlZyHxf6BouFmDV72eox+awAQ
BA1rAU232ZCFt4lCBWe3lfQIrF3YHnR/m4OXvrtrVqmAqcWGZ2AiauC7SyJiWVqD0IOD4zfuHV5a
bsQFfPALDa0dkX6n8GXqlxCok99LHS8taQ3xyk96Zn7lQ6Ubxf2wObUD6/ceReHPL/8KquRML7A2
cX0MP4zwsprso7mZOLQe8i2y0fmf8mJXcC+k8GYwk4Zd4HA9gQyUq+AVqGKULs3GH+x6O1FznhwO
c4vYdL54GOgkmj+gGdA0U1lUgoolqw6XowT9F+g64qLMlqyEoyH0PKJ8YQnmPqqnOj4TfjzuHyAP
RAEUlXVM+qyrMm5Yeaa+ywVBXCSdE2njxGW4HAePt4lS0Mt9oDk1ZheM7Wf3etsHJR9QjQkc5bJF
RTeaH8PHv9UMmeW2MfsLX4fJJ+3jliTijJwW6xV0ftZJP+ErFXfeoXXo15InT7KScbbJM5ZS0r2e
okBW9eXkdu6Lp3ob2bxmIdGEelDWyXDr/nattlVTqye4NBSte1o1wb6G3N2bCYB4/ZXUT0i7y++g
3m/Hqwj3LV2ynj46Iq0iN98tG5OuQU00Dggv/uFSsBFPfjlnu6KGWafVGtEYd9QnpUrFW7g1A7Ou
1EH0KyKxKOZjbNy74uIqchLVHJI43khHEgE2UQas4y4E369J0OnVES7BCkPMneI0vE64N5vKNQT1
mrCUX5MJAB/3g001Ftcb04Mkwrp4eAxpqATNt/ayO9TIR3HY7WXnl/L7p9QIaGFuNiYqjKjaf4n8
HNu92ANxo6lFK+EMBE1/v7m8P3I14hcskByG3Qy0PpmMiS8/FEBVO+auPU70S7gcHLuAZoX1Kj+u
I6yqh9QenaHyFBFFIhqRkDNRIFQDwJal9uN2YHt+u1KHwMU8eCLA0mScOsQidJlpy0AgtnX7sK4b
fWomWs9QjSFkKI+lDpkbiaXktftRv/aAk0hYAGgwrMXpQ3kx4Cr6f4EOh3Iu0OST9bd32ihou34S
6k3lOS7JQ3cpEtzOEyfY9VjT9EoKnZ2Kp8Ap8KV+cVNDSOlu0cMRNuT7AJwo5oHLKntlIc9hYUxU
WCqtJWaTwZb0reZtPX21ApeLoXwT/iNN38gRI0AAoe+vpeLdMcWIHziiVLAZAyKKXdMC60SW26SF
w46fWziPENh+jmbAdUTlPdQtGqz+8WsL6/U7pfCJ5V8Pq8yi6JIzjwu9O/P0KOL13C1+wHmpFYCO
kO6hPQqIj9W/NLLCuwK69n99sA8xLWeOEouw9v9VMQZkoPmNQbiIh7N2erQ4W0QHCe+SMW+KhLYS
ZiSmairuiPAqta3GZE0ty/kWH9pXvD+W/ikndDPuDsONz/bseqUP9i/gIS8SufsoM/J4z/AKURCc
miC8M1Wv0aNjT5az5R+QJOQDm5dpegArsot7wkgIEAo1Y6sT3802PjwV77nA51Qima1TR243euPr
+9ssvs2/LpHlcTKqDybtwWZqH+KylReNWqLoR+Yy3hW7l6CbBGXLTw98xQjFgh+Dz82OguS0o5uJ
BcQsMjEIz2Hz7i/jfx1pVFE5wncMqqwG3EMBwBEd6veoCNxHtUfkFksJS+RZhaveUrLmh6B0cTBG
IduMxt4WN7EDfQW+gpskLjMjZ0fl1mmuaYfujzCe3T2ugG4oSO6hYcjuES5DIp+/3EFiauSQnZJ4
2zCrXN423wx+ixqI5v+EaZb2DEBGlNFSKcNkpmsJE6yZzu2ur3mXKIdSnLw79YTEcZnA4Yy5Dkmd
iIRUmGgEqg9CtRwOhbgJ9+aq35k2YhAXqy87zVfNkapMkWqNLDZpkPviGD0CKXcYaGbBhGq278gu
1d4AFX4OIEsITQLJV6MCEEZBCzD/9J8sMR3ekDEG48NJNF1w06NmliGtB1KD1ydNhqda6VRUutxS
Gii+jm5jlCt5LbHTYpViA9HhJcLqvAJJ4EZYHjsiguC0mqNgizhCve5P3ecKbXKYFJSY0osCvHB9
9+ijoyAkR0r60ezYBA+9wk+OOKW3QWSksgSeRIoijOc5Ds2+r/iPvZh8iMPMDZQNkmT0E1WY83aC
ZTWJ1KKDhO0CqWY7JZAeO67elWmNI7zfEClXWj4vvRDDLvQqOLVBXDFcrl2KfI071uZkgnvptb/t
xFVH981ZgrYYNCxFxc7nQB6yQpx3awmoyrm4qTm8IFZZ7AApeYDd0Xqo+RniGtDSUpANIfrXLphj
7J0QEslAExVziD8b/N8gEOfFJdqTXCBC5K9uD7ARyxZXUEAD1hy5ZNon6udRDzlL5yNxu4gm6U9Q
FUe0tqdSiFBsAN5H2BiDgnGcopveLFOuSIhE/x4RV0iu0qdIlL5QrIVLXb6T/7CJYMf9g2fcTIP4
/KCqf+3JqrOzNOsj93JRykW6au01bCkBCLtcSgc0Cu3OBauEyvMLMhOcK3nX8pv0wU8YfMVCQ+to
V8RSD/jc6cCOJf7ZGqb2NQezpAjemnv3ymXNogJFb02AHt7vlFAOjwveGICeFqd1n7FdWj9KmU2P
dA2nogT99ATzzYDML8YUSqrYJxCewmfZInz+NHeAByw+aXjMSahPGstm0Yxf7m5+WNiJC3vqCpEw
lLR8CgsADyR2ZgcAA610Fv69HUkFeJDm/Wk7QCisieZmHkDTSJllxtffmIyJR8+9DC5ZD3NGeaDb
Zdj6U429qJFHjDJ9HZlgch0EegDIbDnufwwxv2YoiST5fghqWRUeyiwwFZGRaDWAzCg+9qs4tb0V
vBi0ZSDoxBZx/wy72ZK7WkJQOWHO0t8SVpOGuuOk6mxxA55qOPBFiuMEF0sI2ePFM3wVMR/9B2IF
OtIl5YogWN1QVOZOzcJfqiKlWh27O4TA89DFAV9dT3aUrE/o2RGZUfMuf9Zvsj2lNoDKfMNgFaPS
huOGvu1apwae4y2iU7h9T9qRlPpK4/miGgY0+rOenpgUvICVPTQpVbBX/VNjCYmuKIwWas0hXvgE
rwbUrv75c3j6iwGQqdyMgntvlVqBAvZ915mwb7bQptdlPX0M+Nfq6RRdSHvSnBl0o87UMP5/nJYF
wnhlc1QjLoFcx7zwdONzMIwir8JaDGb1hNd5nFPhCridGPBuSPsZaHd8MsJ207IADOb9lgpFq/6Z
YQ/XKpjaWFi3dH2EXRtyTnShALRvpp40CL3EuAusqBG3GRlkdmD5Cu8YIF805hnB8/4F/22+zbCX
MZGZzDPZ2eol2Ogbqf+m+u0pwaPLcV1XTOel1zsSr1x3QwXAwlyqG0j2xH0jsLC+DNNeHF/gtQUi
J+63AZbynWKLYnYYuluQOOJyBdzmTHEhxVduIfc49vKRTLPGL6blNeJopZq4579EkexC7tvY6iD8
ndVA1MUwrDXlKLq1WDBIP6Qted79q0TF0u7XL85OV/WlhvfL5m2zCkkZKKgvOS5uXem5UFIWArPc
Vsm3nlPY2sd62EBOD2gwpC00hQEMzb1nq3Xwu5geSWuQdlhCMiWiE/DL9I7pTaNIuFf481ZYZ+aF
B5oAj8xZVV05Zlii3p1kv4SjAM+udiCXh6lZuhzWMz/bsUjtQzu4mL2t3ljy1wUCrmu9HpqqqICu
n53Ym77oo5zx2YVCU1/eP0VBq8vJJm2OR1KWFobtUud3qNzyahhZwUDHChfW/Av/xV9qsnbK1Haa
ADu2Lm/QxuasPFRKZ/koXj3c2jEAeG+o0GpTtt4hf0su9mhTw3swi0hdlHtbpaXPrADzEBLNU3Lj
rQQzJVJCr42MGXtwTs015E+8tZxzOZtKoXYtvhoJiq5H8OMyByTuTJyxuOL59gP2zimXV2TAGl77
vMdoEmZqSTL1jacpRwKK0pRzry1NMLT/4qgFmU4ZjBBdPdBrhKlGVW2kq2bLAdmsSYCfsJINAMBP
T1LpTHPNFB+6KwxocrRvriVftSi8OcAZ/yhQ3LQG2wURhufQaUPxWwFvEUgShxDDz68tPLIqJHTZ
maXWZihVuy3qb6f0GHgSjUMDsi9stofXWSbCMD0i0M85QMJh30ezsDh+SnYbPtulMmqMXIP5Cul9
Vn31zVMora+Sw9ZoX6s0+KiCPlTWUHTiXmmjOfbZ8Yf2PzqK1AhA7ffwT/x91hkI+GkaPjEAp8bo
jXZaIJIrc+D2hy4rcQZRR4940Hk7ASbn4lwHaauvxlslzaX0GC+3QQfLjn3nEc6gX+I3jY9xhYwI
tFaeP3D1+fY6/xCIFT+eHEGH5FzKXaJ8ocyE8OaOih5Q+olyRLImR2sj3gxv8CAGDdgjW8devvM1
165lKJnp916mjS/HDrNHdVQbCDIuOMPEgWkaAYRYfNyDulls2l4rp4kv9TdFRiuyEPzys0Hq7Jh6
dTTIHDNXvyMMjTdOo5BuKwnOVxc9hjlaOUnXAky2Gc4CnVHW/EcDjBQMHJH1dn2RR4hA7HtM80sp
efCX18mbnARZsSM+AAy/6tuyzgid6HZyvXGe2Xd6R+cJvj1eWrRSFYVzMtDIpNBTPw1AcEUHVvMT
Nhjiirntg82XecORSw5reemjUEuQxu5JCvU5ktAMFkA/QjEww+zto0wwm0FIHQVJDeuAUkDeUny1
RJPCtzf2xJIFWuzpC2AMHCR/CwRzjxgktb7fsiFLXHCm8ClY6a9GCeqwVg8wBZN6aiByivdYe+jC
U9Tyd3E0ItEJLBriDaw3ZqKfoZ4BWD09IeMmlt3x4xP1HOd9H4b9Fultq7Gosp1Kp8KIX8VkS53B
exUHxWYVbpuBgwvFeIEBkMXvaSgpxKqoj6bcZbpgulTonw5h6M7mkLKtRlUd4Ztez/W3YbJh/mb2
04pIrrorV/yCshBlqHGRWh541Ntww2SwKV417PbOPgpnCd3pSkw+DQ6CxSTRuqanroz+2uxNSasR
lI0JxA5flXT/4Q8/6Abpg6JclEy40+ot5YTSxuzXyu+4L+cmx5mfiHKchzHvXLMqnFcWLnAp6EjW
0KbsKLRow1KzpuCrfsEuKavnQoCL2NVK94K8hiWZzORxOjXxvLNr99Q8Rpnqb0Yv1A0+hCkXq49w
8hEY+zph9VwnRjRZUR4qMq37TC+HjKA95BgItj0EepaTtpotE/QWGt9GVsxv1WHCb8CyUI4QB0JM
G0N99Vsof1ZQljRwKVpHkRY5bRDYLyolJasxU+duy1fLpeduQyizkFaP9eQSeB7olWMfMQJ/tywM
pqgQvU4EzPEVGQfzU5dg4GDUqMQqJ9pKRXk1BbGjXkmGl9VcRwhCIeOXwsZ3ZTW4iNDoqb2jId4C
xzBcJtcrZsbtBFUl0GXvAKQ1Iq31MqE6agYHv81JUVPcp+TixticuB+ujRAEWsnzMKRfsuwupJDs
ArQDAu0ajVMp/rWEiMJwj3hMPib2Y34Nday1EQ6tkCAJGvx5E91hfvw7vm0HQTaSBfVYMM+/aNo4
BtmMRLb1kbFFqOiQS5IlJC0HY8DC2CKGj/AqKlTCanMl0W1bgqJBDXIDOfGNrMYa/hKyvnf5OVod
fRFK33dM/5YD+7WDWyLf1pEze1ktRjuj/sN1AKIO7vbKxDR2sk+JwqGeBl5HWLNcC0pAWM+NRQjt
sBDSDDCYzMQFiXP+Us2p+IRQeu6z2PqG1NWrx+F+nToc4pzQrq5nWDSWuHW2qupSLOM0176KJcfN
HBoIz7S39TljMAU0rV7uDr7njobDcCe+AGJXJSYduwVdiM1nHc8XDlhqZHWNTx6KCae2EI7L1pkT
Rey5n3CP9GRvfy7c37mHQCJ1C0snlQCzHcyj52tZQsMfIkwr6r6jTqeXeMXDC4nGHQOKykKF3sFO
jynXwpPFwzOcXk0pQeLDMmZ+Tzy9SLYBG6nPDoI/AASRjjJrlnDE3b4wdxc9aHduXIzz70sBmSY+
XXdmxF9xCijduSIQ0oiRMfd9KMrwZden6gdTBOFjainif4BvqbiWLKmwriVWB5acsk3A+TocRVZx
0bWsuBUzOvd1BNcqv6w1AB1bfZXkKF/D+tQBIHRNIeGHHHYHIoc0ygQFrpwOomv3d6yBBEw3Wivq
3mApfk8H28MDHj5/c5mQ2lLWHKlvwtq+g7CDPE8ln/rwxwOJ10BP0PVV1TQtFwSI6GvZ30uWvkmE
52BQYxiAJ61zJGDKFkiJqockNWXNAQhrzEf/B1m9QrjuJvozmrEgQgfvUZrHXiEDE2AXk5ZDwdLv
PoxnWcqhRnnukwvn9YFeOJysBI3dMk2QwdV+ZCxziidEC99p1xbNkITXwcV20oAIcFm/OH9JxqAa
Qv+D2KeiNwkFT9iR2tIdEfsHAYtWbBmcdwalVDxD7uNKkiyIvypn0hsikEs+8j3SqsWJzWQ8HFf6
Lu+JFe+Z3x4XcUm5ZiDmAcJA9qad2C/Dpr0Rahcq6ZSxi9RVGICVMRefv+yq0ULS7AAcXEGt5aKL
Znq5ZolzDX0isbCmJJVdmJ4koPCSslPTsEER/IP0ZaYr8YyQ/05TOLZ/vvF951qwuYD+cqgmDMP/
Du9NIAwjKZMWRenFD85llqYT4aJJc3oeaWvsZBuTMLEEIjbb9ysOWtz5Mt+RHICbRYbilDMfZm7i
QUjIVW3IywRF/dFe+tzhNDnubM0eMu/41tzVHb48izPir5Fzwhtq2xrTnz5YOxxN5TlFVQcRcKM8
6E65bX/bHx2+gxaCSbWP05Ei9tZlWD99b3i0q/pa4ijh0a6udwFa4aqWIxO/5MmIhk+f2MEOZJWG
nAS6FWhx9SDyyU/LAHD1yU4BvRyldC2142GRWA+uZ1zahfZ4mDlwUuyW4Gl27cJDhBKKbOptead9
Dv4BDgS4oRG5eGDVaCdybl3YEgQELa8agIJ1HAj2Mrrx6jBo694SomOT4dfOrOAFsOjxeZ4uVSs5
oH6dO1QtJKey6N5rGv4vxGmBrw6aDCsynvFBnmNS8I4r6tnFuQQkqYbvIdM/nnqjhpEZBBimKoNW
LFiRg6FQgzKielmn0lPUc3bqaXCANY/Yh7evKHf2nt7JwSQdRliDs97H4n0ISnb6Vi7Bpw1PB0tY
KaebebUBCju1HyIUmUJRYiNldIsqTM8S8eBEsEjxlKWJ0YF3uIL1SY41ZRq/84QPQHq++OnHcbOv
v9LkJlqYuN+BFDgfx6moVAVyFxzuzE8DDKR/3o1u/xV7VVYP26M8ZiIhdAevsTgO8JGeb7P/ii9o
s7Mul1GOzHi6qJzOyfz7lpP0gk5gGZojrmn1s3b3u79p0YIrbxecLNVgdNFqKIJNAFdgr40M8Zio
905uG0JtDkDrxK38hT7c7DJxaouXzfYkeYeaRxQOXyLDGDlnBiucchxvsxEmAwAnqGhq8w7y7MVB
e1ixmwQX7p3BDPGIQ7iWFifM8pAls/iCprTtbcXkiACTh28cLerFCmIBD/gYLh3/L4ra43qE025L
dNSNke5gIBNW7kKbXuPVCiSISKUq/iGtkVzzhoRncV2HYfJea4ahSDlSuaZPLdhazwxfOAzmSCIi
tV7d3TBhBCjym1Fw479pAgKGp1fyfoUGh/EOcVDB4a4k+07SjkAXYQsHaDPtmEIhdDLENkqwBKwz
VFtefbP7m1oql/+z4lZat3zlXuJrPILmDDORs+NoeW0y2aWDw7RNrvAUZRKOnEYwdDEYsHOmunGX
N6nXtuQ8b6AJXwWhL6E774B64Du7b076bA8e1RAKb21iu/7wukt63LnBZvah4ueqSwoyYdr1rV16
17PR1wSdaGV3mf77qhGroiT4cVC3uTqcVNo0Ka387Fbl8l/pI+xt1Xidd4s2cA7GsetwAggvL1Ep
OOhwQrpbpqN5PabLPG99GfVGskAm6/Qo6dORcPEOeHs6Z3CHN0p0a7Bm4y7Ojgn7NNNtK35aZ1Sl
ZNNJcwKu57481fuNXv9V14W6QOzo8NqY5ysk3/rAC2NFh/+wIoDMzUKRJxEMmD/bRa9HwgIbWFrg
nrHp6RciKL0nTwp4vxwPzYwdX18dzUbvoX2PhNLoz+zKLt9ubju5nNVy2mbsh7p/TxQhPj1jN3ML
GJkCeALFB3hWOy5aFgA/VxbOaw1lhe0jyuVg+G733aiMm3Zh4mfuF0vU/gDsWuiHGiX69Xz1E8aa
ZvkRIOSkgyYkWrJ25yAOp1pCNpvd0YDdXTzASeWgjonR/ny2ddloMbhFmDurmMRmSM2MW7ACfrL7
v24uN8FsAOC14IldIN/X8+LEDlxbjloDw7o9Md/oIKm+RKPCJfFffvx6NcL/HlfzNFq44dgD70nU
WWDzSLu7N9WJDBZ8CP7YrYnduPSISY/B71tFR1/Y8jqlOsIvweLAzOs47I1FR5WOfeor+iYRC7Cm
SnZg61bYkfbcZvjvS03rBGtMu1HbwF1mU07DLhc9EyZD16zWUOAZxJltWslraqmCTeD+td9xjBx8
M4MVOs5uaH369XymJfM0FOEohg+gYd8C/GzyWbiAZU2AvMnIKXct7/VKCLePH37o+1uKLP4OUKlb
DCM7qoMi+rfYpXoKK//nAoBQp+uzWo81/rcsjV7AEc5d40T8KIGCrygpbk+Lpf25DUNNIUeo3fIo
a8bRxopizHo2cyHs+2ni8649yrG9BJUDXzBcs90EbQSg+xTHxhCkKgITUdyWrAUNCHcafCaF3Qa8
OmX0NkRvFRjIh/xIMMSzzLDHCYz55UyBCZzxyWlsLn1gUmtvwg6B0TIDZyPf9uqMPwAYXFOd5wKA
FExyDn3OrwusTHf04f5pATv9A+bXBV6En6trvAJ7LIKnibBPxdC763gycb9gD8wkuuf6ej7SqRfX
IEDqu1fHJBcRIXTCB7fz2gENJO2nuvgub48kyWSSyBt6jZJm7KFUYIWgbFJDb0yOZKEsA2N0lSSc
Ns73Fk+nuwqg3MmiaqyK5PuJzfQ1JKYk3r+ZI1c+7aJsHNV9SlmaxYyXYiTeLujGPGyqfk/H674u
4cIlQDseDHDYB8bunJ3aDopO3SmBGkSaRR3QOObkWMlm5E0Z3ST3g9WIOiY7Arrj2TFYBR15eAgF
eoz5O570M10P5ImkvrJqBYBPA1E48MGB7n5q4xCtVrl3p2GDMbXQFSlaVk52gfihuRGYjKDAKQTR
n4f7bmOqU44X3l4huc9lgkTa51nFV3OVZHtNyjbGYLV/gkeDUZJlOB/3uVYA1oMkjfrWZQJ7Z/FK
doqpLcKz02EU9B6tllwsa1nw1kzdKdCxsXF10l7hZmZ4lgVWJKCM2Advsh5VZlx38W0pFRV5EWac
d1rcHJH3uyNVZc5LOx6FZrFjVHEv44u8i1Gsb1hrTA9GdqeYf2ruQP8NrRv7Se8LTF7but2s0mvJ
XSGsizR65iHyCqYNQ9Spd4tL+AOYf/jdyQjNLeyxosYq/77FTl9uceEqA7wGjoW2UcRJ2N97D4wo
52uxYd7XvCZ+F0V5qCdsBb+hu9oKDhcOxS/jB+fHQMmvArCQJ3A91nV8qDexy9Z6aOZ7WPyYcNsO
3pQLJvGhDYoYxnESg3nJVFqgEnGDOK19AB1MJc95KZxTuhMbb9fymz6q5zj3fJy3YyawGniB9WY9
s9rdqq5Kb8wYDj3rgcMaSGXXEvTTPJ/A6TGxgfF+Gkm6BaQPhXQC2ULEA6IWGczHGspQ+4K6LZha
bsMk7kXxpgUefT2dA0fNp1O+l5Y3O0AYGQi6RIyFwPVaAOjVCcwgCtuvUIVzfGdLgFh0TjthdEco
nItfjF+2cjA74/UCsqxXfcIHW4qka8UzIjXjnOBqhUuhgPZaK8E2C3sLCK418o8KXqtjJNvHqxrY
u3L+Nyi5jF3z4D6Q/QdySt7imkYE98g+u2oVaqel2TII67oNC8tmQVeqtU73eh5ALSGzEdXUNDbN
ehP4EHW5qu57WsWE5xr3kWgd1sd3gHn4UZy6tKpTouN3nUkQ2qeAwGcl0nhU3qnY7SMRVSlyU9iy
gsu7DGWEM57yijq7NPzU+4hd6283vdhAcYXE2EGj/s9tEKC6nWw/OHx1LIB/Mp6Pfo9v/JISKszi
QSid+t+WQuRicMuSZ1WEdGZPpQW0J8874GGBQ5V1oW1jaVbKxm89938oYcQ9I1B2FQGBQQ7bKnoX
1ReKhwXC05RrNb/0oy9Wmd5IpvTyCcgsrmf5kqUTIvCd5jK9tMKAspvmAD3QOSEeS2QdZ3Py2ErE
ijARy82jC8CtwZQ1UogjftvIVWZMwE5nz3Un5GZBmM32Ui/QyR8vk0wiVY0B9qhMrV+vo4O0YuOo
UKv3o9gnGftqiWqiiamEalTca3wxSD+7Z5LLQx6QaniW1NrA3fdpejK907uHIG242k+8fvy+Cha2
+mePYufWTI0J3x/7uYHhjovQWqX14vJ74w3Kyi8oLxmh5eMP2v26c2cVodfnTzs+DqEEMdvy03lk
bvL24VlbVYVyL2g1zjufSE2bBc/9Fy4F/ymzmqMrj0w5Rfkx/8jTLbQxJ3dXWiJHUtGNpGIdkm5o
6lnT2KaYuf2raM1pl0Jfgy8oMrya+ClAtLsRY5jxiCGryQ+AQi1oZExl5B504F3WFlULpT4Yuycp
DgU1Bam8SPgXTNL9IekFXwgAqtrBhDaQ3NkEKmH32CT8FgkU5sQBbQWcLayn/m0Cglc4EXLsQZZk
oqmB1Pg+uK95yUfIYsINdMDDuGT6lBMO8eQCeoEcANPEhCSWnh2qMzKbwNNwep5VALhtVCa99aWv
nagnyxJ6AmvB8nUFnuj9y0UKhVCLvpbe8FsiBHY9bjtELeP2qJLaihhhtWdnqj+D/K/O3gxWHX5j
GsxX0b2cqEKRrfkkrw3YRu5ylG3e9hB4JrFNEYEecw27WEscyImgrn6z2TclNu4DihRJGQIYvhIR
0FCQxHUy9YB/kYTkG99fhmtTDpKJvFf0RX7KgGPvBoJN6RSD0II5coq3cHnB9LzmDMA/RDC3XO+V
WKwG3vTEEW6eLOKh8z/z2creilH7qmOj4Z1C5WG7YbM4IQ5yMkp7dBKLxdZuUBoHkharhCpKv3bh
k0+KbUiHF8rYDKLQntQ8V/IdoghzEsTKvJQWxYSSz8gGoIhjGoBN9hW+YwaIBT9RdmmepW/n8t7y
KWj/MhAgpm17OoLkwYX29Wrx/xv1TQrxpZNFhdptbJnEGQhlfvPZyzDFCJxCw5lzjczrQVzHIJxV
Qdzj2RJ95/A42IQpEVfT/rJGH7vlWrd0gB9x08fHSkNuDQxXg425Tr/S+lSFEaZ4FhaX9MWBcDbE
W5hyfvF3f9pT3dsxNzdnHe+pQc1nMkPaF/LHSWgO0b2GVZHlEVx3CorE+7fNqB4s34y59OeVcCDX
aKuKg9efgRza/MypCqDNqGqHEwpRBf9FTJyrZLSGG7+NHLiuyAlvokD5hYraZiXwsjwRjBhFPWVb
JhqITygT4gKoVR/ZBGe0IFA3BqTnCFkqDCQZn54SMhLOtnr/egG/biRteB9A0TFkyUC6diYw3jN6
4jGfiw12QVOa2/6wRZTZe8T5Z9bfm/EsTchu1CSgt+FxKzPzv/6lDyPWlAK3Di62WqzBfImNUAG3
ulMnSOAITmBz+qPKtzWak9j2chq1n5R/UpNLqOD5pHFo3wD9UEXs5cjdPqNTuxSGOVvmRwbzmahb
Lb0qUxuF8kjMSB9cpUG/I0t0AcsPuTaWl+DJ7znp+Ryo10dPz25oAKXZZC/toPMKvgazy82gRBca
tlIIgLHuzPoasOyNejUGOaCAih8N/tV03H6uvKpTJckgTHBnoWzrONm2U9D1l2C+m+2zPI8MRWRX
Dl/Z5hmYeiF+cMmeZU7N3dYFhCF8vnDAwtibJM4xtB8c8J8Ms/bTnzQNh3rbVw/Mg0CiUcd1tvTn
mKQRWRDgRm5Z7qqEi73JmrKcHIXRCFaSU6GPJ2W+I/HaTIfIjCteZIfpEUegG2iS6OSTKaXbRrLL
vURZw+xVKrtMNq8mSehKxS/srP1vZ5OLFVrN6Bhsiu5GRBUYdzSUXwP+G+XTVz0DNAlDOffIpmwX
QQKmBbOLbSMBNuutQ76VFOfVT/n050uT0zcVmsNoNcKiTvlH9ykpeVzES2YBjEW2eukzXwMg8wst
qi9um59MKwfST5mIS4CA0OYB4YC5JMAs0RE/q/5vpRVmHBUvCTv0xMXNZ1vOBqSFLscTX5XxW/u1
0ybqktLcMiZ9e3ttE7h31JUnd9cXJh77tg+XpcK1/bte93wYTqv3KCETWjOF+VhLq1N48pQMEptq
27CcVxsqKXBz8VMHMIlR4LfTnGh2YwlSVQ3guxFZgb6Wjq8c9IlppqUCjnpv8t+cdZtpddBXONfN
mXcN9L2WUOzc2ODufXV/QVRkcWi1tc+knNh/yT4XmrHOwpdmxzS5Nxj1F3Wnuxe+0XO1TyvbcuyF
Ltouz05lHoudlpCtY8XE6HtYFOLsBSi2To0KPp6bRhy0pOv8HriTiXXWRCZzwpA418tyAiBrpdjB
cOv6wPpG3vFtPBs+SYWlU1Rl3LxalRPKO4anzEZXCZwwJtPd20WUYBeXxOOexcd1Q8f6paFtv3zf
WI3z619xLP1iJXjYk39x5x6I4qgsdy81k4sBpcjQeZYvrAHtL5u7G0Vy11SBwkqpfNScy+lrkcpo
+tpm+EAQq5AX3BokGjd+c3YHwVGhIEwWShKa9jq7bFKKfRiTorUcXw90k5dfBp826Kv0FJgZw19L
Yss2vQHil8R9lvLo5SGhT9Mafr2wL/S93hm9J1JLTQZWwaMqPP5mRSfDsjpymk0fg2mw5LZnlemS
xk34N4UVBerZstkrFBqr3oOlwADVpZU4qLDDb6GY5o0ocUzJoIv6dEYIaJ2kuYhN0H9E5ZDbnm/f
lnUKDcXX2kxwNJEJjIgR4MGULy+3Z/ZSk2HvMRp6xarjBohKHx5YO0ywJmyUdPi4izfTcWRCU3gx
/rbmJ2DqCQBc12vlhDq1bcpt12VCiippmgM58e9hBLXt6jEMff7neK2QkePJ6VXm9D7Tc7FLKbwM
MsJ+TEhLXgmjfLmEJnoyazt++Qqp7UBNN5BBMGl+M/TaWFi+7YHNli/WjSsqpn41+SLBBhwhUlZf
4Tk40wIU4b4t1aVZPMnhXvlQU0+U+q0jCFiIjN85Rfuw8U6Hkf7pHPegOWPaVquoQ1g8wAUM4FlZ
rMZkr9NDZI6M8xXeMFw2GRkpjto9XO1ru3giAYOTyPn26Lx7L/7OGdFzhuqt2bbJkvLodFx61zIP
8/jzc1UVK/JN/fvVvv+9ET/yCoCWluj2WnHBLd5Up05vTXVqGfjUFGa6lpIGd8OrctIyu1gfJM+r
u9Tf/AkOfhXA87yEzY3rmnWxD+PN19VfcKg/A/SX4oXw/2UnUcpFElV//FioRXLJG/FDmD5nLHEI
3ZUFbl5qa8OnDJ4oBfTM14eYZAIdAX/dfYb1InJIS4igNgL1tHHV959EguQ8CYhrUk1X/XqsJBH0
ahpNSNbjq3NHbahqnI3PZ0O7q7q/l9AylqFxZFaNvYFPk1k2IyrEaSRfuQLS2rLFR2xw9pPzUCMa
JWHz05F2V8LhVJA6ppNEQ1LUKZvpMBPCnu4cu3TK1LiRJNWD9oafVOl4RDB220Db195yxuAWklN+
GZktN6WmZO1iKHowF9QmwZI90XCug6+u5xpnuRiI9tQ8tN+xLkrxo7agxP/+CA/qx6tI57FGkLos
zkLaEZGI0rS2Ho2mECzj+EETXRLyia2zAzBdesa7fNebPG5ZCplYVuoGC9mUaogmP7Hxjorv7QdN
sVnH98rcH5E0A04dMt8J7SE0eLZpTTg+2zoGQ9eneDOMlfkd+WQbZoD2BesQjuQ+kjoopt4dtZ/p
/kkE6eDuL2hNXmAeqSieH0Jzk6211OUGZmmz1MQ57TiJ2WeWzDkxGNK9km3ZsKXoPkUSPDB4ow1W
05qOlyNSSIPg+I7sUZ4vJ+j4gVQhJJRQwg9Aamn94ySI5ok8jXxxjc1zuPc+9h96l8zsV6quQd1f
M0wz1/b0k+OJszuZly4dbEk7cu/6dKf+ePaU/OBu+kkbbhiTgn72NHOL3Zke8xjNjuSOig44Fu1T
wl+/VewBO5L7lhrjueNPshG3NArIHlTR9aO9ptE9TmokTQhiXSBnjfKiX0Cqj0EeiW4Elh/T2sq6
xXWat65cGhGUk5r7IbYjmfg8IL7Oj9SZlcGPflsUBX8+M6k25neSiwVGhxtEbB1sFXUnpih5mzmX
7N7Z40PQig9ToPt5PRWKAv8rPGnjGUhQ4g6ZTVl587FjEBqL5FD5vk2JuJga4TSLrUZrEfUYt4zh
nbO655I/LD3Me5is1zDAxo9Q5hk3B1BwUrbp6ZR7DGQpNBmiIYd4Ax1BODmrrOv1iCWc1N11pYZa
Ej0NLWaskTTMG8GZnpmlvTpDj7wsbAF82mON3x1Stv1KHCqEwJNzA1yoR4Y8GLHO62lSWM7qOicI
Aah5t6tf9Zr5nvDjrP4wCvbjdl0S0ixbLIwNPrNmYFoBust5EcgxhMNFaVDbC/HH3uZ9PBu5eAnz
QkZgz1rbj3SpgESvfTZtIm8OoGliEhs1HSD57hsEvmIJB6+hI0TBobk2yUNzhzqSv4BAV3VP+2Id
XpiOMvbuue0nh6yJvyiLUiDWevG1DOqtavVZlTMgm6a8Zj+wzsX2VhlRKzZ0Qup5SbTZylmgQ9UC
WeOy7IqZSxL4CfEI63yTX2eX6F2euhIkQI/h07wF9CWh8+upUp47ZFYbRoH93Sssic47yFlJNkSl
kxOkDBIAinnzp+vsKppAf7O+fPGrA906+9WqK/+9ZZJlD/Bfaa5sdZvj2PlER5W1kjeu8HK+geCz
q6eKwiPZ5bBGYm5307wg/PJUfmpg49F4Cbxx6k+0q9Yrvrq8Ib7Gw2ed00AMr9R0Yw++0qc8Tdp5
2ElFNL1aGgI7wq/s1MDMnNibSCy5NEEn93ipIuRGRJXHR2EobRnaVZdxEAI9oKcVkuH09pDHlveX
hCJASz4Jvt4CJgwZuPk3yng9jb5Bv1ssMrW6yocrEabJ49KI6fVRYYo/gOc3QIXB3DoFOBQJvwfp
opf6gc5WmluVj3rLPjN2tll9QrT2XGLz3ikwn82I7DSszhgXAJEWkhd1hTx2XEkYt37RMXSdQLzF
wVJArj+VgaJtX24rNkTccN5QVcyAaUyH9n8Pmw27jsce+iaa7J8vCjKnC3DLWt31pU5PnHj91V1t
7c2R9kNi2c049yWRTOaE7UrWKG/DPM+R1KRZteAglePkQjnyUWYtBEMKCfoJXNWmwD1PtElYe76x
HX1+G3tpmnZkHSr+JMUGn7jXQW2+3M80AscM1yuNhEllyfUV6cjk1eOIzDNuUEFRmVMuK9vyBEOi
YQP3Sx6qVW/n4GEKrxzBfQgh2eDAPO710B5KQCaNB9qL61ZfpnxrtNRpeRcmkylbhiJpwBfKqnjz
WP9E9zgVox4Xy5Q7HTT1MgcjThEycKZ0lZ+kxdGsP+s5rwgg5OmmBvjWLyq3/7kdpzw0jmDRF6Sw
GtdmnPRymiy0uvd7WIl0MpLZUb0POInspktRVUG/ICJcSxqlZ3+biOVXxy8ph9twg3b3gGBG1BVq
9lWzySALmnXRoXsLm4+S3KeZD3egYLhab2UFeE6HW2fzDOw8fCOQoOuV4FyTGOiWgjEEib0/xF+j
4Z3eUBuFXRRx4pfhqoMtson8eJkn5FIyYZ0bvkWB9Qa1Uuykrfj4F6m63FiclM2SebH75gFzR3jJ
rt9IDkGMeh7RjLk1JR9+XRBpbOm6OUhXSj29bnjct9Qumi9OrtVa1+fdgwpkokcKjQBLof09YF6Y
8e0GNQnfCXQHPam/lTMCaqZgqYGPBVfCkbOtcS/94bDhDjDjySWXBhmpJ4r4LmNCDSL3qlSmdOvH
6QHzNFYpf4R/rvLCw2qIWCBuj1ke5CAVPTcc5dXrMYkF2u5D9uZpWrrkKtLVSHcTtEJqGT+DdT3a
uL2P5/Dm6RH8S2DkBTyKqoQe3vgtUI8CbPAMC/+4XV8jHhlN69kIyCsqvWiz5DsLgAEd7Er83+qt
k+fOJc6YTAIrpxn9BweyNT449qmV84qBPGQ9vF2uDCswXFVkLez5RZ7Rf2oEglyGkQ9DRuEUs5zK
R+vouFSfAPisYrAX2yZEF4m8VArEBBLnVXuiIx1u8Ln0//uEWeEZms9VV3Wh1HJDYAhTYym+bnba
RuJ8hehmIps7nBvtqRp8pss4ZmvI3sjgCCMaCjt+ygGwv0Z7ePWHDkrOnKUTT9A33Vk4z8dZ5j5E
rHzR00/gmp1NEjZt2xXdrAzdkQn1q7pKFLYd+u2f1LhVGU6EbPpiB3dcg3tFjCccOkGTm08lpkM7
A0bWKCNUBsqDiWmt5IJc6V1tuAybkpa+XgmlJBg2DawWBOq+vc4S3ADxHJ5RyA9mZPqlWBirFjjz
9CbZ7Hlm1NwU6Gz2g+JbS3ty2vVNMu1clHv2dzjByp2Is0QmkcbVEfNgDub5zwR4o4cpf74pzV+J
pvRIzfT0X4/LEQXLXENfFaoYre8klAy+6GLNg7RV5WiPMROFOSH8VxXZtPym2XZzF+6j3SD9LZA3
W3EUFswS3ojLI8mBdM8qY2qoRQSd8YTFqHgU8rQnR0O56wuJbI+wm0uWdAQv0GdnFzh6moR4gx6w
3WypC0wlRaOtMSBiEInm17392HYVmw155fmfUElE4kPsUfqjpPD7aPH2+t5UfrDAVM1IMXvqovhc
FFfvTASm7Sj+kpihc3PJva615QOVVQIV7cINa28UYmZb7S71FVyilQv9z4U/qxzItm7Exu6qQyRm
cFendDUSCfm5LR2MwHwdz295cTIJHnFaBLkIaDPuWhNsHS+JdIYX6GUc/CBMGOPalt2vIPQ0prQd
cbZJq4vy7y5tqy0EHvG1md2VmHyKiEhRXXb37SFSEWcaFK/onmPMDyY2hI8jv3I7wbFGAzd3575a
poO+9SDiWMPcRZSWitguoLTe4274uydU7P0Mu7nySU8qrQDbNwSNNYKEaZbfgDctxEqVtGWRPKHN
koMpXQM0ngFiXrnMqXMFj6FXsaQFzFKbvcO0abBeVPjleYXIgzCS5j278KI/mGFQ2EB+arfRyS+z
JUK0QfO/HTZSptdIVfj3gzsUTiVTSu+lrHEewjFry6mQ3DUv1nhqU5IShxfWTREsvS7EDPgnXyGQ
ZXIwFEP4wORqczxhV1RrvawfzPMkHlG3jHttxBD/Pe/6sx0HbS7dRZH1Qefxl0wcZuYvfSgr8H8D
dc08WpqmVBx59bOC8UUafiq59N7Mowk22UWhfzeQ2Hf5FPCqYh+N30I6PoVqCBXXlqOMZD3B/nZg
r+urYz4n1L9hAcyGAB9PrNS1jjoKrlggsAKBg2pliSaHXKWmCwyLUZ6Nn1K3/GBuAcsWCRTdgEuZ
IEkVd7KX1vYQzUPszTSWLX70sLSyXWXvC2WtNwEzQS3ukkpQzWfW/s3bJQ94kio2Prj2jeDdMpv9
w88QNVpvJPoqrDWmlcmC7bL5Ebh0OcCooGPpw3+kJ9mWExjQpLEeiIVNGl3fBgGVDikRJHAv7y3L
YFxWbXw4cumUxYIdv+X/6ddNNDgl/AJsuORmn8D63xSR7eftJdIYjApJYZrzqQM02LapmkzyS5jH
wbbwJaGN391cniESm0I0yhYgEf5z4yte9Vv12EfxqCwJ/2l5bj3OdtWtLT6wODYi5LemTZihVUGl
RzBphBQCjcCoDgbUfL7F2Xcu86ngz0d4Cw4fvwI2oxn88rSKMQrtseBXROA9lqs6d8BfzoDQpgFM
v44SeAJBPrfxs4VguQma1q0iaUdYa6rgcseLBllCiZ+I72bCTLEgFM/77cDyk/leEY2wJdoCM46b
sT680QdATQgpMGCrTfcYDi7xV3d1KQLhos49ThXo7AgFtpBTpjBW9GCOpVv76bIeyS2Nt5CgSaEq
JseML5xrabbiJzW/ICSdlAWTe9FOQAm048KzHY0GSdG+5pFVeWp4qdHHyeZFTtDm857HTzkzS6VU
rBLr4W6BhU1kA50kHKDDiWkY+OL+AXzQPpAD3Y7ZHn/IUlwxJMTEzGDhUlq+rcswB3oUks2A7YTY
Etx9eTqRL5CYJu6Qw0y28v50PZXtkKC7GXpskK6m4N/+P/hGHkS/8FiEZcTJJbozxGn1GDNHDyZn
bTzI7FUFAAKeXSpOjJ67ehGqJP/m9mIdVx9YAuMXkIJ382iKOD/0PNnEu5nXaBfBuxMpaw7tmMUn
+RmIOguNMVvHWshwIKSrErSO3B/l3OM8w4d/JdDfq/8woo9kWOcRdmoJXSUN3mBOZG+uafp8WMlz
Z5x2EfnIf/ojGfbmIcMsKKEVV92iejiLS7Mfq2wCBukywxj4T40+DH4wPUomakc4+V1vNjvVvRMg
lDFn7mDlpHHFosgZlhEFZUu3vP6ImdJIim1QGp39lnqmYkxyNsNrr2sSj9igyFshXXk4HMx/SzGZ
IoReT1ynXq37AEt+DNrpptZepIbzsK4o0eTnqFUbebsZMqFq8twWajlepHeDk5vBrSGnumPn9Kje
BtW/jb3+LTaD2AgoacGfx7tT/XWiGFVDoNdAxxXhk4hB9IldVFjgUUrca/9BHuRNDEH5xIgYNk/+
vNFgCPjc1L+5hd2xuLQ9DFQ998lNqVV0BufQ0t18xNkkoYRHvjKtGBufq5mUM9fwD8JbwJjz/4gF
pk+GqN/1dT0fEoOie/jfS7+T/gBE3vBrU18h88zN5yA1AnzqAcLA/4B6ZPVbVEOfb6EzZZcHJmxz
y/vi9WCKPsOEKrDPrM7Pqh7CMU+Qnlz8C6sG4HQwC9mHi2+JGIOjGKSUPfKwVft6cfUoa/k2AQsF
rZBdbVSxvi8N4O1YqG8M2yh1+SNRvcSnrDwpS2gB/50cJoHPzI5Pl/VOmt4RLREj9EEsBlR888NG
bKb+7DWEwCcWjbb7PVPuaHZTyJzOIOK82jDcAqRobhYZzHduHslBFT50c4ElzrlbkgvX9qUvqDLU
bWWbKIIFfmH0Ety6hgm5H1hEupLBFpCwewW+Dn/wQ+LGsYBnDJAFYH3D7EDRuCfJPNueUOcKM2bW
CZDlHaDK8nF6fQwKg2diyz1MarNU/K+VeW9SLXNVyizuf+LR30UIDQyh7Bxw98tsRYqBO5sm3s1H
uRtmJKXhYu8IE8OpZ5Z3VuMREqpGEnTWpJ3HdybFFmMG834io6vaM9PGTw5rLaCyY5jS2d/TVQp4
L539CA7YAgJsjs1qxPYklbLPud2rO6OjRd0q552re4Gdkkwc3hu6d5puTXnY/fiZ1Ha/JK/LJNcU
YNX3MjgGxJgBaI4Uraa8Jgp1wpALKhVxdFPfPwGkfhFl8W3GfhON3VoGJsA7KJKiF9podPBv0tu2
XSBWuqxBEzOvqTtjLuPrnnT1Ek9lRB/Pdl0WJOvHDuInNKjR7aG9i7pYKQiV6xXVFJPhLNl9Mrij
vIRnrfSz5Lpn6/PU7GE2QwBSjng75jtBbvs1xz0N4yxYCvEVRiyDuc8QonqgnSWNtZJD7bh/QBjj
CX37bm6EMVh/i0Co3dJ7rcurE3K8RzhVKYEq0rcx2AhrhkHuotHQd+Mv/kh/ZRUt7weqTDh9gSUP
fJqsPPghRx300FX/IY8/dqieUkEoeIm+0DbtbADNH2U76JQPNYz9XMps4kMDrZpcTWCpL1E/lYlq
I7L4gUDeHkLh83c9ucguvPIA1fI/PHxFH4lbYMxw0Vkf+e3a6fQkYIP3/pfT8zTtwcPdJDkgnHm7
tTAIIribrgIsjUl3T/DQzzd8arrAk+iz/4R+dhZiPToNL5+WvrnqWLf1za0GUWUt66uaTkUVxoRL
Yv6U/dXsVWyj/7AIxRpzssXhgrkWkrk15Dr514RlkhAJ3JuIqJVzeEDuqmfMNHSNzvfNEKLANlxi
mKXBvPlh/YZHd/HfUbtOP1ulYi06NJCBfN7cCD0tT4WXuwBoYL1JT52q0scWgckYNnvDzuyajjP1
EkJmdlBj6IieIUE6y1H0Zj5L1Rf9UCdPbX7ikKRfbCDXTXRONbNYfIV4W/m3LZ/cbJ0zlVN9qZOH
KlDR+WqCCtE+DKMADHWebbQ8juOflxutrgMLaDDsDSH3lREELvlglJFQ/4pWOZZhznYPvqwBivyO
Mph6uz1ZlulOJc3z5PeHmywiadecVx+IJCw5ArQwkMYadf8OuQt7EoYsOUQequ1CORWo0TgSaDw2
uwiVq/4mEyMLgQkHtyJRGcNgwU9Uh1Isot1D5UUYdR2C/Ionw3h6r6Gvfvwi0bPq+WsdSgJKnepZ
4vuKTQHCRDkecT9vgu6lnVIENTcumNmrGh+BYOKEWIZkmdBIiri3Q5dpH2s6aFo+nTHX/W9QdIJk
NldrMvMF7bPp/8HtkpF1vteBK56TVmYrxV3ALun/zvY8nFJjfQZgJmjCZdCRfoV6FIJyIC8tc+x5
zZRgnYQnawhn/XvG1a0p3kbBvqjxqOz+yuKWqRwHzw/YSScM7WyxQ+gq11BZukUtbnlDZNVVB7BY
gVeCxLSg/sgO/C+4p86ysfOvSaqkGWpKqJ+HPgOkEtEm/g6QmsoYEdt23xs14fgmh5y1dRdIi7/g
9ZwOKPKW7iVTFWhX2clGB3vL4BSQv9rUAeMmGrR20USrJwPpoDUXw/m/Y5JC15pecrjPtsEu6hv7
e/AA2EasI9uQBmuE/ruepiaUN3C4fBPt5mZTbCo0qWrQh3ZM7fEsZEVc7xt0MPvo+t0CRzB4lGlP
aHessE+TULbDYcdCMui6iOGQOxEwWQ8y5lZVBCpQb+VxGAAJYjPVCjR0YF0sUUuVKJkJ56g1/DrQ
QNu5rLWFMohqMyg+0IKZh7jwBlt3cZv3ZB0H9Ep3/N3PIcEaq5yVobsh38GYO+v0WKOSZYkSNgBU
oA5dp02TjByC46iiJ5igUXUFE4yfhUcb+fd6Q8hVRnQCmXBryEDLSmYwaerbji67KC8dWxSC/rdF
QkBCbyEus3wuQa8SNe2K8jOZRFDxRq8VIUhT9SvBcb1F4v/USL3fTMSiWVerwJVFP7IX3Ismmrt6
eUZVBhTJig4qR8vy2M8TSBVG372hJ5RIfQ+Rx8qHj1EtOi5iJ9a+4Ely3UPZx4EwAQtQWKq2T76Z
aAn062FOIzXLsO9QXHvW93Q9R1drO9hdbvdLu4la3b3ilUncBB2Cr5r+kIPMeB6BUxNtXB3E42vl
zSc9kf33dsAipSLG3434XSt8cBT1A0+QzApvWY7WPPP8ElpzMsD2v4BBFWTYeSViJUsH+owDSZUt
nzxv8BvQe7JlNFinDATGFWx2nbnZZiCp4QF9jWCGj9T2uOfWGfj9aOSxHZoDm8yL9pJsvqisj2mq
E9ef5ILO16PzSBgHBx/sJ90oMK2bFGaKBPQvetAJcmOBIGwlnUN9SJlKbtKIutH7qt/q6QlhQd4K
7wyuof18tXrzMcVuYx/mdDMzgfji7CVvt+s7EI6Z3k69jr9domTGDVJkycqmWsvTPcpcX/Cjyu8P
ejSyWhFl3WwlJwbHqeao2ZI9vNJSHTl4M6PxNqvaBevrWBr4DIRtXWHVzfDjZYwo7lz/S2wf/+Od
GOxMhMmQTTP5Ye3PGUc+Uu6PTdQEUXXLKucX90LhGUP04W4I6rL+4cWoJHKVV/gYFJXQ82ScA+Ga
/ptEP5V+RsEMQXaAjn4j6iL9/JfnZMYgzn2da4wq/4e7IQEWGrK80bK9u5u9bpNE1n4s2ibJc3ze
8Py+R5LswF4+9L8duCSrU5A0cuOeQQOxoSynCS80a1mvaONXj4o9ul+yVlQsdj8AcL/DKXqWCuEy
qfK5p4qenZC42hyP1PyDKgAUYYRRRvlaYMGvYTl6Q+Fx3K9G9pMes9NTy72LHmNHGeEglpmx6cfP
4Uit5DM6CuJi7t02rg8TqYbmdvRmsy3qtRRV3+5L5KPh43mkjF/+aYqTQ7QwfBSA75VG2IVosBFC
0f+DZ07P1f5L6atw7RDthFuFa0U0K9dceRQA+TPrdHPmVl/T8Of2zR+QcrYzw8LxX+aiRMFauVz5
HJvfX0/OZRytLO1yBowF9ig5DJFIap1nTT4CiTuSIuxkLZr5DRmnfCwcyxqwXYKeqTypCTUwOTc1
YaEdAr5zMLXBhe8KLbT9vCbykZS2xJXoDdGV2qYbhs3O7Cg4xho4IBDlVu3NIvt4Dnf0ZhhnLxt2
tyUvgNKccmZwt146Mms4m6MRLk1+DS9Cm8Gnyusc2jg3LkjHkQeeWx9O0ZjpbxoIejM9BudiWeNK
2UG1KbLuvxzrvbIJIfObFChOA55UVK14oCKg8uYNlPIajHLJdr7rzxO+z0StbZiMhHOVRDkH6K2J
75Eqyc4Y5MGFCn6uXp4vuBy1x45HjMSReFG6WfJEFBBWaCrHUp1xEpnYxytLCQ9jxHL0u5z7ywOZ
UmaZnvmyzo4c16HEMb9LTh7mlB2+fVYqZoc6IHZ39oacGRZIORz5jvRLoTzdcOYexMl9nIC0XEoz
WbXEmqwUr/6eg6ECSUT6YER6eTZTFxzLeMqZODTb6yS/nw03jAGTIobzY0QoNlBffPHw7IouANZh
2iFnP2MjWSWdUnasOS25tRx9puuHMqLQ99ELcjm6GCfGpl9ieNBOdC+VgbbIZtHPiIDKbF/nEEqF
BoR2PZG+h/ZOgywL6R1moHldvoaFzutfWGt0ALA4RV8l97PkAmxlolilCJnIrNC7Rg9SeGNb4Uws
R1qi7dIdg64csY9RCpt+jtyayiyjGLqx6rTGblDfPX071HsBVycdbdtV5O7zFi+5YvdsbVfJt+/o
luD0qeFqbvkcXhIa0q90HD8n0lAuXVNTnNRbWRg9HHzMzsw6eXAUhLzt0mVceNGRgrB3NMC3giYy
tUG97wWbpPBZJqwfmgwe8p4812t2BlfpTJjNNCCbxl9KIQhZ/h4zm0NsMxprgi9tKT5+z/iHoxl4
Rcq8B1z/YIwNHGbZsuCrlRFwSPBqbj0E5NmmPlLyC5EoHjgG1/19E1vwwTPgJ4rOpFsy46BWi/1V
gbHPcALBCy8yP0P99DXAlwTpwW/3AqcPhXhoKCQETILTmHDABk8prugIKySA7g65fWr4tUVZ8ZiM
BtKO9HOaCnKC+3LKbfAmRn5rkX4UNVocONJyB4DVUJMjHbmk0OObi4L2RcUkZxM5LWkPdZd2vyru
Y0/Malw9DhxzEAFKd3KFGJRjf64yAPmQ7mwaxxD0AopeFfv0/e9s+pildy1jlGbZ5QEocseQqam8
8VImpqbAHFieHmntX9NYZbhXZF4RrOMHCIu/LXTnn++YX/hJV2PK7uSamdBRBoa21HxZfiaE3NAv
bDCDBoeX07aLsQbfW6DXbkhTtj4DV6uvkVEzlqxBeU/HzoieBKAeYphtl5d/KBnCwquL94c0e8G7
UPzCD2+NuSHp95dtOYRPphFpopOAG3ul4s+0EQOCc0/MM0pS55XWplvK3yRLXvdtfHoVT96QWCix
+zQA0hEvvUFc5kB4/QjD4798J64hcpttiSVjFnPrweJGt8nVABrs7EbA+WzjWj2TznCJt4KuG4N0
yEL1ii1iOW4RLvWN4j3qDQmqU36lxOqo7wZg0UiM1nnV+vy/GGClVn4Iq0QD69o6Vw/HVBtPL6vs
JmbySfSvz4sVrmTR8k/suC7G1CGEJc2hJDg1sCsNYj3DvS4P0GFDBGC6ttPHX1JD5k8CTouw8UrP
smfqJdNJm1C8jByXcMFijkZLO4T2Jcy5xV3WFIrGQUU0XOTCDlb5TdinzJo73fcSPQfTVYslcEQU
PO6fN8MeUtRxHv4cm2zphG0emb2JTDNunzPTDityTehSpunqzeUuFCeioXzJOUnVP8vq49BnTkNH
bdS5phEqwwVdA13hfQe3r/mzcGTcVUxSLqz27uvElzHy9I0KpWf5lg9Hu5hM7ZD4WTANAhwX123B
Fxzvrq59IzrGjOdhZ55nIVijOOay5gkQYxzXgmFesCoT1N2utFaKrGtxtry5fse3TT9SkVohLeDt
yz5Wol+I9SXEAA/kQHzGy/B/HQMX8trgv5uyHIYOpELlLFKu2n0yqTScGBEB9SqPHQ5D44o5wDOs
RxGY/tFKuHaLCvXrjQV/SgG2psZhphl86XFG676UM67povOuhuWF4Kui03LVTmvk0v446IJasqoC
THSsJlyH4OiVMwrwUNZWimrh50Z3e+uMidzb+QVsnJAz+q/F/444EBxyV9jPbs8WXni0Oqx2B6Dc
E6Sq5Bp5KRizSV0m+LGc4oDHbX8xN9e3ql9B+HkFKUVX+aN+UHpf7NkH7NiYGzaHcLAR4QI45We7
0IGtkdWqymB19mJAI6zH+sEpJcKFWWaLbYnyH15q3fAPA1sAb8NrCUfzG3GgNGjMtWIZhHXN6pIl
AC6PAySpsGDLqBt4A8a6SsyY09hiF8rgKmbV5Ux8y/XSzzXZ3rqD5iwZF4Ogm+1XWiU5bmJhHyJ4
hWEoKraIBn6z35RRhmn38sUsBfqzdoBFYNmSgiRr+TS5UGsH23FBTbyFtoIOshS7vkksqF12d66/
0+VRxqhTNavO+xX29XrPHx2KZYB208PMhH5RqzQ43cMG3f383p851p+eh2uc02HT7ek1PuTB4g2h
UizSrF15m4w+GDbwXdPBsOzklfotGTw8a4qaXkPYlLdmbmgFmNE7e/+mgdrV/r8sK1jYuD9ESXaU
Ki/N942TsyPksW5f0xrqxJ4dJ5s7JPgKGCHbW3SRq2dHFGOJY27QdAYIs9hNb+5IUDbyb45w9hft
3Hl/jyGZE9Xwu8JU+1AFv7A24bmYO32i3eVKygr3B8dyUDzj44r9NQmC8NCtA+HY4Zn/qTGSWDaL
KvxN4pQ4rGJbnvX9FovACV+PvTVdLceaqPNffP5pVtJPuYVzdaq86eUQoeyYGou9s5m/8pUeq2Of
6ZXfUmvfXvBAwiJVRJDEtf4aV4X9D4yHjNBSIWrDxrb1h2OKPfpExVUtSNT5JGyV53X3JSg7Ald3
9iAXEcVv9zSUUxpQ2BcrLMWH4DegpkH5631MvZnySb2KYh/rVoOtIxpIHMgoGeN9PefakD1L8oX6
uLawc4zt+fe16stjpThXaw3yelhkZQQg2zm7VOnE7cAEpToKDFWOEX+sOfMgHJFpqbtF/awyZs0W
DRNC5GAY6EfMXxg9uKPAsRDRBz4x1J0KIIjnry9vrpmT2u93YvseYmUgunXMJnlx27JUMlW6ZUdp
eScv1NCAC4xnwPl43NdfuBQ9MvoGuc3dmOlwyJxf8zDvfU3XbrQeOUwtKrouNrCMin7mw7wLrVar
aYrvsgfBMUjQoPA8jb2zolgALN9v1OMMRVhdAKf2wbWgmeS1Wbxtkpwv0LUTXlN8U2gPMgwmFN32
/atE/EjTJBojRxwkFrGvzLECnhKwvdegsXiINVNYmXfWz18YxgKRU+QU+vMk3BrwdppNxsqhava5
b8gFBdgY4KE31zguoUZOUYvBjia9MuS/q+f3zDMYRfEsuYV3JOi9mLkznEpL3uPCYduLabRQZqSf
X4tv2mLGGMaBtYDGDi6EQuwjSL1MUwzQHUWUxeS57v+/hybQCuPP93hJ9Lw9Vy/GNDtcTx2aQMT4
s0TCsYa+K3gO2NFNvfiHyNpae2Ygfzu0LBNo9S+g9cJ1aqEArqQZaTI0FVG+9mPpYBOX+m05g21i
iG/6w4ca4qJjTbRjqyYhccv6wkMfHjAISF2UzSsSi0+2mYIa/ZeeWgTZmJWHOk6m+xTw4iEd9vS2
nSF8SWOPawLf7kwt6wJt3w3oXCcG97ShGiJVnWYH0X1Rhe3cg2+kZ4lUHIKUNbb8cQ8pT+N1xN09
DdhpI+L13ygvTABPFfoK6sR3k5YDGTtZO0paZbhJuMB8SyNBcoipjy1XEKZs26OZrcicfh7FJzMk
8isu2I4O6hy8ujcTNj4bqH+s9q0qGj44X/LeJ0cl74vjXEqGqwgikdoyK+XTQ2+EQUeQv9y2VPN9
GqZ2jiNq0WAN0pshbl5utnws9/DpCcaq/wdPyAAAlpWV8vmCTtQKqLBIXDb0SIdB5jzLpcnK3O7e
jQCpWkbmn9gzul9zv9JcSxSfYe8SgjMTXPVjpjMj0sI1/6ydLA3gpjCFz2tyZGjdqn2BiZl6xhnY
6NdzwFCt2eY6cXZtSI+YidKvUQuW3ahx/1iPjqKlNO4PWmBH7VFvGwyJNlfIzUUSpnFwR3dLTWqs
d1C2jdL/RBtt0PJCM9fcbg1iR8Z/2t3cu5CAXsjvkbObfKgyJ3i9IxUl671aoHuRav75sBYZoExf
iRaNN9mbYxod3dZ+tcBDzUsDPEhWmw2qhEuz9Fe+6iPFEY6UZpmfe62QHf373+e8z9Nxp5RQW070
gzVTe6r/TbABPxWvGCV4IVDtzxH2cjcGwfeW+U/sSNa1NvDKJuFYPsgVpRw6X5/lHJ9NqEiISCtM
7KPjvYD0ClpH5g/aHEe0pRHx4mCHEUia7WTBeQs1EjtP6IeaQZqacVns1GGYLLzHcEMh+PtTKVmV
yjK9pUEKjKanKOViUX4yv3nUeC+Ny20dqlEPwZ8TXDjeryYUFhIzn2AVX0xzYePnkypR6andnWrE
KdUalX7kzrpx97T050Jgz3O5taylkkJ8YZUanMGbEwWsZQ+iO09jvihX4lLweIqx0ME7y2mGdibL
Ann04b6PUoi3OwvbxlpJCoKr0JyjA1zF472U5ZhB15C6tZy4/8idFBkrxPWtMSJ30GVdXHcg77Cl
4iRPrEvAvkjL91lPj5ZBg/MO5ettE2h+3kH88VN1MHrQXOtXMnwCtKxSnDveUn1Bro5gp2geYvSl
qg5LFa6TG/XykJErdzCukKvTFdf5/9EBuPsUAWvuMJicTlpW2N73BjWhHw1TEfk1sC2mULiql+aI
SrY7UtubLf4ZEsNnaZ6HPrBOePcZVciYTrH8uptv6zDgqEEr5g9zt5++b45rzQf8rKKoRdWeH2k2
fJguM9myEpzU+aw7pwrcxkyXu/H8tlYoSOMc4a9g4Q77axtaeNbhMRUWd64gRToLY1tkOd2yiHaQ
dZsL7KuknwCv4/YMI/xqT7ZeyaFMc4TbQgfV9971GWBV981IODBhKnTFEIjz9ip14tUxdAm2kLtm
uRz9sM4imhgD6wHPlDYxdDzdPfKYc5DWq1VMsxCBd9ihJTO+SeVEVRVLZEzUd/nvovR8dK8DBNBu
BWiFmFshKgCxKN8F9DDN4C5IB3IvduTv9whTROMnve8vxvh1xeSr8Sjpy2xCr95TujaTs195S7lg
aqJd5v9Qqir5zjyuq5tPSt+0OCaJGfqo+213nzdEDkE+4ZM0WOLAWm1RnNgVUVcG8cmjoMRe9b4E
wli0xX4TMhPg+G8oDjp/54lWrLNS/1NRJeV5sT/uMW5K8fqNWaHeJ/75MXsCCiCtdvhvkPzy8rs/
/Px0udNuCg+5W0H0v9RZPy2FiG4MZuPfhvaZFmYJEVpTOCZ83g1zg2wBRMPlXDSv732bbMtOvrWf
ds5Kykg+QPbHPT1SzBouC2ETcbDUV4BV/dQ3K/Xj4z46uoH3Lysw0oJVBkDSQDBSqGF/fyxBK4CW
Cf/OdVjSYNm400Ydz96sC2tgoslgTPejTWHGIj/AK1IybJCVqK6eCYf4TdIUSt2vu2ZYPXkeNQWT
fNB05ZMN0yrsUgZAY0Bu1l7Kl2BXD4B2Li7tbB0LDJN9b6JpEiZv9xFruaClDUQE/qHwRSjVYeG8
uLueH0uJMYxVk5+K+sGXdKiLZnIXwowcQcQcGcZedX4p+U+727FU7/fhpwBlRZG8iFLOrp/tzG94
x30R4snJc7tCEUZ3w4D6R3e/NlpiYz7Ek6gfDYjyFJIy9VmziZYUH9qo8XPeYqjHUi+SdCePANeJ
By1HTnhbM3b8MkC09WpErDSqQeLnb/p6TTAJhUABXaSUSJ0H6hoFQoC7olJOI3XOD3v4Tj8Br2d0
EeUKequveBKlV+zxY0fnf+ivyN0aBoU8a4BvILrXGRnqmaFYH+Rt03bfp/DpjYi2vRP+2CVSRpn6
DUpl2PLsuNLxIpQlAcASw5aFlRcSL3eh0sj9mMJX3RvZ+YcLS2rS2RaRaSdcddKu42KUMfcKZHl0
Tvefr5sNStLKCpqKtCAyHaKe/zJsEpXkN8dnXRROwtTsvSOjYqQNWw78QW4vm6XB8aZmuYl10W9P
rmw8STopu05piksvijJdHdBXPg8w3a6aDPWLQKtwOFLA/GS6IXiKld/Xt5JYtvvqKMMMwl1zC+T6
RHlu6pkYF+HHYWbxQGRrsaRq10Mj4JNX4Z9CeqX0N8mdOQvE54OQuJlpldUXCSMHtWohu5I5/C8K
FdcyroDyaM5rLknEro6B140aIJa0BjEDbRX/N3n7TpZptMi+e+WrwWKcQf7NHumXeT6UXhBx1cca
EoGUFPzCDB3vwCfU5RJvQIMwTgCcKwVDpWKfLPwiwQIKErd2sLsNq9h3TF1h/TgxlEkOd/8Th6GF
wGxH7LvJshBQB+pXpahbt1Whz519pbD8TaIl4Djddm4Gc4xGbMkOEvyg6SIIUFZG19dSXEImlhKB
++REVphr3gk1CJyjG4RskLGak35nktXuPkAUIJb8UBbw+IcSjwq/gEu8+Vnwlxciw5L7ZWO7S85Z
qemfjhv37b7Fvb5kd0kq+0Im2+FQh5U+Go/1AZnhYGcj1MN48iSiIMamp35XGfiN6G8ZMkj394Mo
HLqDMklOb8SnRRBP0lIRXnQ6QsaO80XwiH2xvbe3fj6uliIs+zt6LYvFhtOSU1ua5zcz6oMnVJav
mczet1o6U/tkoADY370nl+ewaRAwugYLIF034YIf6yXUf0MtalhCE+dd/teaHYgbjaEq3VW2EhTM
PrqCWVsVGUmBwgVcq3aTtuoxYv8wK2P9EZx3OVj0/uI3974dA6ZvHE9M5Sp+dlOBDplP7KOXFV1K
ZlSxaOa2456oKXLg6/cXSsryse1sc8T53jTMWZT4CulkpPae+d1fcPUl0Gh3RC5mHPjXpYcWfr4q
iBQkUUHZ7f8LEMARiX4sePawhAE8CGKjHnHLvZmTfnZJNKLm/3azSwBNUhh3f3F7SLqor9n0YCmj
Ak4MoUUlDgtlHYxlq3tAFHVRRZpTZHELKt4Ihhcxkn/5SC1eQzjC9kW+PDwapqVEGltYFAtS6ih+
Dv0BZLckYJUVWFnBlDE3BTR5GyB/9byxQTnBNPqiUhSxjWTpJiySvV4Cw27QofiCmIxEAimAyM7d
6RBhX3PGeDJo7EMlkoggAo2QFb6h2tmohPEzPpMfeIWya2lH1Uls1JrzKibGMJsDDZKMw7vGJbje
jhAWNg0Je7SjfuBS4tdgCPZy2tt/9AZsVfVwFQm2F35v55+L7dHCni+r6jHLZN4DMEIEA7u5MgZg
HiIFhMwGc/QBZLKMdzBPesTiP0Mq5k6kbPeDeSV8eJMj76Fo1mOmt+SGE2ZShyO27J+pPw4r5gcr
GI2DTAJebS05ss1H9Swk2FdapQ4fD+OHcdDjUTgDcSQX/961s4ZserFhlAglFYhWWgbapjMUITl6
RmAldBenHFYcMH0hFGzy5H2qx1l+d4PW863DLqP5uKp4JMnObjoYJAoARR4EJLVS3vMR84Q33r3Q
eNOZUd6xuDqd4Epb84UZoIXX9V6ZgB0EM9r+w55FQYy8UBQN/Ob+DN9WTUk/R3isYvR52PW3jGFr
cgtDstflJwp5PZoZ8nYSo7oOJ1W0LpiEqRZe04EoBsBlEnZ2ETvIvwsJkGj6F849mupOgT7ORycF
OH3P/KQ6De/nR7S1+pCLUXumU2j+ByG0DVaoagnUUUFPEFGqUXsI6hRJ5y4Nf1Dgvd38JuqgW4V1
XrFGslo318VpMnLLVj6MWUIAHq57KPNxmvabNb8Ht6mOdThp9eu/760JtCtbfUxjwPBEXjBVUxhA
5G8ZosxLkkuzHKrZQTt3d+iOmdWAblFTRltQFetr/verQfjYfXSp6hkSsCPNVvMhIXPfBPLmvWsV
a1k4jbgd/fsUd2Hb/Nfe3VKIQeQ2I0+GsQ9qkDZLy0AbqxON4L8tDb3M8GriqMsHrUve45y1DgQl
qQExARBMGOnt3/ZsmHSpTyo8+FLQNA9ugR8oFRikt7EfDwA3mUKfq7wktbIoENqb2L8BxGx82Qna
/QVjGvfE2DjdBhgFmcAYzso1Ls9aHU+nubG15BV+XxqpuK9fAlLFoktErWl43ZZs2CuBbZVPknyr
5ivVcFnOWO5b3ygm46l/xjlPS83+rh6LESqMmhw5BuB76D+GP/1NUTPNHkoQyZT5c6HdPlSDp50z
x+lXVOLGKbM95uRPJCVWzI38e+y7lBiTplDHxdR36vqBNaQQnanYwPkHKlr3cbd9b8WUguudjOrB
K1TtJzTdUDIN5LThcWa0J31lG7j2ZYvkprEtI5fNQGAqkaWnzOtrG9DjAQz5kEk9Jlr2z9D6FV59
XAmu65x4AjTVDB2RLFXq44JnbNk8EHi7NB/Cf2By2yLXZmYW3BzgVgxl6l4UOfUajVbdJkdLYHqj
4VHLMhu4rTEiFNG6Jl2FRd14olYcpuLC8S/bT+OOJuWNERpcjQ08/Tq7JDBk9QbdBecMyBaWoLM0
NCURPIuoRRR08+6nkiUnovM1H/NX1dNxwJEszVxKUDnpK8rojkfXSZtMPieBOOyV2PtPvo9PM8/C
f4XC5FXLV0juGls5yOE+5AhOHj2pCe/F3mCT+W0lNY90FmSjwrNLO190FIfwUJDr80eapQpKRwBc
ViGo/ER223o5HiNwGN/9LIWq+8WuVFYT/nCKk7DQus8V57HnmEQO4qMFNx1I3e6h35NIPJefwBQI
3/LkhE0+lsGYyNFXiJYRDVxszIFi8RqITkIrzy96EmtG/PIGGAHmCrsb1GM6uKjpC4omWq6q804H
VJnFkI91SIWdLzbk78f5/Uooz5hhBDdEyVlWq511cje2aRCiYff5MU2Do3QOvcu7GCH5O5OMTXmI
IPGk2qahbb1jDy/tIwS9aUoVQjQQNJ7RnjVIsNEgCLGSPQIZ5dhPZUUb1/WmyzsLv/aajn3HZqdj
HLn6HUIAZbH8YZil9aM8mOSFT+wrB2N0Kbb3I6lANKzNFsui5IAJ1PnTO4iuXmMYgH1s5BCBJJLl
PYrVc1Mt2irzRvdWQeLFe/mSH8E57bw7+dp9Z96oAJ7zR6IEMb7U3gIrnvstEBkZrOg1XjeRqeUg
AlmkzM97Ei8mHdLJwXV8/+pRit8rEuou6bT+ONZLeJWN2+zG3zjpEBbfoyk7HUYMi/2Zbw+P88Ni
6TnMPGo+0keNBz5pBc6Wcy/P2ctG2Sya3PqIneyvgwqs0z8EjSJRO8wX461Z0Pu0Xw0Jbn1Gj23c
EOUluw8Lt8VpWbbt265h2nlCDmCfr5lruYJTOsKLptyGx+mq1hTL65jNWhPACH0fuPPirRhtcW/D
oJtKzUzI3wXKf2SW4/VhJlEvCK4xU5Ie6oYoO1BQFv+6KSNEN5s1nxTfpFd2f6CBXic7t7Erk5ik
mZTyzdpZhzyUqfZeuP4WgLRa9bJpd6UqrwdHsDxuN+/JW8bvZV+3gEToGI5k86z/GzLa4D5fmvZR
wYOVIBCmxxNEcLhs+X9PXt4aSGQDQyVSuKy9JWaTq80YK96Yv7n+TNB44cllu5TUrrx6d60XKaHv
UWlGcNUY01UdKUbzQZYfz/TTfmFUBEe2k4ip3lo5Tc83Zr/VFXoCt9fTpP55TAFupC+CCaKWxMHZ
Qf+3LTnGcsR33FvGy0akH/sP7V4nj2O/1tpwxRlbZ+oWWAvIhAAyC9wutWudWk2/7KK7KbkR09Ac
/GS3kABDvcG8Ihyv7eR0zbxTah2fJS8ZoId8OQ2K7F0l4HchctVL1mRH7nSCX6ncky3Xg6+VR2Jb
V/syOTqQUKY+rZwtYEk1FVxEM5gS7/2fbCSZ/5kIU8B1Nv0Zv25Y9Ll4qiYPw/pCZvhEbiJc/86O
wIQiW9dwa7OJjzmdy8xJb5RFtR2Qbw4gqTH8o3OzrVKyGL6CoBF4dpjXs4R0llT9mHG6XV9FOuDR
6VvGnDAZKwk147XhC59D3EzwHj3A9kHH/KkNzGK49Gf3ehgjPDq3jo4p3JeQY5QLcvs2Pkk5NM9K
a7/S24WSv9s374wUT5WFXx/oBYxqeGMtVtNFJUbd3Ft0cHv+7MHJsTtQB2JJkLHX6QffnaSuEL6O
uqBB6HxJ6QDp4jDDwZwB3Q268C90rmUacgFIZi5aq4Q30Eyd3vAolk0FnsDZsz29XM3pl0Ra0EPW
/cob0WYMBrMGtHHKxkAEf0iebmu77sUt8A1CN/At0ahKOzIMyapq2SBwYoKpwhNuhT7naD+yxzMe
lPZZItBcdlUIxHxRLz03UL6mI1X1aesqj3T0HQvnubzZQRzM9qmSE9vRZk4AO3UMGHEfoxrtl1GV
ObRy6XV5EiF2lfB6m2SFGMRIoVQx4AwHsVUWSkBC2Ubs7my8Pl6x+txZNSso9iyf7PR18u6RzIm1
+RIPrxAJHtsd4g9stpycARXxJH5MkXaOFXIekbtYspf7s3SrZRj4cn8iHXnB8KxGhrCUTrSfK5xb
M/O0vGg4/7pfyiJX1o2B7fkoNgTsyxVIVRBwuJbtUkxMKbvT1YgJfW6bE5XLv219V6GYF3lb67Ba
MME/AeNGe6uMW3soYo0PPDllovBHMAF0vERnL62s/0SjITJUjoBj0hA87S3JhpGR9Mzb5zQ7h5tT
Bxg7OTTDD+jCcLfl1maVF4tn5fVwnujWdyrg/jy1Bb6gJE8l1SCN0jZ9pr3afHGEDQ0LgwGfIXgR
55v4gugcYfs8An4pZ8sMjwvWAQ9wdg+pwv2djKKOu8KC9WNPKx9nFtUPk6xsgUAD3pQMboCun7wW
cLbfNnGukhQhZGDQCpyPBHUtc3kns5i9hgToFzADrF9YjApwmfRgtf2510BgupvkLwI5l8fD7Bfe
VMZiE8dZstIkDen/wFpFij9EtctJw+n6wYxiBE5jcWigaOmnx/c2NlUlkCS82yUUF8tSI8w1I/v2
T6qMngasRMogegde33X9bVNMf3yfQZ/w4bt0UAahLXbvA1MtgzkDCDTDQNC6/jPsZ6piFG11Shdq
JMfMGbVzIuzErlLc4BY1S8hVMaGNrIbrVxtEKYb0d115Hu36lJEJM9Q6czCNLP7g7dIgI5N8kUA6
YDzAWvCkgEmP+x5MH7AORqrwIGqLxR6VKLbet6Tm5pfO7hNz98DSZj61s2i5GtoTnzsycuMgeeqd
VbvG7t/sR12jxliqv1icWSKooi8v1u/3BqsJwy1my+q+xiKyZSs5tnJgj41FOgf24gjM0JrhvnrQ
kEgwpoamJGxgmC21G9ba9/ceSMGwXfwb+DzwfnUcU9cPfm7yVN+c/fuTmFlCl4PwpViP/VwKml2a
/Mgq9TUixXVyGkYDPFYAVjDv+JVV3mpij685w6e2alJD4+Le8yOsNqoae28evw6mb5c+yUiBxRjs
UoaQVMo2OF+nCIq1BbV1gITCAmUtMObtNGM3BH81UGhNPDThHT5XWJVvG3g8qvy2yG1ap1SQvyir
57UevN7zAiRR6EbksN7f9uIBkfKDz3bPQI4MHUHv7kjouP6u7Df596miKgphxMmZzmZ+3g2/ri9H
UEJjuEGcic5vEgGXuTm4MnZFXjQIWEC5lbHsXlVVYbCV/h2xOL2bvgC0Ny30auCaN7nGpC+ZB69c
fLcQ6diCkMVkfxF9WDgvx+5OFSElTptMhZZBPTdn8qFCZyXPX8lmGRIndV4xf7R7RRfHU0XvAdYD
c1HGp+A1bI6xVYLLlD7RHGvyly+xY9nG3hE0LixP8Lnu21GXYeZKsAuncoQXU6Ah8ASHA4zHzhs2
uLbPcZ+T0FdBzz/rKaIPW4+84YXZKyU1/WEXkXb7/EQlNDF262TKR2lVbERmTPnvTQ2+uVNoEcSj
MXGfblPHA8XKVf815QZ+GYHgSuZjjE2+TWd4jHxBzXO+MmAPGn7h2v6wz5efv8+r5/DHzXecG0rq
G/F3b6MSnYlogwAZs3k+AEt8wbm4rAMQIk3JU2QGgqjeENaibe4Ux3gUMqy8X1rS6/1AzYp1EHMT
yODg5/+JuLex08kr+HkiRn4EinGRDwzDqeVZWMdzcDUW7S96EuWvHwAt5iCzzaJRMEVUE/30n51E
GKLlg/UxcWj+VmKvVPvUyfKX4ijArz9iZqhqxG32D15JGcV72QE8hGeAxqIEx2HCGYQrW/mFZ0RZ
ziUQE8OAtPpgLgiIczQat2cRgqnJBePHPup7bqN5G3HztHLJapEfVBOoGLwaH6kuS67aIfWLnBe9
YWpE1/oHjJgESKT4s2pcjHG+MyTCGAOKRFxwGwKxCcx9u/VxlKKv2pMwqcUIZI97wA93a8Xdt/of
Q/Y1ZnjAD4O+eKPgY6+9IFwZZZB4STpifdRHHFn7eqsv+J0nff8V04sCPc/di72+4iRcasHcyew5
UuRoHhE6ekPIJO69QQxbF9WgmHuFxaSmJzERSMCXRF0DcMpOZb4SwO0FDybn6DwAZI5WhzDumxx4
sdEBELSDXE/s9hVYNYa2P3xsAtm/eWBV8aQUg5WvpTP+wHT4n1KylfimDUGcTsJDJTB8VIE2CI7+
B8lWIpE8yVUxMhf2gsy+Wtchjiputyyz3TZ7bwYNXysNwJPuKdqH/VWHHNbYyTT5eSi1A7kePRpg
7uVBFC0nKVYojIDSByb1OReAo0S+Eyrdpb8y6HK6U67PF94N4/5Yw5S/18H3kms2qutFsvqlT+VD
t34qO3WYtEkZJU/IMVC5TpC35tZu5J1umkw/ATntoxQJVsRkoRKqkEQ18rR2pRw1atqLwV/7bNfR
aawPI9idXym5j2ekAIsK199T05jOycRM83ThYCqzZ8FXh34qx4YGjGLO1vQw/cMBKvmXA+OdjWGD
H4j7MxWbS4GhNzJM9KpCpdC+6o0mAr+JCzKF6Sg/VwV8seAST3aye9AgVkPVdDYVluJb1bgnGxYw
6ETVtODPdlrn6SsUiA9K/yD7k/Or0A/OgnfE0O/QZm4GDC5DaZYtZI6sbwXsCwNdngHDvgHtrQnb
DxSxTUS5npby5LIHIsoEgSTyeEMud+9dwlzSNF9lzMYWbzfrl1px1TpGaKbvQiSeThrt6QyQq+jW
b4jyYBArLftOhYubIUOOOv5vZkeEkgs5cqFGoo7+NAlxZWMQa6J8U/uSEtEU5/aWQ6g1hK41IY1x
CS2kNtR6zd4RWvFfDg4Ce6bKwfLPuyHqL948xFm0DlTADZkw7IWNhZq51WwaVNv2u4B+mr5cEudq
spMmaS2ePFamDf4NBYB633mFdGH8zW+v7jLu/d7nbU/W8v4ge5oy20HEIMJmStugQNnlbWMurQk+
bmFDzTYAOQvq79WIAoKJO6204LEErMgkCH1i6oHRyc2m85+TfncN/NIjhudk8QHZQAPIqaFllg7b
cUHSybN1q8qYPl+1Lo4eQaSMTtP3yLwev4Fhse7yfXooM4S+aaTMB3u77w9gaaNShYagerN5STNg
0Agxe3hxFhjRiYascoDTRisQna1hReId5H7iOZsb2ag1c3tPp/gRZCaeHWarTw/RnlFCD7KZQvUa
4Dx7MDyCnNH7VDHEMF9I3dBTz1SiDoJjawX68aaUP9A+umy/XxqCJXEH5DIstbKW7snY6bfhUrHN
Vqvbb7E3xRvsCadpqM9VMYzpASkgDGSApTs1cuId7v+jnX6SoyAIaU2ESxmeGyY0LUutH3M/K3+4
VZ5LxoW/kc5lEB71onrPNr6M8rU4L8e0zmmHDA3jHbkSe7YV1yJwYVqZ6FMKEy4fInEfItbIFZiz
7P+4Nbs/A2PeNsXWlmxdXxe8f5K+T1Hb4+qTaP3wqXUU/ePMSblpbpJT/Aq4LFdD+6Ly75pee3Dh
XuQ/UGAQJ8B4IcKk/zDGrnA2qtCsidXhPbq7tPP+k0HNJ02eCZKIpfthkW55xoaiYWNxLTdOS8o2
I4+uO6ZqyvffldXJ0TqRwlBOjPa1XCtr+F2H72zejiZsrcvq61fiGSpsVfRT/9e65xtrEA3Wgf0a
rBlV54/sB2faPB3istQvaTWHbITf0K8kvXr5qhzrkm5X0eHWflWrqm2eI1pPsFOzCzzVnlXjxgnK
pBK+Nz/fWLVY96xkllzeJys0CUvvkiUN3I1Hq5GxXG+UgKrIZ/eTW8VWgKnIMJyfEMxVFKrXuAHm
0CoMxEU/cY4+HDRPstG9HC4hewExL6idB1T1fUETrHpbL2BBW8WG8go9GulL+QfZaYqSHfkT0RLG
jTMv9+RicXBbCQ8+FnkUJdMbr6xBrVG+g+lDUoxlg/YEaRHDB062aRzr90b8cAKOFpmeYHE99u36
HNqDjHrKxe5FT3CahtIdPcZIQDu9ko+py0gJIALtlNfOFekneGeLLV5Shfv3enKGpcIlXRkbUUiY
sK2EZihdab6zAp5+ImBvrtEWwDRDYCo2/p5dmgbeSw7uL/siwfH62uA4aNLiusQ1TO+tPruJBV1s
wTM9Ne9EiIhyXUlL4ZWEQPhdSwPNuGJjvjwhgVDtAO3FvN5zupeANevdw10oGlT2G9wysa2KwC+j
vdgKny9+Ks+NTpcl0E3DtPGYgNHqamjuIxgb3yKCBMPf5ZX9+o1lAOmCefRb4SQ+CzKINJ/IuSgJ
ps0MHbWlI5t6DDuH4MxV3mF6eRxIV+SX+nCy4vS8A5sp/yyWuZjX6eJW3shYK8ZsnUPFaofXKtNW
/L5m0Fz84/Lipk8yHnSrAkmfQtOfJhGCgelyYwQF1VQsFDyHYSbrsqX2xNIfuXbssfMMdxgUQ8Ry
tLbPwyOQKL3nlY1Vx6/l1l8CThjRH4FSvu7ETXWi7b7WKP0UoD3CjEmoTpfd5W+2D8ZVjpaIxvcG
cv0vYVQ5MHqZ0tXSd9fIBFEKjmBnzVBG0xmEHH7D9BPZlsUWs6+LYHiDg1CeKSETQRly2NrVw5dY
2ygcWw76t/lNMx1/27RE7mjqWYZ2SbIUmVcTs64p0iaYxFPE6gRULwObFVZ5FIhVl3Qx93GiaH82
berq6td7M9H0TDRX11G6VzJUiuVoauZHpihs1tqHATRO8DgII4D0qksoB12vN9fQTguVe6p4L2Vr
Xjs1aB53seOCIt6RVJN6L5z0WLAyUb3AfVCXsvAj1x3TuILFhQE8oXaFpDXOTj6nVLbGoQPk9xx3
odQG/lIkjbah2LihvDpz7o6iRzDpawvn0eDUHkjklEfPOSnoh9oOZYfZEMdySJ2apGNlpxbcv/DC
lpm+LykimxP29526zmoLN0QgAuv6oUwkSrJh8Yd7NF3ISkgYdl+7eC6P3dhs+E/bzE3fpZHq6Z/y
kRn1nDLUewezZXp7WuYVX0kazfIk5mQa9FMJf0PXrhGUNFCvXWOMMGanm2VL/dfQaG3stEb9ECZs
402fpPlP5fjZL/JrrIpgX/ctkMKQjdMLb1nL6JZzm/fwGS84kJVvfqhV93Lqv1Fu+VHt0g2DFLuB
mfUxyD8fruzjvsTon/kwQLCreo3Bld98zihLiwI61EqrBrXbMfY4EBYAV19YNHwj4XVLLVlnJvWS
tfpX6JRRRROUKRQtBbISRulgAJngi3wV+BwNDF/qrOrW5yC9GlICoptpwO/5s0giysNLgeJxrozy
3dWnU5c0w0A6n93KgnAnHB8DGrPZNEfg14F+aETmx06AhOkKaClztS12HGyvw4iYqKrwazTBET2P
jVPaK/L+ByoqDIsTqqmRsqc2iUfA59QZxMFtstejTg3S4WopM331jQR1Vw9TKxqFwc9M8GbadE4i
5quN6M68IyllQSs+LyIL4NflMW+dM8LrtA4w3ejL/FwEbSUfdfM4IxDzU6Vkg6LRfzVt3sBcHpCE
yAa+o0V3JwqGjmIkGh/uZ6DgF9V71fOQ01Otg/Vbzt/8sLlZx2U18EKpDu2PeLyEix9Tlzaz+ili
SZMsitZi35G/OIIyzerrTUmA+Alk6aKNdPWBocp/b6RF3womF189o/rJiFGoMIPkpUFP+86XkYdB
5cJfmcsTsmUw0jcSmC8CqINpK8zK1ZoK2djxMHwpJA/YQ+aZOHfmGQJyTBNe9rKKjjRN/wYlYok0
VcurM45DlfkiqH1vcDy3AqyK2ZrnEDDlbWZmfnCyIXn/WbiGGg0RshyPc2WfoCPBhVqmBz1tnZl6
L4BKCN4GUWgAeoeps66seExeNx1yaXW8JUBto3uzENah5NPI3VA9ZEvPh4ixw+OtSBICvVXjZGTN
E2lDxyYB0I9vL8I6bp5m4GnBC/XpSQ4jdnREbistqF78wY39n/d9k7mFK3p23q2pZhyr7zKmUPe1
7i1JrAOVj6GiObsPJqRBEjO2aKV4B87SL7D3n6ACSmf0GC7TtH16yJGPZ9cSztNtZrQmN9t00g3M
BfaZQ6MKlXIF7ghhSWDlLG9Pt+8bO9CAbaZfWmatx6evojkbS0jRKef8KdBLEHeGM8ld4OMb8hez
V2hwB/2BnjA+KW21Fhj+5MLqirLjZJpSDEHO0qaXxvwFlO4NHYJzyDpnX0/Vf6xVtQ+KEU+qMpY2
rcSFiGLnw/q39WL0sGnt+S05KqdnZN1p1fFgjtwHqDX39C1HzHZjsS5C44XCChRqEoA1nultzHQD
NCfBzQ27fmVANEV/jLdGJ0mQd0wTuFXOgIo5W3tIN5FW46DgOSHYSFyL/4ta4FYtkSLbtCpnw0iR
YSsyycGTMtJUHRk97gLQ7psCTFEjVWNy7oYjIS2NhsdBHTMK80poNGlkL8pSETjlF01OWgY+rqpL
hzfqeH/qPWiC/PZWS2wJFee/Lf8b44MmVBeZouAvBfF2EofyaFA/prXO0Vcbg7hSq8iXFqwNBZBQ
RCRU0ggmwnZXNB/NYcj4DbAWiVA7Wmh2xhyHrNDrYWzW95xy5JU8HRDWF2bSLCY01Z/y6oYkzm5l
hbsrEfdkXww3ngl2KOFWJdgJNBVfFI5Y63qiCn7+iFFf8fhJEZF6l5hJ5x3qOjp7d2f8h4Dhodqd
gb/i0bGwKLQXfpnhQnagDLyhYwQdDAljBPdRyrqGZV7nKRZ50shvMmS1N8l0LZwxPtuVKJCLavyi
2UIyxXyg+HTJY6RSsd039RhJ4PefuVVt/Jh2loE1jn3W3usw/yd3NmKXHkHbKUMmnstqjVpS/bvH
9FqV4d2TU/LOtheKwcIqk+76UJ/cGcpaZf36B/Bg+qNrYAJjMjsnE13KGHxBFMtX3hRfHweSKmpe
Eiq29K5B+rbMf/O68WQI2EjBTv26QMgrEMLwUCRVLmHD4fDnjzOrI6yX03pTuSng4GqIjUKKetDI
t1Dn0O0gkQwhA1Pdz7PWzBILFL5cVrK11ID1uBcZpqSRzFS/ck689esKa7QweijqEFu5PojKYTZc
OPui+mHIkwO7VMhlAtVoPf1Rtxw5CL64Rb5a0t8tTCIqzZmvidn7DpscbBvaCi00gA+vx3a6mt2z
XbiCFvjO7wSV0qwAKPWiE9xkNPwAuYeusMaMTeVLBO++waFLsnQv05RQmMZBh3jW8VMu76OXZDzy
XUOoCvRypor0X0ENrivNFL6NLLH+3u22hKFwzyblV8fzKt9QB9p3qo7xKsVR9xWOp1TDLVyWFSzO
0mbpvk1cK8VPDLg+3myGnYdZasKFIo4SA/mnmmA5aDshmxNYHheJiuXMWBeKEbThXP8ruRUp+j10
0J2WzyfiAmV1d/qdEnoKZb6eG50mNxQZRCFo9N9CFG/KI0onq6EG/84k6/oFvY7mN0XVqfq50i8Y
Vd7EiWlhPRggrhJnnWNwHSyAQie+9MUEG2SLoHaEKedxifjTGBcK9Hlk0TUwl6SlEmWBYpBOp3E0
DHFVRgyNbAaD7ejtCCyEbj0WUgvdEp+BCgSFbk2VXXJkjVlhW/BSvq4WxQuZp/Hq/f1SqU4UACVN
qZEupSzZn21GUFJ3lOsRdTlWhRfFVFf8gM4zHf5Zp1ROah96LKlnNTXBpmqvaonY568p3fL/k7Vk
mJmEegoLGvFWACXs+Pv1l5TnRpHPCY0nUB2O7PxoqWawX/ncwqJal3xN2A6QWOYJ/bm8ZdjyHmAO
Mz6Nlb1pHPxc7hxpDpID75uqRdUCqd1D8avn/SfpypyiGvtYDPyVT1kv2QzEnxWXfvzPMQmh9vNg
DeEQyg99WYKTWsnBnUJ9QKYYYGxSxa8M1SaQFTn9VZP/eFw++Iyh6fEJKmawbALGFV0B/qw1qnBZ
+TkVV08fHn0LuG2BeNOQg1JA6vj7brbNpFROlIClegvH/uRV5BTjuWMNRs60geK220xFhtoOz6sd
PmanYqfET7c9R+Bj1wRl/wbKyd0hZ7BnsrTP/uJ8cTmZFHmwjbYUf66lU8qg1L3Mf1lECTwpIqE1
t7PiNPuLdZv4fB0h2SeLGkdITy3/k3FZTY52U3kcZP6ZoGLDWucvGNuqZ+SqwwyfXdvJRLaH5JgU
ICodv9SJsAmi3S6jW4g8dl0MwOwIlQehV24u+zSmNR0c2btcIrd582AYkBUbg8ZXrpyoSL5Qh30l
b/6QZuRoWbwYeCLM0YWP0vD+4zoWK0n5sQcREcgR99RkdxGVhsP3aZHyhF43clA8U19N+xgI+PuK
+0TgCaq6CBO56XbjEZSGXUvU8EXXfMHeov0gLqS/1HEoU/RxTpb/qo6lZnNeUnJERc3phqx7PnyP
7USofmTFp7cDmSlhYSLzruHt0YxeFcmWL+sRHtR0OvkVwEWS54N7KST4m+5x/PMIED1Nh0keXgyo
p92Sb1sg2p/s2q3co2jf9MKjBUZ2SreNj1qvS3Pazlmrs7V+JO8/B43PSIoNWrUbRQ1+vUIe1JVt
lDlAgW8sUfA/yOpRKg6ZFScixQjsiGH/GGLrBKadKKWH7TLozFrv/0tURmnb5YVJqRl/eWzkbnRp
5Gp66MApN/JzmYpRwVbJIsjs6Wt3AfWptvKIz5JrnjcdFDsi8Gfe5qlOGDI1z1Uoeebr27dUnfWx
hmyHsRvOmPFk1LYEvOWoQep8CEm1YQ2E4Tf9J1mtw7Kn2NOEKXnUXmTv2dRYejVwzCzidBf/Kcwd
jWF8URTEFm4uz7E+5yDFxu/QXEQG06eJJywg65UkaVh9f2pFsc+thmYoXA0BlUuXnIGMG2Gdhyy2
K913QMWY4O9HrWh1OURkT1ezrsGJlhQyyootjPLDg/CUb0/Tg1JyZFFEzkn5YvYjwvNMIt5t92LF
AHl8Br2XY8UxOiDT8FdrF30aF3aqDDaRUf8WF1YTb1OVJhBU6Qt3GFUduDZSxsJUbYqwqxIgTWW3
+WRSImrnUZumgjsAr+4r3+Q0xIEg5YOa614bHkE3FhetjuGqSuvuWFyc8tOV8kVeqfE43Wxcnq0J
SHNzhkstIFjrYeGp4oMFAT5XL3E1bJaroPBcgF9A0ay4np5hrhlvfL157WMYI85LSEtC67yyKMXR
4C6gtOZrrk26aH+h4Rwk8EjzpKDqCUcJEOsYYQ3aZEsGW2eggtWWkXbLSDMqNrwHB8+9RlhA/gqj
3R7FchibnZbVmhO9DEac5BuoXqUiWqkeZ4KqNLqMM/DbwkmqHczqs8vquUlaYAv0n1Bud2bZJVu5
YgSyzibKc1M5/X6a0nWCodzJrSr6M47mpc+ORWGE44BHYPDNCn7HK7vswcUjjXckMop3vEXgvbFL
V755OK55x8ltWmmlNCEJRjHYyI9yw0Fq6auc1cAMqmYtLkHVcLNn8rEgvHtKoXu0cmFmsxmpxxyp
9jTdFu4q4frA+7GewSAriCLoo09rlJE23sqy1cpun4QMHyeRG8djR8juniNc71lzuylRfCbp0p1o
xKdgFxbc+oYNrHVmDY0FuOOqiJdLmLOuovKA1hvfsxLyPljhsPKSfK52LBbvfFQ+ZGV3bbsA7HQr
VAb82n55yP4rZkVAUk98jD+2eoNiD8pHWBkRsQoXzzLa95dRMbnk7vxXnN0WszN8UOJvKNR7zN9v
DZWilIewuFsIu0Mz1CPNDZ27XgMPKxFEcpzxeykl8eYxJGkkHGNN6KqA8NMQ43s+PGYOKCOzeWdO
QVSE6s2q4UIsbEQ5tQDZRzJdp77nOJDSfhF1TLEqkqc/q6s2aTHfAwKAJozx3GBAG90YCGfVI2S4
NRKacjynnkO+io70F5Yik8D2sV8CXd9NbPdIizPFN3wWSlqK7pbw80O4MofmwZyMXqtxee8grxVz
wyT/fOOcZZfBdFCQSGZcvkv8V7cNJje8Yi48WSfBzS76brPXMHIxMiBMwWpfkX9vq275bnD9pgJ5
Sr7XuLwJrfyQnHtw2dljBCnhZJ7b9sQ20Zitnm7caUE5KNrYMFyYXBX0rbf5Uycn9ezx3j0GRrqu
2NRl17WCVSy4hkkd2fh15osNHGdOM6oDBnR/C99Ae05UVOW9pbYbLKYutqIyuomefUrZB2UVGhVw
FXpC6uySW3wfvnbnIsUi1sE1G3xQqEKeAuyb8S/kP59lRmh49/snqSl8rLt54VgNH/fO1izdW5Ah
k/t9pfn6MvX9ovym43YGOY2/8YlVT1eW0lxq/L98Vs2/2D+jwgRggyn0sA93UK6OMo6NkNcAVpTq
dBzaESwXXBgq+n/6kKihZxE+++9EC3ODiaXQ4JlBITLfHjZ9AuycRX/vPk4kZvAsHj2DQXQOZrsw
n0pjoDLmnHhCdnPERzONtH8BTi19yc2r+GirjcYa5rMCorC9Yv5jAHySKTIGQgJm2vJtJLI2OlGC
AENPOSi9IpXgyLM9K0dMCfqZFvFznK/OdaN++IJpnE60ww1RQ/DjueW9I2eoSfDhnVNTDhfR8jb1
mFIT7FfM++Sb5Sa0tTW14zF8qV1wAzIBPz60uk2bkOf24ozQ66YXSMe6jarZ14HdnWie7CpR9Ets
RnryARL7EJLYNu81u3Kpq5n7l3Ra/66xosPMwdQ7nezksDwnNlOM2AZLObcA+bWOQGdOdL15N+RM
34LraFXvlcBrhh/5XWxQqof3/SWEX3XbB4a26I1EqJBUUFsyT5GV51l6Gj3ceQ9EfeDuiesChKUW
cHcWfvK3I81y9gh/YQnLY9ydiZLL3frC4ScoPf9UWLsbEJBE2w5yDlSfIv+KomgDgAHvq8iksLen
sLEDecuFfEYCOrL/pNF23xtsUJbcgE0TA/hNrRrJsRuxzmAID85NKUCOvT4XOXwgtW7inLTzuDnh
RQHFHhw59XSXH4mNx8vkVzsAzhxrN1h559erFFUaeOFVVVT1Vi4ONDPEm/Kl0Rg8EGPArbXXyOC8
5Dyd5HM6r9mp25OkJDmYuKniGvRn+FUqKnCxhj0DqpyUOW3SzhxY+aCL1hwgEN9Pjc3uuUlGIXF4
QUJzZqBfefxUHB499bbKsaGmVqI4cQRldDSJCCCyFdWNZ9nV7dohNmU/NJz208AN90X2LSOWPU/9
7lNaDIHPSAz27I9yObamC+89WuRDdlxLC/iwxF+oEnMI7RC4hxrPqcjGFZM5XT+tkKuRqq6brs63
IWuCJ0JhVRpCWMyFv2wGsUAo44VemfwOVEC0bNtmAaeJ0ILgkphPDYlcRtc0xO3jYYpEv4bKTOsd
EgrhGtluHGdW1CirXQXUH0DYCq8HXbxRgUNsobjrUWoysWR6iB/4+elEP1Ac7QGr6E5CDWEvX5Km
BcJ/DBvpo3r3/+8VAnnA8UZv1Aq6jVJ3krEB/v2ff0AQ4+M6KMV7mMI+un2YX+UZ4jm7Jdz96LpS
BDLE4j0u/TB/LFyaFTPxd5g3sdaKPdwq4d2N9uAV/ZIJa90ynXBOYuXQxEbpYGFvRX46bLsNlDG3
ehJYJJhMw0YCI/sVnO+faP1KyZPQvQRNjvtWsSEWzUtdoFyBkdCLYrEIsUCv0GXbdIwupB+dQ8A6
/se/EdBAMFyaYzQj0l1+Urm4ZW8C6K69JRRZwrrW8KmmG9lVybCaL4/7Cipqemj4NoMslSc+merH
z8SEJoeJhtK9vxtkl27L7i3Ou2yAJ6QsZDvlTfndpMiCtu9furQyrj1WrEWQRRRAWU0AZ30ryFKx
KB07cLQrEIB7k6DEuPaLxECwPJRpAj6YaXPx8btbgMtHHAAmu2u4fiHWHY0G5mLFHeWhb62XjrJJ
ebyGUeLANH6jih42bIRETPtgxX0BrRA6qV0GJiArJ96rgS0ot/gj5KXbgJrFJLuJJWDb2YX/3HBK
Nf9UBZnf+XM33VxohzEJVhKzwd49lP6znbIq+oXzffQfbETD51QphEm2A6VcAmdhllqXzdnz23l/
+2Rk/ae34bvOrpmR+9TB2IkUgAEZzEe/xsQ0JC63358U2igsBDIfQaQfZnWPrKD+bhMo5kAB+qlS
Ps1KS4T66wwz0Azazr6F8qnm0klAKwITFpY++lNeuErh2AmetcGLNoXxRJ2d40W42RediQvq3IHP
QiSC4agNuLxRCK9ZB4MAaz98UnESjNGSnOmRns8syMxqmE1TP+WsCC4eY1u5IvcNPPlcqtoB9VeC
xxSj8B9VL34F4JOiruqRQUp3zljBM06BEVQcOqSza3LL/sL4QIGctcBN8sEbp3Xehvt87r49F3Sj
yGKomyrRC/yqwTwJU888Su3IBGfw/Dw4uiO/VqQEskXspF9AsWjFV40C/MIT3/6ot+ePIEM0aDR8
JyFWs/RO8EU1nE00FKSrAV+5BeJ4Ntcv4CVbCOdOlSaClcO8F9nXLfp8BWBcaK+8VrRkVR+cbuds
wnWX9elNlKPmT07mSD9cc/W79jL2wX2y2xp6c76iCnhfr5uH82qAUKjOgd4ky1V2Qau3MFAr2krF
Yfxn3poPc8xnGNkrohQm9VJ+ipctMR+wUQKqSWxxQt2hyRmVhSq0zACzHvvLtPH1ytFQZA3IiLZD
XUXKJnqxqVOhaNLCdsaajKYDR/CKB5+jpXIWEcT5asNBM7oWnJyVh+RcZwKuCCY/Kg84JAKopDKX
6TrR/1RJA2HwjAzVa/1heAH5zLMaNaDKavPvg4nwH4hCQ/Zm5CQKUdsAaNWeMgqMSRbncJ1s2Ad2
+SjJfuOa3zPN0wyjSIfZ2er4P+NeYzg0Rgni14AlxO/OlrlCz4zIOg3FvCx/7v9HAsfqBhDCyFYj
SyfS5KSpvHI+TT1Lt7gJyUpMgn+sE3SoFX9nNId5kqgIcSLFGDHRD4/Z5ydYy7PRoKOPagSy+o66
lQKwnU8zYkDVmghcXDrsbbULM8iBpzWSDTflVKCFBPUIzfxi6W/jE8Luw1pQO0uN3x0qWBbtzUPf
YwRgwIH4RA0mNcxg2Bmc+b8hOPJYImrOn7gos5ZsCMkavy0OAg+pKh6AIv3Ck0NNEO/nLmGFqN42
GehdY69B3znBku3Upa45GOWK1n47GM0GgpsvVYIkjugot/4BSWCiucaLejG8Um/qWLsm5Atnti9O
UpGBZziGtai5eMttA9WtINDu0zJaukNLcLo8mXozwHRpizFDFTL5Q+l4ZOICG1ISxQ6xZZZOAXvm
VTEXZXqe/Itfd8CBC/UbOCBzIdkjo1hCmtNUsK0XHlgi+iGKVLBByKj8p0P+KzUAHpN1GbvTeBat
mvT9Ry3uYzgLzP1X/nZfSaK63ZCUUrEiCf5IW/T+xX+DUno+DHjIR2bKGSYg1BO0r7o9mO1+ypUH
GK44vB6ZhohjozDLMt0YoMaEtBaVxLYNnVFxPeGz0FBS1rNJzinC5/BXHg8d0VjMbnHYn8GHMN4t
qGM8KRMxRhNe/4taEnYmsJCuV3WwAPXPVFo1I3/dqr4BZBbLd+8k5VIJEiJxKcfz49oW6HtIkBmY
XLzASErR9GYafFZMkN1QkIxtKpoyhoZKe/aUXds6iNGx/Srr0Vk9W1QawYfLIPgMHrG50v6q39Lm
Iq8X9HamkC/D5pC+LTLGUGdMyZGPOqJBvMYUstG6enpWxnsl2f2vyiz3A9CooDXld7UE1DxxaBnV
Qpq2mhdc0x3LfTHh/AIlWsJx1dEZ++kknBLdq/xo23/nYac3xpzRIKn/IbHXxuWxfqg/AAu871XD
FwN6YsDmDgcylxoVIzAdgdkUZugU+U1KWqlZvTLp3PjnKwL3Xg46EoZI2DOVwNzC96JtvftXE7i3
ZTtBaYSuHK9GdgsSSckU7+F3TkR5JDedyNbcOf/erT2tRJSOdV9+mtg5j3QWygL9LiBbl3sGA9uF
Rr2avp5sJew1J7gmBS02EtvSv027YKaz2hTzm+HW8J4rh9dCAxjMf6IOi50pCiJyQrHYPHfBd7Dc
csg1hzorJVDvKaV6zYYTE/KcovUPuCuomZa0zEiirTMdJ8ChzupdN/NZkZ6Wf1+0SbIaHYb0wOq5
tBvw3Keu0x+WaPhBkhwgpQ7J6KBf4+g+QOXZOoMzswnI4Ns81g18uVZbEftDSNcIeY/LfUUAaiMM
Wca6hOIBP7B9evm8dB0I/9jNY0mhi8ThwowpV9Q656jUvtJX4SyFBuOOsoeItI4kckG8/yG2Puvg
FPhgR0tQREgdGTP6fnwcT//tRZkFX7n4VfdoTDSq0KfCBa58ZEF9LqVRJYhQX4OdNHRtJEup1q5Y
o4HirLlynuLmdgPQALYQnxOLtrjfTic0XRbDimZ09Vg76GJqqbYq7+IovNLsS9g1JzBIWJDi+2gi
SHCbGEmk7lnEZVEF6gqw8PVbqOqCxzzn34w6ajooUK3wWgmzvepy2Q+82QXZs0HzPHaDn3UUvAlx
rlqZxo69Kx+mpC9kIKmPpzTSmwpHv87iRZBYzVfzCXLeFNna7oZdzLXsC/i+9OzDNy9vNY1JxkmP
96qyQCYksgtYsJfE4uklBCzcqFWq6CTjPXMmwzFIlngErB8UsKzSlzY8r9vt5scc9ECiH+Xp4uNi
boLp24rxpn8gXMJdB5O5/YzV+GYeB5cz4JsEO3nsEWUocukkXYlb4JzBNr7y7q+9uC+xiPypIxSI
no4aC6EHmXBgMDwsZ5AMhIVLp1k3OuON8NboN1RVorrbZoCTkMBN+1Iop1CKUN/Q5sjAysPrcfW4
WMyy3qf4csPUiE/J/uOPRMSKOxV81WM1Efl5wJ/cuP//nLroVFNyXBfDZ6aa770hCU+r4faavFHA
ewJ+m/Grg6xNM/AXAWvMmv0jKM18VrPKyDqRx7iff1dC6yJaOcc5Jxp3R59hH/epeinWdadCmvnJ
L2lhSe08f0cXj2n6/pyTNblVmD8OLLRnAlISqDZKVyE2tfudqUGFd2fxB27KYor9BMkaoT+LrW2u
0KUOieq4OYcruSjMnkeTDpG/J5UrI+OpZ0SIq6kRWCmPyUZ10s8fJL46S6Y47LR63oM+3gOwX+Bu
kADZO2bLOqbWl/7GE/b+34dEm4kL9Pj8T7+xhBbx4OyT6WAZGLZ3vZlcy2ykeryN+OI0jKFyuiGN
h4Ms93dcn3l437qLdu5LDq7StHKlREx2cL44wVteBd9MyzOnMAugheL7w2RBVD3Gh9t3237D5x8k
WB2DrOqeXmR7Tn3Ch/mn7Xss1B/0H9a4RgqMYX7kNQtQA7zAmmwaQpa56TAS7Vbvvm8Lfi0BMZAh
N4KoTE35n2C33wsCRFF8hFa/c6F5TcQAsZdcHWv+J9IWAQejRxFRtb31oCfK7KNYsTguA81xTado
lXEBfdAqo2AzlnCER/3bvxESyDw9iMGpWm5go117p9Vd5rty9sED2ZJOXe0nb0h1cn5l8k+lWfmQ
7M1q4D8D4sQ2ITb734dh/rEvo/DYtBJrNjppVjA7v/10kNr9nOMEmN2odLFP3VUXO3uo1OrWEP5Z
Lt7/cjIHxpZAZEPCxCsJU1iDil5JAE9paezUXKC+n5mUaW8smGQrDkiAYbcRiBmrjLY0PjKJWr1+
O6Z96VKPlEF2WgKhlkx1mAk6+D1S5DJ1sNE+9X4C2Zhc7D2pVPH6dHyewN50gNlZzVBWslu6WkAr
fQyeJuEZ68WJLFqw8xUaO3Wi2EEX97OpKJPt4ux7ATZOuW687eULOYZvFEEwvJaWHLos0+kV4B8c
v3bdTfgZ94QXitXRUXG+mkYmQBl/QNiGmvq2sB36U6n8/QvqSRO3P39oHW6cXU03WkdbhfohHnPK
iavaN4aaIS6jaACZGiWdj70gc1x6OfhPxVFuLyTYgqzYvqKuWN8koCWcLkoRBy92jiqgdd9mofsD
KoH0UrjCzyHTmYFIEjFY3DhUJrslJ7B30PqKiVcWeZU/mehABWIKaDvq98Dyl4gN1xvWnj2qrBDI
c0uXbJYcjfzXbFe+e4IlXr3e52uXUnifsaNoWV/kpeqAjEfBc6LilfDiLuUM+LwRAPcw3vY5b50j
7fN7FUr20JwbLzFJ7M34LUqeyliIJVO8h3yXwHgBJdk//oWlv3+Fs0JSPgxIk1fmzwiX4FjrUGy/
Ww9CN4mGUr6FTlihI/HaR0p0AIVn3YKxM5MoYuBtOKxcd499/MC4SX4zbhbvbV0TA/IdMoM4iGJI
QqB5kK27pfYaA59Y0rGy0K4mK3RNhi7AS34oWxRiesKy5Fl3v4bDBwdHle7VGKG6EyPBxKXF02Hh
pEk+OWMhqov8AKMHj4YSV3ZaIfWkRKX4av6LyIL/1V96dSxCClQyikeXKQQ3xks0XOvDdzuTVVJz
KGNTaOvN6lJ0eul4k3pwW30Uh+OlSOxOzAszgg0kgobaJerv/Su/56L6NnrXapCkwpm3vyzMKFAe
Y6SrhyklPBAmqQxmxnjeP69Np1caBHsxBCH7pIDx7jxpbNaAC1mecpdFgkPj6wOLVpXXr4nQB90b
KBI/J9NLL4T5oTc8vNwzfbcYQAO7KFRVAdnB4zpGjoIn278dcYllMenfOWz3rcroBNsmhGSCWC6O
wDuFInSIUGeB8nT9nuCmLl9EBzW0CgBM7wij3hw2CMCugHrUgj0uz383GL/APIemGHLkT4fWwa25
PdymN7QDjww74QEgD11i+i3mcwOZBt308fwijg7qUDz9DnAlq8NbNXj3HZvZfjeokEduXJ2HnglK
eWFbSN86WuaegCfh14OGqBcpJt1JcR8yRKYMCEctkRZrT2tgy+sasKRW18k1X7bQkVGXBUHHOHJd
xN1s8/sqZSf4p15MxPBnL8L3QwG74RkKj2HunSaXKz7FYvg7Qj/Eyft1ugQwqX12fOssx+NLPr6f
eJjoi7uilWMJPRyPzNud8fOE+XCN7TFSDlbOTzx1ZZ1azQlrPaZwMfO5QlGsbKNSqgGgUAvfITPe
h65aivRZM7BiMxl1pmrDNvMRgT76O4Is6rj65aAOu3G1FJxAYnwIvrG3xacT86KTFHmQhc7Q5T1E
cyAxGAboL8ZZt+27Bc1s2afFhYKUtXeKqdcwhaoIZpJPzJeAsYYhXX6Nzm7wBmkYmWu+pGgMHGfV
IeDCLUeqidS5Snhz/U99rR+ulfaai67DxTowtwu7OBh2LEn+VLgMJ6TWWih8qr4aZJL9tcfcb30o
09Jyr9wwDD/3RKgPDYdqV76MpPuvxaM7h3jPi1AqYXwHWkQeKZHMPdND8gp4ATr6ykpNDq3tcIgD
QbpQi1pulnynXpSNc6Ag3WzUZ4wKztiPe92ro2hS++A2mzHVFo1MDtx+6rymQOgPSl+frG1JcGLZ
j9GO1eR3UmAHLmEQEQlsk+cbReGuGFKkIfHKwcct5Vk8fCL69uCzzZ4Q+32W0GQDrv+f+XGU87UD
mzSAWpJ/5Nnc3zvH6K/MPCfqHtjqsCSJFN3jyeArGi+sORV+wb6Zxp7W4sCFSmBmaIvujFCKFcNx
VlCSCs8Up1bWhaFuPDrcYEuh964xCrSi5MQmlVYob/B3Uur0vzqzHICln00RzRgxnKs+nV8RxYHV
VJYnn+JDPxYvTRAGcIQHOVk8nsrYx4mGNtYaFVyV1SCYagEpZ50PnrBgrCocQnGm83VFefOBBHg9
36kq2gc8DUSdqjmJscU4g8kZQ7HRh7TqRg0ZaJssbA/hQeHj1MkB0thirR3N7TTCSrILRhj9JRSx
MkrPWS+/OcR9Tm4r3c29QM00Hvk0jUeenm1gsZj/9hE42hTZTsKWI7LzkaQXzAmtAfkB8o6M1LPv
txmGkWy/N53rroS+wo0cPaFK+LFoJJZVjCHHA5SdczRTsgrt2VAHyLNlqI9Fo1Vgr7BHKDIADaF/
8FUAu0ebyx5LrlTFkJLk06x0lDQF/DWDC+d26A7w1J7cbwy06bbLxqNhUo+T9JMXu9iOgB1bbx+7
pQMe+CV1KJ3r93pm74ct6nGW2p8zTXBdfsQfLwZqW9P0DH97tCAFc9zK12PGQMCAqyljfIZtTPkM
dQ7N7F+uwUUm4YFnt/8G9ycsyXWXPN9zHrbrppFPU3AiBxA62tnNJder1bQUpdnj+ea/R9fVapBR
fYGWrJyfdSagOpQBcoBRE1ovlkGdZF0T6VIOCqo7l2eMh3TeS7T9c+skikTns8Ysfx9Jp96U/ozU
LyyLYjxYzuT+rnI8GkMqCPN1Pe/QgO8oGy79+QMq4FvVHm6SMvpHAE0GvtvO/5kpU+9t6FdPM7X3
STA7AWmOCHdKSO0yxUAVCXTaFXfBzUb5vsS+TqEBOwXQzi5seUtbtXcNMw65zGrsUjntyBqHnEHZ
alaoZudoT41+qG1x6564ZwGt7bhgWyNcaexxVF9X4dioWfubUCaGBhq3WyFHQoMAeSWP4jiTVNJr
x5sjH23Opi3DCiW48ujrEJdaruTb9LQZwKWq/m5IAcbm8yT+vIUYntZc3fu9KlRA98xfC5WNl4a0
YR75oSE7iuzo/BARRWev2vgpcNZUm/qKRSIqTSfE49mOoVyKDQ/S//Wzvlkj38VwQEBpf2TnrrAu
cNJcqS+EpEcQHBpB+D5+M6ubv+Q1JaiOoOU3SFTmI1sjxHfxWwCp7FTtMO8QeJFCwxaKEzKVyDmA
LKW6h7OXVwFw7HZKi7jFDHqpvCXZN7QTZUkBQOdzm7KNC8cp/oHZzKHR8tEhLx4uiOh/d2lTAAPi
Axt+Tt2C6jkkoz68tEMYzeBR+xnZWm8Lg3PAnm72lUo0yx0+1iobAgRCFSQntcf7ERIFopjVaTQA
o98lQM0V3zbguBewCRjk+Oat4g5LKh7ITeoe/jHfHx1mbzOrgzUhl26nJuIc2TPDXZ5ZG6cRee2l
7AX1vtBOlkVYXAft4golrrd98qt635PT5u2L4QrJWIzrhs1NRJ/9yZb37hoEpAOyuQJr2/hE86Tc
sVNNhpq9IXscAqZPJRirCiUyMj8wudXW4eWVCVvcyA9Vi6ahctiH6GSzlg30G/wGSkY83ISPgiHa
+imCUT1euBcI2yXmhF9o/n+7a3lm1nq2aSGPejmlwij11oG7pjbC3NUgmPZ+DttL19adwppPPWV0
Rax3W1TWmc6RxDzGUtuTFcB/sFnuMBf5ZmWkWhidflLPijckumvJ05CB5GHbDIECxV0nkHrVL/Lz
MS5cdWaOeBOssnJCMy35Qkmr4b9pWl2w0IDIHoRShS37mLB9sye071ftL8iPYJmJdFtW/dXDFe0H
vv4O1WnQedGGiCmgjkTjDNl0WNNp7RbwssPZV51XNNfW8GGppiKiSl7Y6HI87x2XLGq1WU4lBE98
70SfaEwmhhpNyNU6ra6GemWawH/PsASmc2/RwErSr3VQjQcSoVxVW4uPQ3djn/ttqUUzfI2TYgjM
fhCRMthBBQEaD4Fh91WkkxfNtd3Go001b3bw42EjMUh9gmlKQcom/YJsb7J0T4x2jxbD/Ed4AzJt
AUbvrPI1TGGeRyo9dWgJn7ZHnJ9XECaXxgIsIH1Qf4zyNQytz4g66r1N6T0OPJ20gK0jOb/jl5s5
362fv/AoXPeJpkniLs6S5v+bdB4Iduvu9VlXLX0SAoVSHT+cE/nbaaNKUOW/VUSBSfnIb+M1r2Ty
66c5rkFELPJrC/0MjBMTTTlAIQuCRNOKjvKELdWvDh+j/oKxC7L62o8jBgIMWGoXfmK82fyi4b30
WlvXfPkMoeUFSC9KGEnWcsDfXmN+ox+zhXYZOAM+3VPoMQztbj7FhCdZC1t0aNQEo+Besjwf7VbP
iUyuAF6rikSStq116+0gQoInajAUNKQOWV34KOQ1/FeovLK5votN9fwjIjx0JuNuiGykUhzBXgzJ
i81thMdlrt8NaM3WcE0iUL8uyTma/LrT06EqXDAIdbNOC3kO8yXCZopnK/umwEyByL7/0GXladMY
2p0rpPyXdkIVBkV3t5rJiCu1hR8NHzrCUSPOQnEKzU0DKb/h3Q9HuWatHFquTTQ7zZMIU6ElNCPT
CXR5+rrQZPiTg47/TvuovzxRtIbbb5kWl0fWByW17JmlaiJgzaIOh8dRkXYp2Wv4MglO1bjQal5e
aVywvsp9ZmDQ+OrvKCnFzY3cpP2WVVStY2YBf1/QTdM1mUXwDeIiWlMioc4O7JJzbZI8/0Mc2Kgf
UzdWj5L1hQJOKui0xkp/H/da04SuYdqimb9y5Q2ozHHnQY7tBtG0EFUNhxmg7KEuegtdG3BqYKAP
xJ/U+UjaemOIJBNygzEbiomxD7+y2wr35874DGwB4wWQsN5V+cOhPrSwNb89otel0KAeKPoyVPg2
caaffgIo8xk7320LUrdLpcNie3bUN/ZoVeE9yOg5fczIuA7xk93haQr5O5Xup3C6Tqalb434HAa3
fU9WhPvqGRqQQxXCyYwhQoUYY3ujMYCuq1tg3N0Sy0vrgrXZ+ipN/Xa/0BhAzNbArgT/fsGZeTXo
w6XgPQHfA3ipu9Y8i+ovBZSRINvWhbaumovIrGNSsH6pQJ9c5RXWiUbmTBvVgKEBPINpGZnIY3m+
5HZfFR+ArjTjyPoMOR+vSBeQ1FJgfi6GfAVavGrESriz6rwNF452OILUgadOX47z4jYp5j4OFXQC
htfnbU1z+yOnRZm+pIqB8KdsfJ3WngLh3e5/hVHPrwmqUgUtnbH/MIKbFOk2mduX04ZVbp2/2sT4
Mmxm9xyCgmADY89uT5kTrDHOB+vAUghTQA8slwvXRI2drHGNS3Fzl/uUqgKCDNi6LDuFdqtHpjaC
NKjwsbqFRTYXd18y15uO9RTd15Usd+KDkgkw1yON1ql/bOIhbR/XHNEhU2JUzzegjdLL8ePLw4hE
ylv9/bkVc48RabURgqZ/yP4stD0+5tCxa/EShItSKYmz9eD4r23SqZDQ+C8kV6jd7L8TxDo+nODo
JlIz1RoHp8Z3QBiyyhqQE0ruxZeV41t+s5gKgGFgKSKJQeKzr5l7B8CrSwnGcpZPF3oQm7xoIevi
S6UYgTbkLerWeDSHeAW4M0pdXie6f/2gYRyrueV6j7T/rHqW2XidPn1X2P/SlLagIwuZVHyhqLdm
7x1+zRvuYfQiRDtyHGtHbFn1W2gxOTvMDSTYJkaFUqmpkpvULAwxQLv8vmoJwK3We6/0J3ljK4L7
kAhDbhGdWKMxyqH+CQMptHY135ik/iqomPbuRdshXJRZe4XjJG1Jes+Q2alwomK2cJ0c80OwXNXc
I87N0VmR5vTX5ypDXP2RQEHJmkVKDyNrimj8jkx1II96lRimmkkCC+EoykBFZ8cVjjJmYRwoWbLr
2VLfaVv4vUVnZ2TUXnLKfKyXtWbXuFfQymyOe3wNWEPGa9HG8jnwvEafa3RnTx1rrPOBGHTFFbQ5
7fYfULpD16QlXoxFwrmvc03WxOUa0Uw0Sv9TvdK7cB6eZzkshxM3m35nP2rpd0pdJgRZRwT5ONcB
G0+5XojMewvKzi4EI8fY8qCUoeRjHWY4Aju2VkVl37xfnl9rwF3DvPlRkFZMTmXh7lmcqr/D7vjF
NrGodtHqE3qTEaOPOAQrEAs5o1MY8OIxD3uQpZ5zLgkoRmlJMbA6fE+lLY7D/hU1tybLiDbBFZH2
VRjTstZni6/WVhSrcV5mxIN7hUKECyGWRcoGJbrfRqmTLQ1+89i5c5GwKNinnAB3D60Hy9qMyjZB
w2zLvqfyvZNXoKRREbim147SRk8f/utPOdOis5fFTEaYbnb0b2or/ffhMQoVU+ObUg35jjvu3NjR
QmWlTYVDsQWvNbyL3GRGb69IySXdS4i3jaWdFWaR4lvrv5SMc/NHzNem6p9WIi4zL9lnaAlJH/JQ
HQFNDzRc6AXsbLUPZaNCfwAjDDIGMANyozPI+VWthSgJfO+TVnDMo9w04f9loNHiG4hTncfpsPmm
5Y2nA5XlNlE4ukt8DiWWEhY5OIQOtnxgC3c/XVgkmv8Hjlvi2rO79AWGcA0nGBCwIgNiupp556Od
mrg0TxLbsAAx+EGlKy04Hx35jSrSgMhaD+GKVxTUgLZBFOqSkrT5T3eYyLOUxuowjELTf0kB2xjg
xLs2aNra+xFIIdAVGYe72imPV9ij6wOvkB0cuR5qmaBWljVs5VTJj/zlytthczgXVqOaIJnggEKS
itKWDBPTWXr8SlygCvmbd9LHc2VNMbxxxuHRFceYiFDdI/RRg10NlDJw45NEspEMiVOIOKT1qIKv
TsrCsBiTSPZbdQ5hDP8F7126qP04o9rHkgrgi4G4oZauKEBaMKj09TzcK37v91IK/SdC8mKhN/aX
+XSFoW5gAekSAKTWNqZ7a5vBWIeNb/M2VLGiUaqu/V2vz0I82IUaXEo1AbBSlbn4j1jmJrMWyuQB
Fm4Zr2A82hZHdx9dH2FKHhJtdG/mgJccrsn52O2fNXWBZoofp4sNROgFORl+3YqcBXgEUa9WkVIh
4pPVDOx2T2ckS7r80f2RuYaQqFE39Rk4VVireP+LP2GPqbw2uqz/dyHY8Ww6oYoMH53AwLjCWMAN
Sl6l2rlmODKdEBKje+KKPEEQZn+aKJ1O3Io4qDu7pjtwz8uG0dLPL3OOhKmXMiioIkvOkjqoiB4o
X4P507i/ndPE3BWTTVzH5XTpYlcdQHgFR4RaeW8zoAOf5n5zC87NQx0uekqE/V4/owZHfT0epGTv
HKAV22Ggd5UkEJUW5C+FR2d5VgEtw0TQlhPxeyOW22ZaJQBWrvOQgABzIRaQvYF85SQ3faJ7nY3K
aq4/ZewnKBfmvi/I4jBYZC2BeTUus0L5KSULWjlMR+BUgBlHlgbE8mxV6JII0Homfui5CXZEgqj0
Abpo++jPLUBBSiwgBf+Hv8CCxU+uxo9MhNpGQbVMG1s1pEzvv9XmRETV29D9+m+4/jrDpEs4FOgL
RCTwCrBvAsFUwnIshkoWufqhjD7zCuA3dPsBd5CHnZA3YpTROHeT9CtqvORmutR23jBWZh9qtKii
3O4rwnQfPmw38szsc3ILqKeCpp4ccYksUsV/IjD4eknIl1i6jTdwFxRBQZ7++vGkJFQY31i1UT52
zYWMCMuEoUuZC5gHrPkuCHcvtlDTly4+NiWXV5RXzwC1POrxcXh6zQytvzd9x8Xz/JrY/QQICOTJ
5PCdjh7uymIeHCBKELAiwm2pa2f3PO9rK2bFRUALR/9u4pNY9fJv7zhTOXbN7crL4RFq0prUS8Lp
HYWH7WvsrEql/LNBSSz85nWO6kiFbBGhiZUeuRfcIFscuPGfgiXnXoUu+H2JIEbzSqfZS0cM38Aw
SeLKE2R7XswCop/M00+MAxHxrknAZCRod+ghQvH6Z5g10PTTIbKFXRxBT/v12jJFNOcEZVKqfS9+
MUfsDWmbucFKKLZF2Qc01IX7QxvUbwNIA9h55Z6L7Hb2g6DKvxFfT59QZ+OUQLfLctY4vIyaKuY4
IOxOFAB4HfXIt6EPjv+kdzlpSbhcMg0tVyLyDq/jzjfmjNRSA6+lD/u+YjSy/jxao+bGEFyajned
c6Uk7OWlolTE7KIxdmlJPuby9jC7HoCzXwy+X9qEUO8e5AvllQuyVBFbTYHX7mkNKHJudi3LDT9P
9FZjzP4vksDKd+rmHtp3TdZt7UegtZMp8cGA2St20RoL6tMLHulSsKhVazwzBiXQf6XZQ7xZi1Fw
oT0R804b6n3GMYoorv2JLBTieCzJKQaKbB29iqngcV5iJXWGn7IrnBXVS/R6XHRZaXSCeC/JeSqx
ux9mUrq8VIYbxvHEFrNF2bFhsPr1W+P8YluauU8Gsv9E90NjMswJesh8poy2SnYd/1XUL8364dlX
16T6Q7Zv0pymkeaUq4ai7/D6DrSmUf7D+PJLP0B/n3qsi59TRVJ/0att0RV9+DJCVUxcN0dzULrV
kcL2+AnEyKEeYwjbQtE2QFPhhRnQY4FswKXLKhgKhD5ZOiEyZOJbOubjJZsj1xWzgwECV8NGYf4V
vTY7Fbmhs7PyOZ8NbAjI3Ok7s/n3nb7fb2gxSla/mayAKoCT3LhiHBX9eCrrnZ9NfCfhrWZVQKPI
HsCFcITwjEIbxlu9it8xmQ4mXkMKkLqRpMZCTNM51xXxZqf7qBbarriCD35mGdTUG58wybjkE51f
UQ6/Bw2Fb0UB2eoxMQqfNDZZnQWZUIQTnGc4DFe3ID0NDBoEMZxF8C00esw+6Kvyr+taz9h064/A
f78TvFnAJ3tXNyRgKpx7zg7E90ggqTwbTZRZhLA1gB2PfK0m/9c5sXaDeI5+lcNYjWHoqPLRnh7R
pJXkP7IdkNJIZpefmPWTo8wJQEPcnWl+XGK2uUf5566/TlFDn8zLdPMA2chPUyzeXKq3djS1SCGY
mujzdiTZBBZXx5YpKnfXXKHFyNricVOYD57iPI71Gx/8gd76L6cf+/lKb9yhISr94dWBnZFXp/U3
4fM4PzSn9/Svu2wRr1ajAFtRGqNykK7dmDO1cPjzbcTNjItkPVbpdB/7reCZjRIkLW6UHU1/f11+
o4gLyTH2RmA33a7vNGZMFCqox2ZAiPXWTMbxAZXBHh0j5hawVDnkROkS5s/ntaBw+rmCsBLydStJ
iM9WtW0sX2Hwh07yT/xnz/XXQMIr6H93zLcLwqiG+oI7Z1THqpBWjNqlCtmWHmqMuUm/iyOR74tP
4Wo2LVpGZC4gbmmri+jHLQV5G6WgDdYyHqmxLlFsUEISvAlua521xicZTWuePmwASFlMQ01yWqqL
hZFeHJoWEsGWTEyVXqm/CKiuJlQW6bZtJelqzJGdWyLwCyQiPH15hmjH9fXRI0we3xolLyLAdWI4
9vJ8Lq3V/19kzvbMCrZalWcgbyvGO+tKFsSegKeIxZYpmd94+XPcmB8770Na13ypHWAzlUoK2vtz
uoDntIWAnKLxOT9+k1jlV0BKWAE+doTPHAQHcR5Ad0WIPrtUxtE+5a/Vi5v/ArmIbZcTHBPXvdZB
sZ4nKZ7AWNlf9lG6kxEpM1xpBHVsPVQO/MIjsb2cROkQGXlolS8dZPoGCG8K7cPmYBF3cBEwdRpk
RDev3Uv+04ok6ou5naATuEkIOO5ZvqaNlnrlQxGumNYhqs0newUzDckslnEEsmOW8hApPmuqZ2SV
YGlbV9NkRxDpJxAe7yVQJAMG5DpGnxZUi14G2/wEBh+DvlGLcepxIqZu35J7/Gib0mUeRciJ/Lq1
G8gUqwIg/79s9sxR4uYgtBdJuZcr4vtQs6jk6NXrCYErQN2iE2CNMoTEawkxU5FuJTV/7FkSBrkA
f5kwT7b/oBLwW8yuQqIxwAfxZS64Aw8UOyu1Hx8Qu67gYVpDQVZjZjYdpiEVwbENkhhlZROuwyTX
O3q2pAfIUj4d8HY7JMSq4ZjBMO5izJuvOR3wLldAnbdNoVdXuMLK6QNg5ZUOZsz7UTt2YLiDjnpo
PtUUSdOmukb0CGMsMNkhdKMnp2lkzXFyhnJ5BUdkFyiCCTpFerIjofIeDw4X7z0eBgYFD7Mw36uN
wsmeKOeJNMDtVz0B8wKwcvPq2h9Gaf/wptk6UAYNBk+Am2c9h/O4xsnnpt8oFcXwjIDJN92Pdy+y
vbt3Gz6sW8TjxZJC1xHNPe8wDsDrd6aBp94voHwVj27qCi0ryHuc22l4yRjKHfcNtZRELMooz8Uf
ZMTWq3naYdoYp1mIexCuoF/1UWqqXb8g69Smzan0FO+g+JdaT5sEGMG2L1KZqnnUNqbQYjnG/dbl
zqHuk2di4Rs6CRYwaeqCWEXN8t2ZlqQb0btXhxjvTvxc5RsYNA0cIYGEzBSdUemCNaV1VSujqys+
PD8hq0J5h39gqgQX46fgFWLUCp1tdl0w+SYvysDdgGbB6gDWzwUPQ1IVqOaaSQgBG3eTRK4e4ruE
r2Z0XWr/jd6B4OownTGGVLktKv6E7X15LHJyvJuUzy+9hA1s9bZQCCUBy8WtENG64cLhw1roJhEu
jXeZqz45aJuYodoQ3dRiNB+FOxLL+EKxnrFYsvJVEgFulN9dHUdjg7LMMdGeYmHIaTbo3lE0W7Tn
gm1WpE1UicpYBEfgHhvNI94xlU6Nuc9jTecdo+rEhXMWdNVBOlYCkjiSXv6Q6mscag9Mu6a60xfe
3WgOoQ74X4JdJxk5ChcZRskVrpzfgWOYBvKvctEsNIM9il8jPZZRdduvhWfxU2qC+RAowk/F4h/V
CUtCHpE2Hrnm8jNwR9U+kKYWZ+YehUo0eO3hYmnJglvTqYmMw67GqWs/KfgHacOjqbocB8ilXder
2XFrGCcKtowGEDzaNYNhv4s57AdmdRLnbPtB5Rqf8hu6tupJNjRVl2c7RDDWIVz1kRb119ydRcTn
Jgz9jaQHljB8vsksdo//V280ti/KNZyRAMSx3ihkmBUuWwCrqUpgesj9ln8Qy1JdU4GcQUkAYWDx
eMP33rh1hDlhWXJqcLVpnsIUfienta7Xevqi5+nIZU7D6QKG92nQx2z9/voZ0bsLHaFA6bpG2Vb0
oaCxjN+nPShvZsnnS4uEBGDgsYlBDg1UTzpZ7Xr0ENr8CzU+JC4AzqI5E7UxOiuxDnND89UdfwTr
F7hq/KtAlrcvB2LUaiBLbvaSG0HQrQT+TWuAVOe9ghoay/wGutp9seVcjqH3E4ql98C2SWZdhGe+
Y9XzyjfY7r3+CJrEy1fH2ewsEcSxbWtmTFaOwKOsqdzkWBOBqOZR9m1k3fFknE5NZUY8g9JMmIUH
rT2/JeKOsn3ddbb7XOUQKQ+iFqWksp7SNMlVnNKpLkEaPBDl23sqmNFXdenme/tpqO4Do29w3UIH
43mQhBMqn65nrarsJlPqaRU7MvgfOVkH7hevM5p8Zpm1CJNSAQq1x4j/Afqfc5j1tUysTyohpgx1
eK2luj/uhQK03YVhzwd5uhCzSZtC6S+e6ePDq7uLsDW4C1tCmkhMLSflxhE6gCvUxg84zhXImwCp
5zcwlc6pIiJaQvy468BK1ERashdbcqZOe9dZtGcGWgwFFa8VdWyQWZH0IVs2tzuzy41d3pxXZB0M
Cq9XW/f8MHguf7ZLNl4y/+FR0RN7yzXWYugVCqs6kew9JZ0GAu4XBLV77hf1MS3Tr0odMjpMcFaD
TAHDGTmNViDlSt85zpyzqTETYYNyoyi831eLRs7mvqfeDU4HE0DNYuFmGAINJUUOhQM7DXzlAuvN
4Z7OqzBX6LZ2q2xNw9k8Uvswu/30kh7YlL2ZAfUS61PhcsK45SBIR4v1FvOi+TnEKYe384VNRc8d
8odee0Rdark6QaRKlIZTOfYaRzltzOzLb0e6PN/3Ql5+E/KHlhTBTWs0J9Vp2v13nI73l0bLS/o7
PJcoWoM1+2D5gaJ/3qdm45j8k+xU4MK6+G0CCeoYxmeyT+GWWHHqO5F8sKaTlOsDWxzCkv3y9Vbt
9wlOUqlD2nMUiT1QQT/r47BDvoKxM5mVH9WF0oMwND5nzD3rCsRLhtKO7RNPRwIBgBnwY2Fv7DxO
ifmWudqNv+kxMW+XOffQvMRVqc1YMBHES5H2Oj8iwwPQ95WbAmYfPvHkdmOyc3otp1Ix6xsgM9ts
xXbe82/EO0SyQ54L7bVJb9zDg2iPMoG6+riDCYKfr2dakVYJROrDPRABXtRWyZu9earikvUR+6Q3
XXv3ffDY4F+8YU9aMceG00veKI5BcQRmIkUEXfhKUAvRN7K8YnC676tQPrdwBcJTU1kDzOHGCpyl
aqUJIXRcVOYXZxmT35zYqk7Y8uBZ7evDaR3wYqOawqZcluCKPN7cxJCZpeLoZ1VMy8hoc3lGvV6A
VbF9xipj2HNErmv0DYVf5sLeXLKmG2bVDWXa286Mqgn6GyeKcM1IX05taVcN6RRSyGx0gg5p3wgt
w/c7x1Ys54u8KrD0nShAQtuumu1Ub6w1+qJ/4eRQVrhRxIU2PrjAJOCn+ArUHIU+8zjz+935h2Bs
86fxin9upTewDGalLt3nGc+8CNBEHXdNPFxpIWddTNz+4jcL3LZHO7Vfdshs72HAxe5ezBVVKhgv
a7vGlXNoby6pdXHxc2mz/o6bJr6vx6wxqzQgLpNMHSrLAODC5ukL3szcGgBmFvp3nvIDp7csCUZL
PXjNHRLzAd84IEJeF1w9G+Z9AC8T64K0zWLP7ax/pTzidZ6SUi+g1jiAtF66DmiWPBw5/8kczOUw
hZzqG0Z0MfUjmJT4VCMhZuYL4fj6yQR4Sn7ypnZ6Vr+z47wMlCD0V4EfT2CVlVSOyHzJgGvcd/v4
Py6NieZoKayN03XoGBpciZO2rDs9VFjseRhj6ZMDsbiBQyf4vmql7PNY+YSrMK60hSF0u2qQKSRa
zFcbKAiXYGGqWn9Dw/whpZ1bC88h2TaxHV40jDhSw9O79KXmHdheBs+fTyTpwTUBYRHUVPgJ5jpm
13nRo2pGbBuJVsvPdZj1Y8fkYBKWIc/OdScrsXjriJskRdSBrzqmxC8/0gZt1T/PDy3a8n4j6aLm
1b/iY8OrrTDlo64JMv0EUVQ80nDWDyaJFYV7ia9FnlcY3RZwUaIMxaJox+68QZtHXSYKEa3sevgB
3VdV8LvkHed36qDgcNKVY/ga/BysXFOJBvY8/UVCjy8VrhDcE+jfLqQITxFMCtZ+dff6kMMano6G
dZscfbSn1Tt1VRlSqLFtz4qoseGI5AIFh2fhaiQFBZMmrVw3bxx94uvVU8+bd6y7Wtu1zSK0Md7k
jI/qBijmBAm4axlopOAD4z8nGhXn6jARXdcwx/DrgMu07FlQEjsiIXhMc28ALmL3F16V7jojbzmB
Y3NUt+D5DVOvAkcGsIxlRB+VJaPL1iWx7wFT0DZkH6hUfWHp4Sp95PmEjezLHZSyQ1LgV/4Ejbwq
Sc0M56f1ij4B50jCY66jPPf+ae06+S66dxiiwyQ7b4jszXiFcubTOocGGkUQWo3+YqttGKhpV+TK
NpTr70JUwB1Wq+CoTslwsutcHjI2bGo2IH62w20Uf9zcK2zXR+ERCvt6+Bm0MubwSAHf5JGiDwdD
UYjDAY0IQafisDnZF3IwQXzG8t19pwfZMrwuiKPc+gLmvQfV6qPLrbMCS8IqpO7cLd3MD36Lko0z
xjS0Lo3+PHrcDXCNvvMxnTALLWRyC5G7pzWse4+XPd2rmxmJaGb/4wRh+nppnlVmeIGKpKo+R1Cp
5tUoCehlhRtS5j8IhLWSlyRAkk6jtMoyq/VKF5lrQejPOOi4BHQoXyGjx+agQDRkXUXDnGbk3oe6
5Vkg1GHzQqqVvK5uccZYpSMXte3DbnSzTrwhpwjKFSJjGPER2e7cIioVPCLkx2/8ZmK+mEafXjlT
knIem7e/pxXBwy0hyBzf/NX0MJvBqpKJFEQWkTMkRpBJpeJhrK4TTIdVpYfa5rLa+B36IQoRifGW
qDPQFYLjOpAzUbWeRHzZwfsJGGL4F3lvgxL0DvDN0HkfvmW+e3Attl0Dw+1t4V9ym77WiJP9FhX6
GLerL5q7dGO9Nwga2gzJcXN0nYKmaeKRGMxaExe0M8uB7KMc+n18cHfoMlkWOSRg5JTiYOZkoMAO
SXbSgmfAbM/DY8XngkY8iYNTymEKXZ66M/e/pBjZpeFJY/FS+D2KQHWunDQQySRKJlF6+cUJbBwy
XZXIW/QTRzQtuBOaZqWA8dv+IcWEMs00Z7MPyvBqPbyNpeqmOY6HQ5dqHpeWl5fAHyAI/y71RbD8
5T+z+lmP2YEwpWbPTOSKlW6WV78EukKBJqcDH/Y/VD4svFz4ZYhl01+p6BSol3MSdUCJviRK3f9j
67pdHmiHbGQ78kvBnOs/H+6hZh9ZmVbVz0ujHTojB6HVbWSe9Xb417iWU+Ukzo16ENGD6EUwarkJ
1EFJSQo9n3cgTWS0PCVVh1+YZFTAUaWtx1uLIaVZa0mDbBVFcUSx9/hqiBv9ZL86HTT63ttI3oiG
F6xs+in4ZXyzVS4aU4bN7fVZ301rGguCesEQsf8+D0LHFHrIYZejNMFu/4l2VkwHghX2Xzwef9qk
huWrJJaGXJSH3gucy3Vvbwqdq3yn6mta41EKK3HDol/uzpCd2YJ4fxltPUpMpgKoW9SV3lr2/gAD
nKfhyk4LbAjI3yfSTyh9DSxgUqUY1AMkneaBLZkc4poDuuxrvFXY/i/VoU+cgTRwmFtxZ27eriTi
45MkPEbstvdKCnTLzjkyYDvXN8hENxC720wcOSemFLug2lKeFPLPzI+biZjv+k+ap7ggoC1myKu0
VWqrVjz6rzX636Qmy/felwmAA8ScTrKZPy59YP9Kksxu2FTl9NeuMO6np/7zROIy5YethkJENxiY
QEzgjBKBb0SjGDStIo6iG2bMc7WtXENUbLIn5+06+IK4FJWZ/OkxsRC4wqAkqa6/0WM8UHmoEXlO
Ib/JNxPCnytrYE91LVT5EGNUpBZ53QJZQXVpSYm8Z3TgQz5mNAhTvRPRxBSrZpJ0yuB9bGPRh43a
Atn31Sj+mnRmq6SHPsJe5gUoHmGmlFdLnWix/hNjSCnsd6xQwuzqg38zszY47wT3PrvRccx+m8St
z17NFxrYV22W2LVg8LEXxyfw9A6CO+mm3MwXVAIM4ZW5Bj9sj2GSh6lVmsAnV03YG4447TaeynGs
vJTdKEHnqxqgf/niA1Wc0Cxp8mUQV3N6aIwSqKs3IngJxEFWqTkhiQtpDN+7RA2F56z5ncAk8rgo
Zxk3Fr8C4/zYZ0vEuyciABiVQlisAYavgGLDDOZhzOaPuVmAJpGzTFxszCRt7YNxi6+WpKP88P5Y
2ze0x/DJU2jpXmvuzQBoyhRfzOioBAaOoetgJGrGr95oHSJ1qxHjJU14RWllcPuHAwO0TkDSGa7L
9+qYfn0oRPJ1urrBGp0VtFm3DtRbSLp7e5ffJTKoCG1N5yPL3SjZETXc2lN6+qwIGGrtUvQDsZLb
ktqH9nc/BhgTIX65sMvMmHprfq8OKhb7R4wgVJ5BixsMqiUZlyZOIRMC8Qqsdwk4WX3+LOlOAxYI
6XHBrNMeY7GwGighUpdDLeQCPP+ZjqVOmStQKBMn5uM6EY4nnknuTZphzjtGphLXKD5jW+hO/ZPp
AhWfx7c6POO0e/d6t6eeYGzdbwWocFko/mE5pEeS+GiBnZTy5xzQwUrbSR+MsNup8bzJUqpEnY79
23vJqdEmRxYCqXrQb/fCKoHKACKnbHEBBzWhSrQ7ocB/DaL/nA/6VmrxidzRz1lcwBdud402HsCq
wKGRwDUDRzIeAhUD+dzh162mXqYN9/gTXsVWV0IGi/1WMGHbZdD01aC2U+x2rS2vf93Wy6fBmcnD
iAfZHRAuE+ThmdryrX/H6zp0VqJ9fBUCt3y8JmH++lrWWi5f350Ma4FM2IknGJzxEfa9ZSFIIbkG
IlP6kPgy4PZ4MGxmlxH0fyYxsVSUgpihmG2/TvcUBIXmqoECNZN/cdtZn7dvmlkJTnQyL2H/rMdR
bT0+frX7CqIl1+6CVg1G2Hl/H5jniT2F+0Kg4+sJQ6HmkeaZtO3TrpQbOWzLo3ph4tGamZkAeisL
ct8wD8fEBiDfhB4iqfx3JXKmDQYlRYac+Nm5XRKn0jGT8/CticBZTrV6fkPkagpGmtgAOm9wR7cr
TCsKZqAW724SnOxtHvVunnL1HOfUwTUqj+nNaRvnwnS2JAjseoCFaSDJGgZdouswrOvOjXVGmff5
wMDW9vJIxMscl1sxVQOG9m+2stcam7zuaB6YoO4TgyKUQeXbSsHI9xaSs3wE1dK9ur7UIjPWkZWn
ab/U8ffw3WDYEVHPiFQ4pr/kDPqDk24K8zCGhtk4Um22nHfAM/549zjmMoPE+fej2WLQISJRXElZ
P9nc9bhV9SndbuvYajPs4RBHx0tbpuQaglbtOHN462WdTBLBG6djopGKsiDHOLq9WmCzsU7l6zLB
9LZsxbJqyIPEoESOIPz7pqPq6R4YnL8Y3IDfgAHWxTZ0ek7D5EuttlJY5hQuzgl6nVYrlZvj1qG5
g9vYmjKAvy6J6tVRi2U/ldxz3KMbUBxoho+AvLlcSSwKJWD61iH6G8EzzkmFfuVg+4NItEUPyQ58
gDpwIBwCDd2bUdYWZVlIp/UTFrgogWpFX2UVal3O3dfX0wCHqrGKN/XfrUCbMsIhTWVPNJWb+46w
GZTiJA+hkDliO+YBPhpjHwPbiDBcfIZWeUXp+rizWp8aDR/60L6+CnV1ay3addiI4FhVSO09JuWO
tnJoUmWeSw8nZo1ikL0MMQcPWg521KXf7DTqL8vbe6AwLMdMk3Ga9hg59juK/7FOEkt5E0vMBxYn
LxCAjvnP7yI4xLaa4dfTW9zznK9T5MttN4OTpVBh5K/Cqhg47WhcADpq6+cJ86xLm4hXSZYuvN5i
U02CQCAdcjvg5u0py/SlxygFI3YS7KZ37DwOu8xGNwqNfDUY8iMEtkDeP+B1rqmBaeVWmAXw7NEB
dj4tlgX2UJ3VcBttrRCEdyia/hwB/ZOclKxoBaY78RZsPO4yhWsVJhP1uNKjlyIyf58UM/QvwWdy
MfUvv4lKOcwmE+S+jIuHLHQ7JNkTo6Q9p7oReG2+J6Onolk9YAgAoOk/X7uCr1UgfGg7nva4IRNs
7VpTHt9Ev2xcLqmWAW0r5nlwqlriBm0hjWvbmV8O6ZHHH122jxWryqMM7kTTpgt02CR/rnbSBKl3
ssN/I2SweWOGmLM0A1Bc2s6pgVY7V8/+HtiMk2bOZNXTrCVk9ijuswVJy8a1p4FaV5l+CWY0wuMT
/7YcIkWfAFa3WBlsjaeEj7nf/M5pVNlehm/R4N/h9qOWupdsH6PL+o8WYvsBJd2h5LCNm27vECfK
5v3OmqIK8Px5zpVqIUgUvfulyi0X4vvaOWSQVoMVTqJjBDgIZbmA2kTSESKTAGRPzDwV1wQRJWIG
4DDkxLffy95fRlUv+irwoD62CjE5mLgQjWeuEcqkTDz51siHMolVx9vPMyefWBwKx0+vgMmwhDeC
ATAAUBy1qI44QX2/VI8Xyw3jXvAQZXWBLoOfJoO/a5cfjpfvA1JuXAvyQeGLIRKifDTK0qE35Pkn
pLgqgS3FDc6njUNLNwdqJaNqfQyvMZO6sGhzVX292DPI5QhWaIJFJTOJVOt1dK3TyE/qr42OLC8c
oAvCGvnTIuh/qxYetuKCXx6SYttTZrW0uBrdINL1ve4JS8c4TMp81YuYjJocha3SW7lEQeL9Jy/Y
PUqTPpOfhCoiwctGcFE/laSzrHluCqm5EMCNjwdmtJiM90MDa102YwEVg4qO7NGCSUUD2Taya3bC
etVWGbnkVvqFDw6I2FI2tBnpEqAnhgahDuVsHmnFgewYoS2zwICS4fT3wpOfJ8QoXUNL7Af8K5nr
Ri065zEdfa53VqRZudUUvy5HPWCUgi075d9okTjvnREP7BwnCKTrHgKa+5/QWWZkEL3JqMWAqa/D
kVbF6e+DWq8Iu3Q49ROsFv84SLg9eAkl5gk6GHAKwKo9WrglyL+lziWv4+0LmM1SyTaX0tCCZ0hH
DHR+k8jlbiYJbciaSNjJYBf9bD3rEX51N1fwLqrmVup5cSauiPwB4j+1z99dFm710ML8Jbm++SMs
SXVooa5RXsSruZ/FsD88UnIvG3UO0cTulsmSA0hnI1nCdLaOBsD6/n5JvKxRXE53mdzTmA6C9AdG
qEfjVSJO5Vn1gtLitte7pfHbWqUMUq4hFE2MgFQnstrwSB9UjIN0fGb3e4IEYFzbtxnwVE5+bM/p
CiAfYR4uV8/z7Myx1t+3myJzQs9eUvRZdSv1hAbW0YY63gv4nJ0htAOKdQblEhGmRUUnIEDHSHB3
FjmeC83ZgJhzgmbeXBuGOMNsWV2yP5OAYBLPaP/h+rcHgKMAN4CfahRsgS/dw0r5n53926gTQ72W
YcsVEbIW6u1CI7rbC1AnUwuDG/Fn7nFkUle07PzbnD7ByHqbEUIcOQgfNVDL752uVNwbt2Lpyefa
XK8huG46L0PXfy0t+O7GdFp/JFjSKD4wLkM1/TYM/dy8w1+f1M4fyPIUNeq49KYkmJy33RjnsaGn
RN4V0kBqUtEFIlfG+BMrLptkZXbod4/PKo6JyQdKedzJkZW+HctAcO0O+/9M3dRxOoPkyy6uxKxP
OgEMCBQZD/hJwp40y6fYjjvYMCgguw6PtbpivhIYzhj71u2OJ6Tn8VoC2vN9zuowokvIdHmxCiB9
LbmCrGGuK/jDMfvc+SvcQ+QqDBNTQ1F9oH6eDLlHtmTq3n7QfWCnmvWsnGiPTqSiJ+yIz2Hvzk6q
DPCMidavVIB3oRZeLcdHm5I+Du6lYQdit9phW+m/44z4L3zgsfECevjRzOvaByaMhZZ2e301vJ54
fSpdb03+uoacgQGK5PqKR63qSnj9jCUsY7uRD7MFVTVFhg7jtqG9cAnXIBncVZSCx7odBSF0ZCxq
23oRWXL27eb5OLYoYoV/DMSPJ8iswJGy+Mw1BqWL9DEi84kVErIynKjdwBEjYjMbR3nlPaI5Ogzk
bUAgmEzD/Gj4wSMVHMi8a1ZK6VuG7+qmH9jHTbn59rPWQamREo/n3SxNpFbP5odJF2HqGZVfz2v6
PQfYz+fPvUXbuyilVWOVPkj/saUCFUznPOxOg5XQMpBB/WI1pZk/aZzs4kGncFocDD+LDQfrxUOC
Ny+pgyW0A728MkWjDl4yFXk+qYb6TIHN3TcfLty1AR+wuAa8zVxUCaSdHEyJzBObJrcHPNjROvcg
BY69C7a2MCS4sxzk0SSDBKL4ABrj/uUXjJdv9dprdn+S0+WoOO0b7pd2++IeKyg8Jcv5QrQX7zDJ
tKC5q7oxmcN7yqX2LR7EvRCu8qFS5vuXWUVerdxLbSHZqSSBbevgP3qlUiZBnEooYUUYMSndLNmt
ndqKPrbJip9igxmZJMEixDNNOAA6m5ZYfNQwRTKnNbHz/YVSmCSD05MLMt4LK2T+iTJRAfJYikYN
QgqYS7YebmxPNg/skO5xdTAbO1AFj+Qxftcz3tIlxt12DwLdp9SSbRNRvvodzaFEIzQ+YmqdYkOw
EIecSPHEMN+bGqLLVAosuMuPP7b+IAAdEfm0jJcYMZDTzL1sNIoaQc8YwW7V/DC1QNn2DdH+ooz3
kgk7y7QImnFqc0+sBOuEC2WRsk2HG7rxUmyhU0LWx8jPrZsfdVdURIRRW4t6iLm+/bw342m2Kca9
rZ229jDcnkI66RhEePY/9hGdovY6PzZU3+6VeHVLp+J2gkZ6DXM5xju2w3JGJ0unXWCekDLzbaql
f6Bk3Gs3lKnGWxZRQLc3w4ifmmo3ZZ6HAGt+gGWRa461D92KoPLBq3t09kWjwwrRSEKsqg7SU8mP
5NhZCT2FZpSRhcUzJhzLSy1WzzoQ7oZh8KUsbvdrbT1Sd2hIVJG0wkEUDkXCWfDp2wnIhn/AObRX
JEH1dWfqQq6iRX5Ib4iU+nZr3OXcTGIdE93ldXLMx/RBVZqliWDCZ1bV3hXakIPvMuSDrPpugEGn
hhfidDrU/0jWGBzoO0k4WU/tP4PNBIbKim31NlsRCsc8EIp9kGZfyKweGCQNKPG5qG9x9nMVuRUM
9zX3/Ykf123D6OAbMnkUZ/GHtwEWmDBEcOv1FjVZ13Tc1TzO1bmklJUMqnWpmquldREzW7sVKuOP
ctQcTyE93e+gDcafXO0dyaGHRRRcQqe7hmT4fQi8xzHanN5pD20ZOjeSB1qVM3xljEn5t0OJm02x
BOkuJxdxR/gZFYdlhR5ZA+pKIZpZwbym3Bu1OJ5ZaBiUm8Jts0EkfOg6jwVw212cpO5YKioXhAtn
Y/LQw/13cPbwL3fWaDzDpEvbcvd6J9FHHyYj+vb/SQTtKTE/WDmmYq3eCr+V25wYGU4an34GSToN
dtUcwWK9MmmxlqYYVrumGk3xZNENG2cMEh5z6oBkCCMTWIhNMP2LRhT4I9unnsJp/2LU6+Oy1wF8
WhzgDSF0gy0K6cOs1n66dUd1OH9JLSVpoK0Q4UxM+87eGCuDl+xvBJuxViKlBD9sWEk+qN0SubkE
YkrXVDVSbl3oQH2BWBYIBppYUoV6pyzQ21G8UgqKSBePzlX1UYcjOfPL2EENNJxJ0PasDIYrtycu
GEwLPcFCngK7xjjiLz9Mbr9xWPDfMEIS3kK1ze6kBm1c50UrzLWGF/gYSF6zZjrRYXWcggCDfCWK
I7BxsqNBThWdjuF729BOmhQGWdhSk5AJLfEmJFsYLHnT9U/mpRbHmaDaNoZdAeCS2M29OJWjleDV
C+4+3T2WsP7c2UPGX+0mC8nub1LC9EIQ4fDCnCAArUczaaJIEome1bG0OdE5gDKv7ez8ygObT0Mc
Y2ctei7gRkJFpGiLPey6UAbi82ZET0//brtxUr/dR7jK37IoeGeWORgwdqecPU05vlfAFZ2V5VjQ
5gWQhwsq4sRPLBfcbChmqHtdZycTobk3NS18cHt9v5haEKdY+eEtGUuHTQgo5AcAoNUHKl2D7cHR
oLAZixpP50kFsK+6Qk9jkPYMEje5IlGdiICYhVRNhdGA1Tb3yOjox2wv664CU2Z1igUebF7K3hjh
ujMheltZm6i7Mg4Q6jJFlC47cZ6CEYN9aQzOKMEbo938bMWj69DWNCEx7hAnlCumVtMdku2HG8nt
MkBBt9r3/JCkGzpwsLfyZxI0WKfU0US/iPmcdSwsoqIdBHKk7Em14+7dNT9MGhqh/kvr4p8U/yz6
EQrbfIBw5/+CZkDXHqJcfmhXlgoyA6ShUhR0qlH5/fCgt6jIrfX7+3KnFu9Y7pqLZX55wA1x/IwH
Wlez2AjPID2xNtoD0yyiTtIWSMYpwZYcaGLACavssOn+w/A2ilX6l5boRHD0Vj9MdeETtpJyGkhd
QfsIrizFLoJwIXGcZzwEZW+KfF1r1RCpkb1uPjixltMPLoFgSgertdlJiLkGVytaRK7EjzaYWm4U
TCAtqKdVRjffPDvWO7Tp/+YTm/uITovzH314wr/35fhOKpuT5KTbcoaeaXGvQAR5RzYk4CbDyLJk
DpO/cUD9AEoiEL+ap6bFokhunRqWG34GAFKcWl+t7DF3lmr0bWkb16zALnMwJS+YmJujoCfL35/q
W7/CrUeig6vNkfBYQddmxTpkijVHnonciMXvkrBH58vxmFAsn9IQ6QEfWnl00yddciVKnU9rBzUA
fLWwUu6bjiLU7q5kjNcbJX5LadhoUC5rR7dr2Ekj3yeHrRsedfGKyMm6WfPA5KpBDUrFVMXrbHBm
Y6s5FULbQoa+gYgzIrtoBIlgsO9o+pPlUIKrfU3eYFUF0VbUJiJGUrDi22xZyBoX0Svy5dW9LeQy
kNviuT1fqQkiVtABYlMBhCGvYn/vVXKG7E/CdSgDxHn+LsYi+FiK+zxE4VH0EtI5fM00rknz07bh
5yxho1OG/RSdIla5/SnAPoYMjc9maCDC+4fRLOruAQptcG9kHI8BEZb8hVpa7Fw68BEQVQhXYSsu
hGKKudNHqG19D6zV1NT0lTwMYgYkjp1iZM7DpIffk0WBH7W8JrTlBBjXreaWvm/d6MmTiOeZ5eVr
0GwonzvxksoFrg/0pum4Lvo/rBoS+3m3dweIC7sEUoJ64wVZ35QmP6xbPa3QBluITWhWQYEhnROF
7OYybk36UAEKC5Fu4cWtQSxHcxejCFIgirUZLSNqgV91K3Nh+hKuv2SvppgArdeaUD3M8sBDOEQi
IWv5C1sFGuGnDZ1Cx/pjcvVQ6oLOjsolRN1qoVTShwqNw8fPuYCQnYuo31TYruSrUvPqM8MYNpn6
GN5ZveHX37QtwLHgD33SJYmEES4orDEv6ZhttZpt3hFOlsqhmeugBd89bVwUZbRBECvtpfcCPIi+
yoZd13rheU3fAeVS2ICC8kqCfTtoheCuOUfl6iNjZ52xzROtajM0hbF0ZG1+4O7L41XH0qPNOqYj
QMAiZobkAPBAje7S8aVfmrQM7A2U0brzuFmCit0YwuZ60PvIAfy6h5fYxdA55s7ETdX+LVc1B2Vc
aTNGUC8nLuxWN8cDE5K9YcYrat2BcsnMgWVOUhHx5TGnOIhoFRJcjaW/x8xPM+F+Oy6eRTnLf1kJ
Ymnt0SoedE32xJli+HbYV+Gmx+icH1xRlXnDCrhbNrDrjoerBF1HbfXTF2Vlao+79btHPTzCw1rP
1BhyMQpCNgYQPC593Xfwm8/19DdzGJ/iDVrAZL0RXvl1KiXnzduV+Tke0H/sXsfZ5Klo7DkYugGT
GSmcuhuikY+JwB9HqYYvbKeA7IA4QatnuUXwOpY9eYIrFUa733OYE6s7xwIysiogemxkwKQlaUWF
R+cFUtoJ0+AJkKyHQXgE7gxB4qbVo1syNldKGc3wYdh3Sy3/zkYsIK+llEvwkvfK8Sv2auN74IEd
eeginwur5vQN9vSg94ZOA05LLCosL9sfKmu04KJ4zDan6ZTccZsQDA6vi4lhE+WBbX0AMmVyeltE
slGTLVN86m2bjwfobiPc63/RINyxScsm3+jOgh2IZ7UpFtJt6Pk66GSJ4f1NK5lN8UvMZLWz0+DF
zQTcMpE3Gqwg+KppL2x6WIjg89V3aC8Voq/wNGEnUji7ZlC/sNQWQOhYew+0rgDLUyAy66Th/jcc
XlfwDkGyMeaesp0mtd8jvMTuAizNX20id5dOeAbobvad88tERw/Njh8PLpv2hLZKuZSDomTdhULx
NT96mAb4m5jONTWq50bnqrPmuwJhCTYmC7TKrY28tZRUSv/uYE+lMvEBLpCfEjRxf7ZH0/X55hW+
G8lhY7DnyTEDTSo4uoUGgHFJ2QVeF2evKuT80nx0t3WJcmr3A16jZUZl57inObHseElQHsgtmHWq
DZ/vS26eTT8yBHrjvkA9rJoBT74CrvURXTGu1kf0xhbL7wa1w4jSSL5MOtF7dVDGTWNSSsKIF0eF
IfH4/q9aYokCqGjcJDLxrnXRCohMBMGd0ItKS5v1Zuvo4M10sHoSE28Fz68Tx97fHwoqDV5xTEIg
y+S+qdFPC+aaAwkPCPtu5Yo5phETDZTbrKqhiIRrB8xP8ufcFSuBXMjv1O0oCZA0kgyVBGUAfFVt
Nast92LDn9h0Qdumsb/Vzoks18sxa+Nq91yVohp7Ac1M0RSzQJ6spe5Yg8g29glb8WWWKseOlUin
l2z0QV4iKuxTMjPxYbifxT8se6gNM+vlg8Li9rYvTomG1Bymadr3a6eWOqJ3LgBBKKQAoEGdRxjs
gdlpP8WQxLGB+5JVFrA8geiMhrQRZS69UBrvP+XGbnvuspRnaJhz1ukIOXHI40kJti4Br1ngGg+0
qpe3NurNAOb3CTcsA+071GPAVLPkeN5dxuDRVyC3TUKXHObKd/05cc55sHN2wYYH5RETCpG/VA1U
y9mcUrXoV7gqdaHS4rdNRuCH3FhyGk+ecjZhVyFFa4wcQs3n6zsg+yIxzvnpixzjfxJRoUkrBaHW
cei3e/sasSUmuMg31uxcjSUvIj/8PyRD6A5ezTa8B5FzSo0189dSNrKWS4PZL21N3tW8n9tYtR6x
k6MGyvYrXl+HpelmYJwFh97UOdyU+CUcd4mc8hGleBjQyPnvv3+21sIS97qxuz/tftvh5mUQFf+w
jZDVoikP1OmrDyoNcKmgRugRvCowwM9VoZe4QSfG4noDxAfrkXBSCnTIKzPXeMQH0iOTCT0DuLTJ
ISH6LRsh2w2QLzOlqWJSFjwg2N2uX3WZCA/BwriqoG3zcVZNG0QxOmnsKaaCTbZA7Yx9XmZHB3Od
ZgJxqyh+C3mcDq4hsYeJJU+cNbf9TWWEmA6n44coYbYebqPN9ebFKWOj1o1oJGFbq2u+bONJRtwR
hjkwzmGvbOa+nmc8atguBku6z+2dkMTmEeIvMnczuTbaDv/NtY5lV/NxT/5G0JAvi70RYUj+J4p5
AW8V2Dm1A8aT9pJtTIXHlEj6beQXQuv/PpDERNgPpw3scBAfkm5sSGN67K6L4FkqfJg87KgaSztD
l64hMM2MU+gcgvIkqkze+VZCQuAJ7+oseSJXPRihFFrjSgRj5nV7S4B0+h2GPK9NlRwKMnQUlMOq
9aliCZuyyqh9ycsEm6px/kAWLVcgeYp3yyWMQaJk1fNE1VMG/5g59DPWzxox2vPf+U2kudcOc1kf
/9G0fMhNxoKaCgqNp8UpxVhkkrNhjxkEWSgtQMLqnnWdkzPxO7eHq2nOnay2Oy3ffNhIURjF0WYZ
HLqeOfY661HUSqWP0/00knHxW3yBtPo4+7m/i6NZnAaSJR4apo1C4VEgbPM0d8Iz4WvKe5Vw50uF
rupFjsfjxzT74uw/vxnhwYZNyDGsNJjyhIYWQhPGMDHzHOh8eHWL6eJ3b74VbJT0I923e77NPP9i
HB8VTpUIaURjCV7cvI3Dfzt5iiWoE7U0nImRwZRUC9wvrLjfL1i9ilFGcusQ5U9rdlK8WpD0DEyU
pVGJb4MPBLoFaPo1D5FnI8T1T28pAT5qfBigwphW6RZ0hdD5i9fUw6rpsGQwz85orl0ecwr0+8bh
rWr1FQpJL5AA1cjBhix+MeX3wvAkfpeuh6JHm9CbP3pJsptMpAMxcj3TN5s/Spg3ZSf0uHwTcS9x
D5Eq604FmNHkTgeD8PpQgkHG1Hb0yXEterrsYzJI/amTqSErVU1lTCRGsoy4KBvimeTFYQOrIq6Q
0IDHc8XlV728YnaReZhM4ZDvQEoh7EkV9zdzPrd2WCZG/i/lKpdqnFZy9iYXQMTowQIxE6Hrka+Z
fWRAGFSKrFZ7IRRA3B299zPbfkSJYB+Ox3/16Xo4c3fz4JlHZfZgcdlLmhfp11n0v67TrNe9FKHX
xhuTjxN2IDNNtWGpcoEQhz26jqcBBbdqwjD7KZMwi45NwSMUHFzHvoj30KSmR7hVtwcA3BIdq75x
W0auQF5/Jjd5ia6dAZF5WDivR3WHiQCPpt7MtzxfBzOhYsGpk763ti8dmWmmZjnRvc3hspp9ip81
2SiJutHFcY9VQq8sEa5opZVEY6/XsbMamj2B6rrn8YiWVa1Vm++KqxT9adfS7UsdqyibdhG91YBU
HhVKTrpTfS7/3GLTQRW34lJkAuDQkMwwszIlz9TG931C7v6dU2/4RGTviVRz9BJJgjRaP08GoW+Y
rJ3kiz4AWZxm/vs3mFZYLD93ghXZGMuWyzp6gPBO4DwQ1VqT5Pl73R3bEDbHMGS3DzJFpmwhKeKH
GzbY+CmoHxUvXGmvk4Pp7p60BOCwm1KKBjZz5G/dAja6Izn7+dVwbldyiAggvJ2MU6P7FubClnuq
CpisajoomXzpoWVJ/5TxZ8+tbF1ah9CCLnoFbGwAyWKdqhJL9VvpySFuasRyAyaJDmhXNUT0x9Y3
lVUvkdaOGAdslw9nMwVXHIwvZAytN8HP8UscI9JAsWeY8sim0LEH1ToSjX+NM26T1lNGA52BJF3i
LlviYpFPYmUz+aye++ExT7LCI8Pcq8Yzu28OwtC/cSJ+M+VS+a7DbX/OiVqD3dnxrtSaCA9FFhaL
6NnQlrnYakW40VCtKQaa8O+01PE84KUksZsTSczO9CI3fOnPjiOlqabgVmiuuGfVDjNTvpLWmpOu
QNwf00WLrfDqRjoxFs05Xtl1dAIw/tgZpiLo4n92qzomKdbxKP9P5UKPFodrrM/DId4jwjbOygP3
5KAUYJEN3IOP1+oYs7kQHy+JMWX/HXJKWJTtH6FcwP5MAtM8xfnWjJDeGyKHOtWCD/LFOYJEWN8O
jHtv5mZqVby3odd9ra/7qFwOCUsgShCq4Uy4JB7hCyLCNqMs1L+TR6RVj2gmjH+8LMxsA3iOuLeH
NoCYDC6KA9Co6tpAkxg+nuwl1ZKpncKzxoG0/q5IPitg0fFNkcT91u/vYVQHW7enQYHR4FL/b88m
9Eop0200nLbF/Y77Lru4W09/oYN/FJD3mS+oBccNGlg4xAwEp9jAUdfnEjzsUVV59Sfi8DoPDsZh
TmOMyhBZO95nNMRg1We8RrcujJmpxGNBJVqwJW8OGgyvfsTpqma9UFHfCcNJS+PFu4Vqnn4NZFj7
SwsnD8rpunUX4oSsvUT30zoxl7222KN+EuX/jL2940HjSX6NUUDsrZZ37YK/bx9CtUH3wb8/2Xso
tPL9pKawGlxJW4gfhqGd96Wb7A9fz3+BM5BpB2LbTH84eCm2Sc+V1W8KaqJToRB4Wh4f/5iPNA6v
GNhLhyvRXoJ/ShVU+o4kve0GMjZ6HhohogWn6g3lxOwXapq7oQkslhJGSAgyCsKtrwvk1ajBnTxD
s+BuxULyMhPVYzhrhbqsx8uILV155b/l5PrJLL6OW0Xn5arUUQQsZCY638qDReufjUI7pwP+0UWN
qglxHfYIHoVY4A+VJdbQyWDZZhh8M2fIf0Sybn1KlHhhC8BFesxs1XCSPgQpm8hQzXNqhg074Bry
ar9KdC1ukNa6XdNLb15k0sF9zqfZAa/47gqlqBaNj1C8jcq4w7AjRpyI5lXjzhWHDxm5DYDuBY7+
pjkBMF1duIqzzj2rvjZnWtGz2ilugdy+wf2bi/3qOU1JRyrUJaEl/QtjIcsbu+yiyWUZQqzN9InT
oGdGcr+gjtwyZXmq+EYQXmo/GNV6R3PKDA71iZ0PhD7DMYeeG7cJZVXZpRdSJpWIqnoOHSpdZZL4
8/lTbZZNTDW98rjw1WPaIMQYyzufHhKne4YZCu/3GXhpi7myQswJyX4Tn3kFQfXBXzWmOf4esf5E
eLmPcc7fAdkw3dMICYbgwHcO2gErqxJj+7SIqGgx3cIhNF5vn8krRBx5beKLVqpi7HCti9PJJ3rb
FrRMD0LMBwnSKpJPemoesDSa61SKFBaDy4bsFGkfr69y2HN0o+X/Lw7xJX0+uSV50Ly2pcsJ1PlX
ImSqqd7uv41A+H/rvvvCHhPk7q7PK2g5stxMKoQ6Od0SQjhJ5yvL8Vl18cXdN7hzM+Za06I0L7bu
fx5AH5A6txF8zUEVrgQDFAmXcE11dHjhpqckx3WbQtt+sNaEz6a8RXkpbQO3ODJQWCflkNzB2I1j
9bVScYbMN3UAcxj5Y3rdD4esOgHOrNXSNwhIapvZWv0xeYMJyyzlk9CZZciAsqQnU3Fhz8nbxcJg
HCDWghGuytqdVuOj1H8xRxbK/Ks09kTtl1nGmih9aywBbinGpqBvQcYof57T3B/3lgTsK90bUxKm
LMq2LN3Tpv4FzQl3Pgl0Uo3IYCA9HEhTB2/umqsrGi0eYy9V+NhhpUV48ilBx5RRcwpYzGRNR09X
hoaMJxyz1ZK7JHo1k3/uha2rXeKKdJuEMLW5G1ngNZBNT7dBF77JkCtZ4Is+JoW+U8FfWa9JaktR
bTAIwjRMH8+cmHTA7ODCS1Vf67DcDLeulCCPcneD3vrt/k9f8EtTXaWTAASO/c2+JUrtXLtI9JcD
1fg8+K6Pmt31yg8lIvAn9eN6fsBr3Br1nN/9gZ3bHWzPwSMjemb5+XVeY0vONU22o/iK2n0h5yQL
xqLcsO6UhrCbxs6DFVeFNNWX0jUKNPTGAbJoa03t/98H6sXIPpbprT0Hz2Qhp3cm7twFu6z3zJLS
eGcwyxAWhVIcdsYTvl/OHDnDLGe+9zliV3kfBGPz9CPSyXlCqVmRjLw+PAfOZ6N+GIixRpOZQzx1
nWcpztEvORwc2Eh1fpNx2IRRykOYTUzUkJm63RRssyvgGBPN8edQHzsOHNTcBUsoEMjNmqnQhgz5
mpxroXJAgJZT56b9S8t4ric+xU+kOuPL4PPXJKXg14LVMrh63QY6KRBU0qYL4DRi7NsZM0BGEq3P
P38+UCOtuQKDV0SGVunAdD9QL31afDxupdKNnVHBgSWgoWjQrlh8YTb8dIkM1UMBjGjev4R+jh7B
tGWYadT/IHKhXyWH1fhlsNlckClfiHSZSTTpkTzhW/szGr+GkdeDBN3QQ+czhM5vvH7AUAjCr6Vv
EMvJJh4DZZ19+0TDf/HURETAkTRPB/Qf4XOUPk6j4oE36EbhaC74rduM3Qfro9EnQOJYjXjGGdJa
PPJYqiD4ugt+HkXIblHx0RJifpj893ZYt8AgSTNnV4bAPhX/4zO4O66XUee0kceZ8TI9aF6WGn/6
X1b/knjlwsv4wdD2514n9pukNEPfbxf87VSjb9p/qNAJ5f4sl7Xi78e6UZquIv9sBm2C/5wpNLdF
SCuIOH4eapk/cyIHcIWfc5fpMtNtifgAhkG7NdExBoBO+yCPoSMg9wh88ZF0A+NdsiBVQ0sXRumq
UlRT4Ozie0s4OS6uKYYnXJPuxcCJQEy7QNl6BaUbzFr6QdnBEvQw5bPSHbNTQdNlHVzH85fsb3lH
J+rXKY3Tkf916d2BhiT0fTdC5dwQTLCWFS/s69RhTkd/XlUiS8iwql8aDsxF0lPW5pWIwKbv+4yM
L6Sza9GFAW1MdsOjZWaI2L9OnSMZpdn2aWRj2JHVSo8v7gQRX6+gJyeDzPGnFMlrp2OPYWobtep0
gzpjgeU/nVkJ/G1PuA2Z5M3ntL/Y9TR3pHchxx0hgCEsVNLKn2VZ/omUFwCaZVNhmaWUjBYn7VOa
ivLjLZLTEh4avXcxAcbkh9Ev0X+kj1Uv9EPb2yxuOSktRFKyI/0iKqbHnSM1JUw+JZxq3eqmXnDY
Zvo/PcyenSjKuCXP5oVzBDdS67t9zFcpLH4kmxcUsnApgWJQpMNnfC3L3azYGYVNT7c5LzxGeZg4
az6jHB9UDWBwb9ZKvoyOteJxaXSB6JF1aHTGN7eO+Tyf1YLnazjEr+S//arbLFDMg4i1G9dfYHz/
qEcDCmk3QS7KwOK0gbk8O3R75SDTyGD0WTWvmIUT/+x6rLmpmpVRC2BXYd/vBLwewlavFZMqmfdy
T5gQAaW4R0FH91bDvXshO2qe0pbJvXjpz+ym7Wlx7CR6f2R9bKcgh8+6QoR11V8lq6qq4ARlJtBz
vOdhhTosMqwo01eKOWEt4rjf05pKpGd84wuJBYniIGzNcurHqVPxn0OhSFJ5PyoUNBZYjCJfWyDE
A1q2wXgGh7+XCAt6YpSR5PvAraArhF1lMcGHUMfkUajC2S95gYr0Iyk3Db8gjNE0VcVi4ImQ8ISs
jXJmLhF/dUcPiE660NhMRJ7aJgMw5j4plyVpRAU11kzsRoFIKxQN8LLw4tU5BMU6oA+70yO3jW5a
rLFPh/QFRu4fA8WV+7RL3xIoQjUcI0Aco67TFK3hGI+qKpG8g3zl7xYaee9CGDeKAqyZzWpUeR7h
VQgl6FOfBPXGAcOqIcxXwTTrnuBBayzKr6YZpoQ/t/l+EzDxtnrgoXy9+aX8LWAk+x+FZEYgdHO+
43cpOcAHXbbgxCHPfR9U92JHzWiRK/Vkn9H9n0LaYj3lBZbGYhIBCk744XiPhv9i8GgtpS0agC0s
u1i8pGltEoVPMXrvk0+ivt7b+NN4wY0Ui6gxxD+Uyb1FbZhIMpT0yYuJeBpVeHsYY0OBzxOK0x6y
P6ZrlLoKthat21y58MNAD3h6+E69PfnJJK90b6FeTteDRG+t2KPKjI1X7a/sZgDlb+SfqmGbZOr5
FOek3XWEmyIxfl3h9r+V96fYOIWEX/xGFYERSlHltcVTuAAWRjyDYI84IgZ+bJ0YKPT8bMqW0bFs
XNDIwtp7KqdX5J74y00nS+HbV8v1Clwh8LkkRLbt7xK2RAC5HCKpgYoTVKyUsfqQcIdcRsKe6E2R
TobacwQwntRyDrHj5q6pkBUIXtwKrJf0X7tODOnz5+9qrRUwmy8cWWUANgcsdAZ1jZGoc3G3KwqZ
pajjbX/OmME9ho+6Qjb/6LTUk2zfOeY6F5a3S0vwFhYxeq7yI7mUe3jZhjtb4W1KN2Hhpn1OfWSP
jDaVBa0eC+pbU7J7hT/YmluxzIuzJRNEYOaUqQ7HraatD4I5YTKgRj7L6wce2E14ADwkb1I3TwXQ
9NRQto9LGnRydgAKtfwfI1NXIzA+a4ADNp+1ROP9lRPQ/EMeEM7VZbLMg2uU06onWzE0T4sW/oqu
BaF2rhZGZ/aVK7vkdQ4hIb99ll58UNxERLC0yvKUE5/Vqk4uSrOSxMNTymp0lE1PiFUNi4VSuuy/
sZRVSh0KrLvsBk39tPjLI3IfeNgwu1Y1JXxUorJDq/uwWdIoSG4NfLNL/SvpF4N5CQjhZZgXA02M
glH6s8x+G3Z+XKC49dMOn/H+H0+DO/HcPPwBtdVL51cV+v8Zt/kN7im9F8+RqHFGKh0zEdhlWUFe
+nO/FcX1/VGx5wOlh/ipzmupVKCxbl0I7a59eOehP70ikiRrWfnQZlX0iuanpLDj2BEEFLVenOM4
q8rkq19sCFxDx6pJWkQPzgme/I+wYQKhKs7tQ7njCf0SScDtGnAmslxfZfpCRoqlHWGblWQE1r6e
gCcA0a7U67ArxXs6NrQejoVxagZP7VxmT+85p1n7vVJfRydCXSxwVouydvmUhPWdohiu+kkSIJHa
3M9L6VVcM6hzgIdhAJuiMm1eNHbcw0G0CL+C927a8GX8W1Znqx5BqtOmULVxCQA1o7AP1kImAEDZ
OELZ6KXrLP58B8Qb4LK8qIRBFayjDIc33kHh6Llp1/b2EXHLoQU5jvWdHaPVuAUYq9cuZrYOolZo
Ws72T6d9EmIJbHXA9c9uwQ5YUV4Yi65Nky8/rPtdSoE3y7cIW/zbyu5m4WF5Pdnqo9lYYGpi8un5
ILTq7ANK5sDLHs+csBNdb2ELMxDRZP8up347fEdQ69YnuHADf9TCZ9uxfpvOHGANGhEm+J+K3Ptq
F+zkOUnR/lR/3PQQsgC/xn111Fz/eojRq+OIzHxBV5zObqbujK40nC2UaeR5rSg27RTiMpf3o+sa
x56YuoTCe2AsyAKRgyX57gzFigEHWV8zSXr+Ms5mEGtIwdL00uWt7JozzKj7tCmD1glN7qfNQnSl
zZDHQ6fFgwgGgVXNclfwOFs6CDAKUruYLgAdenm6CiLNlztKgLeU7WoKN1N3OMqxBK9VQSmr49d9
fsTXDqQs6pty1i5noy4M+T5Bu9DJczxd0tnjSislqZASLryqfeDjAOz96OgOUpx9N/2kdJxyBc1H
Fu3zxxPvqpFk5v/AfoztG/Ar4AEz1YvRz0qdv2eOl27lzQWqsoPaFXEwQak/Vl9V9AxyCPVkKztl
HmMrfiY+LlKZl3/m2Jc+o0mK1LUOflN122g69rlYmkrrFUjTQ/j/6Xwgd9Bf4Gt8eN9H4NEpJ07w
0R4V6eiSuA+vMdMAwu9Swn/QwitEtAMHAgvaIafxv/6Ta5+ChVJTzjV53f2qKCf/7Ge+tchTifd8
O//F1vxSfDQx38gePJmaqtZvHuJ0j7PnMV6hCafFmc2WjdV12Zws/UAjcZ6HKCP9HXnnle9M3DZ+
72vLZCPJJeFLv5reUy6qJkbEWPjtoek6KsJ4KIOr573u6tV+6Bq2HajIhdAlqipERxoEp0gkizqZ
9TLBdv3/DWnD2DhLgYCFsS/ho1G8EwZZ1WJtchcPC7+GecXz9uRcVDoNunbkhdIOWlAQDY1Ly4CN
Ts8AlNCXdxbZKxMjGkxUCmH6YaCK71mce9dvo5Lh2KBQF2UhRXJnkdJn5iFe2QNN0jc65zBH/rqt
RLAUn5No6TKzDxTR6oTD5iTmjbl7uZ5cYjkI513ld+2d4BHqH3+bJWzx7HN29XPkuG6R3SK3W2k8
fU/9LRae0CGy7d5QNrQ0CZLuSlC5jWxLJZ1avfJ1FFDQ8RebPbx2md4NoyIjdwBIeCG872mU1YuS
cOQfgeozNDUb+3oAjLawYk41o7IkoLsaoG/15ZIoyEpoMiIPYLt4mSWkp1cfzUDfBs0cEEmVf4vb
AIS8XrkHHEBdzJM3OCMw78pPq64FcTNrvrtLEmqHVHRpZHuGDAt/sA9sqeGoYo7CeQK/YqeravRB
B1WZ+ABT5eue2JOoo3GyRFQpnR8rd+lPNcvVpG2xegebyt2itX8sh40crD8+J+VkFFBEz2dY8P1/
aRpcQxbtiWfT3ar++dBFw+uH3s4+Vo9IovaMv8WiZY1qohENYOXrn7qWkf1XbMzRs2wQlJXjuOD2
p4X01F2rqnCSbYj4+c1ayiWFE2saM0L+Jn+zgfH2QVMeW9834T/0tr/ev18AXbhKxHMcTfmIiNy5
aqbM+uISsUHq9gjooQk2n/NBgk0Xc6EXjH89s+T4Arv4sXwZ/ki/wAmo6TVmlVkO8Jocufm1ohOb
sDmHfRVyWI3vBiWZ7e6Pz999uwTZkAtQltOjSvUE5gqntYL3/Y4uPct9wzxN0ncqtBaEVHem91L9
Odq/N9JiMsnuQ/b1Pmk4Jbqp+Hgk8UEfQFcoMLF9g+shnbxVZqmLTXJrEXx4poLov0Mz6b9pGejB
Jz5l1Gx0g1jSrFlAZ2gDSODbYu3yusNS0IriT6An0KDFWAkPQ7cu5F+jGl1se0SZdfuB4n+4hGdI
Dnxk7hr5klbGbLE9o64VrjX50kB6nzt7aqK34lIy4ePCFoZlS+dF/EqHQwitW9xMzKM+zuv/ILwE
4h+VnDltkxPe7jiv7rh7egu97TjOtf32Pttpu/CednA+WrB0IYw48xk3GCFaLhu6QB1E8SPEuC8r
F9MQiNWj2ADOHMHNMqjFf33nnCfm73xL+T7PlvqoAv7yY8tgDCyqTTuLObLSa6xq/Cev49el0eJu
auf8LvZ/CNp+D0ixgXTwfmGa0pBlWbjQE7Wr/ikh80EUo/+EqfSapM895OGX/CF8rGIKhKD/SdN7
1n6WARB6xvpT2HQs5Q6HUwmTVe9ayWLzP8H0zpuM+28rCGdfG2J84+4E5SRbYb+dCauBdcGv/dFP
HsCkH8EDqC18XdljusFnIyMKDK+zJDR4o2d+i6MX8I7WJhCK4vKpsoDRBpcmVXromzPi5E2tZ9G3
F+ydLRQml+idseBP0Oanb3Por6HlFedGS0F/43ev+ywUqhe/xsRf6RDwWVKoP1Ni2gqg6eqbS+ui
tBCszg9/G3JSChCAJDbuX/LO2kq6KqLq1LL3KNGhWn52T489SNpghEMYSyRIzSwBdrZDQFKsNyz1
NO4r88z1q7+wTtcb30Il+upuV3pD6wI5CIbF0hT9roJmmybpqMDErkXzn+FoxpSWTgHiInIwTjX3
WpsdWwIzAFNZO3qKBsuxJVcYTaGa73E13CLQ0aJ1kUhsFjwxT/cfAAIvtkD4sF1YQZqgXEYMR2pF
ntttSEkWC84rzw/RSIwS10ebWixbGcSOxeZBFSDyluSsCNZ6wkjILzSbMIe5r4LyiiZeT+zQ/GJw
NvlNJ+ioFaJug2yV+FmMgQ2+GBWOAGszZS1WSbyllecRkaL9VzSQS727PEO48gQ3zXimtqqFUnco
rgNDLM3MlBWxJt0wEi7UYG4N7Ns1FPmxOQ+fEefEMP3PdgsIUOSWKkNVTugAJ86E66rn/lbVMdPk
ezCn5Klu8BuhhAHYHxdy4P1dLgMgyO3oY6yD3UR0Ut9h07Qt3gOHXTQQeB/0C6ls3rzxPVItfvaO
ocWwXIh7I3BNnmVL7NGxhw4nifM/uhK1KURCsMs2TvY+zz+SVQpnnW3Wj8qglo4E+kCOWF9gwUwW
TYHTzGkiuLUYFury0hxAXn+4OQXWzLuABktKntWSm6AvuKw4cbZjuHLvuhSAu9pLE4dKqhZj5ISh
yemyL7J/udEH8hXGNGV9b5GEQbaPXSFmdGstS1hs6FZaDVRG8jq8Gziim7s1HvfhYP8UmemmNYPO
ELO0WQAm3+cFHCdQuGIHqTMQsgcdG0mPKbnyMxPVnC+NjRD4/o/Ujk5KKv+hbGxpru+lao5lNDJO
7+dfeQigO6bAePu7EN6vQIn54CDDfPA7zlOtlC+umO8ur9A95GPZSEIuql3ysR+OxHz58KmFe6dn
9lSsCayoE85W6dRHDZImtKKzFkXdyY2sUzzCaak+XypQ5PCIj/maG9MKvcr/DssWQ6M0Miags61+
qQeIdib158vsdwNO5ziMHEPo3DD9eX/lVtSKg78iER2VadrZTCnSpqL0XCDu7VS5icwyqtoK8tUG
HvqyXdW80ER86IwemsQhx0IKeewVYutFBMEg8kXwx670Jrk6LSIHHicbogg5crGOJr62OXe0wm1I
/GLgu+Ker0W9uM7EplJ4G5SSX+KxPRbRrArmU5+jMS1xb15BGHQl39QjaGO9aNR6JPIcUmjLe84k
6Q9nigTcH2tc7w7E97u0Y9f53XZ7OuxWIIb3Ird6WbYClh4abBzSFQPnPKUleHGaR4y2bxLNYipm
Yu/sqwytZgwQpl+1A1rs9oJ98T5u6pI5u0g/+UYK9kNIVSza/J3bOhL0uDbNvFrJMskfKCT4gpRl
+yfmjMs4UYo4pSkecJBCPyzSQqxSpIiB6Y8ElW58T5T668DTI8ZUOKenqnLealuRjQUnsHp28gAg
o4zb3IW1m0IpXAi21VYSDzi0E+av5/dxZb0bpXaVKhB0qSOxPgXxAgLXffazcBk3mfZbZ3jE+mGx
ZrUPNY//gaz0wEYu1T5xFrKSrtqCzdBoDPvT3AEixErw25YYDKEmflVm25WnY4emTnCsPEONaOpl
V5JOpY+ZB/0tKf7G/tNaVi8ngbNrbisvGHd6t93f81lY2AD2PMfdVOkS7+bybGxs+klx8iu6SZ0X
FHp10pQF4l8Ry/G/+dOJVM9Ni/vz1vxGwmnwwMuK2fqvDgZr8U9fOoB/7rGaTn5sk68w7FExw9r+
p0DH840+oW7Oh0KbZfUbieTDSwR8aKoOH+cYtr7dKCf0BG5DONcVTccZFuVyBzbyL0p2Avh2b+LC
BRNmEB2SQiQsJy/oe2cz/wbkb9e251zBWINeCbktgNneDIYlKepxzWuN6wUAwSyQ9wvTnnxVS+ow
Qh2pNuWIWAEwJIFwTE1Zl3iXFf6SxgIiNKEtY9mhJkqOJehM1eSL1J0eH5KQtwtCmRQIXaLrHRyJ
nle9ivSOGP0zNMC1JOY5YZQM/6VD8WZlsb47SEIVklYlIoGbqm3UdHhhknFIHmWlj11JYKXB8fFl
/p5/0KFekoWZ0R7Do712nMMcNmo9r+U2Apz5qrr0mxeSTuJ5WrGKgHpgXuJgm6nNjvj4ccyygKFi
Xwk9gZLtugPHgVFAaNU9CuJdwkutHV4jpHbllULHagUGAmSPOAuKE93X9ooZCH58dMjyXYF0QLz2
goTDb3PYVCZtN+1WXUOZJDUjvtfBxXxWxqtRZvh0s1tdJLFerDnkNhWsjm5N6j+WdCOaw/cvuNNe
lsy71AGAPcM0EOpC2sM5JxrehsGB5mFTs4M7BCfsNM1tGew9p6CiKXvyK2Ng97wyyfXZ+k0cGu9N
aQnLN3+PjLRpOozTOfcFIZ4ZX38+ymQOGp5abip6jpeZ2awk4nW753gTif1vLi9vrxjzn/idSMHA
Vetf1BvSHEgpM1SaoYewwV80H/CwbOSrFr9D7dZX5gUc2snB6rtPzJw9DMw5zKCBvMX6W9tELass
Zu912O3tMQae2J6dBv2/VEHTWBuaB6+5L/Omgyb0cP+dq3XjePcdFWsUbIReIuQA7y0D2i08ZgiC
9yqWBTRCNp7rB2jA+0Jrf3zZrDQD9a9oV1+Kp2/Y9jzKi2YuwBQz7NitxeyJ4G0G6ucJN4UjzqPm
Mg84kGFKBdaua1TGW9PhKl8lZLmruFoHMZ/6w2s6Db7xcaQkzKNX6wQXS1+ZoGxa2M3PqYuBhuWS
CsxBrplJQfqOGyesxEEoMX/MBrXZrj+LKeR7cmLFxENO5bm2Qqt200k18KpAjz7p3QbMJDPOlaPi
d9Z6WTWAOoxnR2JNe9WfOTzaX5/FZghQgnJ4BtGRv49YALURFAGaqf10IsMx6nBEZObhrwZ3aTT/
KZ590VG30wcZQXh3xJAw7aFT1PmhzAoAWDs19g/U7llwKmwdh+CxbH459uyjJn42aL2juSHrf2pn
LW3hpcS2r7h/v6CrLcWeavv7tmqKGc209kH7iWXWWAasOkiOk8hOqZC7+4+q2p4xxBMi6eY8rfv8
+fW6DbutAnHuWKyX9NJlLzXE+f4n20ERsJYt1JwNY4UUb2aGDFbTtizj0weKlMN9yKjvtJHxxyjv
qC4M3O4avyKTzcAfZrpuQxQ1XAcxi+ji3VgPThCtOrYPC/K7J/CZ6VIKNLfNGym4/vcQCFKjWJSW
8RLxr1qpGrb8Sp4tsP6U9UfTtCpBSTNA4gm6cnTByRBu4MLLHG/QCYfIuGl5IxOZsYPXwnxA+Wrb
cvuEbHDKWkcEGhjFnmbRl3TaTF6VBAK3BEWH2wW6aD/6cKsaMegmObfkC34mHKw/WWUHjxatILBJ
80bpllajxVqeajzTlAyuuswOUA9Y8D0JCyNvp88a0Wf+ZOPvkqkCiG5ac/VWVsALeyBib4QL9TXz
2x/jbbH2wp497U421onwhxYEX81hAHNXYCsbJCX6Ybnmqt49Ddy94XWVuEFM8LimTelSrmd1kUZo
PNWtU5xC76JOlhr3jHKdX5QfAAZaH+39DNKVVV8K5kAXEzv7InU3n6DkurP4/xsuIEkNi7hGkCJT
ZQJfeVWP6JItkAWVu6jUFPGiYouU2wyRrGxXF7o/+QpbEpdo0FYRrlGKpJByPl3roib+4WUpV1hg
zxb8sm5HqM745YDhSIDP/o8S4vRmAZGeRzIyxgBTdzlpZWoIJi9SkHM9Dj8z3pjuipXkRbSUS7Vq
TeMLnvsf6t1E7hI+Gonzhnpja5y3x0nrfBzM1xXr8O80qn4wEOEc5uEqJUUsbRrlnqsLTqMQXR8q
W0IKEthJEniuvkHJj1vP0PGKAtBBcE6jYg5TM26mnAhXNChmZFc4OPysmmlfXE2/FvHz9iLGTdQI
dNyO6LqsawDPdiCUyqkhXMuVdfnyf7uQ/P24gt3nW/9u7+paHiG4cUS67wvvsfywio9CQLCkGGDx
4kQBNcEFSZG28VrJhwVWhMv10l4y7c8CqRcgSpcGDork30a+LxxUZSZ5y9iuE2H8w7Vabbt1y25X
rMNJVxlWya9K91mMB5tVBGwrCwuMNfeMDvaYsEzFG76Xt5zaQxAmkLtkur+BAmt4pt68rEQY5isf
slEzYMemfKOzqOiNx3VKA9fB98qWWuDMIePw9vqAmMkEf5iN8rPx1CvGJTZC2HwMxqt9mBg48bkH
NK3FUV01E0556I+cyIsAoj7s6HMGWB4NfUouRJj2bIU9Y95x/U2viHk0do6wSdFzxQ9BuMpuld43
tIAyTQyTRdmytd0UVyiTnigjUiaHrMG2HmILmmchSfwIRjdXgbLrJSzlpMHRpDzr+P22ey2qCxYq
fiVPu7dwtVn37ruz4Z4G8jbyv0kWLW25Sdif2F/SEXVS0qVHyoSEYf8a7Wngug37hp5cIjKVM0qt
bb97JgTAcyxREdV54h8ipU2LKxPjpPUYVcih4mMRojjNkCU9SCLk9H+lFGIWws2TIug9R6IZIjVN
YA3JH94T1CrIC09JrI525R7T7OwALC1h/WUWPc9YZI9PZfOwFjlAJfSNlMTBCIXuEeyR/6F36zWf
IYjNAuGwhrgN+ggcHdV/JT27xpm+3lJYkRj5fPSnZjR78U+befbhbo32jGzswUTHVhaTH+Enn9JY
7ynfvuc3aOMGpUBfWJF04m9/E+lxSdE7Tn7NADpw4Jxiwwx5Q+7Ofnc//Uva9e98GRGdfLl6GhWB
Ayly+UlJfJntQQp/5vY+8stQkEbrfVSnEeYG85lDguQNld+gbZo4SFDpww0wX7/paeTPO5CB1uBm
glDhOAyMbjw4VacefIc9/F028TjQ3H8eahm10AVvvMWU3I3JYdWvHgPfRx5BGTgwz28IK8o/abBF
Z9mnD/ZRTaj9gtDjGcGbTjNrLN6gqgh0R3awIwCTVQxkjYWANb0eV2d/E1fkrOEG75W3a0CmpbnM
po69dwjI/W2roKa7mO6px9bF527ykyqB0lc1HJN0Rm9/66jF8E1eohUi0ritMbaGuVHW+32uCYjk
sq33VpG6lvdwxgJ0vDAr0NfHzqiVfBAcT9DJR4Z9PIQnSeHPVurK1RwJfUGpxALYcWn71giXGCoD
WWPiBouQDbckxOyNcwiz4fKTcapmocRuX5lja50ZRSZLXU6hBI5nEpJ+yWod+qmTF1To0o/50l8n
T4z5ausyIuk1giIe4DlWcsxL3Li0GeAuFl6Ajv9lVq/ZfeVhkgf1rmJX+GgDLr8tHum3MGOlW46F
QYOVHvbBa39ifbtnGmzihS6EhKxV8LObyhCg6j4fSfBnu2IccMZQ3H+dFFdbJHfHoF3Q2AR0nCo9
SmjlgugnHWTLGaJJIXgfzRG2gxyZTLV8vryTCf/LkKbKgx5MJneLpjFzAB0T7x7Rg1Fo7HgqiuyO
/kxfzINXmPHO0/I/y9u72PW3oDK+vpJ+dnd9P3S+3zW/XzgDrsInZDlHzVkh/FXuhyUTgNY9AxH6
7TiWeMbJcb++fu8gaGWRFyN5aSr2LM/Vk/oqcJQY027MbPNyu1p9lUbv+K6XDH2wSbdg7iDN+ZvW
nHQVe3wXcH2Bn0Pcs2D3CylCMwWrxtUEX1Gz3+vu4xz+lKCxhNoV0wwFNER0y50Z/wt/PKcc7qB9
kndwCNyWkGvsMBBHg/LMmCYW6C53a/0O/Slf0maiz+ZKazb727w2iwUK/inQ17ieMeHBm9sIE5XW
TcVD3KRL+O7CMM3zRMmb0mMzx3WooLe+F235xgmlSKGn8oZe8s9IVATziarvEu+zYFpl82oxvJT9
AReLg76zfQQRBy4AXS703Sb736gnIO+Od4sDA/ys17oh60rPUclLmpkYDldazdDdeq6IPTanR9TY
ggIyRgFhO3s/0yeNqLmTP9TOepau0yHxpV8eMFrEjlB27YwBEH+fWz8pYs9MX9O3ujklwS3SvT+u
ZCHgZwGgdqTSFsRNTUJCutZvlEyCZ3I6hZP/auIbXvyEH/fFJT4WlKrPqRqAZuthbnaXeUMi0bMP
4O+S0BBKfTmjuheVMKqH4xaMi6fJuXglqvIw5kJ/a0Wn4oy2bFGHheZy1pmujbGea4gjfqWJi8lb
8gNESGhgFBDQK/P3kZ1s0IJGuTQA1zStkPcjMdkTYBpitWDDmw+RgMkDoWucTy8kPVHk4bLy1f2A
pn7Zu1oMk1Vu5qhYwXxOxORvHDnb3tn1RjwXuDQA3mFz1ScsA0L4jCx3G4+EG4U+eOqLC249Y5xn
uKnGE391ovzm0cgmzMTbf4YeNhtJa1caGnfvH0PQAGE2ZkPgnDHIZnjkMzmtavT9kE8wou3TICJf
dwcTKdBh6trMaHbC67nmymtQfxlFpy4H8aFMKwJ+dsrBYQRhxqpCeRPJmatRn50qCRbWor7TGOvB
tnhZtZHLViygXX9ko/E7F16ID/dLyIfqdZoq2KVQ8yX/6Vxatft1n+9XDQa3NgzbnJwT+2Iy1GrB
tqDQKsiJbeK4aNOJFPW7Bsuk1gUSD2hoigYke0m1AtqrvbJFMwWLprtjSyXGzXbnbQ1VcRHmxT3o
14TvZ42VekYpJB9vWaczgjI9VXvzOvjN/yIxK957YBw5G2h12dOuCwio9pf6aKjWrQnu4EIcnoki
mT346HUMZphnlrARyVHQvhoCNpyR5DiWwspOj/UzxcjRw3PMIDOHM9KnPBIKev3YMr09GcyXXNnR
6WvCvwSI7fMGs64inIgILLmaB0HGH4zCZ++sTYTArZyU+CiceDY4YzhyrFNjI84cqmlC+tlUuTBI
JtVfr40BBuUfu8/8JIpILkF+gUWdUyj59W5dupFW7FuAonm7HmEEacAIUZddnHYTQaza5y2+EQ+g
E3wrlj9BCghaPT+4LzM783oquU0FtmkB9ayiNa0EaEDQVuznhtnJcmiev6jLSAAwcybLemU3Qupu
1prJvcZnvH+Vq3ukRxcfvmer2JynWNJsanNrzV7BIRyzyLw/7ddR51Rwvi40aLYC7O3LjBFiK8k0
EQRA40H6C/VOAOb4EIHgDoLBXZOvoQV3U/dF8uGwjcXMrbjbqMT8ug3y16+id8GpQJX5W/wRejcu
bbt2vxuflfueN1KzU0ICQh5ISjE1oVGEykwhyJ8/C2832iLS1SLvhnFHLn2AcCYK+lBkhzLyxZ2H
mTUFBfrMryaJSTMZMSjpURTTa7AIr5WUo8c+su+edbC+QTRKG9jNknOz+HT//17Hqh/+W6+DvDB4
tsjXwVlHQGzRY9H3R+xstjaqk0bu51T8YSqHCzZc7b5Pr6fk9ryHgCAMSAqFrHjfqq9gUDmxiRIM
qxuE1jPfpNQ6FAFGkRIS6ZUnRXdBYKvmvlHohW2z6zDhOuEgAwOsAwpayXZUcfq3/kiS40iaNiS8
Zz28SljzMupciImeDhwSgSzGhaWdPpwi4NcyoRjjhGLAa7wQheKuYe/liGF1x4hk0MZHZpzRSmJ+
4dbWF1ICHjadrpYFfcbvvVjet74x8PUn/irMNQR4z0prWvA3KXmpov15+/R9CP1ktrfXHlJhBVfh
npvmYUjGtHs3KsapjsA5HYFsYPPBqp6KGZA0yOLsDJeFdz6QDt349l0I5jJ2kusSAUsnV44Hf96m
fl8RNC3EBjA68HYuWH0/vLH09GgpXx20BgEnDbjHTpeZEMnN/uQ5MSgym6E95LogweByu/rSGVLt
R2pi96S9W3Nz2e10xy/N1DXIBmUMYq6h40VG+8dZz31jWpxxk7hApGdTHmb6TFmpAb7nCEzgVNkA
jXvGy/YikFyjbE48YKXk1rQynYDv+LGY71Yyw1imoEfy5piGwGyF/eHX0ECEQk0lXyhFxS1XSzNg
M3z1hfbmBeBpMfHBr/CeT1bvOYxu/LFpUvDEsWodPMDjRdziALERaiZawxAnmduNPPwDcxh8m5Rc
0z8fzL6e8/1j/aIZrWtm7ibaBqZ5OF0ioCR4PURJK/6AVTUSaKtM1xL4D3+FOsq+ws5llEb0kyxR
cEjkuRSTpRvAmPOIBLrGXoNORpiyfcmP8NIP7mnCkpDknSacVsS0AOPHd+NjPmaqpm93PPevvRwU
yCUBLdJts3s6c4ePMOb9/j/szFeh3/iS1fjg+2WqyLww+ygMpnPKGOL5+1T3OwUvvPJUz3cRNSET
UIMUHHI/azgZDmf9icYXJMvV99JskLmSU8nLQfotkJbZ0Ci6DAJGQYO/VwiiF5UKYIR9z/Z40oWp
ASH0yaMdREssYc+8qHJZJmGjqZEFBxvhIbSM2FYa7RSNy3XLzEFgzdj79exXSYFTZOgcSoBSuMJy
pa1GrmRdlstbCsKhFBNihFBN7R2IpNp0MyiQlW3NBqXMwASp31ZlSbPVTsCf/mKpKAno4WfvP4q9
5hauW0eocFGih0vdt7tTbA4ECCyqR0G+jf+FD8VdLejTJaN4sgw56FAoTWjZa/bsIj9PeQEituGw
s6/2X9up5xb/QMLAnqr9h1QA4V9wI2DjvLGaEV5S9lOUsedisXZniTNiDrHl7qSZ6e0cH5YHLBkV
1waVl6bOApWICadfwLGyMSIgj4ybU+oQKNsTXpCxQagMrWj/UiXrLYfsz88om9oBI0B1+CI8ewVJ
0TGAHPVrSwdnwEkJ31o+3HzaXQsMEI8dMIDb7WVlphd3tx7WwcLEhaXwXS+oiHDvizlWFjbOBnj8
HUqFwgYt38iOtuxa8L2kbbHoht1gDmzAfLVhmX6Bz4oK82avGnqFvNx/enX1pgRQwJMUrMkVZrZD
1r0qyewZHcWO8UmKgtWS+2zL3Dn/jY9Z+XvEE2d71MJ/rbCSVEuGtp/gxASRdveS88tIaOXTKKlj
BYlXi/gGMxHMaKIuqNsPmnZspTPpEFJADRQ478I2SnHVwpZO7W3o2fca2Eq0p4YvVT/jCpWTv7FG
c+HwK8ElAhzeZFo8TMbQK8v0ggoajrJzrFHo4QSott5+DK9XpC8VasJvwPq4hH0Ag61bqgA+kyck
rkttJEZ2gOvEaUgr8s+gEGGTGgo/WIB3opwCHPwx+a22fQKBFDuagR58RJL7V14V1NuBI1v2ViZ4
6jV+ypGNFKaLYEwIj9TUwQMaHMFodVvuaEqdEcy5wGbQan32KUPBCjqeLxvKg3oDwxI1q3+XrdYa
ucICvkVLqJdnaDi65cNXnMFuaiE9VPL1hd+bLydC3XgMFpSiSG4I/e37cQdYBv51cH9X6z09Q1/J
hSQHe+ztt176MydH118n9eEDlXkXMME1ASjJ7PhpFWBsZRFhlGzYwIGpPgtm50QxxXqW82SQM8AB
KFlfs1Ij724rnseKU66HXZtL0XEdlKY7onJ5gPt1wcKewDaxsTgxsr4a2e2AYmNZX4SlqSjOkdDZ
7L19fMBp3is8zbqF0Ssgv7O2cwffkxeL5xhnz8HyXGhhKlxBZsOIX3Su0uEWDpYRkAxgI/O2wvpX
fwN01TRV84CS8yc9hcyqWzPA3teHNqRh3xMtmfw6C3Fzv3318NPDM96+rLehMK0R2zBMRjcC5EDj
PfNd+tEgrne169PkYIUIqirgMDvnk31zAsi528GPecfmG94hUXGECvDV0jUblYWr8a4Bq3kT4tZ1
gX2bpnOmsyw5fu5vaYCiEbv0UAgqt+wyO5p1CqS7Q4lnsbBrgIS6FALFypV2hQXqcXE763l81fHC
oNHAEpSM0h/6ur50VOWaRh8reIRi4YTJBuEaSzfkDZg3NeUxtQWw8eOXoqW2B+rdM2rC5J5/ZXXp
+o2G6Dyx8SypKjxLacpwV4itVPzY/1LAs1/iAYUJupYc8w/strZe53foJRa+nHGuGMt+65BW7F5l
oWluX0kQjz322E6E/+J+QqSYpWe84V0DWi6bX5E/z2LbnKxNkSi2E7WXXN9FebqLRFGAzV7eDRbq
gCkgF9BYNNRwPTMzLiizrQNmrXHtjWQ/jp4Yf9PnnN1N65Yb3YLqdlLkPtcr8dKq9s2HQ9fq8YjT
pf0+VZrly5Cw32m7ED4RoV/dHgmhi9dX4f1T4Mr6TL97L/tz+HW3PRXTto206U7uZYA0Uvrkd7Ph
mA0KeZf3hrq/W7pychZGjHBL3mEkc44wLj5Yf0Gz86Om2NsfW0d7jHOtaC5YrxoUc4PyoXvHWPt8
Lg1HO9rxKWSbJf0QbuwSvzkyVh7tbqcB8JRB8S9nXQgWU2AoSg/uW6z1/gZk5+bszrbTuurMb5hW
TtleoNbFhW/ujgiw8/8lbJh8yxgbNAhmZrox7kcJSocf6WL5mEqAplMQXN4F1pDbNNw1gGeFa5q0
Rjt5wrbF74qJejIlPaMZPQHspIwWAOLuI2hoAKbZd0DMHG7Li42oNHVwjAv9keciEt9FWySpK425
b6XQlqTSWFO56r26ST5WDRkjDrFljOaoQw4YzBJ8XSpuhAK2Io7Jp9UcdFhB52WMl9BNQQs5ucuu
N96d/cjLPXPJbDwH3Q6rJFM6PPVsl0OSUZPdAyalmKZLmR7OMuPursxed5dkvGrJhM+uaKzUYhwt
rgNJWGfM6m7lu/EibkeJAvaEKZXpo15ly/9/0vUrAfee3e1mi1QlccuJgCKSDke+ACl8HHDK3Cdj
I6KTaY0xtnU11RmHPX9UofoAD7/0IOyI/MStx5xAxetT8EP4IxBdcbtk4/AmUwLJP8z1tuCPrDD4
JMX7Vu/E+pZ9510dNlyEZELo9+VxP64aiwY64eogHXREapR3i0OhJxPhb2k/zZ4153NM7Vh7kejI
qN4wFzS0u8t8kuRe4SXjd4NCZlJ/it4kdbAQ9KUYfdwptsIj7qx3xVlzWNPXB9UT548dnwYXov+V
/btPioIyMqUlG372feiuiNWGKUJIt3ZMifRoopOGSbisEjdSsH2/y5b2gP0eB9z3F4IhrWafDwQd
4kd/RGx9LjfA/2AtchxrCUWMk+mjfcWLQTs3ocoJQbrjwcPZw4fq3ymZl+/liLkbxodnrpzpy2LC
R2rrZvsOWxxA+xxpuLTapwl7LsyPnBvWrVC8caL8PtjBIr3grfPgNMp2sh1w4aCmZN642ZBIGDjD
vdIZSfkgfCs1LTYhsDS8/AwTSNwOUE87Q8iRt3IJWcTDFufenfk6/Rhhh726WlFz0suGp7APAjHr
Ucru8fCGy72iF/Uit1X6iAVCIdgbISQUTN6UPD7P8Wrzec0TAl7xghzKFhd8g+rsVOZsKtle3eFZ
umsAMKKYG1SwVlB9ITM0gsEiEdzfvlBkSpvI3tOi5LEntTmfTW5cCF0RMo/E4bV/Cytl0T5YX7iX
ssXcZQ0aRJYJrNMbWDV9gCBkPkc2RaaJ5a8iHYBLdHnrDolCuatABbpo5rm99/msxNneHMkFZdpe
OJD3+nJ+XuP062rLS2lc+F7CAyCccLNj5Mn3g9G1kueawYG8mYm2XXOhYETKZgxYas3gqYEC5OhW
3H/C1ovtQGbAcc+LhdsXUmXDMQ0o/GosromKOMLRHLtBt+S6I6y9eiulHkLfbYMYuMWB463HOZOv
SJgmI5EmWr1bCphS1wk+EKVLhz53f+Jc401TvlERlOxey8laOYG8UkvtKWeC/A7jkKxmiKScQMB4
1JgeWtWtJb3L9exT3g1v6WBUy5TLkNhhXm6EPFHniYQrh5k+sG3+Cmgz74HzPBlBcXmYqePu4NOI
HdJEHU1alfCi/QxVAOuWlF7LDzV19wnYkWqMlGMCeAqLc97Hscm3w0JOWn43ZRX6M+jOr7sUvSN5
dYmlJPKxFXjuUYKP+b59jYTZHIQ8+qn04JB+8SZ19+SRuLpIQ+W1VktPOOh/hK2TWOQzSRIEAAki
QKQmv1TB8gc66VBt221kmCA9qzsI5Dy4UES8OG8vtNQIU2FlFeIIZPhkTFxGrjug9pn0oR4PefMG
167QGfELt5uADh9unklJDppatbLS7UR9Zhsbv6n7LwIH8QQfw5HBTuy+KuJWJkLXE7san492K+Cl
3AS7ZhAXmV5K8OOgNPTXbDpTO8kMGzh6dh8WfjSztN6ErLeOAkuySeO7vnIFHE9y2E1AN17YSQJf
5u+cVv7hhMR7XB8+QYd8faEZhCvu2RbRI7bjWyb5D90dNTBeO5MTzo0KUrDKcVgJW86oMl/6ClTC
26SOQjJbTQPcOPOeNJEuMap4vEBZiAgxztAa82ZRlCYIQwR+lopiVUhfflbXTMqgUhw6ss/PxD5z
H68Pc76nPvQQhFyZbPqSRiIgW5OSGjncKOmbQXORFzSyYGATBxe1sI9LRG5YbLKJXObAQeAT0Obe
Z5SeUYmsNxcKVdXn+RnWXhGp3yZNkDEBcYJBBx5O1gNhqD9MY/ANKuUrhBhrPnkGTZptgdgp5vB7
kzlP4a/FscASg4CULV4VOZ7Zfa/SPUyIPal+YmOcyq3ss5ZhWMNLw+lGeY//387TalnQmwEOIOLl
yJd1qHAm/2cgVVi+tw7c3CpzTt3blfr7P6uTAJ2WU+AxCWUy4liunKU/V29PcXvvqqUlHUDXb+kV
V5PUku/5eQrfHppu7z5lvwbP/RY81W5ygwkkyYEErTg+Q1GuoIbtsvO6v/CGzS+/hXgmjtsm57uS
rYvW4HwHu2eFuahC+M0NcJ53rZsciAVlU6k/62iB4fFaYh56d1IeWDan2/WrH8yUFyFu3zXCOMuh
Sva3DIrnAN+6bZIFsUz6XsWnIyJ9k+D4CfYD1vxcY0pxYFeuNogykJZdpF9zb29jVeSamtgxsejg
U77/UHlCfzM4ABvYLWAdofwQkbsOmc0EqDCoJbX05hgQV0BMVQZ1GLAalsWIzSQ+l7zOFnFSI5Bl
pq7nvJWhDxYdPz8aFyIkup477Yy5BJBkPoVwSOGEu8TokoQe4D3uiz60B/itMg02hskeEflrxRw5
Hvrh8k9DWaRS8F48fDpJZDTIMFQw0P1TNeqL5KpainL9QREpYaVhgxJx2bK2tUm+w6IfOSA5h8/1
FCkgJGXvJx882bdDxJf3Nm0wv/09U16mFkbZ7jP8K4Jnz8Sep7NqL5Xvhr0Kei8sjOzxIBWnRZjk
tlMoTfat5FaPcEaoje2m15RLrO2stkjKqw6jE98fC0pCQruc1WkYLneEt4uuk4yp20dH73YsDUQr
znpHCL+4aFJmu5SWU9FGPtLtBE3ER5zijJweiXLM8ZBB/ZXf3zAvHx+IekZPcvVn+3N8hi+NvXEW
v9kek9hm57aGcDle4/fVds35xQTlimJUZc9Apgg2ll5bWsl3ZLdOo6Sp2+WVkxekpY8lXi+By392
fznRsiPNlTBqH8YrxJNJvV+Flb999KhEzHwgZTJUQVO8ziRz1Br9nR+WVgThFrlFTK3aIH1ZwZZQ
CnsU9h6LhBzvcGAE9oTOLgWkNAzi1pDhbtl/sH8vYCwwUB4mi7v14Q5/Dy26bCIS25VH68LHEIKC
4w662hD2gv9SJyuqzl8dMsC+se9xJml7HdjQrfUEkMcECz/8fJdEBjHC5xXdlWqngusIpQCx7ZZP
ZtUiPTlmQAky94/4ULgyh3aPFucOE0n2jg/OKr1/iGk5lefVEHQFIL5jqacT8FaE4zYQM0O/z39+
x6EitrNI0brEOvepENjNq1eA6SXo/kqbIrQqB/ZQMjBBtVvIPuL38OSTHvBokwKKF8Q2cxrn9mw3
oqLJ8EEXNkj9Cn1elsPEiZryoySf0m6i/PHehCuzTBDXH8ShwdFTzBoIz2Z+ttGoIaAu75JhYafJ
+QBqhK3yI1uJ4HAgvDwdFjePXYNiZLn6xUoNQitKOEcQ0zkWEf/buwk8F/pCCQGzYjaMqCBW5/2c
mM5xYuI9eQrivuNZuttX/3n5zmoXAAOMiKGLQNPtEWrWCjZMuM9kSpRDNtiM2RlrT+yLjUxqjI3Z
aaoN62GQiWhe5Xol+DT6+iuUfddes0SWip+LNf0ERvLUPz7wE73FFBYNNGCbr71LpswtwATW2SCg
r1tA3yTx/hVJ5aYborkxOaXEaZpR6Pkjbr9Pnxp5/VjGGsvSO+/3PzYWwVzzB6sQCDK+zyDN26jB
EepmDFiMRJTQABSw/Wys8j0E3WL3dMBTt/tppXXrGnME9pvAsy1SHTPx9VLCbyEt43EBjb9rCSTQ
wXbH8ym2g99WQAszu4YPe6VYw824nKX4ISfvEY5b099Kv4mYJ1JH0wFCCwel/iTY0Ao9Xb+xE6iL
ME8N9zD4SrfKpDkVxkQosglGsgHbO7gzTERCPtHEShlXocYnmL5q7qu4bik4ZnWWVCCud0hESTQZ
3KC0Iyxnp51vAVC2X1e27Qs0jwrR7MXas3v3+vaM3G+KwzzY4MzKfhWto/bAE6FrRVfX/wXq3bns
JeluaaoltBWSosvxTwQgexwbpLfAkV5wFpJtfIraSa3f5yFh95rSkrLYHdyvajctsnUmDkgRvrdj
ihXQZ4dtuug/eJkjhWwFcKUEZXgndhEvPeMaI6lQFzUYfVyuTbKecbQFL+3k/LeyWPntN7MLxdti
YabpdIvm71nIKpjRs+TnA+v41/yK89CELhMIxK4460LjtjJP72LsYhfoKzU+bSjM+1zqLAPTSxbG
NnkF7D84mF/CFDPN5CkZOXfHjqiTH7Z0jaBJsStdZpL7PapJvSD6gyRIGf/ATnGRXRXo8bA7FP06
gF+OK7OYXo12qb4zttzyK+7SK3r0ASffVb7u/je8+lQy7Li0niMG0WwPP4OC9MPcqqCQm4QeLzBE
I+apmmHxlMh1c2H2xgEX5/uPrTUhK82AX/9C/DX6hpQDge9dS0Ru/PhaIYEg7k3Zqy9dGyWqj8jq
Mj9/DkXdin0LDDHSn43e0U07LPHnHbCLU91TLNcrFiaa0vj7UfzzgfTJzWtNmTqqRJUsCz39Edmt
J55XVjxm3BuFymTPqPdyZM3oiVQ3nCvVKaTIIR2UF+zp5apxeU9EoWcHBmH7CKpWLTrS5meMQdJJ
mYSXpu5oxavDsc/k3Niyl/vdBG0u4VZKrS7GcZLcdXUNGtzoCHucOjw6kGF4oQTnJ8l+++j+DdtE
z1POTR/Iqvs9Zn0JtUTW34L/pkvHkTzytsemUrih9hS9NlcdrY2tXYwJ7S/JSg1wf7MHCS4FYcN4
Bbg9glcs4Bs2/4Zm6EydpFhlFeJ3Yc88JBcctbHnZiRLOnXZ5BJDyIiiz5Iq0DOoaeqe7j60YQtg
NzXY9C9zqMHZxVx1f7OD67fvy2mXRTMrhltGurEsar2XsEnJcjJKnrOdm7tmTKs+zthXDFnI1YJi
fhx6vrGhHazj/OdS1DXB9jye8gP4YxzjP4E/lr7wJVRopc9cdxYlLCn/khp41MHPh4uDdTS+XB/D
XLBTqYsIXf/hd8+HCmOH9oeV9V9Zx1B3q4RwN+nL3R0HdyrDtpL1HvrNLJUQxvCWl68n8zOkSObg
kh3UQre8apxn3NuxVsbZy7BK2z/T/J16WisI0EoUxrV6TDZSpIuMQR+AfmwFI1QEFrDyMX5lmNPI
qRdQCPRmXUOM4vuuq3Do1gzAlyVPfhz24KlLxTmvRy/TML/Nn5ADIeC1Hq5BvxpPoZF5QZdP1JiQ
HPAqZk8XZ0Bib1FucBtfNG25N1jemJckkVCW3KpQgJeyUUYCKt4ajHFlbA/DIuZLKvWvX0PRCEQQ
gR/FvjPU5j8CS9dGKtfpNpQ8oFnv/x0a4WPaVgNJdZ3L1OIwVRXSpIhyTrAimsWuPmwlkdQWKaOK
V5QgljVlpPhOwY+Gos67Mwlv1HTJNFeUToqGEYaUZTHIv2hTyPDVQhZ3NyKh0hGtWMy8NdX0jXip
Uo2GdeTtGK4tr03h5HSslQ6e3F9Ts5AvYN6PVh3PFbl2z6KSaKhvSj9frLxDLYJwM6By2HUnahif
5XZItPHCAMObjWVnBdl9VB005RgVQ9ZJ9IuA5DMRxROpNCuZUE0RvKK8LCFcoPwQ+izdNS6E+Py3
mPiIOYSWloYfWxtRpCmVSa1m2exy7QU+lvCwcEHpO60IY23v8S5Pt0gDtf9ZmD7rE0AT0mcP7mJh
L472WwJnZ/8ZSy7Zdv9+1FruZnpwEqI9o3RkdhOhtl38GQnEQB4WdQ+aDzauepBYiDEuTN7TBH2p
EXoSYxduyzhoTLo2GB77G+TZyTq1DaknerZftJuZCE51qwMEsPbCR+KIGWPBITOFKXOZ/+0EF+Ct
LXf2YDXwaSv9PFGc30Taliy1aSYa9yQQPfE6wS/MSrcyuE3g3XlMvbeRqfT6WO+gW9L7htKcvkmF
tG8rMq/SkcAHc58ccch2TMR+Sv8Gx6Ad7mCYlsqs7vc6zEM6BmJEfMcKiOXB7tq+pR1YaBGi0w8y
SHMULEMdEULbTNKQGZYyHYDLqhi6dupcxNm3AX6dzVcpXYxBhCzBmLVaBAGoj2b6wSkbJMzHBHbU
KU8noDhpbyKukK7CsJa6S5d521D3Vt2jogPcSsK7dUM7ziqAv4zqG6h0LP229ZiDy7Dk6MjfNz/d
fAuih128Kr1719PbmEu6hxjv0Dc1TLFEuMfj0j66gEEwUGvKlq/z3I+8PfOluPJwHcQlJXckBx56
iVfr5GW6sFnarw3XlS01B+FeaB+7oK2Jb2uM6oDxFxj3yGbvlOfIpCGH9hh0bNi687EsK0x/oRxZ
72JdnpX7rTBDD3vrxKxqi7LMTAJ+BWbT/s8Qj5tr6Y+fl6njrKnfXR5szNT0CxzNKoyv35vyzBPN
7v3icvOTMg9aw/Ko1uiu7Wfctt0S6mBTY8m1YneQCp+sif4UDjYUZs5k85Jwq+LQ+zEBpT67aFLU
1lI9YbewSfg+gKTA1hHJoTXv+CDRmFbOvjPZGqWi2YhzAHs3YTEVFC5c13jOhwNyNgl2OVJK0iCt
nxUYD3cmXVi91w2UuVqA12xka9dDLp9wVPjbWfUCKVtYSnoMZO1eTOL5tcvge1iuW6I7ZuzgsRe8
uFSX+H2udf4Sfj/4r5fllL6MhREL5orjsz0q9essCHjASjMYYR4AgOk1DzcSa4uta7NmUSOhjwuI
jdlHJfjucJUt+Fih51pVPRB2EYnRMjgpNIdJgEOSqTUWyUjGLQ8QWK7uzeN065zZjR+j/bPxTy6k
FipVPlQFHWCLZifG/gkFlMtgM+dpCG1J8xLAzsPU+l8jfw57IA0LApIg0bzzQHvxnZMyZ0NAmjBt
5rk5WrhaFK0Z5d1AyTL3Awsq1KzYU4N92DMWPtv3uoSbcQQ4ZnhzOXhriJKB7Sm5kN/c30OVj6ca
/y7wKYJo+euxSJpJDYxeJ3mKPnOlfhB62L8xgU36o+vORTsFIsC2XyQuMUh+rV+F0exSg3jkIY3K
Dfoxn1nL5YxlUfyN/GbLlkbBifPTE5LRg3EMQ2uCjl4V2UUB6pn6jhXA2jmwvR8x9qbc9FXCxawL
imooBGPkWC+905S58AcRlDsojp9gXazBVtzvIb5wzT/u2Z82VhkP03MamVPCwOco068SpEavNyM6
M4ofdG6YamBRoK7byjWSk00QMDmnH7m2UwerSmByILXdPbm8QJGUqW33UAvrRrsKkiFL0XQdJ7km
CqHJli2UbtfJj74w+YwfZ2+vg+V4wk6/QxR8SJlICmoCp4LgQMtopKK643cu8nvHyrk/kBl871e7
axdeespN2b7D7x/0jynhDQ+HcY/yqL+2AuBd5G+xOr9mj/FHUKyuldmf1AJAUW4I4FVGjXUcEILi
XCIC0OM7cQ8nIkS81nuunVTZWA3DB8U3ze5ebnYD+BliyyFsEw3TU6HpdVGE1V4WhrIvbMYUDK21
N31dEnjMSrC9Q1GF1D+wSqDXeleaBns0HSb7gaj0CxcnosJHaneHi9zU1l9r0c7y+EoL82eWyL6A
hL/C7kN4gL7jVAFjmyGeGMiqIDtpRHJizT0+6g5NVTakCa4T+sDq0GQNBE5ndVfkllO460BwcH/w
Dj4nDKjSGNT34RbuVesJU6Q1gzS9xczpKL3c9apqIwwGlstQFosHlOhKOOTwDBu0fjIK6BD73GGk
tL9cOSbUROel6/euG4QwdExBQB0U0EIDaCDCAhNZX1nwSS9aHNZngj0oplHkUPkmbWjFaDJm3AX1
WmFOqKlOM+aJN85LfjXpfP2bn9GnHqEY7AZCM/m2NO99H7ZU13n51Ss0Jle6dsq4epJrQJ73D1p6
3yKWMVjFi44+RLdBIBoGTiekvjEdR/AHfP3Lf6XZEBnuPbYmP6UTF0a+54UbGRpeuS1jlSxz57+o
pLj46d//yeaeRPMvVxSQLFbrRKpaJT3N+cocR1+LgO7Sw/IBLND/od2Ak7b6EGct10Slpai5qVhs
k6aenPvv3nSoZijf8UxC0+XI4IjbsPRRM37iROZ7IPMSEH7GWxQaDR+7Ut7pgL0NrAbbH1JRRIxq
5iB56eJOrco9xhWLss7FVHhLdVunk2d6bmzuA0NflLPLdieltEKvtDfJj/3a1gEXipfZlxTVItyB
U57vX23U6fGrYPb3jE22aU5aVv1v5ZGuLCYE7A0B+hqJdyD2hdcG2gDPGWqj8Xy/NPuqHP6JRiuL
1HW6AapxyegloeHQufHX3j0CL0dINyskCapdq2qt5yZdnb27r8vX4cP2Tez5neYsdttyWgOHoKrj
4KMU8eTV2sov8E5NrnAi1Pw84c+CDiT3t8xNAgoB1BaqIMLnnBcYfgLl0mF/OZcDpSRFcO9Cq5GK
yhoGbjRDhOfUagmjdKsVWUGwG+oeVZAQzeOWNleeElRfBaxoIMuhEEzitQG6xl7fKwSSxqVlyyQA
vbpKuRb7l5YD0GHOzM7XbSszWK9c01TCjDWFJiQvYwJC+JucU9Zs6ILDHIAQBiaRnMJ1PabJUt3s
cvw5lMoTdC0O9p+Mbrzp+RWHqgb3mypInjQjGibFWXXrF7ksdKy69dCW/pKtDDp6A9hFBcWAc2zz
QtfokaMiquXVtvH36axPVLBud/1ZVbyka0xEDu7TwY4Q3bH5/k4QYHt3KkAkG+Z1gr39/9eG3n0z
aAuAOInGuod7upOVqwYl4LUKPTrIN3oJC/+X0SsXi+BxghPVvev3YVvBvaB8LtiysrY1imdb8Riv
1DuA61OY/wItOPB2KayUAZ9EsBQEpqbhhqYoZjtFClog4wI51zZpCWUcSXsf5v/yOWk5cEujlzyg
qXnEp8DBZhJMbPKVI88hQH60G57K4TI+waQwU7yGeVwZWYHO9YusHO0bws3rOaDlbTwBdswbOu90
mSkdVsa8lIR9mXoE4m51XXE5K4x+CeDbdZ5orUq2Honm4IfWN/79VEfS4dNTYd0bY7vByhmvsgHT
7P3FaFA1FV4onN4p0HvffN/gcVwNKT7aZzO5kW+riRk+/hdwvtyth5Nry3GGNHMtFsDkf08Cf+Vy
waaNUtdfKWjhsxklDNJRW06uJOxPCBtplimzGmdoDHpFooPsxz8e1uG56Hpk4i8X6r7ypjvQm8/Q
Us0xfOjspL+wA807kPwuPd7qqob6FASTkXoM1jcvfWxbIFjyYd1SZyHVh1+clos5Lb/apyeQ4dJ3
0JfIlcjGbH8fEsDpfOC9SonQ8vfPKSkmBKXCYSG81kTgj8w78trxXdj2absQ/1n2mDz6QRkSUS17
hlZXFnnO5rYdF+dozdNwDZxz3DFdsbVqgtLPe5BY0HK991V4KIw5MZwXa+yv/qg0E0+zGfbvNZ74
pDw2dqdxRsrlqEmEtsEU3OZGJx9u08eh4kmXf4HKWuP2o6j0RymNx0ejCLmNyy71o2giuJqAKVU0
K+6l4Tomya7GK+1EoUHkrwQTjTa7/A3iabDT83iJYQPSQdNoPJ3nJCTsTchn2kCS/Lq9OhjjZHQm
eqAM4D4QW/yVZjMiNVimhdB+37UUtliWZtMjCVKw2HcwzFnIQbSBAucAqC3CZwpXvCJ+gFVfrJiC
MVrCElc/XPHylPh60EyjOxQrgWlKLstbvzHiIOivukbMv5p2Ttd/Q+iS6U4rx2UrD5X3A27RgSWH
A7tHaPBHHmC9gfSRgccQkyZCeNCv1gGFb2z3/TnFxtDV1oPxdZCKxmRaIGV5E4iuEgkHpHi53/an
mGaRi1B3rZca3suK1USOAcYw5vFaAQu6qT9vp+FDqDVzrr6BmOJchyO54X9JvLCjxmrtblM2KVER
NUF5B0t+WU6tn997hFzFKaQ5czsBgC/0sO52397sWkhzmicq9v2lA109CSz4AqIri/kDMWropY7K
+gU8IN2iyiBuyXc2IscbDA7364VWpgu5m5rPjvdnPuK2kNoaEe9RFOjAtM/99oKPFY1xTj1ZxNZ/
Hdb0a6WL6vBpPwpgwMkwlMFOvdR1sQKKXsE+hq8c4aPIdSdOXLzDFaZtfQd5WoImyLtsO48jxw+P
Ma6EemXIQAPeo5AhLsLgwnXkDPPUgi3Pf7M6SBLSd9KfV/EO2z5VfEgmieGQzglhM3dn6og13PE+
gyiK+lSO3VFTUXNizl9yalSzN88jIWNeiKIjFWTOMrnIlSA1rhTPKWLdZNNZ0cPPJCu8fWfIh1x0
CxityKjEq7XxBf5qZGCU48GkERupUJ5rZ/bEvJL4N7h0T0fv6rrq2W6YIWhwshvNBATpsTcrIcbg
KD9S2CjqscNwZ46MDo15sPMbP2rOcMArQu7wzwlkdqe1JxWEV1bugqPKTEYPhO2ATCZMdSXyD+nz
7yQJZQJMqNnhweN38EH0cUuEcFRETgnV4xoL3IFUPnAiLRh68XazvS27kbQAfnRJhQ20dEx1pABZ
gTdH18RANllzaBL3X23r6W1Z14+AzThQyzwBUOuJ0QHknoHSYsAHTkteX/NZ1eDfZCGb3/4VKYi/
zLJwKs7Wk75G/nVN8qGEY88MRLEAjiMpOxOW/5YZzWfSuA5oXcXYeyTwOGB6TPZgZqlnlAaw2tOr
jMhuDKiYq9OYyqa/D5n3vaprb3Q1p9mS0g0m+gOnDin5OuGlHgEMV3OEqdJSQ5I1TEcVUn/tyX6K
wjY50wHEoOfjiUjO9on+gUTYZQizZ4DR1FowEfQADgzGo3BoeR7McaN/G7x4iiQYYAeMpFwygoSr
PnOCJSBeOK32RKX+OBXwwNJ1o3GYnCahpWMnBmKkFsBwG+hnCPFpAi6mktQ7QGt59KKGowUMLEJ/
GbzBNUsSVnRB4oUTiD43G8LH6CDukVC0GJoqxC6dwVGiWa8CW/t+M/+DoMXV4mKx+RaILDDhHXbf
wlXeEeuc1HTDOsf8/G88VtsLdTQctywYNuU93i6s49eEt9ZHdGnuuHXLwznVps68wjCDjgvGoub/
KGxgFyPk2s/j8M6d3mLOW3hNierD8vf8ueoAVornM9L8sWVBF2bshJwJEMtf5CIMJgRR793srFH1
fd1DKI/TfOiZBeFwbqflXSgxgbVmLfBYt6ZwwlidaaFPTG8WhmfBo7X22iRRt7k6HnObfDC6Iwbt
BB6R40cqtU5GvrIjQuVE4AvrTI3M0d0Hr27gvvNtbMyhuF2xyEmRELtEWGutN77EG216SDiDxclP
oBhONf/jLfAIbDUkW8ksgUz74Po1BbSj8yKOmB3q+pB8OFyKUmzAX8PZE7OLR3jPOmgOdaFUptIn
ptDIhcmFEnZCL0ZdJufYlGt9P4iLNAiXV535OY+PmHOL21MNLictUC/vjNLCFyQv+UHMHpKbxOtt
IwZVVki6yUVq+Z8OHeD3kVnt8o7AJI21MWqtar405WbwEbOQ65pfK47SszsVBHowqh9sILTH4kpk
3h6R+w7LB8yALeTNlfUke9mAZbANDNEKTNVP6DyuLAKyCoh8MIJC8klyG7AbVN1mJ/j7jLSqL/SI
sHPLiyhfuqUIrN0Kb6PKKsyTDnT4icGXYC184rymIqtmEdcOwvFsN2S7uSgxZVt4C9He343nqVLc
jDpawwN8IHVk33p+3riMdZcu18UaURuTaVzKdUnlpvpPaTV2rl/9A/4SeEzJudE7j8gzb4DMRSoT
eN7DivD0kxn5zMxb5sORDGGkG/jCwOs5bwIWTF4ackaLsliIfZnWZMIrx5utWFlf/WoH9lDtifmW
ei2dRYUfnVQ1tktrzkv2n4nAMtHo0CTL1wY/CEjzgzMJ2d2VeHLpEHthZBA2n52AmzULMUjH2SfH
5MMS1yvZ9bmhC3Ig5QYyJTaSkKpglafDA0C824yurBXpxnp6x8Fq9DiJz0HIyJQE4XxeeQeT/jAE
mcWr2ZJ6EM869EjToRSR25AXO9D7tUYVhKY5n1CGNo6oSp9/nHkvRaaizGiF7fV8KPWas3xRNvMS
niKiCxHLFuzHc3j674mA5JbjeO4WLsXjUNbl9ZdFqfPwzYZbWYLpkMCsNT4dnE7uagfY/dx9WIAE
gLbX8cgJNPC9+4VrTn8MkCE4hLlT7h8Zzj7NrrcLpghv2E+idgQgSEL5MhKhYGPkFHwGAS2ZjKw5
n2HJvU5S2dXqLq9aEa8wY6pKEG5KX0dnNiJm8Ps5bsimuLi7ixyyz7GQey+rPrkn8Y1caO3Jicnw
mH6IIPg9Y3GUx3qtGcUHkXoWL/+nLup4w16xwYhmGkG8vLKtUXKGUunZ2OQmLBiUmbhg9hsrSJy3
WjauxH+XJLDm9BqHhK/WxLpUYR3fC0yrgHCMQufL45iyBRmqeVhfJ5I/U5REZ+6mBkJZdoF21K77
sa0vlxSH4Ks9m048uW6wfLAXyT6v2tOytX6QpuslhDLOHoDtc/jylso9Osc2+WXXejUojgL9Gr3m
nJelOFiQpkM5Xfhox4BKN5QlwyLpoiJSKPGOlwOgCP6hjES1UNb8js0hInDrdJPTNbf+vHjIOMIO
tZuFPL6+1oqFxx87WDwvhg2Wh6QLsSOceXQMKhTfIKkEM0u+ihJjM1G0nKYeYMR7OI1t7F3JO8pa
9YtXU/8pO1pJ88T/axYmd8cyu3tAruCw2mOUQBdIM17oramYCor1dNce/Hg5IwpEBqk9DEbuXFaQ
6ZCjFF40pwj64jv/J459ATJT8ZGtWc/N7rgv2rUnQlb/fecgLU4hSGVv8jamLyDwwHbz1SlPn7Tt
LOU0/L6gY1Kh9GY9WQOq6EPubzxbfyBfG3Fq4xE6RYLqomzrJDXrug5JQ7kRgypYzU/OFS63+TEj
7jpFoLUeSxxruRKMmj/FJhLbUU+iR3UX+dx6Zhm6T3kc77VpC5i1cOtAXn+cp66OBG8stZg4eMDG
4R4apSq/VMb99Bq21/iV7xD7p/biX7he41sBtnm64+qGlXyXBH4QfzF1Xt0O8hzET/EqfXFhCggi
s0hZEa5iNDEI8zfw6CUUNKjdt58BhgxZTNefWiOolul6jJcnvfThnmqKyD4LVGn6LF7DKA0spvRh
MT7zyZeiS7cTZi5/x2G6qBgxBPUeq6jU9QrT3p7zfnNtzFDzgiONnokXXnR0czxk+AO7R3uC5Xtr
LCh/ipX/inO0eyGSe3XAs6BEZiUqYNEvMXFKV0/97eD1Db1ao6S+P+jSUPfeBv9Iag7rHlhMTsIk
twjMr83QC4AsSrPs1jBogrS2qqb5qcwZis5DBzuARdGMH37jN7IiZ1+Ev41OL9xTOfiiBqzTNS1g
PZsAGFpAI9mF9/4aTZkMvo0NbF54V62IizZGCy/y0Rkg+4g3hs7dUpsH+I8nhy5SFioy2dExdjkW
zG41CwMAO863/16Q3ZRqBuyL+zW5lTIUtilrkbpBdkhhTUSqQO9N/uTfubQbAAIJUtftauCM3880
L54Y35mPYpNJ/bvJynvz7wW/bxrV4iidlvh9acDVRHVeJfGg8OC5UzIfxmFFjiuaBTYF3pGr+NwD
VaXZkujFTit2NcGD6h18IXLnX3cwq8Fhj6pwp8aXvwNdO7GlGqCtcABZuSPrQFzWmNWsGs+RaZAk
eIw3l7ZLnznUoogrCyANId5H2cq0fdFv+vp4ooGlGh8q1QyTe4DeSLUGTD/osAjR0rfyiPwdwdnk
mw9rzJMHFkJpi9Rk/hjsS6PZCl3YL/zPUkscZ78fJWhsKbDbG+4taHkIGDrrQDgxO2ETkilo3Z/e
gc0ZSst5TZi4zNLwQwo+upSHf/WsUqx9zL74kik6aJLemDYGZn8NhGY26VDJI6vp2StBPvFrO0uC
s0LPVo69X2LqN3mKF8EuEi26cIWe8X++aGCoIIbpBqgoxlWfg1qPIK1hpvOszaF4JZc6llqqQzSm
yZodgcLVWVHKB+Vm1Sb4ZhpYRIMcUfqNkAvizML5YTC0RUowecy3CAevzFoL+Ae6TVG2wWLHk12b
ygOHRG2zD3/vWU+6kDr5Dhxu/JfjdbQfGBl/9tbqSxTgcdIy40ryfJAbdB58YCkFfHOIOZZvhAZD
m+sukbwx0RElMv0lk8vc6AqGT9paqCv1VPBOSw3JArJNAV3a4n00CS7zC+zLFbBNLDe5oFKquxm4
AxPqeeeSdDPNXR80slAxPll/AdBYStAiWQ9eIgT6T9OinjdX7yqoVqku+ibVMcdvughBbSZYvN7Q
XH84Pu4Lc0LuobSRiOvkaOhH9B+m3PEDD6OLmrbv/bVoJe+jwWNqHrFng5e86OQ1xLJGjuydmoxv
E7D8cYYpCt6E5ZrEDupcnsSXIRUktGghhUwLQLjPUPUyA8Sl81m/cvekD6PutrZxT95m/np0RTHt
OZ2YveE2IWnNWQ53R/OvZNal2op+MLmMKFFzhTkkLZCBV9xyXiGGvxiVNbTwKpVM1OLgDc8y8V3u
Et1a6V8sfHkOC1CtvnLIUO3SjULUIkxn70t83SYGRiYNuJoxvUFZwEBbRc4Yt5tZR9kTIrA/p4S6
Stdz2lfTuqxXzLTb84X7AHptfKya656kHK+3JJIBU0L0q9iJoKPIAuh296XVp6uJfXtHxEVEqiGn
KBWxXzYasLX0rFRa02yfOa4V8XsF1e9TfzllISNhEU2RJrdZrVKoRmabj+DCr2zMpCBqQJIXUfIY
VRTyprw4vmbO048hOx+oisu1/NdzfXIpt52ivqxlZiEhGyHI8H43LP4LD2jkXf/7iZAQWoLP/NxS
z3whZGe045i+pw/jb9D7iOpm0pJYzLoACHIylqMGlVIH3ELGcSvEkYsDgfSjZCrz+lHj7nz0lBEg
nMMstdK23G4kvkedQ3jWBJ+IFCEfG/L8Y6ICop0njJGlEXKiK4gRnEPYgABjNbUlDb/XXUUqDlNy
KzDEfVkRgcmgEf/dmD4juVePlwbA3fR2yhSgleVQ56Kmgxz672iU+tF6qF7TFz8V6auretobRgV5
s4+Yv05oaUWMzO6LAt0vogkCt2Cix7FXU15x9z5Ki57cToDpBMcKWxO/2kD+ZFi616RDRwX+Ovu3
s279rNH/7E9skh2q/ny7KtNjumGsLWFxsVqRKxodBk4jJXtI7J/+xNk/BAZLDqeA999asodgTHMv
OGNpPyWs7k+mVVKXWWQrutShemO+RaLoUZY7eJNu0i94XubkywSiiYTmnFBuMtbnj61TZbIztkx1
Nratgz80S0UIuvN2tf7LjRJRUjcJo4aI96UEwGxoDtZRIFq2F3eOLAmza9H5pFFn2/2vUAvJmBGf
Ww4mu7VqFj7PU7UYpWf+GcJNwtQosyPGtu7OFKg8XFqFFAP3AeaQdJEcdoQT0DZPMDi+sdOugZw8
rLjK4vBDYivnUARiY6UB6r5G+MYqaV2gEe273hfxxtIsOeCJLiiV5DROTwGDi1GE7ewX8KV5RI8i
h2B8LY73cxe1FElaBxeaHXiK3QkwjlAp2a5HQGUdCrhiX9MYXvfOTHr8MvIna3ECCQQyhWwk3XDT
rYu9wFgOBiI9Az3lAYVgaxc4kWu0wo+hbCTmmpAJptumGc/soxVHnaT6GZh67rEB2+EMkV69yb3m
zsoQeUCnnmji+JoFg9A60SVWxQ88jTCYi5wQzZWhLJH98KbHVkbkXg3RukBzyDcRtun1jpF/naeG
Bb1TWin3zI7TAPnqbOiPlhoydXLMbw9jKRsUJ7rQ0y5T4rdCmLqj1C7n/fgXXlOo5SO7AachIAgN
kEAAHcKH1ESsZD/7JpMe7WkFgP6emmFnoCFd8SDnpW+jLAxXfL9JZixHL52/TQZTM69GIP1lfwGR
ZTFwctbvLG13Cd2Km7Y2RW/RMYU0Cqucb5/GpTpVHqqdzFSeGEvYOq0JfiNjM44FONZQQEqtxs8y
U4KBfA+ROroJRUq+b9luYch8DedzVwegPwjv1Ekz5RB/v94RKsk7LOdKRB+mFp0DesroypU4himf
LzsbNy4mPjII73L7X1aHtj9Tu7nOWDrB+dtGgECLMKrch31AcGlnU+xwr/4CZHG9dlm8YcGMXzyV
Depa5RzEaBZgHZtISIdvV4j5bC5LR+klj98EivG5PxlW6OUtSp0IXlShceFkoURZh4ScU61GzdCF
W9DV+nhITe7egyQAJWB5/gVTr3D/WI5YGGTGrmF42z9Pa8KUqnRKHHKCE6sf5RsJjWfoZj+6c40H
YQZg+j1ffOyxmYznmt3VCkREttlSVNUq0q/tIj/x4uPJgYGqeiJ6wXnt5rdjwYb8U3uq7JkCUugQ
RX2coFIqpYSiVo0Re1ulIaElvdhqsvBdMOoSKrxXHk2QRn4gYxggQFm2phqXAKJCyAtcc505UfYN
aADM3mk1HcJZ2XhX+QvZW1d82HKRnur3QFwTGLvL+UxY8O8Jj24hOKJtCVjWYOp+d8l7LkkiepeG
Clvke3F3rTvtO1wd9jf70bLX3xEGhWu44ci7A9d9jXZiyEho7k+HfJYB7feHfaakCxpGv6Aknj+t
kC60UIywIyDJTMBGE8ZHU91sinWH8hrUpE/aOic7zvi3hgERYojdYE1/iCw77ielP/l2ZCF9dSRy
0nGT93OQaKkAScSQ9jmW3MSJRattuS4QwazqEmrXmPjIbFNm0jUIGlh4BK+h0T+57tWVD12oku+u
/uuUGJCIPCv32mZyDvNCuuNaqJC/6/VgMpRr/AOCz4unyd1OfMsaggsAYxUQYyUQxSlV/rMa2EHo
Vp7PYjlftopKbVvWoaswBZRpLIfBioSqmu7i0Z/g7s1xVVsRG5E9Q7oIQR2t3iJxZGQyab8p2SYC
ahyRkcQw+Mr2EGHto0bAuibrxOdibJNsM7vLIzmgAx9CAYsMNfKsvVX0MzsMsSGVFVNp0BJR7YZk
K7b/dpx1jma/9OGouINaW0dNNOpMx6KDEPtitnxdSGTePtFhXc5wlqWy6qdYweWsoST6kk7F+C/x
1uICm3UUAErx1ZfUSI8fraBbB41Y6JM4+Ne1geqo6NZD0H1W2hzsw3wqQTyD4qXg16oufYWcQdxm
kwF4EfaSMZAcMAKo6JAzFru0jw47Ag+HCCdwNpSZZk7a23J4eeNLXufCki/WISMc1Fu7rnp84SG2
oUhk5U/VIQE/gdRVfGDXT6CY27Lb0A/GvPUEYOOz3bBes36FDxRfSpyFUubZL0n46Lg1L1pCm127
5hgenOqrud9hG0o9TihfE4oj0CimY3ebe2JoIIUU8MeEflGY6e4PZouJoden1lpCOwq2BsNsqeQX
Mmr5lai2oQk6uUN6vIhqmxVeNZdA/itNDy2Uy97fo9gjlpbJ/w+A7u+EWA61B8O0exh2dxoGDsXV
+rHSn38NpSzr/fgm4EN0TTpqMtqK0k51xoSC0g+UySXYzhJnm6C+JzZH85ic0FrWgsZOa/yv1bvV
53fsUYUURGVshnxJBm/Gqbyt+FSBV0S8qjiEzLcu011ud+sWMoiLzov2iaQb1xDuNvkEPBFcBtJO
hY1nUxEmqsI1qHj99RHtRG+a6TOfTe4GIqjunk+9DzZeWvbo6qX+MdFF0P66zcwWwpdNduqErzbF
7m5x+c+epfcBkfM9K3JCf7wTXwMvpE0Q9VFasmdCiHOHY9Hzf6RTgtyUvk/TlptSUfNW1xWxpWpf
d0td12WTq6vkPSBkKsP3fuJxzGm52KjK7eYIMebDa1ssySxsRnd3sYZVvI2D2dBNBoDFRSQt/Uoi
dpo+62gqDxoOc5F0q3N540kheeAcz/ttPLmOl0dmG44S8VrpzA4Hc8EaXY1GDN5p93752/1i0xUb
P412S6GwlZFxo/J78Pm7G1qTopFRHfxJGEKtebgOLMih+E8hyYeaNOSYUnIqhe/qZ27MoeTy4rYK
5qwQ3Jwy0Kx209nJCCZAUPEmgEzI/QWeD/2KOQiv8vv4phJZS2nO92HMnyD2caQvPXTShOvNXxCA
HhAGmKajzeTjKUlq8Im+vugVHNDzxPOVSkEFVwWROk0d+k7HpJqGf0zabLUmxGIec9audZMlEZAn
BIE4IoxO75hC+yjHbjApPakBCXX24Le+r7XOTmir3JUlvSU/n1WAPqYMx8a3mrO+oqzYgv2ZCjQ1
aVKTVcoafOdu2bUI2i2HyYIAuisgRdDPoERbKN90psu6VMLM2dMLF9iwXWwFzx6efYiS3F/W4aet
QUmmceccx9sK0XKMfntc9jEyQ1IdzxMwUO0gVyRGWVBNQaMvduvjqmJagI6Gpnyrkqt3DAkjqiK2
fFcI4hVp6+nO3QqjerQuC4Rcw3fB1+tX7iMndHKefJSicljIAa7gE6FpJ1gU1/Gr6Y+fiJ31kAls
Cv+EoO723QE3l2tVUXdC/zmW51/NtTnwAHQRpIZ2k2AeD1fcObmfoNGwMDM8lNInuY7mrYFv9pkS
JhpQeErxsWIl+qi2BJTOjx1BhAOBXcijkYXrCSxq3ufD/ODtwd+Xe6lXaWN7wpO5hHv8hGyK5qEP
k3iUMfE/HOybnNb6adoyAdAARc1/9fNC61K31AXkEf8qlPrhobgg1nAEkSc2GD1CQfvaT9HNk7io
H9luqLJgZTfEt2u3PjgPe8YBVrsnrg2O3Z0lLIBLgPO4CKk5X0EPB8gPXRYYIG1hFuzzx1Iq4Kmu
ZTgS06xbyYLsuASEsE+I4sRmZWkVL9sEP4ApBf6ja600y3iLppf1kRNzKbHXQR+hNaWSQsVksySF
MLPSyTSNH+SUQfIJpG9XYkeBpPrZZuZBsHPLsrQW0BvCS+jrrcCk72RWWz/tlYQj/eqv9iFBSKVl
tbWCg41E/6oEcIfZdWdBA3Gk9MUAj+eUoIXCppPJPflvmiVGr4z8lBrj2o54NxpYH0YQ6uMZp8np
YwJeJd1U7NaEN2C+jRMa5eUMkDUeXz4VSjwvyY62zLQDRPkjJ7EafAC+AGywTlp73xs0Bnkp2Bsv
3Efb3Bd4NggO18+F0iqx9VvBDXFbE6p+/iLwujyku3P4BR0OR5F7Wc3LGNFS9AOcZkFtOnsQkXYM
wiqqIGeVDijc7s5zDhe88Lt2rFcyNX0XXu4qyjVBwOGABc6wj8W1QaFL96s5WFVsDboP4sem2Z0o
B0NkenT7ieCp8eQ4OEr1rUwa/LASQIWOXZoSHX6N1LqUb/6p1jFOaFQwfogPwjgijE4b9XMgMoZX
68RK4glTBJS9K/sE8vPwmOMmOXzPqMh5WNq4Gbmj9xwwxxw2SnH0e9wztH4L0a+ZYixniRfiMoG8
nh3b6h9ZM0JGmxv8omlj6vy2GoRs4d/iU6ZpsfXvHUzTNZqKVhwaNwbuYJ2JAFHcdpUv9GJROxVl
Akbg/15GkG2KPkMfyNC6n3rEFq2b710PGr0O2wbZmG6O4fo/iX0HgLMNT4Vahn2EXzDWewPmEvxT
fZn/IqEp1PKhZTfinp+uyxDxT4AvSPrOFWd/CR36qJW1TiaRAMidQlKnuk7xo9oJP6pQ3FRtn8YY
nhkYcYYxq+GIDsu0vwAtlkZvTH99Krob+CkDVYKQ2ffYShfmSVNVGUaTvPViPOIN2ubNTf5eqqXh
HOmqQgDc/1u80AuLc0y8int1TUnK9zl6G8intKDIo68YFfjPQlaNzSze+kw4iNrmXjc/gptK+SUc
7poA+5/sQ9ofInpfzDFw9ptkNwO214TGr+DR9oNeLarYKdF+72g3kUX+MHGLNphOeDz3O44DYwUz
6JSpQHc3QUD20YXB5vaykv17hk8s8AqSd0QguZ+TOwpIl/VxLRWQkeA48dlSFwnXRERu0qV8BitI
WT6Y3Et/o8SYQ1uyx7P+XZN7Z+jMySejUz5DUnbPcr0eJYN3jEE9fy52OmaKn/st71sYBYwM1MQh
Jt7ISF88tDNiAVi0gv4/wTZWepe+stIkSnrZpOLsAqutG8UY0KXbsgAWdQjktawcWP3WJCdRKL9J
5/DYnF+0eijXIEgqHKgXCat7dJgUG0hJCLuw8/GWgfFI7bUkZN1DfyuBx76LdXOEjuNInXnSc9mP
T7/SknGl4/2F7u3ogV6cAyvAV/FOaoBOROmKII0v3iVcHNn++hPfjrH5EfBQ0hiD2SkNQQvrcIQq
BTckgdjrIkii2LffYFSWu51fDAxiNXWSnett6UsYicFxMd5n+54WHKAtJJ9M1fkj1WQkiuQz+L1X
XoL0Z4YvnObVg878DzUSiGR9fiWaoVUoajzm5QyNm6N/Ogb3mX0DLoVCVgYvtQi+7zZg2BNCXgby
CZFy3tAr3hO3kfv1oNp8L+GefygZngl5wLrA6wPiqc1Lytew27XqexRhmRVeia+DGPHOwcrB+fW6
9NWdqR3VcNR8NMY1Ho8XOHwiC9KvauBp1yjzjqoygfYesr+bLI3uY5oHMWNCJaerniRs4pDWggXC
8vt8owk8+PAzkwMKZrvTAVhn27cJSJDLR1/XEiyygzh9vX5wJOYe2iKc1qrw3YIcP0T52K9LZIWF
crdHo1XkngdhQWLt66ODRY/meRfn844Y6r8Io6V3txpUa0Y1nGjJEvCmAX1yZ8LXWGQ3Rn2P0flE
gYBx8IiE9PKyu/9bfvNBACkcsYhVnNVRdSzFAu5b37p4WFtEaOAUE7HU7FU0cEduIVbBKjm8KRO3
NiFsk4Hc3wWgvsMQNJJoUIiaMI616492EUJKU00dtJDuGUdvFsFFLAVWra8ODofd1qX/e2eSmE2J
rIeq+4HoWZv1N2D0Ge/ib1ItMO3mpSWQzDY/Ua/ExDa2hgs9+yOAxtl/qJ+E400vJ3I15vgJEZuv
SeJJ2t4l/Jq4aCcyb20Z2NmhgiUkFM1xVeYJN6CRDm3MfAAsCnhnXbVMWGSzsEkcI8DcTjwNqacv
A4JEKb4a0b3PjEKqL8WPFlQzf5tAs3bJI7hFDo8938fCANumgtN7Av8N2KZHpdq5T/DMFjpTGq2n
l1hRqBUG06p9Ga6kB/MO/pAgSoISfcPGjBO+d5swJnShothWoXOFkhfc3Nmbx6v8YpVhfnzSceV1
+J4BNyCH3c2J1F/+kocck76HoutgDlHI4DmtQZgNNIuzBx/4AA1/PV/jSZ3QZcpewBwDhzsHdaMg
g1vlx/7GppGYzSwc9bY27tsYubkLa2CnevbUZkRE0SAR7uVKOF/GnntPGu/PlxJj9rWSZlFq2ZP9
YdhCncfDd3NZvmADcAXD0DVoaE/jVsUD04RXj66Rk+49/+C56zOaks6JzDKPuW97MBN4lDU656Wa
mElJrcVpmADTFonVIrDOHCjNbfHAQLKFvY1xr0T2ace9lsqbx4EcTbyK5pv+qiyxVl+dqOfGJDq9
+zkG5Xo1Ru1jw8SIFjwm/gJVN8ITy+iGXkBdjU/1NdW0+4tY6U+w3phd9lzlpMwYky3JFLYE2F0S
DzPMvN0fgKK+GZyOH0ZutfNKZ2lWA/nODBza6cu9HbgRMLEQL8p0yXTJYxuGrMhn9cmuOtpJeXKf
9dBuGjvfKS26GhdOF4zSTIh+X6H5fauojO88nv2CnODnwah5X4M7LJvyJpnuZqssvZ7fNb6r5Dhn
/UKL6slIn1x7eVobWSZ2+THir5s5y8kuX3Td5Q6dtm8PTW8wQp0U+vqly6mAiQjEem5ftBS9ylTY
psN2mxCHBdZXZCSHnAu/0WVKJmUUxpYpg7TpwW4SjSIHg1nA6RR2AIlVfeIPNhR15SpXgtyrK5sv
WyQULjyEaHhfDqHEXkcj9kFt6QnQ4YLj95U8awG2b46XuK7HR5NP5sT+ogYhOpAY8qeFdhcUIin5
M+Yd/cTqmmr07mnXtf9KIZwtJMZwSKMY+thyl0HCS9sqZPoBuhrKANj+ffTQ8Yu97Jyj1JmeRJQ4
5rxd9pDIFeX0u5Gm0/jP3uIsYN7icBBg+rCNQw2EoC4hi1s/tQ09LucNq0yfGvA/908W90Ae6avD
bSkZPu8Uf/jMYdpTBHHsccuGDbkzLC5gzy5HecDqKUxkWtrGZR3NanKkhgo/DybUtXPy2XPCibnV
hxhPNK09S+bNKbamLwT9JqzmANAOAhVWvh9uSsxnMXLOzveZ6SaluM5EYlE0C7VUFYwfpa8qDpqu
hUX+6IwDE3Ow3nNevEIYqeXJnAvkPsTv+jtyqvrRs01SX9W971zw0qrFzTgGPxdbvkHv+m9xySf9
K1atxdioTtJa24ggugLLtqAp1bumCfRchJc2+TLVGgLxtz88ebp/hlofByM6M684+ExGJ2Vo/ioM
j/Q21Vh9H3Bb8/m55rTC0HuBV+icmWxvNUlchTxJ6nRzMl0O/71kYqcVzNlK8IrA45qid2HaRXie
g5aq3P6FlT3upRHswmfypCAsx8Lf+yg+jMoRngnd4w3Uy4lzPUkKcUTIYbir11Q4s3vBrzCfnTSc
w/Sd6LFNbmVnJMKJ4oAGZs6+VudgBekap46Iz44ZH5h+rIorUzKDB8bNki6Jpfe63OsPZnDCZu7e
uDn+O876t77p1sMgY9LekLQ4HgNQ5iK7AS+yq9gjGiAgIbKeOQLguJgC1Id9om/JZFun2RI6CT6j
FtxwMdnaj3XfXx/NWpacNR1MzniWBWWLwJHeOzx5Oo1ojO2vrUtVXkqxeM0SOONjzCG0k4NEUZX8
kGJ1BgVMuzg9PZT7KBV6UTyNFUxIeQEfmfUr8eTMX1CZrIAipTfOrNqfncXxDV5bCmtCneyAfW56
rPP8g1XAX8WBAGnepViTLreaBiZbPUrqmTzsGQ1u0zXZnQqADwNp050Qn6Py/f0RokeNyVYSa3ba
GY10DaiGuALp+LG6MNT4+Pb/WDnmBfl8Qupsw43P3JNepHOxh+jRRt1pG7HktpnDqvJotPkuiaqZ
2URDgC2TWJi68yBkBVdsamT7VcoguEFyFi6gEpycFlNdZp5db/qrRJVCqKb7li5/KZHhUBUFPiaK
JiXtbhvGKU6sSDMk3C6CG1vuF/ToJi/DV2cfGXEayEc6WEc+g7jn/1WFonjZPiOEkuJFRXLJgwJ8
GlEpeqx0UBNQyMU3J5/v6kJBIQuXBrkTBv5Ne0QMytCQWuPLlOngb1R0sAZo6A3egeHr37cwKvqL
f5P+ZwnrQJdiAGKD+o7XWCntoTM1edTYEZJ+ctiXsOclbVetDjvDU5bdEfdtJqdR/w6z10famwLo
d8vBET7lZGLPBWZsYkGYzS4SxeFndXR69gyR7jjPWzj28Fbb7Kni6Abe6RU9lqMpZgWtvpuSRG3S
zv9MfGsLS/VjxNWsxE1QzzuHd+3L0nkquRnzVGqdmxzfJqqP5uSuWQ0FnnhsRQ3FmbnjwTfW5ggQ
mbqB5FzZkoWObiXQqQu+KpZnHOEgjdwBO2GeA8X+vAAtf4zEBcL3dfbZcLQ7nj3yzM/AqG2t1zMs
5eY8RMPtYm8WaGajYfdo9ApKrpWgcZwxWCVUcr1k/ajM8nxjZsb6x0nKGBzyzhBUm9Z9ssWSeXV6
8cHWFP9Q0322aj+tT/7ZKxMHQpJ6M2hQIZImb+C0wjWMEhEecicMk/XD6nHo6/lSzYoIvitGXg+Y
ejuZ8hsnMkkK0NFeaRG1YIHZmG9A8EaSE4cGKMQJRrylJQaTjtmioHlgDKkrUEgas8bFuBh8pcTT
Qwve5+OngO3OIwFOv+g3DrCqv/qr1pqITmEcUaSLoIGv32D1hhP/7iQLYTgCXm3rj7jMoNius9+W
WGAu7NBFwZWZoRO5LI5LLeR74T+oquKoEEQpeqO4VaN9+YrvOOa/AGybPNoDYAwY6QLkk0h895VZ
tk/8jdczvpfP4q34DSnJYaXFFf0BMd+uDrv45sp+88ZPLkn4ZuS2lRy3v1w05T8Vc4NONmSC4rFM
eT/tNhy0MufAgAwHqFU0mbOdG01VZsoAaWZzcZcXBnAyucnbzl+wYm7E2yuFLoDsYIGljBUb5pSD
541IUl1LVHy7V1S9DRMr7ABRJIY37kP0QjwNExUTGGjgyWxMViJcP3YfdMRhHy2acoURukJZpCC1
mnMhLQOHiLcCehV/OBCEjKaWxlinFCinKlvLekMmFhWwHQX6SGUdZsx/vHzDZAl9swUrSbjqEeJK
j2Cv1rg5MBgsb7yuUVWYizxzVRVvb4/k1tOE7QFr+8LzH7hAGINHfXe+C3Qiju+faOQxKDiErPQF
IljG4/ldt8W3CDOu+jQneHciTD58vdF0K1a73o62fY/s/S85wBh8eglCxRn/NR5SxKicfbzq76lL
aDetcVpHNHXttaEanhNX39/1ufBOy3eicEK3DxyhynjrrautZk0B25Expvc2pieYT1jXzupnXkSb
BWqlB8nxaeOAp5gPUF0ace/qO+lx1jhuvcMPpzIKYyoUgGlkpDOQiQt5ReWUduIMxNU0Vk6fQG55
kofyQ0gjevXEDG42p+Oja8ffSS7SbGIE8wGenNR7pOR66tgFwHaYCPCv+GapVoXl7yIQxSmGuCtz
JX9l3KTyM+1iGFiDkwVZnJ45wlcLeOaLPmwP6MmwoHzhHJK4dqEN8Yzq7GFaCepQjWGEBpEHglmV
1YxyIBzJBkna/+x3h3dF5htliPxTjoOSBtyCcWiUhNQGgkJ9p1TAr+uGSK1at/94vDKQYe+vLnhl
zISLO5eSGnpkphRf4RZOdqptpYsHUfGaMzYfmg1aQZlPNN7aRwNBYfzeC6TqWo8UMSKgJEUrfNX3
ozsk2U7MgRmhsFt9TO5L9w/VTjJUF/1CXMqqHC+Y/vzYImF5jmZDk5UDX9aQzy5E5CAEkCIgYiyr
/LYDTUjoECaGoRPKiUKvygv3J1aII9anM64w+MLQUffuabezkvG2bB4YO7ylCX6Z8mo7eJVDcEut
9IsWGFYutb1bEyM6Dlvu0ATC0LvGUeJU8PJCJljp3iE+8LJqsc1CrYlsO0ukQYVaPYip9f/9FyMi
AoYGrxvN7qqhOj/A5+XFdymgzSekJbalUL5j4WKH9SvD1PalIEbhHBFipgYaS8BkC4vS44bVJX4E
lKsLD9MfGy41X0LZoUeXfaVrsXDAuQMxpZiRf37iq1jByKsNhbDpy+dWhlgz0tSNyyB4k5uTaAuq
7vSCsW7vlg3OHP0c5z4i9AUCB7Wu0C8lJ8hVFmG5oJ6+QOzezRL8Wj4qZBRwRRbu++ybAL4VY5Av
dnHnt7SKXVzVy4wSClPxdTf6EJcibLUM7DKpOJ5QhCtAaM9fJiBR7Dt4Q9n2gf5cs+csNFrcNp2M
QHdZmgBvp/AZ3nmfqeM+/TTi+YINXFtm3IKHKx2Dtnu89DhVpVIDz66Is6s+SlPBELptz7ePIzYY
AROobLwL6f/A8da0690tuO4ka58qyYp3Q1g9wQ+FxiamJfBEaSvMvvf9D1VT4le4Ms+olFTtSrz/
TkN2AAK7iW/ddhhKeetm+qx7vBXRUfFqX1iz+wAPcVE/vl5wi4/Q0LxcxnyAOfLAZMkEDSqAn5I7
AL5b56JOuveSIVWm3okk/4KwFekswdR9FcCHewbBww7nGurV9F2HyW9k3vK8kZMmusUdRKBybn1E
4jCw2xAFQSSAxWG8i1QMB9bD3SFDcvnTUC3FsAwL50aHdzs9O1XsSRis8mLm+ESnhokB11kRnq+w
5zW8srIZUepK1hTJZdIMp0z28e/ULvwPzxsLeFdtd5TZX1GoY/uEKZfbWtzG3yU+SrGuuguip5Dm
vidMPK8WZb7TEqu0DxCF1gNFOkaBqXhB8lIgRaPeUwdbbFQzuNTfhf84+FPycBAuTbLpP+hDRSwW
SEEN7Nu5+ye7Deg9S4jpREmm0BzmFAUG3l619wYuYIjhpoPOuHHFq72aEFwVPS1ZWMtkFunFf57y
nQXnYJSDYoqF5s0epDhKvA31nLyfxMZmTI3Bo08ef6uqSZaQ7xZMihdoJFYySinWLFV1jGiwH57i
wGTBuylsFVQkMnxxZiBGVsqJxx2ybmi0ueenGJGwHesu/QLJwArWlVv+rf6CTZxdVY/aDbp/yRAc
1cPgkJPJzbiakmHDfOTnxg3KsCPb+ZMwD4OzWWX5h1zlS8sAwBowItOYXJ8XVLKQchsykNPjC38a
Xf6W2/YsKjWGE8u+4S+b3xVCW2BscOUqCpU5kPg9AZLIJvHMq5BrbdbOBJVeXrrIE5XGsjzKFPPN
i+piQoxVR8bT8A0y6j9kQH7+b0fZLwcexJGd9R3tprchiiyRulPKHKsRNUQYMAqqDcfjmiVJw8Uu
6n74bQhHP7XZKnYCzpurp9eRXOYzPgC+9DSthKiPe8bwey3WYIYiTT5N3GggkVW58EPc4ZhEIA52
KZy9PwjpLGvr0wWCPIqCkDkl0HX3zDv6zmZVgPEOTjy4L/wiI9DRIzY2SbxgHXBTDKUZrwuCMc6O
de7K9Aos2CwzIST+Oa4O2d4LG2/ZSpkAWJ0mmM0pEu+qxKtLntEjoeT//myIPsL64myyzbRprz5i
GtMSHnMu+BXPMT6R9apRZV9iAmu/AxYo1yloDza/1E0zpn2Gg8zryAsh1LLH1vwvWroa/38MOZYi
CsKa8DQyjFYWkTDvycYSz0DGfMuQVfH8IXaJFHSLZF51FLAWX48yMpJH6CHZ+FBiFKnxroaGxSpi
Ghx7N40wjB3/xxSyweeMJXUqzPfu/a7w+DhUMWLdihYDp3nEdzDs8GmrezWPQ6SZyMTuGieyCJew
CAvKgldDKeX7Q8jTIUGVa6m/o0jqwC37YbXXJ+WxBMWf0QDN5IvOacrjAXv1M/hNpkrZ82snhMVC
i7A7l9AbmuvufRQjiD6X5fWI5eELHY/rQNspUmYz71DRahAq5ib+9MFp6VcQkijuVD8FmeLweC2n
OIda5mi5mAMJtG4T0Sjl5MpNwvYW7YBvKXqMyGLGZmHgkcY8lK3yssCW8AzMlRB3ZbTOqOKP0f60
NCGrVymFt75x9Ry7QbPkFhZTFpbo9iplgoVdplIHFl6WuR0EMEZuEjoiZyFlwpgco0ZIjltWS4R5
EJqG5T6tP6mWmUoa0T36oYzQELRoNffDN6T059p6yal66wE8T9VgrHqjp3D3dWGLmFhUaRcZ18LD
63aqL20+VUzJxsdAqu/SAbBXVm5gn4LI4rk3eqcY696l9Utk/a/5AT/Io3AtCcpf55g0VsMhN8Yh
ZFCqjb7rZi5FJL57vzcbyVahKKTgWtMziGpQD+FGa8WL1qpDVe3WUC+0cftdySblxkD7SwzMAtks
Df2qIZl0NaaLzGs+nELS6FLuaSU0nt+fORON5nG8o2vnlroYK6M01JdJgtpfcAETZZ9Jb+okl6FD
lYNYFukb3IfbIgfAemoeqOZfqhn6QqgAXSycZuYlKckPDPnwoxNLb4AMUTjhG/1dz6LkxnVRc65p
4Y7nXo1cLDdlrD/pay0jfkmvycuVa2DW8V57tz2cTYhEXrJVqu02oE0dMvwLmFDRW7yZb72c60qI
KPnK1otK8CJ/L3OFY5qQiIhCd/s+Qn4A9KwSzcUPSvMOnOTmyeeLKp7syyHJ9UA7lQU/17xO301S
+7dhxNAmRINJKPrrWZ86wumxVL8FUdeCxCpHur/F8l0T/ZIYlj+6P4qCnghL37AmqImzxHBlCSQD
Em6gSJSHV7aFPgMvfSUIopxFQfEWJKQ0Zg8FS5WZqWPy0GDRIvQhhfTzUHRYVw6079lwUkH8X5Ey
e0ER4QAD2m2lvmBW0iLiPnLCeG1eFgxjuCKA1mGApziGEudGKKyNvgOvsfPVLbsJk5BPAhq1VJHd
k3VmEH+gFqZO9EjH/Q7M7CvObeEHUSSGHQZOeMIuNBZfsTRbHgLcPAl+RlpthLWRB6UCLOXCBQwB
a0qaGzqVB15qTAvYuZVWhFgkvTOxCLNrdxmKp/fIYS4XygEo/wHELau5giKXIlrfWsDRAQcXt5kW
f69fyWmBojvM63PGWIlmL1FA07K/UPwmC3htdydlwb4Qh882W0ii93dHzTVp2dehxc2fSOFzKXXp
VHWRLS7wqTCZiJGNbdd8GHn6ttO0wSSO0W0mCEt42EvFLZS2AtASqafHOwAgW3TgNLp02nH7QclA
X1mdf7FWQtxlle+jPQmhve+0juUyNoqxlWHCVZteiihDgTVb04NSkkVtaG64Lr6mhhbbUgOpWCYS
/bAZyGNIo1rxekQXKIywutsPSCEveDUD3bxNzI+QDyhO18OquhhswORA5uJSk7bmsU804uOjVatC
LrvA9OrKcYJchSbYQIs2o4hyxec5jaQXiBO99dFzPDYlBBdEPFErUDfAbltQowxVhjlZ3StFlrgl
MptwJbSv9pvxkZfpY4AEo7ruZjTsQ2MYzV2C3i8ay0q6W1uQ+GTpXTJ+xKvaAJNtkFWz41sO7cUr
cY4RtzQ0ei5H2y5+GvtngyiZ5F31KezKQR4VvC6uQKtsXIXkp+74h5Ts1O/wgeKbQF7BMfUxnTzb
/S2jd9zviKpM5gH2JBQ5dhSi/sT9Voa5za1MTgaOFePqjb+wVKzAsm8sQLMoclTtqaNIGWbizbZK
OHHkllitaw0a4P+wpApdos/QAgHLP+Dy0FQ17n1WH/WKuvyufjAFsxBWB43b6u9IBljn7Zfw32kt
xkqanm8g38XtFnzkuz7zQnZgqKU50A14sfDHFX2dTZEt4KMyCLhFRqa+trUCbruA5wUvugfpS6tl
uwaBQ3KMBXnzTt48tEzODbMPHESI3clP5FAN4PqwMd3kLQgHHehOv7/pdmFNRnQEYgqih9+dZu5f
+cp0MjGDg26V/JEUlzycPIZ6tMZD/mz+3/atfgHpsNX+pqVpx/i1v6YuF6s8r/bG95DYLUiCLgZp
SG5vmGZyq4Pgj89ZQ2xBRXXTI+PZ2q4y3YDiDoXAkANxDgzG2hQRrqc9btf1av9+iafTxJU9GNPb
j1CCHanYEEQ9uLITseHr731e/cXhfhnRry8ShYNkcBJSb8IBqM1FiMcRrNvsW/Pw36mx8Y94JlVD
oVS1XVY7XoHU7R+32nU98OcQq2wDAalomjupQf3dz2pCI+HJO8EXCC+5cocpnGnnV13tia7l207+
hpkWyXR6auzNMl2I0VU+a8Ar4ZfHqfKPPlArOrcrce+NwteIhmyHkKtcYzcQ1T4ZRGO4oDEgrfcj
V/huHLYwfg01/jOsfiC/qqKKjUngDuf9wdvmN7TDFXdXMQZqKgF+xZWYIt16XMuAh/54S2oUhBOc
Gv5wdfA6ETo+OHxEzeY68dOrGW1Y6l3Ge8xjupYf/FnHPp9ARWCwlnEZz+ufNgBpJCl7HUx6k3mJ
31bnN/Q4iHw1ZK3/WF0EVd2nwqqJAVJHEbY3D3isICYJRMhMW9RYS6Deu7dQ9CVy8INdzemWcDgs
7Qk/X3+Gy7UuIVnPAXhawwekzng0W+vZ7Xxjdk1dJCa6YJilzEojJLKWt8PoTTJ3UiycAzwC3ga5
03ubLO8glpfSKKhG7FWULj3q2wSLhafH4xNsEi0djbQn2Zy1aS759D9beViw4v/4CXoIDFu7GHcf
u640eq0+IFCl8qdXfPX+K4y78ZxvvYSQAN2U/6yGZmussLWh2BDtp3LzkRmLAumi+8oaPiUq6Bba
v/PNdSUcLlXGeGuQmXUWdlRVehgAoz7Xr4F/PIn7i62NJrQLocfxcedNq1cDwpFVFwgvXuG/Fti8
/rebHO0c10Y2h4QrwBZFdTtMY8HrPNwtGdvSg0Gx2N1u9b8BUbCzEu/o9qOUX2CcCl/yMXGcQ3N/
UicOv+O7m171u7BmPg26BVY15pTNBeAFDccwYnmXPYxDoogQwroWf0GHKCxRfC4InQThnNJ/WI14
v+6fCGG7d17Ii/1pB0UgQN6153jwx7HqNg9ULmEIgbV4kYmfub6YYiUcFh3fykIFq+zPE3sqHnwL
4XaVEludVWfAUoQPsIjsJaHqBjLUIEQ1hYfg843zwsBefg3cwNsM1b1TY55v6E1gzLwYeHOpWjzq
UJ3pcip8micYF3MlOP7yUX20orlrNeNTxQUnRv1W8No9CWnpmeEHJJKMYB0v+1fmZVrBOMiG4ifW
U/VqAp+oWmtI9UTt6dj7nzMnWsWfp7ORAFg2+A4/pVdsP+/p29gLFHAJeGUOGzEVDC1VOTxMN/1K
ftrT57tzz12KTzyNX5K8QlVlPdynacuLZHDQrt6eCTjN2Ix9u8YHEkqDOVP0VHauyTg3SMQA+iyg
XL/+stippuiMhuMJeTzUzYjiosyOVZroCtUC289oUgYhnSaVWbjJ38tlVLNc1sGX/slDjOl81Sab
jjKfra1SjgXhD03YAUs7MTKh4Nxd1tML8eMu/ISTYIjPqyrrxUOZ7x8E3ZBWynX1ByemYz8aIWtL
jouD9uhWCz7+Yt5pUBGtj21xxUlXsVULbwZ7M+VDZ5NcbagS1bYMJIwIIICXotfjvgPfX+1jgZ9/
YFNVKDtkFgYd076Ppn9dZSQ+LDxezotMWMXTSo9QPfd1kwobCFB+WcLBDonHKreRLeCuFTHio3Aw
8A3gHZRi6zYAWSWL7/En2SnJW5Lf3ZDyoevs/L2CsoI6ykKYfIRh2W52qGknUdURll9gXTmqPtYb
5k5GUjNTO28Z7Gz70nnoFClbhdg0faHhjeaBnChaI0B41vYG/HohjF694N8gkBPRX7Co30Vj5r+k
F9E8xrluzFfXYB55v5pdtvsSTVXIik5Zs56S9Dh3q9eOzEHWjF2ErrnOK5hQlLZ8b41mxwON8geS
OL/1tRtjmVnY/T3dllgMGjSdxPiqMEFSniDPYWOa3v0BTgT5DjSWZFEKT5ChtXJIhTcVlKH/eFHl
feCRFZFhz6d3tY8WSBnRRQdUawbUqdMjUHWzQUlqUlUzsB/MVl5+aZcyi3xKgrl1Ch+CgDDXhCgW
YXgHvw0zmRH2WUUR27VD7rADGgqzlEuHJim6kcmh/ACojOR4iDd3ALgDILftRdnoOjAMtJ4cwX2R
orple9q0ZhYe3VSH6U/wfuSxCpthFp5OWxovNNAbqbBTeYI2F+hABvtXyIWKDkANg4Iiom04OpSt
15eqix66N5c6fUjfyYTk41UocExjvJ058HR/dqRFl+cDOE8XCGJ0qNOyArnNr72Prb6f8pNMtMQY
psB6U50rUVgDEZKhqlPS7fMNjFuj5ipJ3fqz71P9ewDUvVosIS8ZlYTbc2vy4QNg5nhzYxw+GLn2
lX4JGTCy8vUilE1q5D6q/cDYTmJgQ0uBXCbJS0cltQgWFyxocKVS3B5Bu/JQEySQ8c6yoparLdWU
mBEIJ6Ntmw1D8SePHhtVYcaaubmLQxuSdvU7I4YRTsFp8UHMim7NCJh+s6HC+gNbQW/dHOFIhBN4
u6aoDUMcE84etjP5nK/LUXczEDLZSnbMccalY839yNJfdiiA7h/Kdui3wJ3Dpy/fSMy+mXRGf0QC
i7u/c20+vW/rcSpv3975rfNIi1eCBMVJ8V9IYDyM9PvZRJjWqOYfYi316yeETF/ozTqMKMiZ2MiZ
uLxAn04jJELMUGkBYk1v3Iuj1rgarFKufSaXoN2p8U+KZWd+ZCNJcHh0mqReqjnwx3cBYW88nQcI
MGp6rp79OlSPF6oqVYZlVQKZtJN+A+ZqKTQzZeJMieMATVwKmXi3cd3f6+eyv9ulh2JQmiBUhD5Z
udD4vPY/kahHpdR8EzHK27onxCre5Q86x6rFIDngJq9vNW/4CMVmYbGf1TPK+rZmJLmYgdIur3iB
NKIEJliTzvsrCt383X31oBKYv4AR0cJWBlukRG43a8Nhy9o1bJykRRlECpa7bs8M5x65hX4tZMQk
lRIiVUa+CUG6FLGUKQlzs9IpMZ0TjuapUAylpOa63n5zkWgFPtchV8RQNkU3g2cjuPqkoQtYdamR
3/YcVQ3DOlLL7FTGGmfLwscN8cOZR9d3cC9nWjf30M+utiZQRSh+rV7iIH1O21MIV5E7u7VKsJjN
+YLAPOcD4bsP3+MBjJViTZYjMf6P+OQ6qVfyNTkU+v2/o80+mUGKNmVmydD5DiGLKZBkKznF8Hbe
6uZLci+eKHdDRSLifonPUgVZXdhfgIY+kvGTaEePMiCClhfcqX9wmIrz+Z6eP2xK6KToLFm9rTUL
rRDenhBsDhAg3udTlkh5Wv+pHF5Vu9jkPe8ck2BvgpmUgUla7k+LRL14QhyV+SX1KmKKCemSVIe5
MfsLzkOtGafqJOJx+CJHcenE/kz0C1V0mAX5r++AavgZGC3PoGz80Qj5m0jR3fnEANrJjsST8Hca
HWJb0S3IWJ9i7cWSXVHGRAOw90rbbnESMc/0YTMCSCKbXkWE4ozHIy87Qd21PxD6et2/6yKbZPcQ
RVjAxh6oTr8xZ9Vcp12vjo8YJ61hcbePbYX3qmpWOf7T90spU3rgJABN/JW3joLEFc65AHcZ/zoJ
Fr2hZIo2VIGR2SQpnvVAefb/pzxasHyCAldIvc+nWbNOdUE/h8o9UwsSkM8Qe75a2Y9REAfYtR+J
aX6DtAnpCa+1BFjsp8ioA3H57r5UGsz6Le/ddKFztnMDXgS60qbhVLSYKsDpzZVghz7QXwZHA82h
SE3I8nfeSlMQw+ZxkFQMcz8Zt8fKU/fGj2Ujws2/rViEUy8DjKKVWr8ddj+vyiFLzTY8OtTtf+iC
Y6153cg5dclcIQiWO4IL6OHdhBXcIaJODk23VVbUQU0v3DzIm8rDN3n1G2slKNUB7Hmerd7H3Of/
jA2kxgjjIqWZcttPtSRpAzw7JF3d1g3Z9lFim0YGaC1uLT45mJ2pFt2Lmi155UHwiadUrKzWz8ZX
iC/NNGpG8toM9CO3VM81FSL4RdrITi02E4xsHuA4OPraRyiIV4RjxukmUdLv2WfhiHEgd9T4vmoV
RI5awSikwX68ZTs07gGnPaggdmtsN57jxcPjcBC1eHeo3fSXqBsALiZqSCFJETnyZcXIm6Hxse8L
MPGQQAe7PZXmXz9kOs8jlWWJGGs977VDQKINhP6DIqwcTvHy7F6eIQkXTUIWCgUDkBxr2jkKsQBq
gDt091uLqWl03VSmoXjvjQ6HVrvtFiD3YDgWVAYW9e2JdUUazNStA4hJr2n38LhYRD6SdfMMTNWo
gN98pzqd4ULWE7fyDR9kN5zSDVp3mP9YgkrijzhrXjNTHV9NntC+dKs8eY+xEy4urGbYEv/VrD/z
bj9z8P2s+BPp8c+PueCS5Oy6AD1I29gwkVE0Bu22CPWAlAWJRo56st9e1c9XzO4Mi8HZ6YK9b3mi
BNQ+x27x97NmQvJOakXkxpR+/M8kbpc4R/Zhf+3FmMQHuiiwKiHL8WHeEUJ/2CVltYmC0T8pA9B+
ePO1IHo/YkKiJqUCgQSMb7FWZoVJmokioht0AYmB0GI1wvDwvKzVTo7AsB909ZsgGpyuNQnaynGI
ysfY3Vq3uEYFOZfeq7JF3nTosn69JekobS9KkZTrel/V36w1Olt6gp1i/TZ2yGZdtYt05xR9JRJ1
EQMto15J4kZq5CfRdI6RCH2oG+DIguTJ4CaoZXU30zzZd8q3+9n2YgLDZBnfzvpaMHPhZc0pPYUV
P7Wy4cvNYPZ/JL5AbLPsp0/lQwojyyiaz6xdIt/3HttaN7UMEVwVcAPANGNniwMf6E9A+AdmLU4T
sW/idFYQhhxuL1Bm+AiDltIHj5+o5gqkW3NjIgdEvwX7x3qT6EsBOTz+mMmk0q6o/jxzxaYhrJil
/2SeJ9fJl1+jVfkwqI+uTjQhuS9gLgMO67lLwlj5U00Gtw8I0HiVxe2rgW3/SsUwAQm6K5SxEtx3
JwVFpPZTMDE2381nhnIheX2+QX3lL8W/F2RWJm2+C7AAb4CulLI7bE5cp7BpwSVVJOl7S3X889Kr
d3Uju63Tj5c/BvMJZ3mXiplvqUlxQ86Cv/T68ZrvWMfm2pyXZuymHbRrnNpD2BWiNHhcapobdbDP
2Gk5YWXbxnZXZ7j6CWpTpDcHLMZmwFKNO+BYaE8+zr2StBif4JVKSa4OFbA7NzZ0vxRRcNdcsFXB
L2IAD+DC+gxNRwzzJMiA4awcVZi04dm68ph7YSXW3eRg3GRW098QX6zC/XROsaLlBFfe6nc2KqfX
+jIxjE0jvg2shTQmMsLk82RSbGenhms6EM7l23U5FZB9RtSsUbA4HfC/+CjS/3Pt6GlCUqgdup/u
Xo0fzOWMHqlsdx17AFf9VjJhKrtyXXdWg19JfUt8QO4d3F3G6MyNB3iRlFpgHadthZpMDo/IsIdS
587S7Gu8aS2wf5Ai9UHT0YZZCFBs47S7s+jgvkUshrpVtVN7/V2fsO4/IGFfLAFBqlxTZB8Lb9FA
3Z2PfwciV5//wgUqHbVTha/6dwM9A/wbTMN8NlRERTdKPtmaTIZzp6gTSWoaT094tTX1GmH2vG6S
IMNAVwXoljTVVKvUSvB6ITWsL9hG8Q2DiKnpPkrNCukY6HbRAXWN+wkPl62BUnQ2dpS/5VgIMInV
IrZvosIrMaySkiYWkWid4gCIBgpl91s+wO6irdgukYmMqNRilXhOv3FgztGob7CgYlFlaQ3Qi3iF
QcJUas4MOH4FC0Ip4E3CLjDBzfGvpKqmK5FkdDuwAU3I7/S1ta5FwLagu8NcJRoBD5dTWf2axyeC
qnyaTN1bv8XQibYpKInuEo5zXIpSmsfzhv1+w1pclZ/sc6oL1kgj9y41f4kXuXobmKCkDhi5NqpR
sDIZa++PnYpwrGTnl4PrIGqOZiOu8R8zl5omLP9F9hrTP3CDdeCht15LR5KuVDXJ2fWRKoKKs/Tf
qvV0wzsEZt2kO2WZJ36k+FVk7HraHFrZoCdw+aqw8KrKnjhQtNEvqlDbSV863qg7RYNeZQBq7TNN
34vhRK3388evrdeI7KWlXJhBXzBkYcmqYnGer8UZ4jPGUIwTbKNFZLBj1vq6llFC7pJ9wdkosfmg
3UUNWh9ppJ0Scba9Y+wrex0MbD2q29iydXzMkCYb/MbFHQjd+UKX+KVU0Mtc+rB7s6UxA6nqmt69
HE2DJ4G7oUJnp8glfSYDelLHOcjOtbQ8VIAvC3rFSxy+bckOpiVYa1rFs10V53mn36oEJp8rJ1Hh
T6eZkyGm7X8absQRONcLMRHKiSODTq2RBtCJ1JrAmAg4cfs/4ERNt78HRyoYT5joju3r/DKixdQR
aUhqjV29kdcJSbV2b/AFDiUYNhnRcXESy/44hx9LouNV5XbPRRiupe2SEv3eCm8gwoDybmbxzZ7P
A3XaorM0479mSe5oH1XyOL6tprefnTdEfUGAFjZvizlAJpU6a5aGQo4rGNxl9/1UspC/JVaakzjr
v6B/y/iGilbKpp6qLkzi5TzgeujJQZZwwlvuHOYAyD+oDJkkLuSoB0jQVWWsGyILmDT2uwQ80HvP
reoYiMFAnTlYoePRg7UTxr/+mIkQ7KKfdVXDe0X3aLfOkT77fM8PwRztiO1YXcQad6QzfJJnItoq
CJXUVY0sSPt83J5pER3oTCD0DnA2xLBadu4i2f08KfV0McbKQ0QY1DAu5dp5hEZldSjchIUOGlfd
nKllYSilC6Pe2iQpM4m4PHcPEuVQdGjRIolfu3FvQZtDLdg7K8EKmbFP1nWaKnzBLt+9sSWoNSIR
YBiSck+Os6+SsGSozeu2VKm7cCvHL8bpRXuzHpcl5M2pt0Oekgf6/ROeOc6PRSBcc2FDGyADGr2A
1BX1SwYQ5yMzIIwI/6Fe2CXFdSV0S23L4DSkh0Ta/ZTBZeW5hNGKeqIUU4xIZa1yPnpEe58UoQLu
wBbVxiRwYdTMeQkbzip0PsHJYcVnRwnzsVLkivJ3uHnAUrfsnBoyvebpezELicESQpqSPxJjDPs1
ZxcmH7Z5BB34manzSN+P1nA197aIXDexmUbfwzCS6XJNNI9I38tRnZ9XN39M61MLkBT280VvLLhC
jYWqTZWTQtdRV4Vkgf004XMG+wnDXWcyddRHI5s9wSIDUuiGNstlBOh2E83Mkuenug1uMfbZFHIb
F2ApGAi9rbYztg7+Uc0nKHiVGhc8wjNj25WpfFC5obREBduEt4yyc7poBCp5GU6VoJITqdG/ARcf
DwcPJRN8pU757QqVrb3cHXauBJw72XNt5ixLTk3XDA08/K6RJ9wV3OwqanfULGQVI0SHE+BXaWlZ
nJNPU2hHb0tEvnRJD8k0Tx6O4x1SycaWPf7P9WMqjKxggeG+sH3rSPAtxt03IZK1JUfEXCxS/9Rd
mqf9hwO7S7Xo8KYzmx8s+Y2o4upDsRdwzkdrpf2Nv8ImYuCSziyVATFGWihuy+Y31Cvxio/jcU0N
BiYntHEYyVvueOc3vQ5WeyJ2gocFQW/VJi69hiGZwrEURn1w9pjsOzmBKDHBcmrZEIK1qD2j2ueS
dV20nzLBMJHHEG7+vmi5yd6kVp3iee5oF8Mv+WTubUvf79D2lfBvGcUGINlZWpAgD5zO/03QpcMG
TExQB00OyvLObeZn8m/zXO6k9eiOx9Y6ALjWcvIimUxDk2jOzpT2CG0hHFraB1Ur5auu6xqf88iB
GP+bXS8i3y4BQtorEtXJ2U+wxUAxnmkHm5koruIJYjHpanNGP1Lj4P40nYrzf73mbIqsj0WbmXWj
HWgKVt4IzpXX7IW6+lB8T/lp+XtZm0qkxP94y3WxfoFBETX+6H4yTRm7/KcKLdyxztUSIaH1Has5
2lNvywifps14Y9D4W1c8odNz9/xBqiqjQC9iVn6Mh9wcD8rW9MvplVJJpCKXMziovSCvdC0rso+z
stw/EjSMgXs8WWDSUj16Orsk5PNwN7lVjaKJTjOgYqxdgshJCkoikVaHH6FFPAdoe3so1kKh+L34
2MO502qeSUdnmdd7NK+ML+oPTdrdewzQ9p6C6+uO1BG1Ze8gYcxDnG/5EfFNyJ3057pi5TMNWapa
e9+LF6UKs8G5rDPA+6d6NeFUZO2ZLpN1k9kT41u8Z2B3VJk4AuLUDPUZyEVJDCqSXIlUXOsXYu4g
KlqF+PeQFL6bjDwVO+jTTlxMcoKW5OARiJoEnAOaRGP50J9rQl3N+DGXNz3cHpWws4shFHOhQ06Q
arUYKZlctgfOuYS5grN6Q5K09wkhDMvPH0YNV/a9FoEzWPrUFd1MC966sWN+ljfmrSxCeFbrq9WX
8z5A9FZCBl9qITbHO6KUMSlqGSYu97NPqHE7VqRdLlP26J1ocDd2tIXcijxol0XtMdOIiTr9oyu6
tiChv6Eg/YI1Og6XFSRoth8E2xmaQnuzO83i4sOFaL+c8ikPbB6t+xEhx41NiKr7j+JyE5ZsuFTJ
WPcA4ugHsYIz0ckC7X8+j8TZdYAEGf7tyBQ91V2iUOkCKOpj1CndOnx5rL0BnVp4Xis81kO7fVj7
/VNNu5cCq4o3G+dfZhyzCmtQJQGN+LcCHkPM0haleQO8nwoPvRZCLnamkCcxWbtfSz5u03k0m86J
gKUH6yOBLDKBhg0lGSdTdYZbV8Y04R8nABdvaa8SboVRJ/e6QQxE6hWTMvCP+5nT45qZcVyHbCti
4ZDQuqYgmU/KJaJBJTnT1JKB0AxiPTRqu1cnl5BAh49HAefAWQaI4RcHvAMi5o1GTheLj4Y0l4G7
boY/KyuYXcGfD7KD7wLvLuUvtytMKZ9oCfHnEwfY3Na9ofrGgQUBRTlshN1tap8iYjJ/tcpzfXKD
eytEzlBJSJ+/eIsf+jsTpjSvO5HocpMS+J1MjwX4yKeM3csiUcg071B8KTmQSFA56ukBBN+mq1BH
QTlz/3pW6rwi6cVnYEh06RtP8okRouDg+MDE4Bbb9ArM60GORRH6ouFZSIUqHQnfDKOnqd3aJPPT
Y2qNLBEClkYdZVHCj4Jvjng2kRbVywdu0RHrwLbb2htcxsbnxal6uvCDIbWttwuk5vZvp3YffFr3
nblyYD2rk35WAf9/xlkYEH9szEmiXoAC1eFx3Ec0fnM6695K3HfyAzGuL0+09Z5e4jBB3DKZjHFF
3LMPSXblfSmynmMBYrsgwSCHEe9NvsFZHjhdxx0C7LRuvUD+f5CgwoMSipDqqY8EAm475S6LqAxj
qj2ZKZe/7wij+PLqoqkVXrtymZDnLVllG2c19sp8fdkNXO/B4FPwRFmaiQmtYqS1Wzk3nZbhzUtE
T+zcdxcoWakopQdYQO/Fr2T29Me+ieNqOi3i0USyuvQg1yaFBLdaGFM24gk0QzqlLst3XzHoeQ5j
M38Z64x3odBaKE1WBt+e70BZKTyL8MIyHCokrp6XnwNKWc8vCIqYcuEM75T50TdF3cW+F4LYhNy/
5DR4ZXbOSDzU02DYD09wAwryi8DbdaB1309iGfNlQruHfH6hnYvLrqUa5j3tC7XKHvxnhQeAJ7hN
RtSx/kGSty/zfyrhVdWTxZd2dQVcj0UDzQMANC2fUF1kCpxFC3ZALfFWBiQqgqi/UTd04knlDeFf
eWvSCw+Aqpk3pyFz53qdOICk7YXhZNVO17zbJlEW0f8uztNSOpCjFnyzJdiMzJjQCLHXdvXOg63d
fylUmS+xcyzkAopPjn/Rr6bja+ylydcuORbSnZKwJSw3LyiVa7+ssyw6j+2hf/p2F9dYXOhFAcGG
5Jb/PCKZpVgvZK3V3s+8ClNz/bo9iifiS96pHXjCXj7rbw2Q0YAnQGd2SWznrFAsyFlblJzR3MHE
WDiwfBquDFE2IhHTzPPF8+AfdbusqOji/CZoOIoBqpgsaOJKl3dRZFnfkTJAsje1Nvaz+nWwrOfv
/xctQcGGBHtPpUFH26Hg8wE5FPaErHZ+AgkrWy78a95Cm2LSyxTcWwVTkT5p9u0KHgIpxFIbLGNz
/q3pQnksuE4dZdRvijU5ptnptp9sZo/xosmYWbXhcyUiV6de9BxyQLSW78NtaS7VhaaG/SvPrbzP
mRhUO/i+ysLhTGb7FjZ3JCqt3viKL1mrFXX8WyZ6eO46y5aPeVHovdi9r89khPxrwVyvEa0C1x4s
ws/Yba6hACU5V62tIK3t6qXqJu2b2V0j8Ay2prI/Gx08mV+RRovTvj+A3yYkeqiFPSVNmdf4QqGw
AQ2iXOnIf7hDQOQBEhFvqnbcstyV2qgbcRHs2FknAsN3wrAgQGjrPOdcBIJboc+sQkNBxOVd32UI
tS4yJ2oyRdkEFTd7Tda25RAennPHeQHlh35cvxq3gjLwsDqqSdsVx+Fv/bwQQEpKP2Qqy1q7X96q
1o1nIuuzzVBGgPWZnFGzCGJ9HCwqwZNbwWXzYWkd274f5oP6kv+0mEjUPPJV/7DKywWtaTnp4+az
4X2ZabHf4X2eWZ1Gu68IMxKWlVu6UYMuQ+x6I2to213slO0axDWo1+HK20wlnAgjWLfBft9BNmFi
VIpgpYBy/Q753Gj5l46lQdXrG9GEhyWmaDenUVvAlmAMeL0yHjAPa0ISAA7MtDLy6iFqlZja4EDq
W8f9qGlmBtxhrRAC6C/DiqgxB8uSzGFrJN0bFijVA/DBrSDqATSQqSOodm39WTNWDn1HKCoH3NPc
WR4ADegn07vjJHZiutfzxm6t0z82t3PSD+qum9q7hwqQlaQ/t4arYPHOAzYaTDRo1EMeOdBbXTP3
wNKb8mh8XtqvYkopUztO2YM79qxskYm3/5CcngQpH0cHEM+GktbWqbNFhoD5HI/CO0Rak06fjojt
93XoVSKgjFihgLTAKLq6a29AS4ZLWnYWTw+cri7vKtLX6G+9c0zD+NkYwMjvZOKyJCtzKmBc6qTF
zJBN/rEPXZOypG2hyg5MKh1BND6OIZWKD9zKgbDNRUdnzIBHhwxobsG14RBeQUC2svUjbZ6CUMTB
f/lqELSdh9Cho6SMsbu/yW8A2PQJkOvMnWxRnsXNgpfUbSQ/o7mY0pU6axCPeYXn/B+k6A0QsE6o
s+rFFrxGE9BtIkols7x1Rsl/qTuwyxDwGcQyayR31b7Htt2XbIfdgTcDy9/FaoQvvy7U5YWq9Ib/
u/ScQBjprXvvz5dM2tv3TXn87jNfRaR5UjMDMQBIElElque55nvpf07529N/6SEDrM4CfiDoAXDi
Dr16okg0ODGkcQi1JIjYaTSiX7TY/f7cpokxGBUqO0wP+Hl6Du/LnjFzSrZIyPWm7WsFxSFLioOQ
qnxImBRc24MlID52q56mprX+MChV8uFjm9BcAvOpl5TDCgfgVxbuLF3OIWI7GjDG9TB0gbQAzzH9
otBwSQ6MCMmQzqa98phgYkzG9+2z3NziYmOGXicX/ma9NYKJpvjbFIby3yAo+RFCcAnYuRuC40qK
mVbh82bOpvkMgitNB478r8KwMU0I0GPvCxkrhtSWlGwdPJZWXjMDvTK0n5chRHHCicjjVtdbjkSu
pFOqdZ5lWKsBBtkCc3k9VNdr1pyDUYdPiIIbTBaxr3qospT2Y3eQvNPDLcKohbcjBY/hTAcijMFp
4txqfgWPn5bUgAYggiG1x+KqkG5q4M9XrgL4UHvEdE1VoSIOK9GmwnVERni6l+GSq56r6h2QTF2S
rstDyGC509Iu3xR2fx+qL2vaeyelQ1JEBNcd7/iJBzqO2ocV+8mlEnjbDVqkWddwQJumyYK3O9Dj
cI4gSuZOdekxvAj0+Dz0X3eBFOVvi4LGxBkQJxzGXSZ0iLm3UgtotEdLu/VTsfuFtLwawB6knwhn
2ifPW+6pmaTz1mLBqJ3PXwk+H/sb+oXcTfnQIKHEZGmiBtuJGGmk/IA9YrXRBruJ6QNvxSIBJjjN
F3hIPmqqMnfN2VCY7GsgDUNA9oHf2Pop0eOTGdNcccOPnOOah1rbNlmqWsphAW2PdYEdCOEohJLK
e/X0S8q6ppv4crIyTM6VrX/9hE38V3rMm4m8yUfnOi/VXh3lib9faH8YKHduqPDc0sH5lUAEoQEH
0QEIovcD/J6zyUl3bA+XAxGQIwjFhWpY6Cpw4Da8VOHZbQPSYWStf4ro6HWM/4KsfgXDCZv+hSyd
zbvrDEZ3oyMAb8cD/7KOMJWfLYRw5SG9+IwlNfGhwhvbvk/0jaC8THAg1dbo575SU3MFjmCoS5xo
4WNLmzXdhvo+KMRcEfYVpsFvFWox7vrkhMq5JI+Ztm9Z86P8VDqQOAbNk3JLGBs1ptMBS1si08Au
+DlIuj4TqQwZgeMjeRuRuUEFRniHxe8cM7MjPEuAB9Wtv7uI/Sf9M6IoKsiDEWKI4OrHZ2liARZt
2OhkIEijIEZEgGYh9sy+Gecxjmam0r8LB8WQva+p1SnXgPMyssBdJymQi9rDz7QYqEIxXXgqFyPq
+TF17DPmlNwMiE6fdcCOMy3rFpq5mURZqvWDc7y56JLx4FGg07JhnTTRTCFT4ZuDRn4MsEvUsKbc
HBHFnxZpgKjc/VO/Kh2TFwooC5Zq9UgajaNlCv2SXuY67ZYYB9bLJIqABWxshzDklVDAwCOEOABM
qs+Iy9rE6m3qIjj+b+KB8OSpsVTLH+WBqFGg1mhOYRbQmNQY4Sixe+WMRdi4gZUAOAL/4+ik2Z11
LqpN+qDtZVRY+q2owSrlcTUxHHPnr1puCdp5E7djyHWYsFfYk2scnkqcb38GtQ78QdYdy/TB+tGI
PYeexCLJfeu7S+40SuTwKrU98f4sf1eBk8e39qy5bb5BP5EUPATj91OSaEsO/gftTGGSB2rSNE2H
UW/HO7HX5puYQpsNXHoY9serQ8Qzk3ISLmyMEMzsYu6jDIKOVLNga0xkNtcHzNL9m9Plq0Q52Q48
SHEo8IpXaxGwDaXZ6o3QqIR/Ck3d9NDm1CKSPfXyWccOZa8RGnFju5wjYpGOL1jGf1PMCXuwlG3p
aL9Gwqf/GjJkDcotARdIu7OYfwlqMrpR977yOMmvBhqY9nEvRSSi1XzubiCSMEORFOj94mD02elp
EbvEtMsVlQrogM5+U0lH3VEuYEm86z8uCp4yj5q64duDMQLee4ADdeZ0uQIBzQPLAVeb+lFlAf4D
qbQn5tM2P8so8E7NrXkwPMzI1SYHl14m/sUGmdBGtiiFWh3OqiWQDNTaWTGso+nnF0E6wyPj2iyB
U8HfGzroV4MK87ddHF4jbriPFHhOwdArpR+V+Io0NPqc481rx3rfm12ZYEQge86kFi9od5NXtXBg
enOlcjT0w61U/YhEBKAkmyCrcZPRAkvZPBAmA//LTlhmosGsk7BbWtl+YHqf4KrCC850ZtelZVeZ
kfTzjY2FaH6XbtAgXoK76LRaasosnt6jazIBlV3uul9TqGTgUIs/Qk4T1gmNh0HGSery50n2SIJb
sLUSAzSOwYeDozn8v2yXFu9PECU+inQkKiAd1qucczujlAqSnrDFoA/Koht9Vhj/KTF8gQfovBBH
Qx7bYBYY+gzRKrypIY1nb5p78oPRTLLK0oyRHCtBvm/ni78TJVInLcjy4ubfyKZOa3QKLMmVsC4Q
x5TmCC3nGxWSuCzuuSEjPhD7hs6mUc5oUnbN7rSrMmvz6gAiZ4SAZ0Xkc+MXlJQwPkexWMiSB79Y
rUmfm2v3R0JTIU0HjEZdqfXWdcrfUkVXkJkFg7bYJpf5Zr5mu1sdVo6ExIVO/wJTPt3/cuIJuxUh
chOnYw3tC9YfECLWEjZtWvc5JrpPedAAGWGMXhdR+s0VmofIrabEUZ8lGL0UlD/04fmncJ5qs1kp
aMzJZp3W8vaYD2vKdeqpdFEY46saTpPI9R5QVUKTXUbsZ9B1Llslts6AKr8F0pzVhCBwap84/Gy+
IuydzPrpaw807lwogCEaDnQTXyZKpUShQVpnZHh/Z2JXGvrBXdFIobB4WSxBn0Kb8ldfHqeHS6yu
+F7I7YANrYvIkIJKO/yPqzcJ2v4CIAO6bHVVeCvB2xs4bv/3ENlM1lmtvZafRErOIVxg6z2VaupE
ggjLnigd0PUrkVW1s/Hwhqm+lHqoWBPXYQcS6QXSjfH40uFKLKPxz0WQIeZq4LjZKmdI7N+8Pg78
5/dr+nizStm18+CQPvSmnkD5FcDs/mWHJb0dwEOrFLex7TlCtnxHgkZYx4P35rdCucb4D6kRBLrP
xgvOP396UXlTeTvYY5qtnzbWRBuHwhFi3ZpG8hv89QOH7MgvtBY36gfo1YaV8jibg5hmq+FHbCQS
W/22hIRPq9VpJHaLVsAy0ie9RUSBmArSGxZHSuE9h0HV49VQctSSldwybk7eBPEWxfyvO2j/7I7v
JUJ1zQ/t8d1nuIugSNDjhgmOD1OrNB+REzZy8uY9uY+mUIrohLJmkdpttt3xrAfZPN4B16fP2YL+
RqpQY1OQMnO+Sk1NH/M7BxxZECajjmuNIooHQ8L15+UHIOs9EE2DN4ZOTjFtE9RlHqWsJ5WvTBm8
m4RbQ6THGl0VbfNJFAuAgAJP9a+jKmXQ0PUxluRKN/WOHInV35Plopl4dNdf1ta+G1KI+lZAJgCH
7S6IsCe68jyzO+0MEBikCEY0SNqfegzbjoglVRklSBNJH2TeeYVxMykSP6tIo+Ldmve43uAYz9WK
c1/UuVpv1ZKbSKBO607iuLkqMabPPbCZogNcGIIM8mymoF/fowNzv9JmbZGseofT5y2/CWO/ZxNn
Vc4M+KdkgnEoYZC9pnUZYgLJl6oZOUEnCanZyixvgQXlz1JFkzfmGrrPJFkc4hONXswQN6PwmNtJ
VxpekQLpHvlvywwIOb7lp5J2s3dyK6dlZi8QJmWNiRzdF/2lutDRTlAeIl2LxmEMtB/3QrHl+lwX
Kax/7TpQMyh1G67+qZkCzVz3NVED5/25VCFJFcex0f8JiO5bbbghj7C0JogWcXosgzgx89OqHzpt
aDvbyWBPJ+eGyXfhhHXn6MI3z1Bcc5Y8C6VWN/DUF4u0Qg5juDNw/WnHvD+92Un8CSOYR1e7VN6g
FwuMzdlGEcLtaZ2n0pLb5LWsTQykbVq6TTspTDKaNvrm60X0BpmuSvze8FX/nnDggS694ktSL2an
Ipr35y1XeT8uvRzKRKq+fgT8qcBrQ3IUHxFtWeE5T71B7QczuD/lCRj39LcUHIdI8KNzKNzZSzhh
9HKZ/yqMcHUzdA/biJM7kzZiWiS4Mg3rrFq3PWkPi/zZZUSmb6Llis1uvO6PWQ73wo/eFB7Rxy/6
k2rbbs0A/TUm8PljGKGOw4BBsZWYJ4UeeR1TzREM+DAas/BuOjmYNX+J3dSl4qyvfo4eP/megIcv
WX1nrte8lYBBkGDQ7tfWeH8QSyfn2NDYAcqkdKxw3CJXsphg19jCv0Z16+t0G9JnRymaisr+uFPf
gd+2OgYdHKBH9h6QtK7ZGC43G8aetmTzVLVCoSwMTDZOEPxfksApeASGHPqiSIfXTxaRIT7N6ueY
GXeSkj429xnLpJsHZIeIV+wBZv4HpmPDu2OD9/5DMvbijTIJBLZFShaL9Y9ylclHGW9XGUjMtIRa
ggjrTqTo918/OE462LBkfXtVZhwK/4OP0GplfFeUvvIoQEyttUco8QntKaHb8/devNciEp1pMrak
hvF8Bu8kwSHMwBD2FLq6XQSNrbDiarIw8sfL5FZgEL+bAoOK08Xdnpkrkn1e+tIMMKxrgEUBukAk
Y6mSpQmPVSvvw1YmplZ+b/HGaGAZgBad1tVuLYn8w3fiLIixRbHpd7+PE5Z3MyU1mvAmrhgwT0v3
1CHmec/f58fL9BLi4oHfYvMIZNRGPhswfSFmjwUZ4VFKShf8ioad+X+jpm0Uqg1ySbW4ZYk1dLXD
Yp6rH/B+CKWsk71O5riaEVyQ7YTbaNiYv3Yxf8KfSe+4Lbxw6kjyQD+UEY1KrWwEJQkenF11mnIo
cDJ4n2t3V9LzHhNsVjMMvu2htbdzyYnfhpTc7K8jCw3fBtIDo1cyx2z5lvDCvULYRBFM0NhJ8XPe
J8VoCqUuihdqEZ9BjBD8OJlvXvXLLBvyoO4EDZJ0WnDe+GzpUlCb+gx7DaPzFZ7velp4snSmaalV
P506ga1u1IMwYk7d/5SszqsEl+lRbJXRjpq8TIHZuOxRP4FqNsR2VzD9hfmCFM8Atv42h0byCMnO
Smg/VYkrM1zGXh1XkDvf5lTsoIk5UvDh/sCPdwpRfwmuqCv6C/dSx4N8KtVCa2HQcfbSR68newk/
odX9/WumaLiv5trB/eXma9YAV9E3juWaANBvtNkpY70ixkf3GoK/Ls0k4ngGV3eUUoDur46JT7I6
hDUf38XYnwrJjEgEAwkRTZSLqJ45Sp2OdYA0X0gAPMpDhfljJTuZ4SNim3LnPP4jJCdPOcO+rQnD
qLzdLOHoPuqVWDOFnRsPzEFOEb0WJ3KVXxCkJ1nLZNy+SJK708+jj6NkoXQsLMFK5rnWy1PfPpsC
pGQnOM+r6OwZ3CTcqpTGZjW1hVqDS2AYzumG09NkmE0bu/9rJhIlRLZri/1cZmZo5VKU8mvnUX2T
6lnzg3G20WL+dvUH6emQhMwPF0I0oeMXuFUWGl6NoY56RbrSDS3Thi1gAIhliUeRlpyb3cEfCWqn
LKdKruIdpYSDzsdSSoSRnPucyxmzfM5c+X45JCKO/t1GOxWVTci6orQ7autmGuzeXGbi3S21a2Nh
1Oe01Z6gzmSZ2vAMHcOnQ1Wxdq4DJP8xt+BiCiici9JUFOguVCAbr9Z8erievC4Nxn5ME5bE8ZK5
VMC1sU6aPK3ZJWV2QTc4C3+2P1qiL95EFL5xeEkht/NcW2iC1iMI+0g4eG2MXEXpktDCyxmSjatq
EFdgWCXJC5xXHUxfS2+lEQnoaFNpUiOJ5WNcUufKBj3H4d4Wjymu7Ca7sAEd5K4Fx73Z6DEbutzu
1KYWyhNPLMW48fX7ID8hwiL5gHGmj4v8NKAd5+X1pn0MTMHmEeV55ZJzrHSq4hezDaaZS1OSmwRx
whrWuqNK0A0/Ga/HV+t6n15IHJrTL/Z4Czak/Uz32nykxVih49oWteWHPlIrED6IUTiz5NpoBJOz
8hEfkhVjrOdJbtqHRFfAp35Dk20z9sZzLx0AgksKGRroEAHMKThj79NFHCL24OywVlpxj9Q9CKkz
qS20eUAQU5YqA16YWmM+sGH/uII7+39lFaFxRdUDGIlUHs3iuY0oKrOMPqC4Wr6wADWr+sXZ750w
aJt7uO6gR7SpJKPetwltGLc9Mdyp2FDq4uQ/gONDudEaQ2SOitoUrx6Mmw4Z2Q0fGsKQt101u1Pr
eQtgJY69YPIGITync6J+ZZYw6fMmIyGbHFpx8wAdWo0XTJ3cs0QzQiAA8mbmN1SeTTel1OUFHxzo
yQn9f/fZgyU6aPADqg6O7OJwLVzIXFPtSNBzP+y5Y6upXUscSd5b+v1ySoPEd0bAczs+UqCcXq1r
I0+KEK/DcDuBFOoKyy+BimhX75bOReOT1CxZludP4s5r7OebTW5dck+errPhJ+3+0JtRhZ79e3mo
a0TrWWbIdWBZJicedNKXmb/yYaPpyvMahDkKHKs4qWPFUhQm3uM/UW2nEM3Y7Oi1iY4D703aCHc1
N1oE42F2P/Ev6/4+WCMNAtMWVsJYdS3+r27awAvLRM2ICrDYXkImfwBsewOxK88ZptwMA3J4qMDF
xj5P/AKpT6NDo+Z1oab56vu79JgTUk6uW7eL8gOJ68VkmOu0MWB+HsnnqpVik9uWvnzfwppMooQl
g3p655XCEaFN0hHMCyKCT81MktwxmdfVdO2KB51l7sEs8I16F2031zTAOP8xv+MnNkTl4JP/9to7
8nWOoNCWbKNSX3qjpTRtBEo28LNeum0QCljuJCgJrZYD7MYq0v3vV88l+ZfJm11qX++RuJKPI9c7
YupOUoUmtIVi8l1DwRB5grz9T/rHWf0tXr2YXEfUJBmut3KTCTCoUgfePVP6AT6qTSh7n+B5a27K
JnAPaNk7KsBZoTX/3PwySs7QYDAx3LOAeRZHmWlO5dweIxkEZYCyDbnzc8vhpekR0VsgEMvoX1ka
ZZ1zqW0Akvu9Z7Axtd1d2hEYy0A4STbMjmGv123QQSPli3Tq7ibYmxddPpmVO0734acgnZFSFgxx
V+x1siz0OdCxk0In5MC13TUo1KHBDGkwmbOxRVL2+86b4ybQgtUdGVbr6IQmw1LCvDPYKv+PHkBt
9v2rZ0UCGmrwTK2NYKB2RoJIv92MJmKUxcm3syH1pBFmjW745UittARusDqce856+S81yJFpje57
hR4P4AnhYghwHV9ll/ySekazJhg3KoRKf8UJUxhJKn6sQv4Zi3ax+FjB0El0zHEVZd5o6FJ+1zz1
/4knl2xxzpwORSly2FU9lJX3nRQ1nxjkyN9FR8le2qVBlbdR/F+GUh5PBKhF1UeTdExFpUqc/+HD
dtYV3FOw2GfclTQ/JZLl9/FHM58bUtN9zCLyH6CX0hNAOskwYsLmlBxiFLXp1U6xeMWuNhq4K6VS
IPs29D7oCP9euumkURFgPj4m/zsNkK89S+c/+IwBGrqIddABOlzjfBYm91xuVoD9djTfHtzhUrzR
Vk3R4h3jKhYI9zOXfRNSmT+17PGDHp1SiAqGV7kFCQxfwj3s2ckFKF/stiKttDBf1elN7K2o+IM2
zafhPwtKSEhYwWjj7RGkz2XYEdFAXLmaxjKdQTtInUDlgAmM5z76o7ZT9Js0aBHbf49yHTIvqXQf
vxkABHflWQUuOk/wvxlWyJFGvPbYjz98++TL5uGrPmcXOMje1CD6wynfp2K+yq/Nh6PjT1IJCfE3
0gKqLOqEHicJULrMVTq9SztlvUEyocjOCGa24CHSBGflKAxDFGG3BZ+ztO4O6Lj98uWI2GlvwuBl
bhU4pOVTtc+cEbXV/3W9ntsjYXTw042JntsTo18TM/CSaoPSFYrq0Ltl5v+xVWPOrmbuw06a20WF
zsTMyerCSBwwlvRFI4R2tq8aL4CP+PbPfy4v+C7rWXV+A68MFxbL1e+sovgRuUiX1Oi8mdyZLgIg
7xKPFxQxT3NMFAcmoeiPX9krp6HG7rGzyaTGu79UjuT77QGXN58qPWV6Ypp6kJjY1aWXyEjGPwr3
XJC5ViwoyEanKThjjcaauYJewpU4bJ/FKPa3QiHtldbRUQUb0kbSLEQtxJ0Ibj9OMibg9sSkTaG5
np+yPOYO1+fikZsO205wMnAA7TbAr5aOg181zSfCZZYfrlLxFdHsZKjpIaM4tKBoxlKLP71pW82B
8WQDP2Nq8ejac2lmnhRNdeDfbmlso6PW5i7lHCT9AyuQJFY+RxwjX1KMcLh3sTja24E448sBCl75
FtFJD95o3keLIX/tR/8bJwYf6ii+sH7rb2qVraf/nVHr9WRjGjvjd8v4d18e1msC6MPCwklQF/af
MDia27p1B839h05IvCANXR4mAlHbHMyfNfEy994vOXz7bTsgYUINISVitdXfY85VBNVlyeugV3KK
nb1PUJWAFN0KAw2Lr2xVMXmyg7ODRUIaA+eFXG36igXfKtyb/IkxULeRIH0/ehsYAx/i+dAyUhAj
UMK0arFreuAhvHNcsxUFSCWVTENf63M9DssopLa7pgKkVxZSDU2ybq+RagdBamQ2hfFj9N3YRlpG
xsp1k7IvimtEW3yxQ5rHiObo0e1vIv9yprhY4EDLweuBwDGHoCL9kQV6CeWLqr3pJNODQWfY6+Rr
6DwwNoNo6U39bH5DEhaE4ccIWMoKEGoyuZ4hiTY4Nor7+eywsDIe5TX8FCs1R2a8sYE9NodUbFIN
Cmb+qKL4IROviBE2TWYlxhJLtIcrI6ywxtv6Jx6z5Ei2ZOVRh84ocp0c46S30zXkH15uCDxWGyZU
Y8xTkKTrvIkSJufNahg/zN0GOav1p/DW9sUr3KSbNo8qhafUcRI3vOw4p5+e2Nr7awzS7bPXtgXg
VpwCSq80pfSz22deV/wnMPcNounY9AG6aUJcJnopv1DgNAd3a4SbnF1fs+53uKf3VhcFMe+rTlZs
70lR1+D61BkYif4+lsHo3g+/DWR6s0d+zzCuFcGJOOBk+QBhvZXhEKddt+IuUdOkE8Ua654nfTMd
kPM5Wx1vdtKqoGLwtkmqJSrw6JzUSkYLP0rhpV6CuRCLKRQCIKExkhz2rQiuxEaIjUD/1Gn5H7G7
D7taetK6F3GMnZWgemWPlkY3qZB4Zyg70bxeu1HXWGCn+524g3hDVrKnCJqnQqDuaY2gReePItUK
hnPzf4FsO155duiigtgZcY7CcIVuwcd1Y8v89s/qZTodP9+JYUrpPKSAG6w01Jdt8l+8Nj6ATWK8
CzAzzal9cyFIGdzPY0V9cEVNgaLQzbxSW5D/bhfUXURcNmj7fQ0dQuS+g9uQOPGKiLlexwnEOVR6
zPuOCOuFA5zjjqSSXblrsDh3uQ1xtUT1aKf1ihccVjcuFvaHFnUzyMGBIWoYxFhA4LAo4wmYkgwq
4ZEEK1z2YpjF6MI/6/6QoS3C2pb3/EKrEcgjoRoGlrDK/w6HkNK2+nYIzCCQs/dTFTHw1YrBuoFX
rjkjDWQlpYz0z2Mnu/i6lKeKjDAvDIpzQrhW2nhM/Zpkd7BiOhbYXTNkHQb/TTGx+DBkZUKOz179
tlfvmp5gUv00hmP775s+v9MXIbtHKhMDeAWsS/Qz5So9DdKlMTbTNalguv9y8g1g5QY7wJvHZBKY
ihY1G/NrFmkyUgEWDpjrRSp/Gcp/CqQJsdXb6RlJXJbLlFetfDrVKWFLOgayRc4rhMIESrKU2log
BXg/XyhTjH6YQi8FUrS5OhAzBjUdE+aviTnuDpcsxCbL1rQb0SeNMz4/ZAlf51L+6/TzOlCOqLBM
SsIcosPq8f8JNvmytTf0nskgXF0Qbkp1GvTw6MpVt1NeqobmCS2s8MO1XJel+quiWsNXMGUM7dG1
hGW4mCffGmjOmxXZZA5udoO38WgM0evp9wJKPV3OVL2YDjhlLcYZC2R7Y28b8V1DqowpT3YOZi6M
hVWu9D1eX4s2R8TkxbrrRtVa9hxY4JivBrtk4shiEggZERwN4gF00kgf2282bm5Zzc84o9mCs1xd
gWPT3Lu07kbYkSwa/LpxTwTrLAWv7RvM+vOHoLkzRNVxQO0NFvfN0Z571WUpMZ1pGsqK3o0Oebzl
hlj1ISB68uO5wLCOsKeCgB+6N1hBYs+mm19J2s1D7Heqb16xdGEPvAZ6a1VRxm7LGSN3pykpnfc6
zaNFQZO8z1KsraSU4wjh+GGALvcURSLTwYfA9R8lV1azQpAGbKi1r254eaS4W6D4W/NZ0rwu5ZeI
3I9Yozp6in0cG2OPj6QK+1umeNhDQiBpWjpxAi9V3ZHSy2bHbcard1Tcm8NnyDtjwTNwkSaZ4F4H
VkGguJ2ovPlNAvRKgoNcYdD3Atrokf69lL8Tc6emlfgXU8beLg3liejgomP84AkUarkZYE4eqbw4
/35O2H8mD/39fHAWRsKvVJMSY+6QbeBeg4wIBBUiZxqLqp4w8MG12CsHPWGFmdmHcIYXzXG3+i8w
WCbjfU7eEtrIMz3TgZkeSy07MXWyvChaYMq4Sn2RgThshpP08beADfA7A/RtaHoXVBTLV4Ba0rB4
zrttNLoOpCHWjDKrfy3kOQ7awLbCEJNPmyisaiF9JkqkreGEiHN1BKqfCKnoZf0Z5pcdLNZnfYaW
EmvqLdiMAcrFV3jt/p7GJGQoUPm0qNVRcrxOB9IMKSVQFSu540rWWoxu33jKBEZDREm9K5DddOmn
a1ftyztgjc25OqF2te6iSK9kbEUrqHIn52cboALjIBSQM2wES2AVGNs47/5kDR6CR6nFvqyDW28l
n8vaQDKF1t2TGSu+dliU/Ir3TVrOAh1TQuI9A3tzkTXyi27Cl5Kb2z+P7bukh0tzQwHMO3ceK8+b
0aD2JjnzyE6TiNbXi8LlK3spachj0RNVQM1Mv1iC9xP7FEgnsXONnq9Y3uJJlM9xfqNfbiYfCCC1
I4V0xX4jQP2zPVtwLGuw7hO+VNvzGjp4x9pAIwdgyIbd99XrCkQAc46HTpZ7PSFnaxW3LcRNUf41
axgktObzfpqiCy1faNn8M+usbleBJTy9meidCdigUVEVwoOqPvwZWkERI/LCIBvbPe5OzT7RUhJt
p31nYT7MWQXYkZ2Y588QQJMiel4ebQdQEOc3d8pkBRqiR0zfRpzDnVp/jpaaviwl1aSA/uSJOwfv
Qn1+KqU3gknC/W3RE2Es0hl28DriSa/gcGefv0IAxnhhAxJp5MaUg/j6XodMHhPEU3OTO6QKG1h/
vuIE4BK+rUQK3eHck5JE2eNs4/6MO98eFTTdsjLk3mL9iJnlrSOz5jeZd7iFCgbn5x5HJ+E4DecT
OQpOpU4TukbI8vo0E07O+EOuVqMv/aSPHj7Yki8+1z5J79sF9Ne2+nRnZr3+nFeGf6NQ/ObjlWti
33u+Q9DDdFwe3wlHqzJC9U1MUMogvECxFl9CYeQzqf1hQj+iz32RbuwkmWH4TEsu1sQEG47ilEJ7
y98ajAX8MCO5O/p7fvvPjIPkasJtXyBO74ZUn4EP7pl8u8RvHiIQ12yPc4d+sxlnzqTf2kwu3au6
brIaZpckcML8mmDZcUeAQhextDoCAg9Yl4AJf3yhTFpvln6gNcQNys63i9U4mANEI0slN2Lli0D6
3p4+uqV5q4d5dOrUhu/n07DxJHG9XZkJmh/0qOzidY6Rk07kjR1r0GgfaPZnwbk07Or2QHym9SNb
TlDCLL5YpHjQ2WXiz9NaRtpsQhdoNs8weerAQx+4fUvgGU57xT48617J2SlYiVLxJylJvsZuWs0Y
FGsw7MIt7C8aExoD5k39SCwZCs/SMcgoQuw+AM1gBX7qtm6wKTEFl5tDFXMxDyxeG6KoWRmHUFzV
JU8lKFI8r8xxnkLKhuyu0OBXmOPB/UNNNNk1RG2TcYAcM1ep+B00vOfsUBzF3AFtmNfvBTvRuh63
SCsnRs08M5z9ae0MhYBiCL3oxAkzEqo7k+jr7d3rSheMLXgFnQ2x8lTxtkOcyuf56tomMqTHnGrG
Y2iJCCPq/Y9VemGyfv/yWXf/T6MTKFSX5hfRR1Ba4uknzuAirLe19H5hMq83Ngd7uyLn4pm/ILFJ
ZPp2jCLtF9hgVRIK+H5LIFY68IJAu1BO9Rl7i2KVHOZpccJTsSEZ2XKQ87/08Bs4jRGu865DX5c5
hv43tRIim7lLmeYmRPRZyelRldjkwJmwDAvmTU+jaY12RQtsOV9145B86NyNioslcYS9VhMqQFyz
Kjo+bFI7591Z37fCp1gilsGymZly1YIWTmBhy5vqbQwA85mXk7TXSfDi9WJDKKWokjOefNXZKroE
5bn8+67hw1tD8bJb24R9PxukMWCgmaL8eNpcjrFEcE9kKEHjuakQpEYT30+MncFt8sQs2r3LYIv8
CcMQg19bXW7FUCSXJXMKi8eg9t39Y2Aqe960+/32/FXlXYy/lk/BjJheawdbjzu3idvm3EzvuOR4
kcIgwIFk0qj9VjdadUZtDMgD+/JAJnB3sI2FgtDGcucx/JwPz1MecqfASa5zgrteviEaeMxTUmKZ
AjDXIz2LjbVx0tNDYoKhuhGZ4WV9n5KSfKXv8qxbfIQ6mEn6EQ9/f9Vmkfc2zqoOo3mIFxMD3CFm
HqVp3r7ljtYphhqHAPA2PP1amx06iF1IieFzQf2lMMSzdK9iANdWqQill/+KO1Wue/NclDAPoPvw
fWWO9Bn3nMXlYPMFix7K1cLvzWOLrEJ07qeXhcAdkbWJKq5/AYQmzpGThwGXLu99Q5IAiLUTxG3W
FDFAkbgJwUu0nn8bg2X1h7+W8l4KXv4/qgm8oHCPv6cjQcJ/LSxfflfEk7i5LL4Uc+CjRzGnCr3W
/+G2ztkym2WXIc+oa/N0WVymX/hdtzajjvMEyFxuACDCM2ugUys49mG/rmDqDwLna6rlXA8d70d+
IakfnlTNW/Y+97QnZuBx89EgRTW7zxorBUu8OQk9AlrAtl5EbpFLcjNM0sb1DVjlO6iRzdPp3C6O
OfuHF2jdzqorGdn0diP+Q8UzmAAQ/Xr3I65178dETyRiSlJWjESEx4iR5UI+M9xNNhMUYBHTYNdD
GH1P2vpWb9lQ1JpYUagLDJeEiOhOLQYLcstMpnrYtgyfw+KeeT3RwFfBWY9XROKK/2IgpjrLd1QH
V5ziwPU8TRsKgLbcwOl1WjCssa1mAKYhxzzq2T+1WMPArM3OEL4AnVj96CI+agMqj0lVEGP2GoAg
NFfqVMt54yzRh2D/vLc7iad7/8HjMY68eaAkwdJDGShpM4x8m6gtZsl7OrOrodplxhhaPbaPt5yi
7chxtwUmhILWWhzEwXtr6PGHhXfuprzQ0QJ6TF2+UYwzdiKu1/bWsxfwfjFFK1J1bbfEzhtMelQX
x3Pg6RsLx8dWzDJRF27AFEoJAInVmE1PkvK0r2x/uUGW5Q7F0o8OesaF0zzocTIWPuqUsexQyHsm
en8czaCnP41wAT1O4Iqd2TlWvtdzGSWSuTzy+9fNanIwv9lN1Y9ALyAjZp/+vjWsfmW7D95phC35
LjfXPtrAZXUwSMOSOxqoIQO2JQVBX6ex3Y/3nPCqDMsxjau33WvW927Lfk1gHcs8QJC2jCQxxJeP
szOD5v6uHybjfJU3NF0UUhOOKSASnUp57q/Gj8fULtNiqRulJsNQw+kGg8ImcQtfWeOkTvJDqbUd
c3EDl7Vn2fR9/tLMwe8PUY/zWggaGsBy/yEXBI8s3H9FWrFH8ODjqlrUpnM1XvKOaIlOjDPtd0p/
s5WFOS47WRuhhozSwl+5TR0JUvOEwreEQq7k+c60XYvx6fmwLPcPsOpvuPs3kYZ0/p4YwbZDdxje
64gtVg9FiScknMTT+qCB0OsQOEoD+dRNct27Bmpo1iOVzg5Grb+XvWOVrBQiGzlsmKfnbLN2NCPL
A4TNaVnhtGBhUNwghOnHIhLM5UXVCZbHnz99XHLhtP26zm1JJwfNq6oEfJJEMk9dOulzIFDFhyjB
EipjghHmDq7gj5F0rj9bW4EZJY71C2RLUdbe3P/bCrmPjI00x/HFCY1xu/JlLlnPWA2SS4cjyIvO
YvzL1123jnHuopcLylPnI6BjkdCVq87VwETeb93q2SHFja7aozM60hUYwIdSKDZhgDdezpOQuLG1
aVH59BMY7/xJI7CJu9D9xJ5nGmxQBNvdfTUzXf8F7BV+FFqf985QSD9gz99ry9Q9TyoBBIF+TeQ3
J+wIc674le0Xukf3ok0rClcna6dxZLiDa+9FxeI7GeNqqCYJXwx6V7RzX2Vd10ZigjbFdfZAKHxd
v8kI06bCXohTxxp5wCvy/GeOW4XIajOPlL/mH7wRyCJxHGJ33MvV5Zgb2QvpsiXT4/48FsA65IV2
nhr1B0KE+XqV77bsb00zfBHbJ9lYCKQChZYYiDkFjoZCQcoK1Pgs0zsL8KpMjXoBN/kwDs3eOCxY
GNh3Y04N/4KeDl94vBAviwnB+GYwqLQ9zP/lEfo3gO+HXSNwvPIRrSsDxrOCSefporn+dxEU1Soo
+XYZ8S2H3JzEFy7n2+swR9aeI1m6c+UXEcaQjIwqqJSdkdlITJqB2DpIm0OIVYasKtHS6SNW43WJ
82dIsBHJE3P46RsfOO/Sw563pkWX7y/F6zwgq+SkIwq3IPimS10L7I0J8xb+T3yTk9qgP35ZyV4P
64DbJW2SuZQN1RApfJ5v33QLXkv5WuCFT2CgPFTcoP8eLkMeFY/H1O0rcF4rGfx3Inan2YhozmC6
Uu0HMIJbffO0Nttb/XLID2lACwwIoU++N+a0YaLVVYC0wURGDjXIDp+NdIrhqVBk50dfIz4YVrM+
MQ1RAzoZsoc4lBYqCtHcXD5dLThe3+9HXAAD7Se3onPhwz0F6Y1plymAq7fmha27hVBj4bg+rzdj
QfU08byfrlwsB77Ii3XJsx7sZrTJ6nTSb8GvQxI4uAsTP3jhKHMfyD099ix9cHvFQ1OTqfUkd24O
AdXirWzxNkaHnuXzfRziTyVi8Az+lGKIuL9KcZVPBy4Lo2scfstyc7jI1v7Qklf3cKEQ/9xEZrWB
SoAyAmMWdKEn5M+6p9bXK7p2TZQlprMq/9/duHA/gUqed8KXU9MEJib8xYwycL06ar+wJZDDoGhq
jbjQKY+EEE/BDDn3gdlnZnmLKe4CmnxI9eRMDliAU2weApkSExGWAgJI4wbcWTpVAjaHegAtYp3F
eXKQuyrAXXNA5MhlslW9xBa9HySTSxwrHa/uK29wFZ0tMxISyyHQU5m5V4TtUj9tSJN9svZd0GpB
UkyYl8wOOyUO8eM6QOGnxe7QcQ+lQ4gbFKKyOOWg5sMPcGq6i2KsnxmbcAer2KQik1Qp3sI7zsxA
3/ZiptTnxLhuV5jfrQYjjgdeiqMkOYxbc3g9bnQLNPN5+wmwn1kAOxFY1OZw2uViJUNYqxDVBhxp
sDAt52xf4Ox/UrIhMfTmwkgY3CWdNJ0bGO0vfwrjQFs0x6kLv2QV1ZDLmuqveAykLCa8Tvkvv6Qw
ZkZ9rclqtikIh+0DDspypbuTy9h6iWjU1jVXthvJS68y2g9dcGBV+ONjCSbK3J8gz0K2KkhcHWHq
O8qpE9GQeE6RZem0P8iMutTQmNSZUD2KMesnQEgVZlyVoMhyEgnoxDN5qiuysm/kyTNZZYEOTvS+
YfK/sj7LJcw/gZfhy8uv/EKzJqWX1ivtcZoRywzU8nbOG01GE58YPqgbGD7/bzaJGTrA1492mWuy
P0/6uYnHUPhgUcGKIJgoqsqGgFTWGyLfuMsw1Nm05eJlkW/Xcz8WjhqGvArol8vfN8VIL2/tadC5
RjrserEklkWiw62rf4L028Bt0q3e2zgnFWqAygCioioDIAnuQ0av8eJfzcboIudYIzx5b7yP7WqQ
lDE2rBoq7/BWSLdx/eJ3gZsm1pVVPD8S074SGrehTYgBGQX3KjNa9pKJu2YGiYzSWpr+TDDPhF7r
LoG59oLmgVZ2viDYJNAz2umzNz1BuwNFGjoDz/SaCJRepAZz7dyJBX63W++sPBGZkNN5snPRLufl
xL6vQ02cZ7z2pqW0aVRzsDbUK7VkdIJDQdZvH8w8H0dfy5eVwWBJAOT15EZxhRliC6OmN8jr+PSN
Z6V9RK61NIPVXhqSB8pJ3yZnd2nLU8TVk9wsoBAaHxii5qyC0dnGtNil+AV938HwVGEWi06zfgdU
TgHzLrL/o+OrtxZU37Ihrvr2m/YlhXYVNkw5Ozsm6rr3zyzYrF2tEo5oqJznKz8RSg1etBjchrwM
13rR9QjhCG7WxZhAHlUSk+7EjItNFcPObFmvfJVHLoGPszQZGLz3ouxMivG2I/FeG+gjeBPtot9P
t5/95NU2v8yPNWXovkXcJ6kdr02Pr3ecmMSuO1w2nR5ln7+TqYsA2ep+mYCqGCY+8tNIDUAen1Nz
SF2nyoKh/bXxAlqpqYSPtHCBpz32Bt+s5igMf5id7A0fdKT1BHjMNAYN/O3o+tAXGDDNkiTzbYYa
9UMxX5UYNKuC22kovUoUUK/nSWmpUD9Mbt82L1S63nhP7YX+cmzh+zWbveyLlraLeAsiR7gGhFAL
J1lszKGGGOQHlHI/Zth/oS6gDHKDStmawNQJNYNa7Td+PBnNmFMXfnUxLwedADvOd0isTY+/Klp5
+QuVAf+NWlC3HT76mLDDsfzvn7B5xaFeukKP+yCfEayuqJJam2tI0UJqApG45/CtGkJeZPivvHdW
PN8cnewN9RD4MtSeSd2lhz+/vcvtkoA1kDpTjxUWjiah5j2MUOI/V1uv9V/KPNrR3w4VJxSpCvOo
xy+pa61feOOVz3fc4jsQMtUofLU8ezPM6wsKR6jh6wxhSWACsXkSYrG+X7moYAN27jgS3eBMit8U
uLjN3nDPkKwSJCA4Bfx0BXuLcvklU5ot3N77Qg7RTwYLC6WVYhh7Hui+WICyKw4ofwqFZimtwSeA
5MUEDi22nW75/YjtZ6Iw3YYkgAL3h/egc+/k/MFijza8jfA83bQj18bMN2AhDxYgSmWupkRdt6kF
HiWou/2dbnWe3aS47sGz91Fx4Csh3KZqjY8clM3cyNoTrJLv9Z9nScsG2JDkhRoxHrWQzKVKfVMe
jlIYVUk+0Znnu8jP5W7Dxz3ozvdf/8hk4yiFT7hzu7frplzMIsDQVZ6uv9gbopdR8N9gyyCcg0Lh
ishlecqRQtaptBhmx5FJGTjDjWdqwsAdrGpht8b43lOSR8tW1pqQATLHbSz+HoWRTGWtygfKJyat
KMSXZDuWpxA+aQv6R6OI12+7p8fzs33CmQTsPJlJ6MGDLEj1GqhsjcLdAYRjWLFyYhAnUJrVfq85
lg+l94F9gEWdZDIH3gqC3rjKvHJKiX5jTqjJTAXq1N5NDw3nQ4Z0HBVsipkcw8glj24oEPEu+m0y
jVzWr7X2tgayqsFF5IrhIl3LYJvsc2xTykuBvF06ruOJ+4i2wPjwCs4IFtsSsnUM/9disGKwO2pw
trFoze6M4CjC4Izzp0DHZg3aXlo0a31wk2Doc59UAqoPV2Ps6DQHrklyqh9YhFPGaJMGVW8jnbIr
mHIZKT7X2Mn8NtXhkw5p8u0wF5sCH73W9pYdzxvJxM/H82e9b2Y0dHTRtMMgw0U6NgaidmsKdSGO
a8tmr0+bhU3D8/2IerpJ3j+BQrqYJ/U2kMPZ84CfbKhCMNWdakMKK8j1C3FhnAul+AP2fVrOuNEI
oWHb6kEhT3B8yLzGvNuDvnC/l9gDfB2iGt8kv+J7DcyHC8BbumEMLtWaszvTiLKMnDQz0Nimq+NC
PRzUFn8rt0v81SKnIouXkQlwIDJxIt4A62us/4utIruz7RlnTSgUWVSfFHWpCX5yz/FjrIDHHr5x
EvqQbN1FjchJTSbNPzGFNbdhW9W0zNDjKVKBVT9szterH+e7Ta2M9/h3uecBdHyBKqJVQHBb4dzd
sx1Whf4LsVdN/uncAxjZpyot1nv0AZ9FMrW6wI3raN81pmp8Hz3o3K3ApxGCFQ11YZof2qoHOxiM
Wxrh4WXKs0E7gXdwd1yzdaPSPJ45NzCKCD3Xhkpro08cuMSPRpmG6JK/Agkypf+PSmBDnZ3Z81Hz
oEKdGags/IfDfjA3/w6S8NSw2lG3yVjeCnrXrkCzoQRfOkfT+TyXfXUMpPmo0LnqlsLVJP39kLlr
mnw92Y8Pa43uq+jKbqngsjZxfBTKP7D9w26nnoX7omjH9g7ntP9SDc6wn9NZfXRffNZ/2zocIkfj
0T4zdLAgY82cAPmSasAN2TRejE/QI5XEhN4NlsC2zDcYpw/gM7LHabfNr9E+mcLSlMailZdvNpbd
R1504bxH4Aowo5NSG25OgtMi8AtA09vMvcZ5Us2AuarlG461g78KryYThnF5MIYl6Ct5295evCbP
dEBi8lkUTubFV6Vy7jFoevvgqkTCy183vVfcVM+B6CleK4TNgqOMylWwhqQOFxA2zEyP2VOtLx/n
wK7hWKn51LvGwbnvoeFYOrDD/SA7DaYRdlfBTrK9HlTZbffrbMkWoBtVTQ9txV9qsXRoy3mfJgIt
DK9adxc6eCZjiESRkjSrpVvR62Zv1YY+3gYfXJVbdzcD/sQBTffSYxClb18oix54I2xoMSg6Ptmx
Qp7L/MoYKRKJiQn6jl6E7M2tNIGQfhPxaL/tpRMlbnq6m7sMeZxwTE/Xq852nND8ok1XFDfYmVfO
97ENebRlryXmyHTSnK3Qpre8+wjs9J/zLj3lxaIDF2QjJAEfN4Ot/FdfydFj2JhIc34JuALL6h2N
tCqtUaZB/aVokXWSYIrzmPJjAaW2NBD4I+sU7rDmbflKrUsAe75BWnPq261L8D7VVTLeOgPWl8Pq
0OwKTFoUPJu/Mx5kGxMl06rjdFzfZ/YnDj4oc4V1McEgoEcxhTlRH0Nah+XdP9+wolxGqs3I4zpO
y1FbgoS2JqkgH2Owiz9BZsySRXzMMCfSp6Xqi0jdsXhBdebt+oestZpvheXNMZNJShbWKc5Hwv1h
1PrJr/LZJjWhLKvkBGYWvx/MEiLIV+IdTBHZXhK5qD5+pirrCJSEviIwH0ALwAVMsMs9VnA9mPf2
6bak/7m2AxzVe0IJmKkHQj6dEVRje9ZNcU97+qr/qP6LSGmC1g73YXjqkPs+gffBX3P3ms8vZGVe
jSSK5XUgFjDtysfNYZoTnwDaG6S/6vgI0Ehe1JvyzedPGbPKWuezu1pTIegdD10AyO0rhh4bi0jD
OqWb2gNb6kom7QF0jtWzZUyvNuYysuJ9mrklUqV5VGk6CdFPcJDwuib2oVW352LEtasY1lnFbzv6
psnNPcs+TjO+XWtedGw/LeSHsX53mElkxTLQ6Cj2WTGEdyTprMR6taN2xf4/W4d5snXirseocba0
/oOllVILWNbK24qBz1FpSkgiWP97Yo4E27mXo6UMNeNYixNngONz28tOtkBdl9rISu8jqa9eMVMD
NcUlOJJGMFCxYmUs+BGSPoyapGOw81+4pLCOBJpaHyfAnEn6B+a9m4LYnlrebxy/tpLr157J2CDk
4Rna5KOYD/vnR3twDZK4MhBzxwddtH3fb+Js1p0uvwrtINrR4MQSms1a7Wr404NaeCtsXAJxxYvD
CBBlZ0KG9xdX0p6SLzGdvPymjALZ1T6wf8wbZ20h3PI8KDnd1B7hBlBOozDCIOgO2IRuhtUJcLur
KC7bbz7bAq0lQzPXcNcAtd5qc7PxujVUt5YYd/LD2ji5tisgSAZZR2gOUVEKoO0CqG4BVc9plhR0
bbuPPm/WbMMH5xJW26tqoJvn1c1Nk54Fpv4ygOANk4D9lXnHBe4ZuSAzm5IKm/AMr16wmxc4L18k
P6oyGZV7Fv/ONTfJp7h5UEzmNH8YltTh+x13gmf47yLvGY1JYXPwF2Jwd0PKNs8JLYGKzYuB6Qb2
hKMJ5MKsvfbJHW/WS73ZpW+n/+p0J7z0PxSRSH/s2UMYszkW1vUS0xuz98GPdfC137QEk9+B8gmF
ORWVzLlCSPTH8lVk9A06EgYT4VZAv8WwVAWCWemVWEr/uKBviKv2p+kFmoW7JnyHB3FXZOfdcFFd
/eDqyVlzcUKGyQjuFMOEhd6xfGLM4LGm8HRLzOKtDqiE8YtdIc8K4qySZYn/YIEmXhuC/Ky09mKb
p7BhyYmI2CMIrs4GkwvYmITVASmNcVcOZLJ0+P6iAOCpnHxk/bihXp3x2/uDiejhyJEL8sPdN+0y
zDhEXGieTEseFF5UHXO7CT1YJVdHoGZ7xkbftJSZQyKgLtrpvLqcvNVC0Ter7PGzq7D35vK3vp47
0wIyZvEr2LiM/JqVcYeKUVoUsZZCVswfhYCXMZnemHziVRyvtLKQeId+Th+XIiKbnYE4pHxnNQ2h
799mv+/K2TErAM7qyvyYVEyrHjAgYSnIQCMhB7Isxm5OY7pq4a7wYstxTQyuFAbclo1z5UY3RnyK
i328Tn3ylQdBC/CEApSVC2UJs/s7FZL18jem8Y8xhytGxU9Ghfz0ifkI3r0lCep7EAFuoPbb6KlF
fW44mL/SWq1JCC1GFftoqjiD+5flrtOpKLT+VSu4BkeKjbXWvPUxApBBCWNoKsYb3rhwJwlSFY3A
tJBB3hIKUWnZLSX8BjJ/TkV8He6exP2JThsOLE/L2BU6Ah/+IZRUDQpC/ALPinXKYuzaASmafg4c
x7T5u+IMiydp2I8Wtk3ilEPTli8o+ctP/iEM7hm8FE8DvWzZFVX8O6suuhw3UIXEIfbZJqWhwzy3
NUhj1mVO3LtnyB9NPH8xL73MfF7SZfI+eibvENPua04b6n5FqGZ4bSlGZhVnRyCpIsSQLRjrPAcv
8wby5L2eh80QOlY45vKDBucxGZKxBCaJDH+5xJX4uenL0nGZFNk6BaC+3NLkBXT38R4fsJ0ApgqI
tmLY3w0lKDm56FwoXJlJGhBnKNqps7fvDbnWnexdBYT+ed8AdLEvIH4Wc1M+iQPS1VQquIM/wCHB
OU6MylfphaGA+j/BIGFiim1JuEA8lm9kmDCyalQJSlE5BfhISEyL3x+R0x2oHzkRDFTrDXBqG17k
rsg+xV3e0eCT+hXBlY3inw1bLmNcBchNvAeQYiGSd6DvYCEIzB1NzBOpGMF5g6J1SNYzGt8bQQkE
KaRsYjwmlD+ylX9PxSqxfHiMgyAJ9zt8PUo7p8i8RXwoz4l9C+x5zBgEaqic8pF1AgqZ6tbYZWkN
sjYMjG3/+/KIE9WuJk2++tcFKJxmm2TKsVVjRH87IRfmK60f2vkEGT9z1qQCJTJ/smxv3TBDb+wC
O6+YgUICYlEWc7uXCPT6n+fCH6oOTAC7i40nhvsrO1oYtdwLJDZe7eGmWetuf6WzXlWoXQiGyRAc
PogRmt9ZNwuRjqT82u/WG9pv/N9gy3x/K9jvSv7M4w2aB2oprv20WbtjKzubz5XpZ9kXsjfCleVX
HxvJCb/R5Se8L8/eTgFJ+CWsxrXwlnjCXJgzzzHgGdp/NhtcWViADBT2CqfvY8Qt9LtoRyDonwNg
qoqchvr3i/Wud9JVhdB/j5plN8Ls1EHZNM9IyYWAxpxJPvBzVwXvzWMbc7U0rQfA9vjkRQoD45lf
o1CcUzg/RSbsdDRqutjO9jk24ZudMz4OLWFvpvCMgoLkUyN+X6ldxp0NCqGE6hICLL1Xm85Rn0mH
UnGzB9cP/B7MIaarmyxK9gSyDA84bYG1/bSXEDT1zJRynSiY0mYS8svZTpdy8sWKgNLEjEXUE3XQ
vSObvlu59SGhT2nt6MWlNV+iZrbTzjdcSCNPVPunLgDbgSnNABbT9M3cPwWo50YGxzzrtMSyuEjV
1FLwHhlrQsl5wNrTO96dHsIa03PbSjkn3Ww2jnsrFUW1Q0mT74t2WD3E+cG9yhFFL/1Y9OzvRD2h
XuSn3+jpM4J/pqv20oF+rvURm8nPtFmsdUHvFFeQRLHZ2UefP4yRZcG6dLs8diYQQff5kvxKOzqb
wDYslKGO/CG/H15vcWm9F/2lVHYtuWJQkJT7qBgp71wofBOFf5ftOZwde2Ku25IBIKBG2OEJYkqK
+GlTlWJvTm1C6oHJMcYWhUvb44HAGfQ5EZCqGx9CrmHDYBpEiSb6yzNLEi3R9r9vZRvfmlJGicKD
b9aLBGXPE7DkM/DgPd6S0kdh1kM4wkwKpCkwT2ZwSilK+XrcSx/WY+ejg5j12Hks1BdvzWmDpr9X
rrXfE3uzpBQdsCrtfkNb6yeXx3ucV7vpO0xE1HfD56dBORHdZGiwZILVGqzMAb2o8uORrFErA3To
RCHM9WdYkqtyOTSkLuVpoqqBLM5Cek6HxcjtU1Ct8zHBUwrC45Ip6A9zOw73nworc7VngpcSO2TF
vWKRJNNhY3TPoHYlO52bYpKratJY2/sss4C+VNdv/BC9yh+zgoiTO3v/Bzm5SRxugJvOtKixKOyF
opaQzxT9d6sLi+scxSK7FJWYps5JcVR2/3DbACVxJO5sOsIx2cfft1/loECYiw4hj1kVZnXcy8yF
igmC6k2Vp/hwnANp1mtM0FA5iJ9hOl8WreCRB2Dvx2lQlI8WI28RqfCQ3z6sq0goetcyJC0x60ky
kqOaHfHkKHWt/L7V1az83I425jeNaPp6/sKDfcU+6CwovCtriyzt200V7eurZ1Kc2Xp2/Ci1ne7A
Af/0/6WaaLGEKmixr7gNHXYW6l3KJINB0GpZtM96NpO2CJL1XCynHFP6t9XZ8POWk0rbL3uR3ufq
qGokVkP4kD9QXud+ugoLigBm7NBEHB1eVcKvfz0VQqHq/akYmoAfq0tc04litc0zZVHn1rQ0r2my
oXtutrPeQrlH+mElESJphzLKQ2O5vKR/M/41X9AW4lKwF3uTJuHBSFQnHQuDIxLevk/o4IZjWh1T
wOIiKSfcwloGw8j8rYHzNvz+S5i0F/OAn7Jc+QcsEFLlSt5sTUx69HqMJCv6XFpxXus+m0Cj9oH1
plCGIPY7aNC/8j4+ULTyyyr4rtIZ2q/Ff2amRWuDANymx9OhvZ40o33xXzCKJgHfBILtOZfKXmUM
aU6pKDqARGc6c3g3eMUJpZTm42whxJjq/oYADV8J2fuGGTwKES2eJEUNsXt+D9cJzm3ufFKKhE6Q
qUZCid8rp63GdQu6fNeAF0pTOPWA3s0JuacNNmuoo29sr6HgqMs+lZ9yy6EsZhOCI9PckrXn4TjI
dGHljYGMdTcvlYhqgwLODcWlpIPZrtuzZvJCX42y8s5aIO2cr9dX0CU8+1JUuHqiABIDfGXy3bQa
CVkX5hwAW6cXvVH2Pudy+XwOVqRFkgYU8i7Y8knh5caldmRDs+9dpxxgVC8c0che/8Q4uw55KNiE
mpKXji/7guWQYZIl7hGcGT13vKi8ogTf6N5bAGdIkawyKQ6yWg9OrngyfFsz5ybNnGlj3wWuD/rC
kW1/LbXh2imsGHdasr+zT9oWafejyjeiT0vCcFLh0wKvY9tkXHfO7Y6Ed2e6XxNdeOwpsURLzVuM
9ksN67h5g+i+8x5btYCDfh1vO3eeDIgDOuWOYDfbFw06J3Z3oKB7HpA/YCToma3eOoRjRq9kspTW
sRpnz/VjXxMa+hbvfL2FKDVfoOjTa0+DLgUVzjauYJYTs6g5kihe0ZA81De2Ef2NsGCCb9XsxUp0
m4Y/J5zMKbySH381p1tl4nCt6aKUkJdd/YimjgGZtfW3Yxh8yjKoi212WOv7Baq9mqsYexThf8wL
z5uJvaWcRVUqm4s6w7+UJXkPI4LhOs/JzOMmXvVZtRneIZkzoTsKYPY0j85be+pVJz79wsf3G01l
SkScUOFFZkwHlwvRknzD/QBtz4UW1368LpwXTJvCQF4pIF0Ua1Q7M3bKgmDv5fwRpq427HPApOQT
Ujk1PQFUQLx83+7h8mj8bO4gWs4ZyLcSYFPuMLWIi+mzCcthNAdRTP7lretVg525wZYh8w8v15hn
foja7CjY+Hm8apcxG85XIsM2wDuYt6rhFf74oYgomMzTXpFCS+HqnjjHCYQ5TPNxJAhXhCC182As
7pXpCyGAvws/F8iigX73etgoqAZgfha53OX5ASvSz56rjXEL633lHX0T0rgmAv+jI+2sKucLDv/Q
CmVbTKesPtx28JXEZUcpqF+zZpqHvQG12z8TmMunqmbS+gO32vFNleSyd7d4fxjmpnkYW9B0uFfg
g2Za0l9tbIcSXoVmTxHOms9Pu4C8UqwnRsF4RcQK/bKZpbsA+60GCcFQL9mZbYZ9UBJKZrT0CDcv
BTgYr2vXrpeh1SRnh8f+cNPnZuPsdIniqwclxqpaySEfpzkY9V3IOmaVgoA4FR8DIzwUlrBAPfRQ
bBIUh6FRfkvpcK4on4cSJuln6Ftk7LEEX671Wl6RE+dk84y66zCW8JNoIKtSokiGVC99NgqvJ8UO
UPQDCzak0r8Lnc+wCDVHw8vrD8kFHp4JGgVNf890Z+HRcMLGHzARxb1dz9lJVr7Nu3EufnB0wS7n
eN1LsYm4HUN4EOtiyssaXIDqAF12WfWTWuammAuBrF5lnUhoFnQHL45Nc6oyqOxo0qsnEBH6VW5n
4GgR2ghqN/6Vi7o5w4zYV0zM2wdZheavcJAxEmpZxL1Zi0BXYf4hyI347EMO6YaTFjBQHGVKMbhG
mxSL5n9MuSrzxeEuaO8b+Zri++w40lDLmgfj5Dx8ohmZrKpX1DdPWjHeNlSvxGbWASk2T59t89zn
iTMSJrft5KuCPf0FbwmwSp0fY3ID9EYK5KC7uIkvW0hbvXuuVbKStEYZwqftId3cIr1E+knj+lhY
dVt5wk6UyrVypeSJu0wXig23eu0KKYUBUb/s8CuptzHUMYGCx2F8Ci+bsvI8/Fl/5nBv+W/phBk9
Rt3s/iMAG1inuGIeBfrmE4mDBq01ge9ShzDz/HZqa/GzwstY6FV3GwG35997D5KKIyLZ5gYKGvcd
p4a1WfYUcz7WybpsaII/xjdcvBqDvEGuJixuC886Kv9m3H+X/CDVTrLvvtFWwH/Eluf9JlnaYeNV
CT5xpHF91T84pl4cWmWWyd+e8hGEmJnc6KVjkikIWNqqf4OpC4a2Xv7Dpt5NYF+msuDg3cJ967vK
ouLahFT3+ZDI/HKDkmXElrjiP0uJ5k3QTYhN9rndt73suxVz5Tk1k27keCHK2ZDYj7aF3+jCzfek
Cy8zZCSCMtcUfHeFb83YQem39ogufQAHgN2f4XhlSNtSV2n2r51GU1AYigSJywEoOg/nOII2UfYB
y3cjLr4WzozD1K8kZVOD+ieUrjwpWgQ7ezFrV6gKdtKl68IXC354JUzTu2fTDagF/KgzAXy2uiTs
R5whi4i0XAvrj2H5IxZxOso7HepIt3SAeI5YIs84zwhDHbM6VD79KNw3b4r+13AooBOeDk7wZQKE
d8xqtK+EJAZKMuQK3MNBTd2ihQm233Tmadj+kNueGjP8wkpazrzCl8mGDlj3kxWn0/rtp1GMvWHw
TJ5OtJLZMhgnDy7Bew45p/Ij/rN0C/HX5Mr66YRp5HlTJ4GpqcdsQERmPxFnJsMv3fYXmS+WxWgo
pfPnXJ8bbV8Svvq5TaA+6d+HNyx0tqWn5TtsccFHFHuoCYueWakMf6mmuMIAhUaR7i76rlRui8cH
AgnNcPma7fKz01VSKznBpPJlYHvdvFBK3/5ZRnsgYyqaIT31uP9RTra7TxI8qzlwUSEjujz2g8NL
wP0jw77y6j8G46TJ/aXWf8itf6xwSqutuElTUWV5/DeM/IZWmIIgVUNWa0+Kyw/sf+BgVbTWGrax
TAiIvcguBj8kRErNbWLJyUaIsYhPtQO+ID+wzMrxllTNixb7VLN3H0JzFoVDe/X+Y79/S/0E1JKA
IEfISql3MezYiMoUXb9lTieXvFQtNjcxanqdg2OA29GO3j0kzrWC28mK0qa2V2U8w5k9N47DF9hD
Gtlq6hC0BFe9Mzg9yhI0/NVMHIgegnulPSTDbL5unPef0yiW9D3X4/edrye67jCCr9Xblc4Uhrlk
9TTssjh8fZxv/2QFGvHCu8fcmRg4Xj61rEmNETOmsC4g1A4oe9gma7GRIhbgRugQNsjyLif8pBy9
v42Zfy8X60CaIkpC2rQrrg2hqfh9ERzbphKgO/EK1CxiBUYTZdCKQec3GwNbkgIk3HyraURQTAB6
az0WDt1biHmA4PxIcy3gsUwwsPMN8QzPDVzzyJhUZuHs9RsqqczuA51VvHIPLmQLuqOl9zpoK4B+
0Q8SbhgnZESy7m5iFs0Ka6TUHPh/QjaXKnAwsWn3TFQWDpdp+E9pKBpjqDVwc4VGj5Vmc1zrgkST
8O4IStLi7a83QzFkcg48moHgmgh7kjCW20LltcvbkKpvMmQplAnNV6s1aZkieaYlc73fNZ+VLq6W
rwL28KzO3QNF0dZn86TnEMW+sCp7e+ccsIQJpoV6ypurwirPXNFEzPxRZve5tCA4YBCk1x7ljkN7
0tgHhMifSQjyiY88xTHD4EIes1FJyW8ppiqMh0OZhqJdvdDuboIsuV6HNBJBS4hhjsB0p6Gqy2SV
0WanJowF0RsWlHNvMNzHgAL7aJwV6Srq8WLN+aLZIl202PLL8ADS3BWDhVFAuVGnw//fQkZb9vgt
PmR34BE0UiJdC3XpQpb+wYlznOK9WwDxlpHWG0ldKEDQ3W0zQPzeWaGVn+3gtakEdlDWrIDNgkWP
0/O2zDKFmuFbIl8iAL5JpE9LA87iOqDDzudvTLVBBvQ0Lqa2cOHJbc+oOXlM7qU15UkMO2G7ROFC
Oq6RABk/e5HeZoGm2bCTyn4EC59h3ZTPfABYqlGCqkU15zJnL5bj9TiTi+4vk1qsOHYx6mW1l/u6
uIvPfdB4qF9EAGkA33iZ11fEAf4wMyYE0dtgyWBlYkTW8QdnGkgLSjdhfxcbkpiNioI1jIzUTIQ4
8qDCfkqLnDX6q9WShnZZ4b3XvOvxsEJukzDHMMezIxP7PPehviN14sBxuNYiQIyHfnkYVMBId1qn
MnB7Njyo9CZn9KU9fj6JvoKKgihuJ6VsIQYFDlWdjhonwnRoxfPvYKkbOd7BWgpdhUd+LMnt0wzc
LzB83AWAZKtiykrzQR6fRcPaETaYpaPFpMLbY83+Lq8xUoRa7y3vLadJufmAmWeyYDWBga/icKGl
NVsWObl05Ki0QYtWv5BK4JFCnvlP8fVAkJSRQCqC33F4V4g8k2ShJe+x4NETdMXTKHI+vVYsX4Po
sK3Bfn0AVc20QhRRYqKv2Yrs0iMB6b59jmR9bEZZSEo+eWscrlhB7aMQp19iTGOE+gkVYYYYUYW3
h7blMAVadclfQm10z+JFOI5XjjSuKzZTI+vIZ8FWmSSYC1a9eSTryCrKI+8V1+i0J6iTpHLZ2K7N
6JbPeV6njnm18oXHye93Us0zssHb72zm3ALLApZNz373e752WwG27cNlTwdFkoBjU72FTF0/IV9U
+VjT1MYVdxY7v6AWHEaqL7rzlz4D0BeNvEJx5gf5IhJzgvPxZ3HdXcoKtpVaagPqR7wxKmN0dPdc
KC326V5FhPFr7vYjcqEH55ngc/JvCuXjVlLaOzn64k/vsxT8kJKCZyWEY8YTx9vxlD60CYshk6FQ
4krBrOc3ies5N4d9h1Z916KkyHWHDvgsJ5WJmYm04ZQZsOsISVdZ1FnKPmwX0ulYJ57nQLP/rsdt
lyHu9UWmf5yM7l8nwBjKlcQ9gNmi8eAlATT0J2lkNmax+Sg6dYY37jQeqqHQzCffXoL4AluT0jvH
beL42xxy7RZa/DfaNKM/4BGRzM8cfRnrejzEupQBE7gxRlIkst2E8DLdKilLOHCqHhqizVYbms0w
SQMN8NMzp8/ff0hJEWlMWYvVKlktpq048c2ztiC6q2KTna/4ARYNTWnCskMPAOH4tKjUchdaxiVH
xBnCHeBZTNWej7eG+4MWZKj7KYDBHa+qzeygQGc664Hq5ViQ9ct/xzaMKpClmDLhui39287pEOoK
kNwn1NqfgyP5yWLXduxlFK0GniQPtAQhBWvn4ypSfuUsL1wRZeBzC0YKl+Cdw4t2ekrwfCEnvd8q
T14pZXyEfKBfoBwN4tATmA2AqJWSbNBu1uHr90xIjbMEM4mSCbO9y2xjm+7wXR3EPyHCQVMj03p+
iS0iDyo3e2/7GwF71IvSaqfk6vr2w3HA1BicRMvv2lx7EgLTIsPD3ov7TBwDNE8SJFVJ+vVhuMBM
mcmRGSOAZfFU5pewHaaCQYLYUM45IYHpCGONAn/l5HuFsdgbmgCezD5Jupy6sIdXfJqEYKbx1YcR
qyksh84VkvMyUXGs/XKqfXtGRwJOZBJK5IMazw/OdXQSTQsM2gkB/6RexfHMNKmxigTh+9/Cmx5O
z6z6VoAFXhNmO0jrYpQYRlP5lan/PBfjmKOtZF1MInjeyhjyeO71LW3P549s6LMgh8KhhGFMQ0pT
WjK0zTOnjVVBIeL085ybhBx2oesR7zeQXwxdSCXytwyQZDy3kf7WeqwOkXtiDSq1hJsRczs18u/B
2SHA+c3DVW3Iwtrr17ZkOMUAwtplVSSiKOyyxqZc8I3UStxhKPdSXdHofG0h51FiHpWdTpA6eDtk
EU3f08zxPcksEk53YWe/WT+xnTsDcFCRsufTz7A6qMCFSWT9aswJdJOIhiERjFgX+tHaW2El/Bf5
kuDQNXg6b7xewrr+k6xxeVMVr0mns06Af/GwkbhCYBMvaAnph58ejijtzNgEQSiGae0e1nd0x9JH
gMbPaar5ea/zCyI6YSwIixelkq7z1Tq0voFcuh9GZAK8qd/pY/+uBhPy60pwL9gP/6w5dp7+mN+p
c0cmkOsLOUzXBXTAcWJV1rrtbOq9hq60HUcjUD7x69hz4joVM7qmLpYjbVxtsSxFtj4juaDA0joM
p1rap2A1Nn6OmnLkrh2v1pMU3JIvxf0sgiuulckY6T+MQiR1BDbKgzJ6+XJkxKgsS6wU3OmfimRp
IQ5bfAC2YWTA0X+LXm8fPvlxYa8iZFl6bVQD5ckylaRF5DmROxnUDB6qUr5OiGc8dbwYAYgRNNHg
IlsLXbGvq+3GkK+C5rhcyX+vQN68AfqCQX3/y918WEIBN4dyv2f3q+Yp59ZSVRITcahUj0N6pNiC
gmZCLHgzNEZRMRX4P7Ot8u1Mpg1hEf0hSa6rHqDZFBicGZjflhgxszmBOlDndn0pxINuQxGSYE3F
k+RDfG8rL+++vtrmgDljQdU/a6B9gi/3ldoovCP1O0GdQigvfT3oBd7v3zAPFRHJ4gutVW91aIRV
w64FSKKZ8Qz5SSlBsOvodb9bFJbQ3bFCZb9TH+wtEd1CdnERxOrHdEYnTDMJbIzjEaNpsmejBV2Y
xvGnm6EUrp3KHtJR237Gz/zFyfGXMs6Que9oRhMEEbrh3JVloQARu6YxhmENMFA7IYzyZW+4fMzu
DMQN4Ed/B5K2a2GFHMsmH9VcTkaQ9gWRht8o8CSu2yLrKMvEzVlEHHoyLQiRWMn38gR7PPQmxImE
YYI+PM/cIa0ox4ubJWUpGg0qbmwsW1NMOvZ1B4SypEfhrru55N+iHWc4CA8NOevlqYrF97blnLH7
0e7bOslZjiSowoy7LVaROCNWPK1vX9hEwDU9hBRpckIM6MGvyOpx3FXkx2obZWwuTP2uHA9iHvwm
iRDr+DNbN2i/DQG4LXSqgcGDKNTKEescRyJzzi+r7Pr1Gy3PXKgdImo22V4EYJ5NN0NW8a4UJUty
yLxidxwcssqgpeG084dU/hj8Y59G6YRJWuMry/r2iQbPi6+LuFP+Yb0XtnSG0c8t2z0kVyp/xQcM
lxQYNTzBVtStk8agYjldRBLEfGCKIxmL3XCU4xPiqdvHy6i2/HhitHVn0MJmGMwgs3MhKQ6QSS5I
+K8HMq9pxHaaqEvOvcsnsMX9Ek4vKETWBjsRdMuCitbm/WCmY9Z7SqwiMFR/p8Kbyk6zcYIXV46w
MRmUMG2Hd8uFRHDoOO/UhQpJvCRpGnTzUHBPo6j1tyTnqZg5jAzR+SvKP3j7KD8FVIIObeIcoT/P
bG8zHVEfoWpVl+Xpqw6Ovb4BoiLBN9BH0SQu7uAVl+E1cc3H1L3tnCblX6/+yAP6t3ZRVxdO4sp5
lGmkxpD5U8LQZSZ/uILAgLVvlGNJe/qdfWUFTqx04GzLk0PtZz83xV5alNX/yZfUQyrXwLR7LRPv
1xIkkzSOHYvi9n9AcbujXmoW+BiPACd7O+/PCcqiSr2cnJkAGqmsYO1rMx8YHbV5E82WoUQTDsUV
HToRemnqBBkXiD/49zn5iG1inQE1lh7cHOz/cH8+SwhrfPkOCAugxcp1Xv+F8YJ2ozBINsj+TVbP
E+Xtn6eGhwriGVF2NMY+PuMyVX3QS1oI5u8G/is7cfcl05VuTYe7uHphUdC4bvnVZip/tTaS2g//
Jp3FRLoI//zMT+r4sdfA+uS6t8m623+fVT4gSyJ8nCbdKsUSYyO/CwQs17QFrWL/i3cH4CiDBd9V
H0G44dePRiSGee+vWtR5a5DvoGzO1cyg8c2M/q8pK67qQtkDiIg29E2ZUs/DBQRUmlf9X4XOo0qk
JoKFhpOx6EB+ACtEI4Eg0F+apP74RluZw16n9cu+l0xuukR4ll1jVJQm+UkA9bvvOmgjhk4DQZ0V
EwWixpA4cRfuBxzieBG6vjRJz3VLPLpdSZ2W5NoUHkppOUeutq3hfU9lzCWopQ+N6ccunYEcOVWs
SJBw3lgPCTD8mwVDsAHE0t10obfbkzFMkvM+WklAdnySIL1q0J0kWLmfQAOAkV3lpMWUvB1L3aTa
w1Rd9RA5A4Z2IkJs26tjiSf4OtxW2Oj3guK5SJ8lLlyfReduVVSAHpTtdWtiA/I6Fr9uHmHCwI9u
XJ/l5Zoh1Uk6hC9C66P07n/QnyT1exjFpCHA6rioVcPvm+E7KCuBm3uIecvfMW4gkeKHAIZ/N7XN
3Wq97ggmTQf9uH2kyK8JYXsRS2K0U2n2wPm1dXMW7Kxf96o6QNW6u/l0QnMv0EdJhOR52DgliUbH
G+Gm9gpK6rooaiZ0LW7cHHZOVarWWDqu7DdBbrzAPOn0S2VhB3NA/PbkHEMcu92gwAW8ndeucyB7
tzCcayPap3RlreiZ23DJ/M/bfvJlDuBpT6Ly3Lb6wiS9xNQWDcdYsbeACMdueo04nPaX4GwkC6GW
XhDF/aAkO11bBin2+NzA2JVLjwVflxA5yPUAy7e2kSQch0f6oLhJtrZ/bikm/IW4mNk4IsUhCS8/
r5iw2/RFiijoRysr96lmCoQy8iTWK6qCi3g/janBLaC6/DoEgdtKG7xO30Pme0zeWYM0cp7FZ5B/
VhsQjFJBZVCWBLmLtESdkEIM/2YNzn4/kE+CSTRWsTmzyVRb4rnrqKeBPqk5Mg4BXKCPacoEXRac
pJm51F7piwp0U1BVryiu3BkexPH2jvszoHaYi7XOmCrSIv0/I2VTNXHxpVOI+jRsc9uo3VPqcMus
8H1jeNZQFTihSHlmvVWs3aqpTbETrLG14yl2y10vXP32bHH/YDekNkIkw+xWkAcLVD8fEeHTGfxc
mB/l6FnuilZxERZw4Dnh/RLlFCMWSGjQi+9xLnNsL6uF0ORGBARpllFl5uL8BxuzehUrLyTTaShQ
Bazifykmb94Z1qWh2BZdWbAwh27sap+Q80YS+3L8YLzYZsrN2gnAxCj9fDCCzTloS/9jKHJYXwCO
7GZvqh/024KELS71raFMCJoUDn572GpTNSffxwk6tRgYzY7eBZ/PEn3xG32v8Wlb6Lv3JlgCV6SP
ddakwAYuR50udOtYV/GMIDOOwSJ9zLpGgEAdGXJK/NWyZFaw2J8lajM83Q6K+dRfmAhAuDErBLSI
eDK18DBAFKeNy2/2ZdgNtYbO5jxSMRX1S6QKrx0fu+eIwG042FvbRETnpXO0DhAK34RFlCd8C89S
qvAlQryEcbE4rJfjodQ4cTgRqmUxMROrmVlWOZ2UMwZtKAisNTKHt5SIILILh4D8pNI1ojYf+qdV
qA4zpDEPiIZkRNoBRoOzHnJUj9U6EoqcgNU85Xmwrn9LjpIGNeu3I+V35AP8udxhMeZxtBG0884i
0OAv/x4gJ1nIhi5PoUgcLnWkQlXy+zIkA2XI+j79y4GcWf77tHeERU2vPe6xkY/+8DzHSdHAEtM2
nwD+6OYSblCZORMPAsT2AQxKb1jLdKqACg1sIyqdEfsUXxTJItab1B1/hKko0HeE8rMkw303ZnsE
F/TiORQI3KXWctVawr/9m8LI15rzP2fExcte+Wtatk6Qif4fMn1jamq4FPjLW2MzwbTmVstLVJPQ
SmoJFq56QDL0VjC4YCpBJfOTBads4VD7Ct7QhDKIKRuflRL7Ul6OvhtuLox+scyZ1hb8K+mUD5h1
aLrYfiHV9NT6sXZMzfSBA6OcEVlJhE6iU/rBVh7WsWWuwIJg5tRAbSOnIKn2ZCotEFGD9ju7oE0m
xQ33V90LXdQKL/0++MEw3IQoKpx/5wVEXuanflqb8J7WSy9dN2gSBFKPB8ROg6QGYaGehB76s7x4
hzahW7cyEAMSuxAnTwmidxmoZ4ERykx4W5d02l9+qmNRJTeS+wKwJtLboj66EG1rsb66c5Zjzmdt
GunKouHXDHZ0R1ILTkKCKe/ZjhGovH23saevcKO/Rq40yfrzk8v9DzJB1u3re/aEvRiNovrNwIek
S/nb0YRIqkLac37xMQRHZCZNcqRfvcbxj6VuACvblYajSwsLvxju2ymiHJWhPOgOmD+axraIgPbb
kSbqIN5cTQHt8NNUVpgBgJwwj58T/YPI0LjrpoU2oKZwlXGLqzXHsAsMTsIOlvjGbpKBcv2ysKcK
UBXNndHdcK7bjRY/QEULQo5KmukcMNba178nWnB3rGKJCZ1bVrJh96bZjS3mPJTv6ZT7RIL0AzF1
tlCE0rTvPp+QVIapjApZYQaiBCyFQZQWIPc/9QfoucnwVSUhkhDmz09v1irnRyuuRhEiiHe8SBls
icCPrxl74e6AC1231WHv7FxIdAVs+582Vll77JUKyCoiqlN9Ql267dBuxO2MxBoxs4vF9xPiZWh8
htoWbkU04m5lPdjFpLqHRssNBQCIDDJKTHo2RvJgYMWt8p0zfygX5jmjDbn8G8XvEnqLACGXuYr3
nyfFtT3hAKv0oVOCpOGORLhd/Gx7k3bv5VfVMxtnRy9N1zanlofHY+20eQWucIQKAmNJIVJB5cVf
jeKSYTIYn3RAcvNdyyrNqQ5BrBW0kpsFjIVbY4k4XfibulfUwClJZlStkwThiDu85Jvu9D2vJ1WG
10NTN0KjDlpOTvtJk0hCJHjVt2+YscKFSwJoDoumOhWL5XUA8UjHPxUQQrsZuOCEyijhpgNXlfG3
Y3WyKG3k3p6mi0+2SBhCIUEVfnrHyiIWkTFG4NGwCCZQ6ZkW4F9eqrbWAGY46EM4VN73YfnUAWgE
17InQnl12pChIbQslRoBoe/r+vq2m/kzp4Suxb5SFU1yez0VO571xLhEKsvdarMzHCqJJ7O/JDG2
6frcquYQuWUffvvNn/cIu/2Ywz4j1JN6tq1ebrU8/yhy1TQucg/4X8tZIbWHgU1VGTqkJb/LsC2z
4+tYW+yTHwI3SFsGKgQi/oouacMcTlxX3gjTUbTqUc2238ypbp3/oBWEiJqxXpzEnHZuUbOwKYt1
KGQn/2H/tLnVLBF0+OJaGsAqVO2wf8xwe2iAR/ZwZ2G4wflGDfBgngVqOe+4tPN8j6STcSQJaHcE
tcUQsE+7Pyal59qF+C0HrAAc7Xq2Cs01Y3bGK70gGn7t8+vbNSiNAXlWIXQrpNr8zgIc36jS+OjJ
19CuSuV4MTTryYcMJ0DxnnAtD1mzQTWuNK6Ir6IsRapxxiM/+/vZa4Zi35VnQN2phFUvgaTc91Ys
+aS1PgSHwnezuaV/wCzRMMKFrNXEiD6yl5bUA1bOsnk7C8hOX1wfBl9NCoPG7iLvXWMM8r6Lv8o/
z9IJFIzP4wG+2LNA/bqlIejj8aAmUw76fMCAtd1UGOGXIqZFRt0Ab97TpNX/ppSxR9b3Sj38fgpD
fF/9lSkTvDZvrCFPY5meiuUzeAz76biYrJdXcf5XA8rufpbwNRL1iWhteMtP9sLJWX12rXG0TWSx
87tnf5Z2sl8EI9BuZ8s+uKWMmoAI7E0eytaZ4aF4jrPGx6SgrFcNcCYsTOq2EHTF9dIiRErlVGuk
p693mj3a1h7tgzOx/U200TiiuXOIU2UFWriN/VZj4O9vJrRbMWLKgeVoZeY5tFdYyL5YZZBjevci
UzL8JhEvKBOYODeR6Rs75TA8Cru/gjTyp6YLqUNEuD1UbXMA1BWvKI5SsLpOXD8+OjXDsxn5bYn6
LG6muj0tSw8rLLE9jZkovL5v7iWwF2AWlvZb42YKo1KFwzxZ8PUEHTbcSen4z/LjP+p+b7pTHhDX
KnwPV67IZpXTGVQmxZ6yZkrEIWYiX4LIcNTiyDkcXjs6UJQwuSPNcSG8FGikx7cA43sb6nKXZRjN
ijjT7YBrNMYvQZME+0uXsxSFEA3OZpFXFF6cxR3h0htowuzl5sqsb7EUY9s1MlpeRgG6E8jzJiqm
PIeuLi5I2U4JxPv21OsiUGgcyO+0H5pMyQ+Z2MXrKGi5IkUQLPXz9fxJeKBkC71pY3BOgVTB/HXN
n4bJAigvn4hiuQKTxbKBQqqm+J8HzG8lGUWtoVXELk0/j+j4YpJfkc1sGpYCjznN9b7gwY3zGVxk
DqH/R9rXDdQuP/kxSPCbRDPfAD9rMm6wBjUcA/j6ayqX7Kpm5NLL/ommKxVuIFKZuz89pvhpe1Hs
whO3MWLzXEsu2aA/g0l9k+s9A8VIFBxH7xRCGZO3m1W0bz9/NoO8PTr3ViggXE60+Bu4K4V8YvP1
Ohawd6TBAi8Ww1RdyXP1c6ffRAtBGA029a/iZWzFo/ymibLySHswAWQ+wx7NYLQZZJsuCNncghZK
8JsbhAulgoR6hntdYW29BJq2DTBB6AMVbHnhgkk056zOY1fW6MzlW5ZF87ipR8V5X88yexRiRsmf
MF9tQijck+oDIS+tX3gpXxsnJLTyepODJDTP2PmmO7hlc4w9Fhu0qTSPPeWUxZ1w/HiTJl0lryln
+xvIzNY3zoWFp9IjFWBixJJCDpqdEqaDAjD14tJ8A+uMaLYcJi8BGeB3H0v2bMoMFAXEoJl1cJny
KlQfJOpjKvHDOXNGJYmZuL0ikI6MN1XDdijG1mk+kzdMcfIPWA82n7tXI010hxxp8vuSLzsNfNOV
DaTjnJiW7WkjVsfo9fAyHfwGfcrYL1Ct1j+CaZi9blFnOycUj8G22hWFaduaaZlMx7IH7maIoaGD
hDbHg576ynksuiTzqt+aBYC1j0J5hBk2blT8/S7IkF94eHSyiRuWNX0Syp6e+XzPKZZt8iTrNpfb
xsKXCOpPTmjAjGrWGUWs+E6HZBPyDv35k1wO1DtFgnNqSW5vl8bW0KPTqks/OLMTr8EqrXl8zKFd
EiBWPJu1L0PhTF6HD6MW/TYQsAe2K5JdRECkgKEJhCPKJWvJC7UZYUGOJg81/sKXWVvxx7lJAxCL
A8hs5/Qoj37IvBYyeAoFnyXbi2Nv/VUHAmK+7n17JWrtSpAJgRgAyfefMP/unESmz8/5clY5pFZi
N3gAT+CSIi+GwxXSCLyIA/Lb6u05htTe5tOhxaDorwh8jc86vvk6VcU+Sg4hXESbXZHaJYup+5SG
B9H/Ajet2pg56aZu2xgasWD0oMUlX2AK/vq8Xc9RaK8EGYHxbTK6x91G1AjYKbOGBkGj2apO4PaT
rCvGO1onLKKspg44bqirrHFKg5MCu2Obz4h9g7cPeWyxUt3Zr1/dRWpo4q2EEsGqZgLNQlr1Pmwj
AVmHtUAFaRPiKugSNwotnGfr6ckkEITDZVef6MpZieTnWBVd7PcTtttaKze0dOiDxs9YLLfY2LdR
8mYASpvVOsvWwJhxOPJCKNnoJTkExAh9NA8mcO2gm6y+AmPa1uFqjj0dlMxWTmXkXqcbF3uSEdVY
sGGGqui5pwhLBlcniwyuqD/inzatg/IJ0tXbehgC/AWnAuyrVL1l6sr3oAnMGjt9y361PmXVHDfb
OjR2WSOQMVxiwKV5w23vRlOwiyaf6BC8HTMCcHFAPys/uoSUB2qhaSDNq77HNPetCwZcPlFgWubw
zDA70fJio4oBBiKkgdjBSKaAb1xe8Ur8B6db1nqEdR4dogoKGuFfRFlOU8rgyH0kyANywIGrw8oD
4WQp3Rut+d6FqhpLyBcb1tD6HM7tH+p5r1GuRusgNmspI0qIH4CTCOdKvBT8IMDFKs0DdY6XPe92
HU5iiQg8IGgIIC/vRzNJdKHiUCdw+u1onmwwfSpBpM889PmhGIH3Li13sMEZ/0HYg/JzyEim8NJ6
5Jb0VYjp3kgl3+wblDsb0qYha6EhUm8zLDlWunn6PLtgrg7aNHDoj028JSFuaOKowDNefRw77RmI
oZQfSqocqEPWxAsmwXJe3c8RT0BnMCPRDYJo4rKqcjEQpg2iE1eXGxoppLzEpMYpvT5JAuchJGiW
4u1kf4f7qtIAPvuhbw9cZ8gMOOEv9mwR2BT82h+Ct+4pqmg+520lsaYonEFaWgi7WacP1m1pFAzp
a1YJ/Jx75n49yMRk3t7qYPG7/rJNuI5fMWX32X+lYgKeUdSODZSXnv+RYfXZxeVGxYh7aTvxIZNk
Uk8+C4rwOpDRFah0O1kYonAEbX8VAPxnL6csdgyctEFQLckNRcg8oqNNzrk2PxIRKwemhSOfEXuj
WljXwVnswagthQ2eCm84MFm8Vaya9gk0/bpP+he2dZrUPi1mvmcatf/kf+Dg8KO5P4fII23GWU6a
yrzFIAlUPbioAovYLvVXcOGwjNn2ToodHa3bI7tosWFEJU7BtvK5Wlzz60d49BvkaqSNRzVX5UYd
ua7mLQptzRZVoWeeTOvZ/W1wbxcjlhfCx8nbDHwKLCzJMuqXtu0Gx02007qSi6al0P3iXfGKQAiL
qhN5I/A/xa2Z50Bwji8AyJ+fCp6yJXPfh4ZG6ALoh2jmf2tT1DlIbiFI24BRIYQLrq633cGZB0mv
uDftyTgHscu+UTUzUd18WWiyCBhvK43dUH6NhrnNW48NKGsMEDgisOo5alwQvJUEuCx84ZGgN3vd
Y6fvObbsHJnP1TAyq+gdwZUs6ilPh/tmPOWTEOIztRSjx6x9e3gvhMGmaWimvBD5W/AJ+YIdMFU+
QPOkXM4MAf7Qi2mOZVxu/VVT+swwNxKbyQOwOsfsr3o+R9tmUkYn10X/q298d/UtExL2CyJIak4y
Lj9ERRm4JYpNFN7SkhOpZggFAUDXa2XNZXkW3LWG6YxSVidRjUUgOta0t9HH74k0Squkz9o0Kq3t
353Q5eLqF/nvRm+qWjXjOrJ/FHb9anCX58R5kjMLiB5bZYJo4f/+nPDulZOiRWSldIhRqA4MdCkj
wG1gsFcbmK6/KSg0GOZsgy1zrsqAMmfCfov8I0KfIWFv2DgFAY4ad3KExnfHXyc9pB9LHUpafd2r
rb41bmdZ+iVzhBx/lYSEG9gSWgIZNv+G52GbzUpJKw1OOIYutFO7FARrtwW7OMWljJ/nBKY2JI5R
94Pdku4z4DLf1FGwEligbDzw0Lsor1lFHAY6syQNn9/H6e/DCSI7MBX+5/1muATXuIA03gHCjaAt
xiG59e8NVAMVMsrQlL+LH4BAUMWwNFuE2alDBQQx0pcRpUM4EmC79bs3T4qNj6dPGW4B/AjKUxKn
P7XCnN2mClZe/EdTobNm7jPHYqDDta4/A4PD2DGMpRcddasc1GzhmgU4IZMVY43PS8DVEGs5bUNV
lP8zDYWTk6vEy0HrVKOcH6GjwrVv8o5woPt9UMJJrPt+xc1OZenwuWcRcLjMfIQQc3onhqcsTdED
JYAb5nKJRzn8SW6AqzwWEzzKMpI8wensc/T371dv+gn2nyK+PqThvPyFpa99bf/h4fklnrQI6DVc
01SmfXaok61nr0SjgMjtzY9RfI4Cbsw9G3Neqb+txOPFzQWo3S9h8TWA0Ai/ccrFHiwkn86+OC3O
lz0JYJwzBuyusqQYCEQSeFEXSzl27NRMCu/9Sp8LnPKRiWwF7Fs+92DnXjwatT8ED2bbPVgojdsw
tPBhlwJoD5LAjBBx2owx9xC+MqVkfxX1y18fSGqbKPWpWMHPgl2i5f8YQ5c9h/Kwdm3bgoSZV3vx
E44tC5HpltHB8cB7kyTRPiCcw3mMY6FXbmIppF6j2479jujWf6QLXb0ahnjdW6RXIfnFNS6yOB6k
0i2LzlccbZNyjB7K5Zec3SGu6lJVkjXtPREyuPMw0tbu0miw0xYPuahts9hyFjcisvEdu1oCAYC+
NKlZfW94xiM8SBSa9/qRIAl5PKhWEGpLpa67rWde4ummb+2qTAhtx8L4fhd0cMBQUpVP92PkSjb9
ujzCrwdy2VIdf46FvJHof39u8/52f/aqHuhkpE6l15T+SewmlDt2OtDgBuLrv+nHR4g9ESTThSSL
vxVGT1TZjA+7tXMiyHydClAFWNtOy+hEo33RWncgb3fCHvKpJ7CCp/zCyPn5bcFcT2KWh3HIWb/v
jBuCY21SdUQ3HsId6zSxYK+ZnT25NJCnlRaEEGkgiTjyXeMTDVPejQs1C148ZfQ/ql7U0prarIJM
wSRc/FSib1RDEAcgHcIBqk0/sJ1pURLcb39+Qld1c5PIA+X+7YNb0UrioZxuCFm41cvJXL/8xj+9
Jb7jxXr+mB7JPLKMeN173UIl4R/ZTIUHqKMu1cu5Xl6itSvyQoGeVKYOfSw2p8Idkau1Zo+wAOFU
M1hVsBys7oHtkzI9Kf/hg9v/mdlFkIsbW9oNOVp2FckWfHWhj2lHM30/sVgJVLor8f9pvtPRAFbo
6w9Y3CLLRyLLi2eYcDJQXCwMV/GNivYGhPl+lMg2PzV/e+9eAmZnknTvq9stWqngq823aKeBB7Sd
/nRdixXpgXldRbMZarro5XKMRHkQDMYTK/MiBljIcLnbZPelDx3QPNsU5qTU3meUHdx2mGQ7zfWK
ijA7WWzEYWvaHd1cRrn3aLG9kiHUx9MWUAUys0b+ziO+pEzgpI5Ip5v04blsJqQuiHSqSdAECReA
Q9D7LaBOgvTOEOZ2VDZOak1UniHk+ZevoBlWNYw1r58kFEeLHFJZtA8ggp5LyK2UWlxfw2w7GnPf
KxFbfiFYODnj8Tdd+wcMbD2Vk04NN0Zdtnw1apWKDs/isoO6Ll+TU8vj10O6Sn8nVu172dxfGGVs
x78gRyFF3tkY5xqu6F72+cjr9Y/mh3hnj1BUIsJNMYSSuTTTXCWqb/+cn3L6u5T67v9f8zvwb5ye
rgNDAJE7nkAzQAolBg1QWXix9iZQ8dUpU0ISermZ8nQ0U8D2h+Jeyu2WmZJ+IaAPZJ2I+sE4V87j
oci7X3WN6yZqapk6dgvyfGB0unIThIkDvwn2laGTBuiKD9wDZXDpnIDWEmZiBllP26Y1nuAjboM3
JlCaytTsIkpCV9TRTA0k95TRRh7O79ZdOGimj5moSNrcuONT9FzjHZvREVk4+nPOkWG4vS4GS/dy
WUibZBisbkoT8kVQDmLCRLiT7XQFZgRu0dpNAgN14BfxnNO/QbIj8adPMvrCzIY4DMgJCDF0EYVu
B0uEG+sDQkkH85SDVk32FM823Lu+Im713CE6CPhajZ8pZnbs1cKMPQnKjTmu/zl5BmjtRS+heWMk
5Phx/NMuRnj+Iy1e4XeBY1gKbsCiGtr5QAMyr2TAAPj/CmGWA9c4MPArhSHEYQk3lcFDoVmDSX7O
A5YQDHhS2VSe6s8y/I7DLus5J4LWqZvaeTBswWEyLM9TuPwtqDjKVkln6S74lqWv1rwzWL428E7x
A0QEJ37t7PMBPgCxVqpWWgTeKibllymWtbGl9D4EWh5RRyVCpAAUe+rY0ECn58sxKdjonRqjQII7
saRdYTiF/nUF04PN4d0n3h5bo0R7x6NELvrmoWAEh1kAtkZY3oIRGKk9BdTS/0Jtl9v+foZ2EVCd
fbh0DjjjWOX3OYrB/HhzwrfFNlzciUlMeIFzdXNsHsPff8CtC/aIL89LynmFkASZmhl0f/MeT4Lw
Ss9v4XDGlqqXQ/Cg73T8YJxg/TmwaArP6ch5l+7JHdJq8ODLL1bjhvuGE1+9LC6ttKm2JEHOBTlL
5QLcpqNmxv+mM/osYWqbm0nvVLQlETjRmjWn5NV4QRAZ4Y1RwSgdwbTz2Fb+n9ko1fOSbPQYd61B
DslB/YeGx8LxH0Yz6AUt7dNrD4f74GAGZrJAEsRhN2YLLm9l+8PW1FQeITkcAyMG8fjzdYfKKj2E
DesJOBxfBnjGGQP8AjsLSyXfKqAqGhXynjZPkv2UpWizTMk9ykQFTVl94yTxAipljhtYvLkYGS+/
qBeQ6g1rQtdgnm0A15DVt8i4DsrDcGHvmku6/Me1E3krBWhT4BcWSbuZIltwdR6q7p3pjNVuT/8J
HWNOq5N0oO4mMd5eQcmh7zENnrzBHPTmIrF2EDsRMMxKoxHs8J4FCjtKcPiNl5UbqdUGSORZpLrJ
9BEDeejUAA5BIMDTr2ruvSLRujDJZTgXnXUq25Z+ZeKKkQq+ZFUGSJQAQQlyM+GNf/hhiY9CpOR8
AOrPUsO/5lkcXJbMDwQoTc2wqvasE6mgBi6o/gnOqNguc60/EnXem61+z7SmirGjuTo8h411hpO2
hVVJbxrCDfFRjEf5qCK6lXvXSPGjMyjAwGF+pnwopHJE3h2Y5Sfsz2ed59K9KRC0qudRwBJl5rkK
qYaGgeDa8JLZI192wA0Ua8zM95Q0WnyaJ0uBK+uNreTHIeycTWUwhpREu8byKMPbJOeoxDP37Z40
h/bHKM86E482eyOKkRpQ00P6lrNkKjL630mXmT/5pNjYpxbA6SlzbSkQAlvHssBdFZz8L1/tXn52
dI2iOJ5ryoejQbS3zsbjsjm875MmvGlYAiFK7WqvlEZk2IgkjQkrDTCM4lDLCqs8RbH9ftZRVrIh
2KozaBokn+KT3fqyVdRXv53cs72sPCC4ZlV4T8pY/lKhIkedUDiEViTXb7DMTqlxx4itjG6SyUDV
675zIxGHbZ7EoUC9f9Pow8cJRlBOTfs4u5u+4v1Y/RljU+YlrSwmkVTQCxYyq35gH070CvEc3ogC
vEVrNQsS6pUdgLTmxnphDLkDUqwJkeVwXXr0Q8FKUw1kCdjsXgIBoEJUr5BXcZGcUZvp8AzGb1Dy
PeQt8bTyH/y+cgpUy1N/y5c4n5pAO5YKvgZsbOF8zs7lE6UlCXPs+P4eewGrisuMz4tvvu/so3Lt
gwal73HIKg6MRMMLss9eLAdZFiGF5OMl7mo4YeXw54j4Q++31K5ydTArg3zNiEY+B9kSWoDelQyj
8x6kzlsduSjHVw1kKv3hMMymIgZLi4IqIJyvbLfXTeXSyKPS7YKt31V3TzilsZsFIOeDGmGD7Dk7
kY6oAnMu0jC+FgA+RfXfeYl5JWJC9h3jJwUqSzbHUXJapdlC0+T1yNhhfaJ1Nz72Jssf6pV+PdGS
jwsFfvX5YP1gKpFqKAxu4kS2Bw0cj9ojD/8OvCxx117BXdDq88Hp2ZT04t7oHvdCCNsIfWNj/U7p
zrNr9qoPeFhJni0MS/hnDxBt1U3x/HduR6ArIOiNenafiHZtw+3HXHd8Ub5YRpzAASNwbA70OCH0
tqj0JJc6FF7cZfcGW2G8lLV+1llrO4N3V/Vor7h0dBMU6/izVqSRX6F4ouQMJxg30xR6ifU8CA19
ujgjfHf69SRt7k+WQIdSgDFM2XLkkoRUHABehqwGVsjVmLxG0fJ9rbc4EfSq8ZE3Xi11iHF5l0jQ
6LSS9lz80+0B+msaJfjioR4SA1aNAToBP/ST7xqOYVjGZb+fqLhFHUtxHmuSmV/UfEr3OuFOAOc0
VAZVueqhot4zFV554R2G42oHbwDJsc71r9scwoyMoaB6wKTnWFIIwBdZqd8IMCefQdYH/vajhXjr
PpPUR8UBYAukkE0DPu6PcVOM55dcKxsLz07anKalR+1GEaftpJJGzZ9ul5/ntq3F7cXwUNx7VhOZ
awACwPpWuqucUjHMgrmwPFB+pt4IjpKUVGAVIVHX28D/ppkIhLJsFaornTGM3TmKt27qEYux7rzW
wrcPLWSqkxqRYd56KF8ZaqgLYnQk3npZ4jeWYdpL6hsj7mpWEK9O+DLn/DkMU2lRbwF7YdJ0y9aE
e7wlCmS+GSIJS2IQrim7RevJVftuCtxo6Ek3Fmrm4qKBuPH4YAQkCWQVJF2OGjizA85EKQnbOGos
ElP3nXT48n4LgOK8wqG7JX+zhnV7ksKi07GA/mvzC+lCH1aC2q9UW7RSN4RrtzmqfMmHl0Y2UElO
CVwhxOJkoNLcTQz9quCJJ0qZeQnsSnnOpjt8vkG/v8TrmTk7ukrbwaNecm93eX+zVVPs3ucxRzr5
i+aomU6e9/ke5t/LTLXjOUBglUBK2qfgqaGeGpLcTFk/3yqyVnI8GNCsebHdZX1lhd9pUxklSDXb
8SHMs1Cd+vuQ+dlQD0BQQBzBPefxu0VaGJg+96SWjBF7tEhMlxFP506o7BOHUOkVxKdNFr8EZMNl
bveCoz8GStz/xynyCnb0vHzOeC2JAW+hcpIW57brT0vWi8HEd78n1B5M+BFP3Ee1Pxwcj6DXYGtr
r8QSJTrFWnBZBvGlup0XhTO/nq0bWN3qc+s5OZ8XgAmxCAj/zA8ouB1daOmF9RjInCcDdRQnow+n
Qyw82xPm4flpiqIX0vpS1kl4sOlofZebkSZduuOyLxo0UOUaywf2wGOGH5PPnwKZGMGcpeHU2T5h
nda9dcLqO2kYapdgQygR4g4A4dIYEPMFl9YTCjcs84m4n+3YjOELdsJAfpPwy1QUvDVd4AmyVmBl
I5qu3++1sU/DeT7xNZ79b10dm9Jp9jUA60D1zZB3CI1inXn4+XwmcT6txS/moyp7Gc8f22mc1mc2
H2nglBlmr968nauj2rAgwLQwGJ1hbC5Jha/OLSkwYYnmF/HovK9d0oaY8Ap6Q4HInnjbPP5CHg4P
84NWNl+262Kt4ppDzGZSLzQANGCLXpkq4mzmAqGGSBXgiyQ6BJskycQ7MbqHV8BYQrCpAtvPAXA7
+1O/zN1peNuIYPrjOWRCrGtakFhn0SFs5ipnSvZ2fYLFb+EJ+Qt98JN0C1GaT1P9Wwd4MMLMuTlN
xGfnE2s81IYouQb2sE3egd3gkh09H7d5D8gLYb3eGMc94wVM4bTKzys4u60JrJWWHRIRvoOnCg3o
zMmgpl0amdj02zPYM7Q9oUoIGTpsRjejMAvwGmc5GaN4lVc3zXxE9NtMOshP5S/jZ4nClfoJZ/Qf
VHyG3S32j2ipm4PPi5HTY2JITemwn6ckb3KVf6KbAkoB0TqkL/wuuUMSXRdIjgU4k6qClvkZtiDk
4Qty9ayBghBR93ILIUDQum4HXm5UiHuthOQrC/jblt7B8jrJI1T+9etgaeZA5KpWVm1vnlyZKhLu
CvROnbRrU8vJTle75oF+nHYdL3uY1XhHR5Vo8WZZrOJQg5n1R7sTgcDuSq8FrWn47gIy9/M6AAEC
1Z2Lm++SyMJ4aTu/ytrmUPa1gnyr3bnYk58jTK+lT8JC+KNiShHLTodQakWFUPFofPouwpKbGvHb
3lVWjurxj7Yl9gFb1jHf55XvdFIeNQPCHwj+WFnvchfKWMRrnAiCJT1KyFOU/pe2fXBvyuwOUmJm
f31u40/1Fi+VoAmN5Ra4Am17NAFPnsHnou84Dsv6wR8Dnkxwipuejg8YSWBFdXGqZkSu4kWyaWnD
79068GHTGFn1w/Z0BC7c49mkU3DrZvLg1mRcxhlEaQioYfvaMiRVLhvLm0VGSbyVUg/e6U6twm6i
F8qEgCKorfzlPgybEpe505BWBjapI3j3fDNSXzf5DVcFRm3zi7qaNfCNJE2Xz3xrOngA5ipK4VGj
WZ6eAngCqYuq6GjOD84/qR67LMPTBnpybE2UHOUg6OfhpEMnC7GoW6wU9FKBwjtbFdYazo0dLNS0
O+oGJcXLGDfnnU6O8cqn3RDBDVZAbbeku6GsATy8nY4j63gU0WSqHmASjmchH4F83XWovZkdfZ56
36x4JJr+oYNLpxjyGuC5+cl/nCZI4ZVOoTc1FHv20/j1NVhwfM6r5gcUF3EVjRRqRTAUe1xRDlS5
etxqhJkqkbahAONgS3s+8k3eiOOpJzzduqB+siKZR85OcKL5fE6VVwAtFumRjIxLzSNE7G9GTui7
jn2zHfTLm6ZPmWs9yKLeO1q9jxaRwKgVyfhuetthMQO+YQoyScMwrlaVYWENd8P3QoqWWRinhM3Q
PqsMlxUETVOJQAJhFRixlTtV25LgvNYU4atxTJ9RPy5z7gtvH2rJ+JVg1l5mj9kjhDYdV8SXLB5X
FaVCdBo5PTQTn6NFBNXtD6SxI1cNxPLRQ/R7m2eT0SVxk2Cn5F94OieV+51gJp4xQr9KoG5hVoWI
+RHTTgodS7/Ef3wXSjo9KQiwKzH50sYljVTRV+PvEUCVwlSPwlhTFKJvDe90WTN9cL+Q+GQIHjc1
5oOt7GnS2zefT5VLcQu+DjGugSvcbdr5wP3aVKuR1x4JSjyfLYRV2C2pQkevv54hAt2dnO+RxXmG
/IlDqUlNwO0r30LHrqzKfzdfw9+mH1w8OmBmaHg1VnPbU5InPGtLjEZSfEzHH/iC+n+LKEZyP5OU
1H5zh+W6AxahnFUbfL41zZeJ6q47Wq1j7VKpDuenHlKIROC7j3Fvte+WFYGEDv45IZv8jWPfdC4U
MLjOqBMc+2A+cf+8raW8h4jSaeDqQptYaSNO6IVDWXub/lgIWNqVMWxQUOPXqXetH2Pxsw1rTg4b
TF8vRyC87KRR7axXnTltCkeKEG+tPy+dJVZaJTxRMSyGMjQGyh7vgCTZmeg8d9NGwInCD6Qp/KSV
oBZI2w4BxDS1AZUxuoI0FSecu0CXFeOzo4OJ5GD1/mkFTorNm/5UUqhHPulw5v1m2isbDrQRwnK+
kN1JUd/5usvukLnKlDTgS9xV0tJnA49aBlDgeZSMRlRVR0h1Kt1qVAU0uLVKRhelxDIIRkr/KriU
GA/DPU204qOpk9QPYsS6mWqJ1+J/kAPi8bxjJRK6sahzkCoEigxETJWHtWgplTI22LIPPPFRL1Am
3sDKIWVLtnA+V/nrXWearZsRz4JFShVNkO5WDBy1FfsXUNdy5yDRcqQDHKYYwjP8r0Z7n0n+CwC5
1A8mh07Stfhus2JsKC1Vn0JiP6K5fVCFzZ/ue5qfusoLaGZGrfz5jmTcLSCjhyFTPghveKbFpKt9
Cw+XT6UqvqDjhmTvjtlcAelz4hCacmi4sWtNvh5wbEO6S4kkIU4HMdARD57GuYqh8Z7Z9vhSMqjK
RCV9yjhO0YML6J0rjQhX+E0mh0IZBp6wL9v8lJos4RzmNsfM5CAenb70Ho6nxsd7MmlOyuSwGwfM
rJqqGDMSFtq1xV77xSiyYczd+rF/A2mkZprhc0q8CD+6Ocf2y4XNT58ml3yc3vEluR9Lu+Gexm/a
mJmis9hkqIov0pkg/vlfzmIsGX260ab+DAaqmspNu2dqF9vXn+OdZZekTmSm67sOM85YdcLyOZIv
SMnuU7a7xH2AjXlAKn3+dNHFd0HdLa+qoxvDJ2WNMcP3X8x4RPwk9ZKfX2pIEKDJeQp2+pJ51zpA
CzoDAUIJUdSM+OTdRweUsYSkZ4bNKMjmOjLR7zt7l92TX+ff5eusKEpC0W0yPjP+XLrMZnfINL4G
anYaP16H5A46GprwUCneZNH5tXd4UlpkVUbhyLyUZgSrzxKnCa8dfoSg0VAKUBh2r6atqQnAT/JH
NocTug9dcFxd5zpYCPEUZ+A37H4BTivydDNm2e+aC2gOfgjm888+2UY+WL79JGwEaFXfT/Xb7AiI
BJN63jYvKLxjob96Hwiugb38yb/GLfEwLzQxkEbJ1YKvLrAiKVfxllNmA+xBGeUSXcR1tg63zfBk
Vt3WOMPkTEnn7uFsn5qE+KjsdBfKqQXXfba97IXOzDLDr3iJNrWRMPkG6fU5yvp7K6FANEY0wbLx
wnWSmG2Z2JWeEtTLZBV5/5iRBcOLv/ZBxp9ERXwrq+11kT5V37U5u/9/FAiG7hh0gr06nYVfR6MY
fsmGN9lO/fTsITrhjpG7So9B1dKCjiE0MutJojTsN85eK+gBsy9SGVFwNms35MlCmP5k88HHVDdP
IVyzEBqF7ZklKN/EPjhOkaJiwD++AKK75TNkzTIuS8yGmKdBsu172uiSXHInNuq7VsnxRhUIfroD
EPjfyDUyldLzcKcYkxiXg8nLkFhTJ2Oiarp7gMtnhWuJoaio2gPmznm/NFLygDqVCnvmvVlEoGky
cWTUSXVKobqHNmOsddkL+Ij3d7xYEcyQhLtHTEKieBG6URunPzT3Nej8d4tIaUil7VIBVf3JX+/a
5swYnALw+7Itds3qMVx1T8AnmWeBnvGebKTWzNR+VSuf9S9ybzrOafn17xwVpMinL/XjwmaOPDod
QnTX7w62t0EpxHd7DsJArqrjB3JVyeW2dJou7O20OLOrG8MEFK5+kdC2Ocv9/FwKJ7Mds0d0UxnW
xqjSI6VkRmf8GGcKPDjkmAgV0/wqlTEhchv8qRykpCYAnIjP/2rIaKBRBMn8LfFpwzWS5UxCK78p
Cp5nx3vM3UVMwUSwFcFovi4FmCc5daPyBYPvpi835VxjFiX61AHpmimjXDTW0Dejgb4XJMoYb109
JyFFd3/KhssZENL/sbXqRdqVeCU3aH8InIpPJAxmmP2ddxhEvmtUcfx8UJmzn9q/tGz00TO8iJpp
cftPiflUIhSsPfXC7B1QfgmBLyhGigtPotk7I+7tZREjbJFgHiVCnPLQzZT/k9UlozjwDN9tYryv
vnhaEnhFJ7yW7dZQwJeaGJLfzL5L92nsoed82ewC458R3752dzeQF3y348U3OvEMuaGBjN7N45o9
B+0Ojw8+Wqhg9XwHnR9VZ1X4EBbHucao61hRnRefC6mlPtOnlxTt4xGsMLetorBvHMAUCn2h7uWy
5LnF8dhq9CKO1oi+ytNqkRWB+r7ZXImLtXE0NwuU7DJP5XLByawHyJaNt0JueAalj6kaPycS1Qtg
wrSbVgDeuf+5fklRn3F4vAyXhIZKBh44GzIwsWk4FC0HrCMq9MhdkHsLTVfyTx+lzrHP/fIG3ycd
PMYfY9wqwkR6bGoGAwJKQ8J9+Kyiv1kdnkPXCdRxYPzksJBToqdvKrziiBWlICjVfzxYdd+dY+X+
BpUxqQE7+CW4W1ftS9gBqqKmZkc44wCsuhGyjG+ofkDkpBBV8W6fX/IkuYmqBjQwFrkDCQPvy05u
5Tcnz7n3HxVs3wYWb/ab3hHBfISCzrlLpoCBG/sEC/zlYZt+bJMR3LGQOdrxAodpaEd7u6sjI9iO
GPSevQpLB6t5mi0mHD+semdGLJ1ztii3UefDiWYF/wv1wyhGeEmtw1W9pXx/rClMqqEA0BSCoPqa
i95qxKnqzxuKg/RLhkmcpF4r12agYrU5pyWmeUKyE2sJ2PLcT7Lao+p44lRWyK03tgrmSv2y7zfA
583nXQPL/vMoj/EZxhIm6Iso3cfjsWmIqWXAt4cK8t0LBnfBGEEeN/mC0sJzzF2cS5JCNSMfd/KS
Kx69+KPQ7OP17K9XqpyrmLurxzyIX9m33260yFoy5yPDlS9tsIaGFrdmytitQE+Q8El9N0EkAnCA
ZdDTEkTqoyAmkNOYalzyaktPFZCfBZwijVEKKnlzk6eTWFBLKI4jZVPZGIqW5F14GwERPfk5hB9N
+qAAdsBNpLiGC5/zhrz96BGRXXYFpCuE18C1U1eLw9nJPlpwRpNjOLx6lCV8STb3iN1XzY2kUtYR
TFQCCg9Q/W5NP9avtg8vWBjrWRq+cIHFizCWNCoZCgKMDVQakduU01Nfg51PSK4esJe1VdL/M1bY
TP/sU3DPieCOPhSzOYjJcJxDR8g19pm22cI5tJ83/EpNP2LrFCKV2XZW4IOfUxsMx/yP1KRrNz5A
fXwpnU4aeARtd2ltZuJq6WPWs2Od4RBXevMiLu5GG7aodHcs69Da1JqOld2a/bjpebFlxffcRiaY
DdLbo9DcrTbCv3ERYQxcVlrJiHYQdNeJZxpRVUD1pBhkODTIKDfPAGk67Iuyli8sxgys35qShgJv
q/SGs5McIdB79okirmOmNp1adbSBAw/7HexXPh+T+BqCuP9sl1y10XJj8dI5tEqiz3qkrp7Hcjuh
hSMIAMfb6QA9BaHTjMBBSaYgdpctDLEGgZuRKAB+6IWIbQ5fMjD0rQw6pSeM36IDgJraty7Yov9l
cHG47VYubsd5oTVB4MQRowj0D4xhLP80xi/XYGRLfs69Aj7OokJlFJ8YsVvfROE+8KkkWWoATzGN
mnlEUX+hK4E65uRFZaSkkaIvfcDhwSGnuI5S7qbBg/eom4uWwSTlZ4GlVBmNCUJSZBRSlbCwN/0E
MceUnbOGlYbXVBeCTQIO0/hnHH8Uv7YWWDf8L2qws31MNRbRH37qDvG/qMsPzLsnRac/Ju0bGRRo
KdKocbmtnTHZ/0GCI3iUsqCNTAVjDMa5iKh+57lV6yZorxvee1Yl6B6xkx/+FlC5YG02F8ljU21W
XOz4ME8mef5dlJfcUDXebTrhLt1ENXk4qimke3JGPiuanlZVuaHZvPRsVwlSLkahACTSq4x9Hqrt
GmhNCk5B6DblnFjJ5MdkJfXC+u72Kw9lJT5GZ9d67TSVK9rP3+PTRMuoF7FQ6Bw3gYZTaiYjk6eD
VbuyqiZjVwPhqcxjGBYKFdzAxZANnNkiWAybllRB8IizHgksBVSG06YlkuS3IfxquNcw9D4Mky2t
ckN5aLpC7HudZTI7CbOvZ8ajtVcKwB+vp8M3EU0pf0GKnCMAAliPDlSxlg3G1lmzOGMPF0d+zi9W
XUq4yGiTxOy0Nk1fx/5nOtUOKL+FZ7x0O8YVjNQklBQNnIywLbpXvFovmScWVAXV+Fd1II5rPDGr
FV7GKqQNvOV7vcbm9QEnQXz1dRucFE+/zIGUCNp59cb7LgcddWcOnUzTBPp81MzWcf8r9z9W8CMM
wR5ZotaibxyisX+fGvOFJ2KLo1yg5FLN89hLpjIh/iWyuzFij3t4xTbSh1piqUM5oorhz07KRx9D
2ePZdQK8OJLj9dfJyG83Czim38R3FwSbVqMGdYQj+lVMxsyiSe+RHh78nbo5fPwlGfDvApT/wftW
NewEkpBi5WhXZQfcg/tk8fQpol+AmCXPUuEQLZEySRDA5Cktpdiqy9SfV9xtthph0JfD8Y+PDhnC
I+753fOtIsrzFfxJsCqDYekYLDEXw1uAhfj6qYQ4k9tV1VGCvlG2nniMNLjr1F0fmLXj52uennBa
qjhK2mOrrz6sbCqKs97Khe+fOg09NU5tDL5WLyfEY0wMOdkvm6DGPRMjOcxdc8yGpKzFBZ/3iYit
NEMAwU51/6AZLesgAQieWQktbNRYofDrJhb+R3xnAlwSgM4cpkIaLI2tovTymcvbalKURn73LwjP
+Er2A2uRbmMLgY++0ov58/3ZNC8vVssJCQM3e78Dt3IvT5Cwg0ObztHYfcGuqa7wOFTmyR9A5K9p
thvh0q4rD+hSefhCj+S8PCOL7h0RPozh+z4wO+vslNZK90GBgmUJYRbRUIExAx7Ojo7aIoCQah7a
GPSejuv8U6xA06jG9Qw+glbs53wYnLHS31BamVYvvqeojYWmjKMC6q0EguHP/8eK0JHjAhPSFI49
irPR7zp5nbjpTOVGXr/vtfpdL07uW+zGG6HV+deLJIFRMhPm6yiPR1nLlkrwDqT6gUvCzqwBqTC2
8liBiuSlRyGTpgtxwC/YRET3zoi11N8omZpBuxrTKa8RVBfUcwkbOltb4EwFzSSooWH/QetFi/GM
c3ebF3mUKrb6pugGL4lQ55dxdw9aPwFFmCzoq6MIRHx/BZzGElnxQGyHqF9E5aOQjMZJulj1r6kI
JdPVotzWSNzEjkNbN9I3X6wH9o0zCad6O2oefz9HQzs61Oj4ZqG+zxM7vWcZC6kYLe0qCHU2lmVj
afg+735NDQ3aS9oZD9lo+hzLavbR6G5rVGLZS0G3tcBYRt8WgK4DqjiKN6H8XXk5JOxNlcjvTYSi
hF6uLUREIkS9HJuNW841eSnP3TaXdn1jjYgyBQsR92WBrIc8XpoXWF12n3wqH0+R7550y3vxQ85a
3fWzOpIdXWqwVOoiqiTNkPNNwLrecHuawPoB+Jkr1Zj1pZ44fo4D7QJ1r9CINQl4igya9IPMMPEq
JWz4xt5ypzF5JyxeEpnXVNgSqH5g4WwLhbGrmdlGXJqZBJO39TIqvcmboGPpoF6yw35g8UqEo55Y
NZNA54aiydR8Dl0/s+g8LPY4Q1/OLh8jtIf7NUCA4pFtao8RbwLGA0krC3rudKLXcrCyEQQQQ2oC
3Q38UiHOAd9NVdE13NGTbOnHjsFZJ+vcridm6+v8vdsmZ8CU1nsYxuQTKcDr6Nz/qBOSyAVp86BB
KgcXbxmtr2RBHQJ0bBKGPUDaRNXewjR4lLb2sN813KvfagRXq+pwfMp0x1FPZFMdmq+6I2Uv5J6L
4VtJDJdKZlDMqdfpgt4jIPCFchk2tg27K2GIJiRND61N9FaKFEzrUB2TfKcgZ6JbmIyZ9bjTQXrh
ChZ5gaLUgXLcTlrq0x5n+QVIpZpHQS3bV8w6v8ZrRlmjDMU61TjgYI61XB4z/Mx56ZtVvVonMutj
ID9QsOWTfcfx0iqVy1KduDc3ia5t1Vls8Qys3L373K8X+0+o1o5G3C4TV/OqNtKxnbiuZ1d3Ndw5
UmnxFbfvJRilIMiqaU9kHc2XHjpQxjxr7dL9HVMdDNCdMGGWqkrWpLWbXhNthVlRbR3fxN/bWemR
wy9xjJMZGl+LxkY954nwYcXmMTH7HkBwWgB5vlXfNYsGMD8GVsZJATppmudHrxlyxrGwW6oeemVL
c25NgNHdpM/0urEiexGMUQJM0JL3kHBXJHq+zKctC1W6FaH5n2hSPjD+X10bMfmTS2cqmQPh4GEe
sq6/Zs0i168dPH04lHcL+FFJ3ssA+RsnwtELbZ+Dx0hDMInSQnuGCZ+6gB4yJB4G2oz1fIaF+2gX
ApDlG0b7rOasVE+0SnOFl6GYYmq7uxHm3z0/BsdAIIMRKW/lPAS6djnYTNYXST8+icYYajYYjLEx
OA3o+77vt3hWthFxHV2QDIjiiXTBk2DpcdYo8vvLD2hthr1lzkNwF8kWzP/ad+nGkxU3Kpk72rGc
3i2sk/vCEpDx5zg+es74GQjK9YSb0fFGF20DVl5q0YPdQ0YWDocY7ztd4ZBDExanBtJRqeDwnqLZ
ujrVgy9TJJE4O9KfL0CYx3/MF1QNJb/KVt/IDswZWwjTvNBcvPeqIbyeegNrZM/G3Spmr0Fvri+v
wBMLdhv/9zFRpGSotrhDoUtLq20UPR5U3BInsVAxaXI75itEZZI4I2Qj6aX24yUmLpz14psfY/Lb
zpksQ2LPUspKLSrtiPu1b8KdKRM+mhVz2hDDpzabfUdxVqrt91vRWcjSYClvQyb1uiJKaAT1PQWn
2CdOX0rKpuezx4xARX6parcvY8yqC5pYtE4BGfF0UMc7Mv872hCUmbpTfb94ywGJJjhoPpbj2Ust
Dt2khbHZC2/rJ520H9lyGdtk1Njp3np1nXAe7Sj+PlKxzIOF0A8oBqT1PlsqP9Ybe8KWCxTV2f+D
coBoE8pIM6tGsQ4sE7FnMKY/Vwg8eGRhep36DCym7Qs0xVUgTlKoYljHxNmcxfD8roL8WQGBH9oA
sTz7WkvV9dY+vBva4W3N1DZ3EuI6Vp0NMvFqi0QDgYEBl7U5JgTW4wRFOBn6gcf3tD6PF+lg9Mv9
I2+JAcAQpm+CvIJR0jRZOTLmcvGcNh5BmYptN8RHIQWLdXHO1jD7FOIRZhO0aME1pVqtmfOuE6Xp
4/miip2r7Ej5sPULWv6g0Jc5ks+sRmdVwoTTUgnOpO0kP9K4hQvcdnclJB7UrT6KJtsDmOR6Etea
omJCgYoMuwHRUOZ0Nov1Y8wBBnLZlcpbSaNmfTGmy3apKa+m3AnGCHbHtKU7sJrBgzNMSHhVa2+M
H63mkVZ6Bd1xUsKjMkpCshRMkhy1i4mypGTJntepmW84lBZyDJH3hexBoL13zFYnwQ1IE66R01li
gsYycYaez1wMpGby++raTrRW/tWl77Q9bCFAmSM8X39xOPU51YGesfLqenflJVSF5794T/wr0xR0
smMP8SdmNESS31LP2KlrgsmpdOCNCTE9ep1tzTayWZdXDDNUKbgTUmFUBoSHlp+5wLH3VNfaL4eJ
TA/YMOU1ywaXmtVqWKxqdvNOhV97CBedlOUYLGI8WqYKbe9w4uxuDLaS4WsSkIj8oLZFDj48eq2n
6Rxc/3IZtUNe8LuO3IsXeC12ewTpLkNC6FEtCOvlDyqKlgy1eI8LP19oKDhOqqScYjLPcT7fuQS7
n3ndPtSCa65VRC5szEM57w+058ckDGAeXIPhBiW+aHjEZsdyPDPKRgadirMS5KCEbkxWReVBf5x0
1LXh3sjzD+n5xConFYYB5Lzd/1RT39CjJSQyNUyc4esxkHi+J3SB8CgQOM9J8MyTWPtHrNctAvys
Lz+gxm+6G8jd6C48sFbtx23GFlQB2dWFZ6QZ7psEKlWaoBYt4ae3NZq+JYid52baxDNdKBoIVTq/
7+BmouVpz3B8Ahtb/vAyMYtIXyhMwrqKBBnDwTzWoy6RcvVgwOTTgxi8SygdXbtl3N8wFv0iY4el
EEP/cq+cvlbdGpQog/EjlP1bYafvF8XQ5TuGyqyPYYdEyccgEBc5cGmJ9Yla6AQnTTLaOxD2OqC5
LVr3lpKnV6LjNAyTvjS37OS/i+i2/VeZIlwAO8MEwWpLUL0SR1ca1TZX831+Bn4dUr9X6g8JcdNH
r1LVr7NoB0dIsOAh+PcOh7kG+jpa+jyX6PCAO1U3dM3XlG2fSmDY7HBUlcJuh966NRjXTcY1eHI1
Amtgn2tEcwBVtLjOYhJrPJp9olGjdJf4rJvinkrVWaaqjwQS1YaP3JQ2vLV9UVDCl/Wn4t/mHTdR
eSyLFDSk/w5T3SC+ZwaYVWHXR1Reayk2XXorl87yRgNOoam0P2E1UJgtSmbuwcMxN8jZhfiOLuTr
XFrIZmy5fpknnq0sXo4kX5vxWAtW1MG+QQ3qpLBh3+Se9Z9ROAqNMxsSh1PYJrtvdU8u3DoMUWMq
MxwCcn14lCd/2jM7b5REuV7PmyYy/R9/zNVXtlcj0TkrHFIt1Z9OjWkl4XJmkr1IAjOXYD3p3NAE
65YyRKISccToYd5j4lASl2FcNmf53Mfn2RJEpk0TRRf4UbrFUVSTEkhcHNqkh92nmD6oZTA5sKEG
o4Cux7Efwr6no1KCffql7KXDsDpdw0ApcN42uTyNZrNFMzS14s7vuEEqd/X2aSGRdUeUlgWLRTku
Ttn6UJffs/6KilgMwbwRMUkMatmFPbsxFEvtQLt/rn9BGYVcjk4Zv45GsFWIlWc6u4/ZBY4rZ/EH
0mUKe5Io7SdjGP2Yq+gGhDO42MPRVhLDA2h8xBrcvyOh5Y1quTF8vfG09cJxP8+JVe3t3n+yzD4+
c2QWgKcG3kWcSrYvNhRYWGSWiON0KvrA18o+8X18W3EbpuOS0++Y6D0L74w1MYNSrgPZ0lIhO7YB
4kkod3sWlps3hvrR4YVBnMwZMNkroS7ZbA3BqlAHDBQBiFwvOjiaR4Qy5AUrXjGNGcC+dXouJ3ND
8M0y3yhrINUPdgX+0586hP2RrLDprwTucdEqOshYtPp/r2DOhj2INi5oCpBTLIP8Hykwye0v6Sce
fI5nAgikFJJKRt/lXYoM7dFTZIO2y4zpPFJJKH6Vk7Nq9DYtnSG1dsQLWqr+VPAKYVBfRJ53srSv
TTMAXTkV2oymOJ7FTerQHTzd2Xb/uX0kwL7YZeTasMIAtZ3LsH9JsSC8y5dI5s+P4iTkqhkZZQhp
N1XV5HYmyFaJuw8ZiHuiUTuhB0B7969sHG2rgG/6TtVp0z4bEVjiokGsbkkt26WJWOh10IJoDCI5
v98xiOb0i8kvl2km/SPjWTWtkz+QkGp3DgilruZBp6QrIq42gv0IQIsScyAFnmF7ytTT5dK3uGdU
05tR3a1FokpNuz68zcPekAHSElvQeHyvfb5nuKiDLwzbWP01Ns09Xorra6EQzB8guJdoWUeYZaBb
bvDZVpgdKgq4nm0ugRL7ASBf0PpOaSx55lbAoxcaGHF/dHJ1pdi5rVEk4vYhPYDkPjBO6jlXVpos
MpAq62/QdN0SS65faeHAyEyxNz/JtZuLsNXXs6ujElOB0xfy/XWyby+mw+gpJE3LCi5wPDEQavzy
lwc7uklToJbgv+UIxStFkMLA64mQAzeT02T7RB0DJg5zgFa+065dMg6QfnuBxEgxZXq/6GtLwZix
z5Pnl/tOfn9PyPaQYZInObgbhFs/jJBdwiCfHVcZjSR5P1xIlO4Mo9iqfHixHwIMWa9JjEwOZSpb
akRXBEE1YtRbgexF5fkO+Dx3Pnvd/+UeaHw3XQwsSSW3Hr8Y/vHyEilINelP+uJ1y9L7LbmtkFbC
9Mur4LJUFRzWGYHGzh0UUZBeOsCrVz3IR3UtVrA6rA18rHCSDHrXNyAGs6z8C2wPBnvmo10RTTgz
zf/WqtqAhaM1uePB3BPRiRdVC/jq1famiCqEngAMjFeZS1LtI4vK3cUF/GNuUFbS60mOtFSaMsC8
P2spm+HBNOsjGYUF3/hf/jjHndH4xb+ZplcLwfTOlm+Mvw3kccMl/4LYaF0WTbXG+wEWAJxR8Zr6
puALUg3VWkykEUb1OBjTHLnFSgl0iWedvvczj+58fepUixY+v4ucw1io89iXrO1ZhHPEtwsiZ/EK
WeEdiJRyoPXleQDZhE8IpFcJlZGtJ8zEeodZrOsE4B1oYPisVXRTLafhHLwkddIeinU46UhB/kJL
764BeIQPmnK5ODKA3JIc8Q1zhGS1Ekc3s71/jxxuFZ9Zl8YxRdLtQKFPyI90fuWOetEddLyA0bpo
DuqgBSJqyOIovhsuOXjWPtVjSOoIiE417VVBVa6O0jWx08nceMxZPmEGW7nG6x+fjYb+95J2fbnD
hrsNvLxPEaTn37DIFyy/Qg0slls8Y+h1hMjoEpQAhN6jHtfCcs4I6lLBPx8b1zdYy0m/j/ck1z89
y/pXRXtTtiihJ1nRWmZgwfvruFZtI6yHPruyLtpRRjgBfI8zeci0R7b5MeMMCseZFflxGxrFd8B8
dAVFRZkvvUnSbEmxPPu3xCImUcguE75PWUYla3qhqVBs6wNfVyDPkNqRezkkjLy4gqnpigc3FA4y
aMg/CvgYbWBSU1s9qDNUshUg/hMndX3+U7O6/wcyMgC/kM5hSjKZnbgMMtFtKYfXxtPXSH+OLAsR
uPRFY6FCXGxuhGvpHOAfpkAvQ+bh897DLfOsRhzLPbGbNsQyH7CfUA70LB2jXVgvsAEK0AQ1+xzb
rBSd7DX2g2xJoV6YSTJOoL6aHZzrMQzJbd2trlsI8qE34TK2PhLYwYK+Eibw7vcM3BWO7CaPKnWu
70oN7CoupxH1v0jPXg91xtjfXmvRCVfv+Te5usOWLjENVwaKMCiOv8hMUOQMMXxWy2jCP3QnZTuz
+H/9cOIlB3fQj+ZPyVcjwEpiwrE9FQwqOU6agWSl+M1oLqAjJmpA48HDyhdVTYTELx0iH7iIvgt7
v53I0n4gS6AYeWjpITev58FkKUkraOnE1XjfhbAHFMhF3nFk4Sl2XGNryMSdhcg4SfGxzwCRjpuv
2ztVH3mYmG9Lx1r22x0u2kObVmksOb9mokgE/cUzCH0nXjKWdh1Q+0u/nhLfkgHLVacx8BHHGU2Q
gO/qvfQj8bA2KfybFNchzcmbrQGPOqU6mwKS2CsxDneihukQ2HCO9msheqYFLox51Ke8sS3BNZBK
azzyVejrfz82ijskXpA0Aq6v3N0xNOdg/bl628RgguJ9bcQUSs79bISe2tcmV7DmlPI8mZlWty/o
KJ9szWUG77huEHJGbX7WtiO2ODTJB7OFpGRQJ/wqJec0nZt5t79divrCSxC1oT8Sv+k3Ptk60tiy
/SxuryHK6GnXlVSwF0ZzUvivIRBF8qcFscjJANfYjw8wr1hw75/CzhA3sZewheUPMhq9BPKDjaj1
/AC2ieZ3cCB5kd3kDsnkzEhPrpmN8Dd+31O1dxrSMnWjuO5B7fgz+St3lgUdeQlkyxh4kK1Q2uHz
Fe3GevrMDMyRhbjA7id83XnqLUFsWDw7WL2ppSscvWsXjGvlPSmCvF4U/d2nn6PcqvEMA/exRWfn
5Fj7kjzuTGk3/5Fj7pqMuztXlyxG7al9xAqZQSvA3e1lSg8MyNCKveszk1Q9i+fo/lqaovbknf1n
cSUzchztyO4J1467xyjrTj54BvRIYjT+uSVR5Pc53TNX93uTNUQ/8RpWRX1M3SJctqMmqikOCJgE
VVogxQqkUj6AJs+AQd1+ttATyFFlZMdyQ85UMX9rYCgnoaTEx5Q2liWJp3fXKAlHpMBbGu0Bctp6
xlh1mlWAtiIPlq1iEKyBfXAnW775aY92Jm7MrfVbHYBjObdnOYss3Mx0fG/0aHpuqQRhb/HNbFo8
iFAEgHZZzwb7ygSGAYe/d7eu/kWiZvuUSmsO7c0wKq9XFx4Ay7cMxFUOqC1JjEZYLVJ3duIkBSqx
LQ07SfjwMfhSlpfyWwZnEixmQziXICDd78ImlpOloiWsBgUPA27KWsqY288GDWQSwFxmC80p+X7X
vvQOR6AyyIPo4ZRowoqedNN4ElWPyPocUxOn3E3JJg9gggkQH+BoV06cm7tUIZgPVBdRYvHMAWKF
KRvAQhmir8h5JvkGED2VIVtVCGUgxAH4tIWcmwV0FOHBSoka6QCsoHEpwtMv9D96skoOK96RTons
/TueSoqbyMmKJflR00ExI793/6AC3PWWzp127aFsfjA/djLEL6N4zE2WIcZqa1Ohp+vPkn9LL3+g
L5Hn6MUJhkcvGb+BYnkqlG6OXMkCDrn/R4yy6Q0sc9HgFPHSpX6kUj7QaHA5phZY7CIx6LM7+4Fz
NHiFKQKDpJEAhpOX+XWVrYsVyukcHcqfVQ8gvXFW5W3FfoXlfeiOrrnh6J80UFX/H5EeEgv5UDEu
6MtabHoiT76pOSBidfsn/YqIiw0NigiVhRd+PQFugZrbPomXYgAj5ABRf+wCp1QUyTfwBusSxpIh
N7VKREXS/WYv2EA0AW/lq1j0oIbsW6EznpOjGQgPIOAI5cTIsioYBt3xJFLS1yWdklskVVhaSAG3
rG2Yu/lZjiX8+7RuZkT0MaEDI1fXeoF2YdyaLftXol4o+u2bsz0FOYacoxrMxS2MgsQJJi1Vi4P6
nf9UqLx+S29RHGd9uLS5L6EXSOxYnXXtTcEQ4i9Tpz2SVCv2rcJ6WcCD718aUIjDKJed+NmjZx/2
h1M9uk7ki8QpXwfAUD2KAf2MJK3SfdqEN5eO50f3i9AEM3OlXiP4r/qwTeiDkq4I93JKOrY4bPWm
dyK8WAj+CQbFPMVq0xGgP6ecjxiloz/VKQeGO5o5HHBE9WcbvGUihJpMU5JbI6oedvtV8tA0J6bo
nfsiO7ttOI1Pok+85DwHpq4DHposOnwl1aU5qCJtSeejbj/qJYyQQGkVouQ6gcAq/2NY7T3w5fIy
+k2tvmnExX53Ihc03WoVDXlr6uq+byLpYaP3lLzPLIdQx3VVLcSMPfA9ORw9be58RuQ2Ul47Yb1l
hL7TET5zVyoewxd0M+NHM8Rm9Q0IC/Ng/S2fTdArje7zYMn6v6QUw4+iJy7CYwYxRdglOMW6uKSa
1WvJscZKmDd1YVgICfLwZNDuW72xrRq2pOI+P3BuKsmNPrSukfjUk49bZokOCBg07Hk8Dte+1i7H
8ayD42ypN9L4SnpMuD/g41S7GmMGAehqwYEcFWI0pZVubvrf6sAmWGxm36coJw5LGsQtTYEAHH79
RAD8Kt7LIKlQmtZ90/3pLsSHsZGafTVJWy47Ukuk8xyTjs+Cgd/fHJsUirk74sK+tZMY8pnOJ3IJ
dJJYXGmkP0H2EOxXlWg950i9dwgBTB6H7V9lhrmm1SWcVT1LNRga3X7yQkGKGd0nWFjcp+wrUe8x
34ZRfKmTALrE4+YKGqtGLqk9agWckIoLygvJ1DAWfgSMkGESKfKTzqnDrfTHokhCH7PhPYrG9LDb
A7Xmnv6WP7tG0Vj/U1MYoDxXKyCWQgV5fpmuG+4YG4u6JvwbStsAdl2+KYyFe1xlFeQJ3XmhqmDN
qFfVcQh2LQNOZxQW5WxcvU1Ql3gWDdI6MttzbqzhJVmzPo5u4SCnngRpke0dMIZ3+iIrgWXYipnI
3kTtmcZYj+e8JHsvYEWjFoJWfBAr2hhE0jsfrS0RG6Kx6EpPbDQ27fEfOnnokr84qP0bYofDw+PM
oiyUxetJ55eLVYzoTFOLnlcmvIwY+kK4Cgh4diO+Z+aQD5329RZxIuxyJm+5LJPULvGizmAYF/3+
bSZ5xGlJM+pyZ3Hf6TDoe9rw4fpdu1TjL6plY8gbNPGhaVaA9LWArwti3A1024OCSeFddfIPq0AV
ntUwjkpoztPFMBVnzJ29mjdd3Hoo30fVA2Hw8VWextqz2DW8vs6RHrEKKuEWYLJnc8lZMNOiD6uj
Nsnis2tarCAYb7NJBXtNbRWeEUmTPkdOTnOpqjAMG+dmY/KPhtKNpIkgDi9tD3TiG6kXG0qsjr59
xmA+Oj1PR/XujgaICt31I6gYUkVArdj1j898oLW4UGyRo0EuLAnk6A3vjQUJbmsFOpj0A1o1Cpoh
uxO54Czw0S+R+GqktxQ7XpaGzPQNE36wB09o9DDzsGPdlTjnczph1FrAQqgjQf4I63oyC1MrIgvw
ewiGfzH2SSIn3sFbIxTnFbyPE4F/u8/NhGP7v3RAxAbIgAFnRwcOGCVJUYBXR385ECFWYOCLcxgc
jFKmRjRsL1f/SGKBOvNmyr3uD+SgaUGfm4saCSKIOw7aTSUs8zUaQz437EnAi8VxivhDWmHsIwK8
GhS9AnqzdjnCKbHokHLHharvgErTY7jG4T56UuL/ZYlagk9FHbLu+dUFeYakYDiYLo0qXSRM5YS1
CjVLw7scBLSS4WZvjbxMn+jkzKuQsmyOWmNzRnCOMaSZj4HaDAXpbzqAJea11fzwfJLUJqXem/AQ
noRfO3b2xn2U68zomrRBDguhhMfLseW70N51WvIj1CNO8qPbMsSPs/qUWUx/Nx14gGc8O+p3oscC
gKnMBd48wm7ZIliD92U6o0NmTPpEUU9Sn54BDfrKDUUSxGiplcGFvWL8cMKpDdF6mAAdK79vHvpZ
4mMQ34t/j4JO41q3edyt2bJcj/77MxIoSQuuajwMViY33x7ygnp71xrOeEz+boIPO39LGalGpKbV
+2WCjFOmbtHNg44IGYwlTgfKzp6/+3ur7oKOKXK4xNb2GjF7Pteu1LCj3Im4Wqyqh1vlVUwhm5rH
Suy7pJ4Il30mGBSwlpPsOZffGVDLKqjPfBfIlMN3YkQicHLlH6eyR/iKArucI5LlOJgNpq0Nv3nb
zDRndVWx7xA14/ftg1IwD/c6oTOluUbFpVg1kbjevYQXKq+/RpW3+V+nOkekJkey2lPKXKQdG7qW
DEzWrC0Hvioo1TJw0CQrN8o8MajAFeIo2h5cMDL5+Rs6XE3xhfaZZdybetyawanLO51AwdXacc2y
Q60ZSl2Rb+n3/O1Iq3yq6aXArYvxMcwTxRVjNCkdz5u7eFuW6a7EviRM73fhcueRuTc2owwOt2Ww
WP09CN4xYmjH4/dmxdy74xBJ81IS3X5rDcJ40ssg5dZvpcgjzBGviYQrbwTiqWOqRT2PNfea6x+l
hvCwJeiOEInvgBPuc81XzS+mf74Lw2auiaJcOstK9j0PSxZ+X0l9/CGuK+toVIfKE5zJcpkx3npI
lQxByJaqhyMqfxN+wWiTJe6iQzYvNkUpHcNKdp1THrB22LMrP9aR+8Z6j0hMrAFcLbAiaMvkZvHK
X6fkMZlpPVj9gvEgfgWu7JznUS8Ngz9kbVQDiw+U0D1bEjUlUTvIWQbxzXbHNe7XkEKTV0sqBcKp
ES2iLiYZ3zfqE2AgbTwBfeuT9UFm0rgozcfVnyUuuUuhVw9AmiUDEf8QYujjrv4ujasM3R3BlFOv
wgKbfhjWzQj8+WhxAAO4LBwNC059ebPVZ0qJCWdd+M4ZRFUqd0viiE1QzfkEp3bpq2mG5iDrAAgb
lg78T5bwoRiRxxiWJPEdcGyx1Ki61zeGLh8psfG8inpEucAx5Z/dtBaEvY2B7JPyvSZo2KkRV9jH
mA7r/9eEllxUgRO64cIFoMkH9Bt5znQ9LMWM75VaGwewJde3YuqQbWlJUXP9AP831ZXC5TwdwXlA
+DKPNtDUSrJYnyfAxQ1kx2wU8dYTw20dIzkdFnat1Lu2lHbGVGib3PffWkARMAOeu7AXHkwMCULS
ulJ9Nhjx28HQkMehQiY3C5QJd/X5blqauDMardHT+ByU1blxabN7IxBNbCECAZSdskJdj0pVp5dk
E6q8XVv/aWpayfogzGM0Py8egL8p9aiX0kRLv4VM9bpMqa0a8fzq4HBexTtlMqW7h41GXEjDI3b5
v0RUQ2lr7X3b9FPFcbpEvn4SnwCUzWNxUiKl7U0BTBcWehA3hN2cci1Kbe1M6svVaOCUnr7aPLHc
2s5L3HUqjtT/qjDXK/2C0DjKwiWMnfym7m3orfnL330A1pjddfzUbctjFva8zjYarjINr/Ct62ua
N+5xT2GNdRb7KG5ouiOeRFtN/bUeA9q4ZXT4YzVjk/ObQ/eKaa29N9NYCRDYxIWQVfbRY53JSMV3
+89wZRfni1YcuTOzZ6uvmqULYUfH2fkeAlzwWOvsOXVrMfyalb8msoDiIVNPPSqPlMkjTR2ZcNH7
yXK0fBM1POa+3YvN1Q9NdVqLgpqkvjKyCk+vN8aCSsc/C4S4SoZv+nkr05GNjnNCzY60Aa1PgrEL
ycKolrUp/YZNFkZQdKSlWUHZUpaF21FWf51e7FlK4U2xC35I0Ti2I/qfM2nqFEFvQVCkhq4pkR/6
ALgfgQcir59/hM6aLymmSa2y3aX8z+dsvXweRjfhCHcCT1cuUPKksViyrMAXxXyBOq9gfxWbjpBF
9piF8f3qqwu4He3GBwbpBLq+Bpe9A4GhkRJfakiPEXINSrROjv+EdhMP9OZZmJBP5mMYEVbLq5sl
iDoEAwwPZ1nEiU47MNbh2GU6oHSkV4j20gzbL4MVSLr2vH0i/2nnLvR2ZwqxR1d6ywrMMfp89oaC
57nXqtKOsAfehMlx7TnQFqQOsV3BukosFEPUdA6trhXxxMOPOe/SHa+cGyCEeB/+iXFjmWxwzBqj
XrdFbEOhcRQqZGzjVPcInd7/ntbaQI9ufmqE9UOlhesZeJl70aQLcQvalGrODtONi2vJoKbdSFha
/L8G++5e7NsKiXGbn1DcpwgSy73Wlj0eEQfWvU26wTSOO4zoXyGhWI4yxg6wC9tse6cZ4y4+M9Q/
4ZOgZnyKa85A2DiZYioMHE76avrJl7tkzyYquLy/Uu9YSY1mJ617fNBF2np4S5B6nzSF4Xwb0YIv
tvFhUVCm/g6D6QiFno9OdlYAfJmXyErpW3v9mOXxaYWT0nJmB1d+Yp/SqXsain6ckwFWbLfe/6Xn
sKpp3dO0dy6yBZu0yMXrdCxidvJCAhheHGyteESQXcfigcJpfKcGk1jT+Z8eWkgy90H6JxAr8soQ
bdS1KYyLN8BcTTC1ECLbde4m/NQ0FPHhKf5SbQD3OLTt7X5faVzhGBP9tjanryBtyV3QMfY7gddg
LZv03FDxM7Yf/VOrYTf8U5LXiyscn+RTOsiL4RdkxYaDMV8OPqzEqk4m6ye8folKsXxo2jEmxMVH
0BPqdwNQbdQy4pRK78QQ2XKtYqeDjnifGPsN8CFnOe+bvB/DNCtRq1dSW1KnNosJSHdU0fd4+AKB
/zInQ8lCP/YehlmZQ0XLvaN4qDg+AKaXIMPim0LMrgJy0olTRYo0yw46+ASACL6qgmtgQND770Y5
6H4k9Qym/e3rNgnrWwQCImupYB//kfl10Mpys8oh4mGIRl7AftmnVwtSIhk6JsgUhjJO/qX0UyAJ
/E9ayMgYASYZs0v9vRaR52uJ+SPKYl71IHFwq5VcpdWPpgVEYKKsd5XqiHo5RqCyEZwAjmTvjUTd
ZLA1ZK/aBKFY04Oj071XZc6qj5VLMTcv5MrIS+5Hg/0xLMa1Meq3vBTqym0S2AMgh9jhdJ6e6klv
LAtOgTtbdkH9mkOKiSHHVcB9eN7CUUGmQhLmlpvJQwsv0zGnH4Fgxr6Wsg1G4I7ucPSShTpAkmgZ
Gy/Ztko9zqxkK1kzomfqJ0SCUMywyQmc1exZL2DgeG8IA2W6VDgpRZ5nuAxz4N+ndUIug9hr36Es
XF7UQx0notDoSqgLrQx7054r+fdONQ0mQ5gIrAiFeCX4smU2YQTSd5meIKsEfUDhfdIuAELZuZRh
cPixG69Kvrwoo9RnnTLB1UPXXqyF8TCLBY2xhBCvVwylkuxW8NUM3kTDmtbNi9qnnZ5iqR5Do0HR
+O+WghMM1jfBR28vaaFTZy49jgzzA0FQsJMNc4GOET9NM84om/GYsTtfKKP0Nwh69BtZz4eWNOLm
iqNi8FEhnTqjxnUYEfWu+QHXQV2cxLXRrSXKu1NW8Yd8zBiBDKJ4qrnSuuCVc5pb86PZhVyfjk5h
Sgo8p6rFnceyXydFDv4kGzmCPxojdh8o9c/yevQj1XGmmhKe/ITboQYImQVQZD7GmfayZK/Eld86
7HNfldRL2rqCSYWHuOw0ppYH853G0cricKkjDDGdDsj0vzJ3iTxgGocQPtqmF5A7XWpC0BeOWYTO
huMGLXXBcFfGm4VSJLlPFsK2sLNIdjXqQznnhfBiYt2CFhG4MCgM8Q6ZmW9TDXWvlsGKou1v64Sx
apfCaprHWBPyfmnRBkzLdm+8nP5qGuPaxrI3gzauglUtQ6PG7GXOSGJ1wbV58DKKHMqxCpnsiQ3m
/uFky1Wv6cO9D3W1y9cwxuSPYtVoN9+AleuywQictG13VIJLn/eFfYsPl2zEHEIkVTPZTPQkipdb
Uv9Vs9V9LJl3o7ccsYyoE0b/+BMp38g6kbTELbJkSFNtSUBgePZPSYAhL955oFbgnfRYQ1U6rc9F
7aBcwbUOauMYdQzE81A1hUsGETQi0/IZbLmkT2XCPHsAJGRgkGZbn0bgKI35yC87ojd7oTyAVbI1
oOpCWl9RSvAczvSRx9zqYWoSbfRBxBameXdwfLUc0NpdFFRlbaqTw973/vxY32cIuzKCIz7b4j4C
ia/6cFNpuM4mbRzaH6OColTYq5oSWfNHFRvg9/ngyCAjMWOCWKokZ/aTHtMsxQCd19inVGClgek9
sDHifg3BFm/6pWvrlAnx+2PXhrz8acbuVR7eGnPSSea5jqwunCGySJ9yks88Vw4N6cgEoU4HVRsB
68CNJX+n70tjsmDxR8zJOCRcnXzlul0ptBuoITBJelaxIBP6/itS+Q7hln3LV2IDHFi/jVmbxFYU
jpXfx0zb31UhN8Yxh50LTFpDzpcvIIUPO1+igytjKnL4VKeFrlKgEd0VvbOEgw4vprz+v7zy5UDC
/Dyrzr277Vh5w01rzZmJxAP4Iah2vVFoC1seeiNKm2eJpxMvXx95px0HW69E9b20VvBJGchpskMf
oDCdkG5pOpxqskPJ5DffWeKLPcbH06G+u6+aavTrhj5RwWxn9wBCMsUGVxTOH3ruMi/C8JQvp4zT
tYHYTtfrjSDDijkMvTwOJkjN0TsjEue0q17OQMd9mcP4XTBmYuG0SzwU7jxRJmS/DsnjiVFdYI23
XeSKsIdzM4K+XVpqzIvkULLHTnFeJtzIKtbgA+8B8TUnsDe5ScedwSbrim+hZr6oh87sKrOUARsm
00L6XZoGabXVHqoIa6cryv2OF21bm2foCjKmMIN944TffDp3fj9lXF3ycESiAz6+Yx6DR/BlsBpG
DVS5UiLRXlezkjqf3XXBNQtFbef5eNBWej12s8Ct2NnKH2a/xaY3/25WCQLtBULi0FqHQ9n+Dcuv
cGBXIM71V35iLYBULVKP4Sd9EkmsEDDPNg8AMQbelmBCiHm02mW2hPblUe2ZmGh1flXKZDy4qmTG
PBwMlJ90xGNDsgZwwqkpBN7mHrKJgIbYuMsICDBbQTc5DM0pJwRxEDrYf+eWahqFGaAawEgHkgd5
drFwsvleG3JYsdjoyXjRMM/4S2yVba/xU6pWQBeoqfd2sWHdm5pldxXkEjLJ+L07cJxCY0hL4YD4
xuG6OZ0tBWazuMoZk7rYYiEMoqy9iJXzC3RAciSwSniP8QxkV8+t50WkuFjnirSKj+fplg1T1kn7
RUkUqkRDliLOAHV+Ai/JrJw1xhKUjGwF+QsQlkGlSCwe7jZS4Sl/BILMfxWEguwc96PMB3OFcPsx
wKJNe16veRM4yPS20o7f6S1gRT6vR31S18e+/qXGi1tfnWo4Lq/tZaKzWjefG081ehVLKWWBi08/
XRoizvkllbfRjJ+/25AHURJMeVa79CevM9/uzf0M+xb04gQIMvP32rwgrH+Y4UjvdX6jGEUX/9nV
5usHRbhkfQcxCRniR5UFw5BLvlVHRcvosqRfPvIAVpzAf6vY0aSW5yZEHoosBFRdIDpbvCE6mUOZ
RLPhhJ6gFuOfvWqsfCpNa/UZo2fSYxUGUMKhhbZWQGTw5Qq+brQLAIrWMMPo2mOfoMNrfVOmQO55
HvBcdRwE1zdnDgn39Shkw4mVPY2FR4YHelyZlyCo9lgB+TJa4LBeMo2Yt9W8qv1u7MRSMB/PiOx8
r7DGiCFE8cGYBIK7k7DS7MF1Lej/yDoLGc4bqdRXO9qOdCq2FlnNj7OrE5zz1JoJjFQmqhPl+nF5
7Rl/yvBlHrqUr6JZNzPpcIlSvUkiCwV1kgeAu6JXktzdhKP8rt+ym8yI0quCv0xRfnGuLD+qvyH3
lAxWdIrdqXNfS0yY88+6aqVZDaIwcrKOSwcVlb4mV6IyZIZ1MhV+20qHgypVChEo+sQBbSteNDux
HltrZ2A1wHXDAxdmkPo53NjUWOJXdgcQS3Dn8MqpP1nB6CJ4MsyjS6RnDDKR92/Xzd7vuHHirvdb
qiYNwvxvuFINB2kiCdYG+1eJXS/15zmQeG4kYC3qsuoUYzxgn/k7Lqo/yV7Wd9APBcmNGFz6qZF6
fgv6kV3yKNlBQg8mfcdaGC9WosdcPrqceJd6PMB1lpW61/Thj5eukiLQYSUgBufPZfbpRjbzYWsC
aPdtUf9pc1NFLYE6NzY8P90yrsRpIdqpsKDiPGRMg42/OwYQkkcuc+7m6rTDml3l5oxPclLbsw4t
nzvPgQcFQoqLZJpIE+b6TA/fwz38ztt2RGeODnbe3V5wGfRXWOcZAoaXjBslJ9tivdTYhnwS/RHg
FrUF0gL9FBGerYLilOqBaGqCFV29Ppqrl2PRwAvxh3YJcj4d2Wvt67wzjFqq8CUbCRapj56TRLgr
QW0ecmfi5sIJZWGx5czdBLdh7azbx+1nzXh2BEpJPykJLvV9r5MwsVzsM//gs/tYTsXyuow5KfSF
QaHdxlcP1Y+2hEY73sITZsDlaYT8lEHS5N0uq8RuXB1066XHtLezqoNGp5tBcbS0nmrlumY9Q2k9
f31SUSek9oVRJF5yVlXxuOroP8zXTbcUEJxpqWi1sg6sf1Ofu8AlDmNIQkHLE1n0v5pzVpJ3CeZg
1ZgYOYiuBSjsgnbD+Z/2CvlAfOO8iOMAeddF8Lpx6JlFZXhc7bqS2oLMKza/LLn4FTphZj9uWdvi
9g99D7jQd3s7mfWFQuv8iBtkb8/mu0Vrf04AagVVmlvOUVfkZQjaV3+6jEaEe1S7GK9/xo0H/M3j
+Yn4vVKLlPF443xoYWbou/USVg4XBDu8HAaaApQVVxJkpv3TBhGwRrhETR1NpfRUZ3PfZuxVak20
TPYwsJ9GdFXlHfeiSoRahBqAzWbGcMIs2MWi+A87WjIMCzA7Nw/M15ULcuQG81DA11gGMiAY5E43
JW3VzHplweLgjSuJe2t8b16oqcqFT7cIgo+7a6vj6tjMbg5pQa/o/4oaA10kq0u5HeLtaxSLGNQq
Gn++acjgHdIuXTmcsr+yU4N4uQOb2QxQ/zdBeKyDJNy87AeOtDPbjCl97apYQLsGADTOgnAjs0hX
8bZA7rQwMk0aEGvqB+KB6G2XxtWrK7SIR+voC6vxzPraYTHGr7TRomoRlyJVZFMnE4+8rI+SRr4I
p4C0J9LwGIRVgA35wMxKonDYWKpm78AwbUscb+4mNdIRG1gEo/Qb2jn5l9E7CqHT5opJH4I6/4gg
5bKAqI2STkD+4/2uc7DHY+TtZLdQhynWtXyU/Lvm+nGAQaU4/IegQ+LPYd/aPJl3Ek4FGxJ24dff
J3x7LN9fRjV1doz2uZduCEWxFTPV4MGTyvNYHytWUC23G6V9JX/ZVGeNW0LcNNnpm6nRE4F/WBJ6
NyS07YdqHCiPH4CQ2e2SDuiyxT/RsO7l1uUS3ViA84wtXczjX7wbj2y2bGTCNc1CqjDlbgUnI9N/
/ACqoBT8ukWhJ+FKq5RtBATLBthIU1qgQMH1pQJ4BoUC5AKzD7RcVbelhNSTKsxaIHyj053Nodit
ON4cwlu+pz0U2XYi6va/HtPEGAgJGKohrLO4R3sFJn5MymZ6/l72MUGHuCxcQLrCDq4iB7H7ze5r
ajs32MpD1jEDAmipAjZ9FUiC754jwINw2sRAQ5K++Fp8VG/EvvG4879MBHKrSkrz0Q60FinQuJan
VY20RNLwB7VRWJxcyPWnSdUCn/uScMvrYBrDvyD98sVExc7BoBGGYA/nbgcHDkqqbAYz7adsbBpx
CLbKUFJaKJZD5WgpcTEu29JjaEuqNC7KzgfaR1TtiojTO6luXlk5LPtX8IwFXTTnj+Cq/Ctq3uyR
G7aBxG6WAaNOS2mRw6KO+DHH8ugLVi0QyvU+1X0mbON1A/gijzs0Sd2Rbxi9vWbs5FwNfALmd9+O
nrK+Sb3R+im6y1d3Y/sINh/ojuymbQ6bQC5TjJwx3PeP7Fs2CbPlKzVTctwri8jnnsHQ5E/b4qnd
MbLNZbMVklbky/b1toF6iRTL7Z+9SqzlxgDooUjGdw7iUg6WlNToRWh/rke3IhZ6agsaq6Qkncxx
phCl3faJXN3TaxvIMubYcdPetLR+gXXArfwYKV3OMLr5xYXRfGbD/9EHOsgwx04aQHAGcdJbk/x5
1mf20Kr9WMSTQQn35cA7c3CvfbT0gARuOEGlFRB4PN9DW83fLgdzsfEpKYxAuWrREi1bvYbvtl+u
m1ojdji5BIQbH5IP/UbnjDpDLkO/Liy3VreLHxsYRKBKd8Yw2ey1Cwy8jLH3iitykOoxykRS/G76
F2uekCTi5XgtVUVirvSO/w7XKO/CzLzsd1FzMTxESzW7Q/4N+pmrq38sRwg/SFOxtS5ArtThjmcN
O6mOPFMYkgpgVfZC+Anb/zgXiJuawYuI4xxuizMosR6BX4kdIqJBvcRgITHoZxZvEbmmbB+X15ul
dnyzP7hezq7+/dSS9VGt/6BwlZLoIcohTWIOeyPBg3JLuT+AfUX8UXO/GBh/VJdE5O0aLm/4yU5f
f2gikbdibgF2h5M1WJMa1Jbw/8r9QOmpfVXW7zYihjnvD0+YPP/1tYvr2acIZYSqUwuVadaiOKJb
Z8jsTscnN9L8UM1oUsvsQpAoRON6z7SusBwGamjAc+GV8UQUt2FUsMzErji1TqJvu58qozRkwORP
m+CF/ykT7wfet4jCVEUKxeiOUQzCZ4CZIPRNEuvLvG3dlX8zQNdzGSOkak8quzGMh8bxQkuy61/p
M1Rk/tBaBRrXB31h6cFCRQebVgmRj3+eBWSPEMO17L4MNOBYoY13Z8T2HJkxlMva5jmijnVg8d7b
cMEE331g4qXbsVqITmYcmDmCDgRLwZ7pmMFq8bKIQnmUCayuCj+svRRx66JOp0kV4mBbZOjv+7AE
kYzt8H0e7P8blEQinD9yg9wax14NHfiZvAMjD3LLqCY8F6fjnmMGd3NZ8sr4PiLdl/MNIVnIcEss
UBG3mdEFU5BcDKlNWmBpnoCgy9AmJSkeMtiDL9xkqtWyloYOKviX+wI/5rkunW55LYAc2QaNdvhf
aUXIbiKBKJM96DgGEMaO9v/Z44kGYCgIi3ePAubIPq+PtKJ0Y13nz8gSDni8E93wISrqw6buD05s
6UT8iD6nurum6KOb6rclMQ31GMjBCd8KZ2c+NN7ojWUfiIqTYVR1LGtwNKGfdxe2JKydclk7g53H
IKpABkZLBJuDQz+QRfxlSwt8yGflGhWDz4uZRdM+9LtlvAxWpo5Hf87gMHOjyLO9T2EiZqVAVSh7
dlSjqmQx8whk+10jT7WvuVCJr8V8qcfJel5867JKccapddxkFsK0IJ+IMQkEPxilLBAG4RD+QGoy
Qv+ieulXgcwMn///XfUd8KyDoqwm6spL87SPKSd9cs1iqvtxNS7d1r8pywuylXbObxXZbfs4zX73
wf3ELSQ0sVkbaR8983sz/udu0ArPWj3CpAADKZtvE8wrIhh9/djycmTuDT9w6vNihG4GFYj5/Aj3
FRTxSCKaBtciwpgfwhPcNtSIoT+kp2lPgW8QFex4pfqSbqAtc/tpk2pG5JLDEzWLLspsCcEPMIVB
GsCpvnSEwSc56gc81qcL76MoQtfWg1vGMIi+xR4RgIImPieGAosVKESsPC00N30utGrzKNbGvd0O
hDEZ0xMUT2pLadY1xBUBeKtawLXIwcvMattR0agirYjNJqB0YjIbCwSNN03RNLeOeomoV2x2AWTO
UNdnZuOiSsGGLJ6at/DbFn86ZJwW1l8JHP1PVqHKUxBYCl3RDSdH0kmAmYrPok6hbynFKlccnQng
qfwOee2/ezAr6RMKyH2ZXwrV0a5pIycx7O2/OzPmuiCceyJfLMjxeOkS/Mj6SRpmyLIvYu3xxGNG
PHXHnFr7hQ30nVoSl1ZkokJTLCTIfJxa28QCYKRcd4FuxEkCVgVI/anbPT1aBZ2vpMLWDY0+vooL
PjdCKqGm10Xp6ZQqSObWeq00OfSIcGg0Z8u5gkHK+T+mzg9rvheCFFIaG+o69pPL98Xifc03WRZ4
EcBHZBlsOaoEe1sHT4O4GVQAF856cu7LAHmNI0sayBPHo2fLiO2QxOmDPuv4/nS2bHv4mVc0g2HG
bBUjWAjmjjXJs0sePIMMsJE71z2SGIaTY0G7Y7OCELZ/Wgig3QAQClQsDLFXjq2XPfHuzcgLdYTO
82lzoeC6Y42nCFLoJXCeZUgqKsPsAHoM6G0FYf8iKxhpZCkhQncq7Ff5Cx5kf2ZX0i5bwbdxt65C
aC6JqxkdHAHHKv3M5FVJ1/r0H78UN38VyBoqllN6Wn21B6iUnmFpTW4HGpSWrKCYfIy+uCE8G16u
Sn2S/xSt1jEjYDmhcqPy+m15X+Fac065GZ8hTQhfqvkgEXBgxV/H/r3pLOIUV4aL+y0orufryhAe
XgZBlSCgMRqSf4jiXmA7hCeD+HgRA2l3AAKx6d7yGfhjxpDl2aw8MxOrJRORRjM1jqyImNWM2XKL
6yLxmcX+tNR1nlnxllsHidsor/LXimsQqZzXYUvel9sjTT+gBrb0Q8vD7sLiUHJce6sFrT6GP4Li
D8U02qtyOTOK6XD+qk3Tx6K1Dq5AwrjLa0u+I1lxUljvpGAKJwrKnx+8FtNDgZjDYDus+wlLYA4G
kwdwZnjKFFoGtlL2iupKJ/BeFlLTsxc2LTTYEtSMmgeculc/BsEuKY41nku+LtaXt73xh3tEN1zg
YslnR7Ng8j5rpZNHSiXBcOU5FwsJduibhLVJeS/pCcOobg24KHnw0OPnaNgDjkna5Zd26+z8ZCpf
C+rQIjUx+YuB5b+iWT9zDXtf695YhdJQuHk6RzToiqGyAP5NPu1+XTjCnkhxkoj1hts04U8N5huv
kdO2uIvdd/jTl5lvJSuuzO3Y2WiTOE3F85HLI7lMonOEhpqhAD+yAePtPXkiU5u9QWC1onxLdV+l
qMh+8J2w9I8AO1IfICWynOKcXEDlzVhaBtsPrfdVt7BnQ/uxsz1mHviss7205/azW+dJx6D5sM62
lAl4W64cZ7yOm+L6BJ3CEgz7LEKPLnq3/qKgE2LIo68A1InMG4+J2xpkfZeSxLPmy5wvzEXRLq9v
zU+uZNKwu5A1QC9BqKL5+8X8pmvsMVrlwZ6KY5UtyRPbrg7FposYco8QGxYL0IBv4ZfnIIVNoI5N
X5Ac56t1MccBrV5iu3IOJvkejvFhEKpxwUGK+LfCEqI7W9l9z8/6NRNcdm2lcf/dmsRbj5hKRq++
Of3e1mYyAr2vk+Q9RKLTwV27Is3y63x3E1qEzJV+n9n44FFtQTXC9iM5VXl3/+yh0v3VpGTTd8nE
l11TLX8EL3Ih0XfRLnQj52AhrSRTizQX+CtXOyWqsFMJXHfuiW6+RqSnTKfoVtJcig56SFt6dXYi
GV429uauQDSIIz8JYxBSLnzI/Z7RX1WHwGh5MrkJzpfZYbrt1iETpSXnSBfiw5AYUo6AnO1yDEnX
vUKSTzPhQh5/e93bzcYcArDcMJVHRgfjKNOYTqt8ZW5KMiNrjLQW0ekW0qUokxHMv3+xWRmU4lOi
IV/j2ITolD+6WnF4MxxU0NvVSTE6pV/8GBuvyvrWz+oEzxC3OO5D2M93Af/NQcrb4wvxrVVXX/on
ZB882Cb7xfe3VMFIE8VeWVPUECgZy2JVk7GGUUqf8D6Hc/+0gEeHc/AGIL0X43Q3lat6semgJAZ1
xAUjdM7LetYyXzCBzMmQmTBiPXOLHhb+AElB3LCC0N7fL8LGXiRepAfvB0qOy/J8fBr6oP+Y7Lq1
XfT9zy3yQ1IqhOUJyaTFP4zvx4yksPytSCwtd/NAkKvOzzvKD6ZbH6BGtSKF+tUu9pT2f6IdCrRl
2ZSt0VYtKbaHzFksrOn1vrQANTjhMZGxRrpzAlv/YlnfFQGSL6ibt1SNCD9SSyVUEqJ7shFIEbES
OnFeR42TutzFgQdcYXoEJuCQRlWzr2pjg13Ep5kmL6Ivtr2WLcHlMrgX/idqTXOWjAJr2ECfVN9T
D6LwcrEYZtDPhLAe0aoQEs/uzlGrAzz2kIXZ9zTkEMh1/GnjObZprj/s7G4N64SwUpb74RJ/cD3b
ZL2m2qBUyeavK+VylCKD/2E//dgPSfYtkurPR4S4ag/0axyX+aajPKuCYAEGshJ4b2J1htbrR3Sp
5XRjPWoDsRWFz4sXiMSMeL7TuapUpNVBq7SqPUFH85OhlFgdauGQtyjrc7dK0l+swMEOQIOZdmY2
9lGwyZWxBpVAxeWcJY+SeqR2pmucxo7vL8fuSNi6Ux6X0iY8hpa3GpNknQ6rHJICIY5wLTaqrg9J
vwDZJGowKQ2DG8obMHv6ox9ufslGyPnDWfGxs2GS8hG5VKhfnE9ecw4U/w80AFIIgqIWWPggi8wP
PnYi8syCmSCo1g+UrlXBk7U9XrG0CdjTAoYvTHZs3KqHEF1+JrZWvzE42tJ6ZDWVOJJv6p9je6LT
uWaqZqsuA2vUbyt2IoibvIOrdjYh0uyGX5tp+7ZQTV0IjCezUHgpPENGcHsAwNEkvHfa2KLHub48
K8rTpHM1Lm7pKTg5LTt6ovsyWj1wNExZkWbIoiwolpndE0RMXwGLz6wBI0EXlZeH3fGsQ0eeKBQR
LCYUbm02amhIOCJpjpAmefbyMTB0NN0T665/Tv1kUVr/xLhEfQ26SqcTHLwlKQIEejV9XWbYSyfM
zpOYpxnLVLTXROSLIdyQGO3hVcDjEQoDA9H5HkVJfwBbMjYwtE6al4PMvOhB1PUh6RVCxmUWN0af
v39JL2CHorgUU0CFOhywNe7wrk7FFe8jK6qnIGt1hpyULqkOlc4oIM6kTi1+BoGorJEODPSkVqNC
JnNtNbUOq+y00G6vVgLEg4XqqGjOgEoMNG+OeMV8ntS3f2oHq5EIpiPVSnX4K8x0IsCcXo8ixGTQ
Ixt0qtv4eF+55+kuVihAO4OXdPyM3/MKJT1s/xf+j00xe9E+1C1LWKF38pJnW8eJ1btxC/1IEMu1
LM7+oNvp1M7+GS0WEyFwOetwI991kHN80+DnGH5ZoR2h5ivNnSFpgMinfKqCL/0ex1lgtM2rIplw
DS/pBZHCoHne8Ky34GWgTGIQ01drWbr6opyjchxBt6vTnL5Ue4WTQHzeUeLN4ZzTKGDnGNNpiBUj
y61WojJQ8XSWkpEROZXo1YfydogpqKScoawCltRiTH/VeN0ycmhV1wiuRQqYtoJfK2p8xdY0Z/5K
WnZnO2HRoG+R2jHAiOkuDXV79fq5nBqLSzLWowYXZXCcwtgPRvQlpLNH30ccy1ChlZbFeQjJVuAd
GXfTD3M/ItLdAPdlVwaZmQe3dlmmkX0vnMet/1bSWomiaE0COgPfGs/ee8NnPro3JBIhgEwMUTzv
OyU3fi/v+twE/mEJE++pTGmIWkiBp4v5S74APUb9l2gOV4NCDhIR0IyMocyp41O6mZqpYamh7U2y
0K/gxeZaCo64buwvH0s+s0XBWhRyCcMRZcidcY+RmOIx3PPSzmlf7bw4CY1522Mm1s4uzgHIABaR
YuYi1hnzugQt1hvNYmMS/Wsp4MzS8/bV1AAiPTbyJ31IM1jwnLfNr+fC7LGERA4XxeFv3AXBFyH/
nnogyvx+zOAp8Ip+F7yNOfHTiuSYFqLrwDESXNlTA/d6ibCkZ6WnQh4SnUoosU92vy4dEy/Pdifx
nm0FXAQfxEg1/SQDRpOVd28XbpbMcVIX2Zh5qYE/lKVdntxKlgUgTs3efy/p5cvVJVSdlkIjardU
DRRSqtqgoeWMWfVyp75bwPZo7YJ+7nMI4gWY+dpYSQ3K23+9a+6FK7ZC/7G73sDz84PisWKV9c8X
+gXfWJKrZGLJ0Z2Md5wPqB0KhvkTApUV3FIivosB+IGtnNqtDUMpaU2EwgHCxuvQwE7xx9nO+k6E
1rj6oqyBYPmcBG6Wd4Q+CTSh8juZCi2LVF+n2BVS2j+f07i5GP7Z2gObv+sd0ZDpPr9oFyUe9j/G
BpVFIbaX6jmrGlMqeRvBlJF2TRO1MVdMvrKngvoLrVNltkxYC2f9PLQFnVsHPIgTyRuRMPbOfolh
Gf6PxbNrb2kxZuD4vWiM+qrpbLh0kGUAy2zvErCYzpzEl3maV9dZNRNeYeZeuDmkwPZuzT10TE8M
aaVu9waUkJQhNDuapj7pU+ao563EW4s2DqE837YlDc5a0kHEixtTk/3WACxaEESfhkggvWZS3+qD
9ILNMQjf8tW+3PBPXN8tRmr++cly9n6frfA1TQdcSCV1dyTz6fJkdDke9wpZFhC8y+9FvBVi2d6V
1ZE4jmDgu3HGSkuqAchXdhob6fEjrTELNBh8QHw9qENV1guMA4cRNK3uL/sig3Iksvr8z4/vBhYd
OZ/QIH4fz6IejFNKtTVa1gZ7zb/NpwbL698qOpb2+tCRvotxVTLGHI3xy9TcDrVcM/aH7F510vpf
kbpkQsm+QqbfMznvwGtLbCbyST37tkERv6frGZqpTRzDBqQ3RmH/+sTOl2fQFXrz7lm8e6RygOsF
J3ZOoBEsEMtDfbypyXQVb3UJ93Fn90Yp1G8k+hmNG9Sp3IbsOL9Y26uWrYcRwkjs5j5SPPIc6vCA
8nXIm+Nu4CNMpGs+yOVtOYWCpwYWIy4nP7F5dEPNQ/MJbDvCWbKeJWvOoBc31ddQqcbLo/fo7Cn1
NlX7rZ/fCSdZsvsO7rdlcwsPF7T+HT+UcecIWeEwnEKcVT7elpMCRXn1eb8bm6QNZ8P1LWyZyk6T
LDtNxCFfYvek37ChvUpiTRWYUoMyLlll1mtxaBQch1BtStB/WgNuTlvVtt0sFRR2ILjH9PtHCtCm
xMZR7mpoHJXRqfAR4/2KwMl63/WSP4JUi4MFudr0ipNIANm9gfFQ0HBDu2byT4s8tShTjVQO/103
EbtI6btoo5UQ/QDBfdr3rQjvco5X+t3b7+NRdvhdWMuVPJlMGCVI5BKLG3ClY6umW5Q2jKded8SD
q26xj6t4kMj7cJWQCBd3rEJ1y2WYDg8hLn2zoM/Q6DRMaiiix0748+/Rf5hfNxs5+td9k66whvUc
e8cgwJdDNoXYRVn8qQpCnmtEyzvWLqK/7orcdBdPY+t4qzE4zg6wSaVWplI5Vqf2PqL1axiZONnc
JlMUCEdXp8lIpKAPUOZ4Lz9PIGLK7WahH/0ROHOFqS4emYu+ByDNznpBYLioOhkTaCmC3nHeANSt
MPvh8977c8bZMuXxpKOLAe5tzpVo/jXNM1Ak6uHhVMXLUJpOCHoAnyWpEOE9+psGhWIik7nWGeYn
+DtoZVAmlB2uPbrFtu+xlYpQ+ni3lWRquFMkIVc7r6GEakJ0Q65fDw9TxgK4oynr1J/Ftzco4cP/
aibBXUFMVsbekHaEz8Pthm59u8ajC2LwJEH0sBsvyeRkn0LWF/P5D5Bou0fxy16K6J2AaHVgaNXr
j0wzrVmJJpAyvPsxv+YYb8qk2DSQyyt8LYP3WzvTKyb5J1D++l9WKDnI6DG5HdCbyVdNp158KMVH
BaHT9MhzrBsAfuzYobNFVApnzxD1/8uuem7Y3gQ75GfKpDZ5l/s/Xtbj/5A47QxYuJq21R/z0HK5
oEdUYQuhcZvQI5GtU3sBq3Gn7e5MgUfgxeenXjyK87AOw5FTQuHfYE++MrhYXXWUw6T73/6teR+Q
UGKZ4lrpZojMsyA4KaPwqCMPvIJW+NLVdN/ZRoeX31/HU33XqTNsluLg1f9Fmdqzfkqol9fuFqKW
bo99t5EFNjVUkLcM+H7MHSh7LtTnyWB83SkkEWdVCCH72EfZlDolmAKJF29hCnudre04UnSWXO2G
XvDnstithXK+WJinr43PGBf6hyaWCMdF+uH+ZPo6VFgsjKBJyN1/kuaKbjWrFz6iK0YOzofzh5Wv
3Ibo6/ve7mytQqmNgqjBbAg8YjdEXde3XQJzDekU1TG1HqCjPBbRSs+WDOouQ//83D6xedkYiQDa
UCH4qiOTw4TZ1DaCEBKvh3QoANe18cquWHb9BMXnR+tds2t7Wb5ilpOBFThfFh7fJit0NcAFyG/k
BiQ3phLbhKWNcst3CI4Te8sTAGxXfdu6MaHWhm/nc0r+JFiMfi06fF7NGBM5VvFHnLF0BQRv/4wo
zmQaUgEaIzQ51OkJhj4u9rz5FxsDJEaSAXgOFHcYWpcjlK2FO7zWHulsnnghkeQmt0jLuUWilAp+
OSj4XSJJV9PyjiQI2PEgeDa2Rr9h/a6B626c50GNDTBsvH7pON3e6V2ViUBN3lOqikZCw9XUb8eb
nzo6R2sr411BAP3kkusUxcrWtRF7aqxmNis8+J5eOoLK7+4zGPbdRXn7b8g5sr0ryX/dbt+PKPGR
tO+LtJZmwdES/pTQrqn/YeeH0QR55yXLq2NecrjT12yWB1gqPXWuwKrG2LI67U9Lv8zQmOdRUxpS
HN7lI61s29bjGQ33l4b7LDyVaPb0FbRc54k+kU1aOBnlAc7CYSY6MclCZrAgrA9LYUAMQ17JYT+o
hxTYKPVhqAgZ3K1f0Gjty61gybS83+Tt1PxNMjcNezPHeOGiwJRuynAzBIpznKWyeZUAwhXgzhCc
d+ekYpjGR8gk9K3qmjCm8wP/U8fxqHzgYEZRqTAbtYKKU3ce151Fqo+H8Lcy9/3xL5U1lAReQUAf
lzSJso0VDg6b8EA7r5hpDcOhuCGWlPvd5baGyUBmM3WHaiBRMS9Js0ylyBJKesP4JcIGGselt6Vn
9C6QLyh938qhKad9jELjk44B1I5ha7mhkTL00mFsEH69ogD1ROaCzUw5jlZ1ybxLdCp/c70VYvTs
nxfv3+ftLRbzsjVkywdM7W9jhE0GfoJ6RnQQDfr7GzI9VsYOUtVvLGF88Ob4WdHiGP7hIh77KEbE
JA29dL5Rxxitjisnf3utXqRgImuEq5QQ855W76tbqsQ8TBki2FHmPCoTkDYRuubOKrw83q1KT7Ej
1mvkCuYSPok5M3m9uoRwAQvR4z+8FV6smSqSc5+g3htNvPkamy1uPFeqSV7RbDIAvZ3MnmRDDx5T
Pl4yRTGGFAroWxj9hzXvpY+dZbyRUsz1enopG8UKBuGfsxh1s98XN8YsiqGAeuZZpTHVijs2YnQI
IF04qIwoQCgJi+xsgAmSX0v8PAOraYqgRLbfwTKQ/hjXnwnf9paT2VgD8VA5Ab5tbW8h2AHcZUCL
DxcTyi2ptEY2ll4H/nIJBBR+rdnLfCS97lkkVt9W41mW8ijQXs85KqhCRXLLJ4pGor8l4b577vj0
GKGuzAbA9Mx+F1j7TR9GEm7h1vsF8bteed+G9QGdOtEoelBvmB/KAsZeg4zzk3yE0xdDavYJdr+I
1t+mXBS9cb8r33P50+ADhH6uCsb5NjVNaF5VSIlB30k7pCKALZPANtSJSUZAslEm2KOl3aekxWLw
VVGJt9Fo7a//nT7lLYrapiBqGJ36KoG+veJE56ezO3JyRdl7W5eBubbiBayBEU2OyRRWI+Nl12lv
L+JwXz/vnb95N683UDXcpYpzV8xu5cZWUatYZ+U20BHGvbvvZ6sf6XcZIhwl7CSpUepPGsfKjqdn
QGUQMkDP+EHT0jcOWows+/dPuw8t5Vy5ShGpbnTTZBixp4Z1WZpcPG/AHneFMIcmoAtSlEiF8U6V
h0vk+YkdVxokxqFMX/FB1XIY0/aAjvIOWY2qYH0yh37ez2WYfUrIxobmhmwci1k+Nmb0pZC2wQgY
VOMnO1j3TPOv34I6uSw6Zb7s8s1zrgYTHUl7SEwmQXhAr3fdygXQQIWXonB0YfeB7bRcByaj/eBE
KJVVMG+SCKp2qfkeWabBWcFyxApDrcDe70rhH/wmmHeNY1ihRmMlrYiPv3XdOMbvSqF8NYVDouIV
Z6kSQ2AKn1CZQWA1JcdHIHKYg1vd6F8QEKTSopmxRT8gC0Ou8mKWWKHRDkXygxTIc81xbh0SL6g2
TpmzNYqKvV52we82J5wZc1tro6xNwbqa6+J9anWrgeFsRrQfWuvOXoxwsqaDxWStKUvfhiOQakEn
7WIxjr18Sjmme2sql3NskB2PpSTmoXg0Wy3Ez9Y/+116G7LgTcUURxUOxaDtX74i0YybIYichArG
AP6ukD7GOvKVUkbIyngQeU+W91UM00Rtmi5wsNSq5egi4U0FbJ9g74Rj2QSBAJR8m0MMS+OFT9cT
YmbrGi46o9nDwwQjeCKJsOO86ywFpNhjxVp4UwMXuHEhQr3RsBtp1UbLJVLXOmF8tXCAIjNQg0z+
7O4wMgBLPA5NZ4Ux4tBuHcOBVjpN+ud+ZJpn92+Ah12Rdo0TtNHsSkGw3XgprIZrbljFcA6JT8MS
32JYMdgraIPXFGLJRp1AWT+fqWjlf2rp+8acXVajMAUHIGFvXjoN/Lt1YSJHp6OX4jAqroxRd2g4
MV5ladPQdDFa6V83cfsR0t2qy+CviHAB0aB3e6Ncjj8AW7h8Cmhu5jydyv7sJdXKEmkP1pdMSNdA
XNQzPcu13SveQ9QnuEbKQieELAAlmckky4ypnioVC4c2z/xdeGMSXpFjDX6FupHPBuifQBv6KoUt
MTdjOKf69zB2bhEj7ZyOzZH/2tC/0n7toitI61A4k2CpjQtnBUrOoIZrRx4lDh++rXRqd+mFS6QW
g94dtayCEzIix8Lc/nDk+qZF7sQNjv9e8XExv7v6ZLpJSK57SencUHk/IGkVS91mGZv4Y9QKcR2V
YKISQuVDhSKHMIgz/FQ158KQeLI4vckGI9sfSII0XM3tD3eCL39+o5IDcy+ZkoaKKhlkdcD6T+l1
rj2s3KA53vCQ/BPaSC4Q/G12DASIY0kUW+lwM9s9U8dEdWQFpOY+Cu35494KLx57nuSMYNSUHwk8
qsU549tmsMaIkisVsu7786lHJ3bY32pHYGrZCGG+XrnCfcvPP1vb8drRxQQfeBexoOoav4dZH+zI
lVOoyIASOCNtwRtv9gDVQcrggjwMDUn5/jHc4Z+0Z6qg6pRY2IoLxeSJncDmtVrKkA2R0TNcZT7m
5qfm8KCR9rI5EjqUdnXULuVrmdtIVfvGN4ZlY3FrRUtYSlGwg0JQxwFvrsOkQ6PWmgAkxNU9wPb7
JYBMyxcBgr08YTPeYxnsG3qR8wcZSAB5fH7UteCz5uA/dvvTggtBc+C7uQuhxR0LKfWXQ9h57pGh
yIp/+ZU5DyAHzyu69cBOrcsXxLYeJcQShz4RMyYVp3AoKNvtvX+UTmCqWKjJoNz9Z1dS3Fml42VY
DmnpPyRn4kD+ATVwu9GlbveGDspcOq0JbD7ERL21HBNwDgOw5FGl1OBqUCPeFYuEMcLBFPxreQ4K
i18Df1YulnZHNBm68PjZVtAQKcStl7GFXC5Jk5M0HB2hqjjahAD1kvJVzrErSxTwP/yUtA21iEpY
iaoGKf84kSzVzM6CIHUzuJSrL7pO1nek+vy9Hek8+3j7eLR625hVTyt9TxEcSI/aCgKroDw7gXnS
WUJUzQChKUnumV+KUUBVgtS5zAXCpUORdvPKdnJDbuqEIwvJVs5KdFaZ5OLcEQbgW4KcwLmfOhJe
/aakGHgdbfSFRY+WaOjx4hkCePGWQPzIkfWtHrGx5kIU3yTwNEcuIJN6PgMqXFQs9CfWU2ER407a
bwsmpxm3LFPHuPIRMmzZ9hO9VJ73KMlgHI3w6DT807msy0rkGssrdkW3f5gY48zpszqIcOI9OwhZ
Bf2GEyo1io8NZPkyYOq484shLj5aH5oQcL5IQDHTjLTPksWOUgAEC2eLGmYEWPH01r0ye+JfX7Tn
IkBXBCa1CtHPnLGcZF5UBgTBnMwJL77vdVurD5TTtINS8TaDGmL2+SnYjDxzGG5p7UIZWPXOPs/P
XN9T73/jwgAhXvCzC7BCamzIE/z7FwAAK6erjQxrA22JoloxgpO3z8PDJ0Gg3fzCFk2H9Y5PfG16
/8ix+ZTQwNdHiR7uaB4PcvW02PDZQwDD69t2zlQp7GT/bPhSrdkA30xVDVgepT/peNROgrSNfF0+
8MQ4EMN1VfZrcwZXnzHNyMDwcR8ZPTHkVPTHUHrj40MWDJrTMU5GAH5VWgR0rzaPYZA6NmBcebrv
cLEethUVVvR+MnrohExWL2LLNdRQZ4VSufGxxTrrlHOEW2O+hn7ajXDaEqpquM7Pzkxe3r9EpXbB
pVZvpe7xVahuSMzr51B2K+7YqxrG+riUvMqpcQHXd/C6vRLkiXRzZNGWHCF0sYfO0HREjKT+PhoQ
R46ar4nINej3cG2ymIKukJSubKcJvtdTP1T55HFRte3NTd5mP+ftVcSz9yazvo9GrhC8/xWrHyO6
92WB0ZCSs3Z0Sj/dzI18hcykQQj4UrbtCLivmchMcvMU2sJZ7heHaAa3NzdoQoVV7bRSpbSfW+pn
B5uvxZpyAlUSL4B1NqNuJVQNB3AuIRfNtJc7DvTFcSBQJy60cck0XWfFSnw3WZhHTMpm02rFZEZH
pHgwUeCriF5Smui83XHu+upwM2oKxHLAa2ESMzJ5+F+ooJDtinQkqCmPIZwWI9CR/hBXmsNKRcVC
hos/wTkgL7hESMC3ymJNMCWJcyUc10XmhyZYxjWy2byqwtz/6noVASfpmQeAhlW4BJtG1Vn93NxG
KOhEch8shtlgg5d2vO+ih/e6JIkIouX3p0crMNC4rRHdJqgO01jpbfN9TjJvFWGyaP/Kzb5yBaaJ
0ijA+7DZTTXvwaO0pX6i30Ok5o85zUOOjC2/f2PBN3RWOjXGq42883GOpS9wvfI5QmFDfrchBxyV
rb5KsaBKTCqVaoLYsPnS20kUP54pET7571tw8MTWPVA0UrwOfY2Np085QFRLBDNbt2C77DO4IwFC
gE0+I6MdYCQB7pAKgRqn9NK3wpHFr+vZsCK9icTd23ExVyDuBeEOa1ut2tehD+dkuCg6kkIkvicl
e7Apxz413QF6Xg1fCgxYuTxC5+kzaUyqp1xEx26lPQHfF7dZgpnvdmOyBbxHnqmDTTu7gsaDU+bc
orBHTZgAl79M4HXr54mQlQoUgxOR25ArpKelezAUYglyShYzorO3O3+xr2UV2v8zEOdt3CewG2Sz
YcHvB6qOqBhSYatBedaXEzXStg/rfI9cjTHVvQ/xzmTYRpmAbYII7ZK1gMdT9hTo7USiJf0rbbA6
U6Z3G14vVXIEW1jiV/BkdXhtRc+3Rc006fCdx4D7SjMqVqPT3mH2sH7d2yPWVMm7uytoIbuNTf48
13PnEFJwo8zMhfz5llgqvw9WpEODXmD//ywvZYq0LV/LlkF2RITbYd32CTLFia/HMg/uLfemBqRp
5ohYt05RLN+9f72KdpY7MwjYvrmjgZJzgjCTvXazbqb49Q15CdQh/I/IpWpIqeGDEuVS5A6R+6U7
gi2qVQay81apnSvaygnWS6yiCk21B7Ltp0EOE1cPg4tGSKLqqjYNfPsO3b8ZvFitHltqI/XJXyLH
NzSOtiqFKXnXrkCh+JjKf9zPJWD/Btr0srkyA5fu2IgW2o9o+QsGrgqjxVWQvt+Kw5PYyyZY0A6K
T1SKbVVJVZ8fSczAaRw2I6DkIpig4Ymb27a+dSwwB5dwFlCQSLFhzx87vaJM+fJsdMXP3JmLmRvw
uWfpPxIi5CViDuHJsuRLFrvEG0v5wWh3z62BRBcQX+nitFvo94tny4nQuZUm2yep8tXI78pQSUDt
F2Pkf538MtZWWcW/cEa9vlyas0F31xhRa3y1J7lzcP9pgtwJchxgpoK7Mz4zZMFhb3+DpZdtR9J7
gtpOP/ymdEA4zxyqMkoQRgBnioMu/v3VVu8WZa16FxrVYyMvWJydxr69zFoB2dTsmBf7FcV3c5iT
HsNmAw274b0gCRxlg1FtFnwkuhEYJc1DWZYgMp30X/DtXLqqvgz81648iiDh0aBf5QUcTRJtsRiw
W6krp2WGsexjZRdkla13HYtBFzpCmuD+3hnaKCtlLyC0roxghHpN1MlrBE3hCW/nMfzCQUGMxW76
DZxAetKh7JBsCt6dtev+3F+TXuYXQXdeDzPVL+SgEELuTR8PwRqTAWuZNCdqJ2gB+1gCehff3vvC
sWsVqBK5XV6a8L7KF1eDq7F114zKCUOP0YT60rt4qjfocpRLmVuTfCUrX1W4VUQszsQkMJTC5TEQ
xrfQx654susRQfErBwQeegftx80NbRr43ayDtj4VTqSkTz4JH25epVeGAlZzM1q/8sMEa/jQ13t6
wzxgQUQ4zI6aYfLt+VM9z9/djkEqqwtcd+JMPsZmBVHh4BfEx9/F5aBBD5dXhf2bRb1G+n4a+kn6
+sUdgdTiRQXTYf/2XhUkIS/IP40OKDQLMjmZeV08Tb91AdF5zAnPn0Cn5zHapFtUjL+NtVYxLhmY
rIBuG+vYnOwna3CkD4H7ay7N/njCbnBWZMAA42dnk9Yg2i5HYYajtND57HzgSRYDuAP9K4lLGyEd
jWe9N1VOpQW2TFjJKbNXA1+VnoHnQ9PC64rLFkpO5WA8v3AuFnonOQJASpXSmd9lWBmJN8RIbDQO
TMcWvZtvMAD9pu8tliM14JGVxH7i6MLhf3tgLvgTjBAulcITmDUYndxZCnULharn4AVyYLFUmUWo
gDLcU0lHYX9Geiv85YALu4xnGWMck1HzsgY4pOhk4VhpAuG9BhttfRkSNYGWsWaV8E6k6dmT/bAy
RrZh6ADoYngWDf8tGfSIvop6mlUO94k7Fl61Y4XKpYmWh8YoltHs8pb8MKGilBj5+yxa90JKhJvS
MuQmHyfoAF4a3ioG6XjjeSyC17N8kBFeXnQKAux5K+uU6K4gqe/UqGlEj2LANAZ0tGpR5hDrmepa
Q9Q1Td3ylEKzuuI2hEylVD3oKrZXlw6QUkXjoZuKuoLdC0tcqZ1MwmW00FHMzloqUDzLZvNNJ0im
wWB0BQCNlhEX2Z7ot7W4BXkUbXhm+jpfZaPWAUx/AfaQoIhZ2Q6h3SKLkUovtjsUtXTD76ctTdbL
RSoqTtrExLMzaEg4YUffg91NQjtGwSRmZmgbI8L9533ifOkDe8EhbeK9qo3y/xFfdiL56Qg1Zg57
SxpqRSXstYpXz9gHswR+hEv4LMAC1Ji6x0Lh5lZRpotngzZ3DjwcmSVB6qgSGA7JVtTvgRowJg+v
l77tFWbx5mvREDVxAkjNEtMSqU+bHaedSA3jl8EvnrzsKUVd/Sim4j3AjP5yF64YFB2Kti2jGZqQ
F8iKqMw+2ReaAxJzczsLVcytcaviMAe7M+53Sre3y39Kr4vKDZhH9CBINHdTrJV2GtdwPj9emmEe
sywqdRQ95sPCOkR7A+dovL9F4OJ4/NVN+YeAMwudAaxQgp+7e/zRd8GHYDLOvAj2WS9KoNj+HSd6
3ISj6eFZHefqweIQPPTlfhdsNXSeNwHrvpwrQpGepAyFrGtBhN5bAhe0/jSr2rBGBeNvxc0p4jFp
oCN/TZ0IGu2ZXp9N0vnmDsdsE5b3Oj7680aQHK033Y0GyOdODWD4Sdy4x8GEMLuJtX6vN4Vj66qQ
Hh/BNkpeCimj8xVFQT445sIBiUTDjlcWnrqwXQy3aPGjEYtV0qLg9RzXR3h6386VetV1aVL9wUOK
DedGxlClfgJDFOFqInTmlIjiAm3dGgmFtEUG28SwxGOvAjiJqGVdUl4dK04sLeaIeakEKU2w1BK2
nYvkNWiD/q8MDp0DHHD1T9sdfOOxSW62ZnyPwVdSEFiq7HAehQrG55k9/CFysS2FWOY4+ya60uoo
iIHa2NeDZCwh4cQBwNzcBS9Eb7hLYbzavqkhP0IcGUp1JM+PwJQ+Cqbekpwlf1jA3rdR+fCkrO10
IrhjpbrOVkLXkC2Z6awGoG2jzx+GtxAD2Ce6F5D9paWQ44/ehrYp0TZ1HILSD0bGAeoHv37ss5IM
vK8yEc2jl4Bn4JYAQmA2Se/hokYwQdjzy5Gf0zRXl9kov2yHfyPJPU0GHTNDphRKgSqZHaL/dXau
ig2VWYb9UI3M8xbrJLvPRJ2IIDFy3UYkJppLkUs3V9f5PA94L0C2Y9y7DDDGXmmW7HjgSY6O8wyn
te9ywX4d3ssBp3RRe+KYLGd1CBRl4tya54BNK/KyUgetl+kxC1XGfIpK1auIdxZxM+MEMmHUyOoU
10PYLXdhalfh7A/FMRN3nVsnyL5BW7NkfmEF6Ud0+VjZcg22BkysyeXPq6XjD1wGOUQIIIBZJGoA
LH5NvT0lw39FKWdxLF0QIT6m+XxPrpPo5cq8U5jNuVpue4t87RIRxaOvmTRaESwdMqxSSpLddib4
EmfSd4aMTdigboLiDSJKxTwsjBZhuYOfmrxF4xv3vPo6SK5eFSequvYEGxCMKZTNxeQau7LxQj+R
aACkkrgmjdZ1qfvF4NBhF+uMfZOX1f49+AOLAVCsz7V8IDDR70oj1Iba6KOxKz0vjYI6+4L/Wnqa
3F3PYXwh3g3kWzZnPK6M3Qequi5wd2DCMAx9YyXKxFk/6lRlSg6c4uzwSGnkPt4ihTh5wk395Q4p
t0ODjIOQA7uOrJq7W3EEJ/2QEQUORQH3V4njy02vzcH+kA0+hOCLyf7oil+LOlTQUDsomHMUMOaK
wkyHIjDmKQ9rTpfdk+rn0aO5mfiHWLo+ast5B62vFn7K23+h7/bA9y1faM/jMbpp1k9X2opAPDjm
7HYmWVx0NPrvUv6RWEb7Ab3zYId1knuQ2RAPUsgIbyGJvfpSqKY6pRaZ2zHJapt7kEc5YVqPSULt
tZ0lhDNJyB9eVla/Y/eN2zMpIxTu4gHlX9VNNmnebQ/I6SNfDs/iMo6KV1E4pFRR2kQ3XdB9u+5N
8EXdPFKv4uNEbpaweRv2xmA3dUOOwFx3ad+wN7bzw4Jv/YREJpBPOU+VNl9CmKIVEiIl2fc+8hKi
Yw+H7tl2gyjihFlpI3f3XcpwCKTrhqo321k82ZqOJy9xSyw1VtSa5Y7HAk+NNMeZhZy4E1B3WqlS
RohyvFNAG+zBpYFKKSwx5hSM4Fa1cq6RAaD5GXnweC6iFK218Buuz9xRtxive/Z7OvKDpDiBE8VL
/2lJ2+vGwu7YlFxCk/pDK8aHmcnNCLb/Lf85K09aaOKIe1o+/lbJz/V9YbLY+BTkZq+Ton21MNF2
ONzjYAOy8LBQXOaDd7lWasQQgQBXbBpSfkYDbg7Uwe1vWVwCiirgZLNblbjfUajxNcg7hvBGhqI9
QwLncH/Eg9CML8p1pcLklva5Enj+JM3+YbRs9Wje6Tw8ZMncZWg2xRQlph/MJJ9ZKuGhCRpRs8Xw
76Uzmo8yvMXdkrPf278NUDDsFOX1cPhBYaF/5qpO8obIHQWYL3dxSI9lNaB9QRl6BhYggySZF06c
QTdGCbO8A0D8wAOfQXmn1pQZYKydFDKBoBXnvjK8eLuTzNJbRgfzFh4apLEmw6tk3sRts6dMkVXA
IERiCJqrCl4XtvplN8F4+FTXa0IzfWVeBaR/AWeLi1YxQqy+Qgc8IACqNn91b+J4Ud2pNV5iyETF
MhIL9bjm6RFyAUSf3uHaCqLLn26h9v9VdSvIX7nvXXRQCk337NLHuYAwqwJlympjkmIF5pX8b0aL
15xnLiGiUpDatIFu0oNVgDqrx5N/T1l/vTrCcl2LnTwHswgT/C65TcQxF4sqi2opNe3HJTInhBvl
YSYlJdLCMytsowZAmX8j72OkbkfcoLabkMLrxTLg5GS+4VzG86CYb7YFAXTdwX0Ean/nsI+v/1dV
7ddxjUnll0nBwHCTX69aYW6NwJdcJ55Db7Hc5H2acySO4X+AijCGsShyXhit4okq7P0RS3M2l+di
Imr4m4zdlmndPUq3OXdLVTL3N7m4mFSpfeDheACVudNen8zJ3wh0KVgfXZqTiNqUcB8stZTj4IPb
gpmLTY2gpde6q97qO1xTw/NKjuRJ75Wl0BjgcuxagKR27w6QOd75KvfPFx2zuSc1YiDdf76h11y5
PoT7JxIztdT7K0KptTRYDTgJrLt0zaS1y3xXCLRIXSgeawOTBJSMQsBH0dzEU0lifbkr6OQgVbKj
tpROJizbHrY8VBpoSwgSc/Y4QNwH0yKFBEWELxQC8UlUXEO+gzL/bK66VUMVJaY3tFAJVK8HvwIj
+G7COVw/K55+dHSAwVMA8GAy6cXhssE3t698fqvOCLoY/lx9ezVKZTmEkszmwszDlyRGhSM4WjVv
OqS/huB2gFdyJDVUBsKN1F1tR59O/4422qjtNrLeemJ6kzo7SOb17ar2TZP5Hvl9mTVuRr04xNAd
U7a6KQ8o4S3LSmbfk1ufU7JZhsW3pdxi8y1zNzpki6/xemqiUHWveOhnLeun631hTNMNUowpq+tx
PMltdGj9K5xn2UJpWJs9lkhK7SBm9CZhau4GyYsUNZKoO9UdgUYs0oXTtss9qu6uLLDm76qeMfPe
j+JiFO31BKQd7fv+Y8Y0Y1Jm8sazbGnM1UtifoOpG3dPRQCVmiHswx5uRC0nln6KCkGuMTDQ3dDt
UG2qpGNfV3TuJZSsabVKJYm5hiEAVZ64v+0hRjCP5vzeWhNojXLr0g8CCott1ssD1ucxW4vo54MY
+D5mmzGPzirR85P+7bXrvaS3AEF2cyAD1pwep42fiph8VgCwfV3bi5M4OfrTsVGALRn0bkCKcURd
Ns/YRitLF+oX8/F/I+ASdLxLQHuKiSAMm5ZJ3Yx0x78MGo0zxmSh8snt5p/M1LevnUteGJ8DziV2
kolZjPus3ezyfJqKvscNVqg3Q0kcnLwAy49/1/DeccZkmjT6XSzl3juRzGPlct6wnAKuhFsz8zMi
lwDbw3izql4qPjAsFGQC1xcpEMk+/gWIhBLE0JCPnEH6W81oWMp+q2bp7wJN32KkM5waBIClOStr
b2n6kql8z4UDfMcL4ZklGrNf6Wrfh40eMHAgw7sYAQ/9N95rT56QTmlOT3JOEGulZZ4RljKWNxzD
FaCxYQkOWW1rlLq7QBLaIuQq/C9b2KbOT7EvkwkhCYxhcBjudNrCxNbMZYcXXSMDzSKtlnL2lzhb
J0D9xDKZVWrIdZKr+kPkJkZEpUhWY0V84VNu80wytMn8TL4jlDTVYN2Sjb0RlFX58l07mZvveggT
7OUT4bks4Uz+f4WKrXuSILLdCGyIn4UP+Wj2Tcw21mM7x4oqKyHYy85VXU1lHiUFDKYUH6x3GHRx
vGu0a+L6XD6L12hyIqZLzdqI12YvMmZx4Fw2gY+6NZpy8aWpF8mE90jlhgOoQzmSE4h9sGiu8/je
EWt7t7hYG9q321YeujMXBAZIGZocYMx1sK1Ge61fHDcCL2pjIbOgq3n8TICs2iCQkA499GRrz+XZ
52XNUa4GDQd7a8RGP3Wq41jJOz4yJrl1xGZzlKBMk0L3qfM0BKvWdo+xjQswBOcv5/Zn27VWW/Tl
VgtJY1tytPsF4vlvhPTFScW3HkdL/A/HlCDDyxbc6CR5ykJ0yKfsduY1Habjb9fO+idCS6TPVLnE
SNBPazpI0XoftqqZ6JV1GaPPI5eApcu44vKwDm5mbmANgBWGVZVnMkD5JU9omoMc4so/DoSuQ0an
pzpq4wVWghro3UwTxPdCe8OgZWrva3ttRg4ADbr9mEdRD98LnLbRLnZBuYm7DK200oYyktXB15BT
3FBlWSom2hfr0BS3mBAnJoVnNsnTGRGZpFvVQyNKy/HwwYYkKKujRafUTVSvdNQ2U2ZHQhyVyti8
DGAdVH/Mq/fEYEjPlSHIXdqL9vn4DZq++obRsCMAKIJEspGvgk7QKR/NjioPinvje9vDlN17ccYo
mchmzDoEDwNRh+P5X9jwOh8jD3+pmli4e01beVcTqdyAEVowBaVb273wtjDiu0JRjMWNopkSyI4w
zji22L9rj8CxZDYfCbLNCzcw9+SGkeRoRlVUviWBHhiXPNge5K9f1/XQxQGx91QD2X1vMRK1A7O9
Datii228Bc+5UE/UW+tRj2XAo/jUa/qfp3DN6NzDnh88TPDjUkZ7aoDJBxehpwzRR+Xg07tsgBsc
NUPpLoRuBQFWsvgxLrt4oH1kg9A2vVDNHfSYlYBIMB0MveAErSmvmsF0jSqQm/dUbh2ei86Ngk/e
RVcNRH6EddymWmKBW51ymY5I3hNXUgu/YS+HtV/sTdOqOdRp5fzhRKHSvPSlyxHCAScOlGJKdoH9
LiPm4n/w7fi+JH9pGzfX2p+P5Abom6bkFuGIAreaE1QcqJ81lQpnM5bk8w80bpv12vSqgG9vrGGC
kaav4pAQZXvy8lGqaCcuMftEqN8RIFeYAdmQadQdoIOg7Do8GI7qLjexmOkENW3sVXWdM3xLgMK7
UPw9JWyh7/S38OczoYLjhHtDll4n9k4co0iJ+U/uxURH6vBbNGNm0swYEfNi2g0djbDiQESu91oA
sgYfGmEK00NdwKEP4FhEPGMNPF5f0lnhGWZOLM+f41WqzGQqwk3+oM1JB2sy+FNCW0rbuPd5uEYd
UskRx2IlsCXtNM1cuK6H6spIvNMdKmGmvFfJZDUDs1VYPilQ4VDuQgU0gMicWoBV13FQhdh/+6Zm
LgBVZVkY+3yAcmJAS4N10QK3+DSN5iivX1UApmuN7UcUrnAYO/bHfuzQHmXgl1oO4FvK8FSdGBl6
xrh4Zv63aA8lhwUbMHfQ1fw74JFHYdaeXM4gIUrW6DHmi14Pyt4M8NF8TTxMBWHFi+ILiywcj0M2
TLFKlHuaWSN8bGq7vfdJ1Cv7k8MGebRrVKTav0QImTn3SwZuyKlM6dfPkf/LnGTN5Vceh08Lx2WG
jHp2o9Ni1JXVP0uJDVbtC8ZHVIT1WQJP14m5ykvzujRT7ejvquQ3codpxN55icJa5wGErSZTFdUz
olH8N/SsiNBREfMauJyVTiGQ053hQYdvBzfCBeFPVp1k++VjwuqvRj02XYDyBRGx9nPR3Nbu2UyI
UWFpheG5KF56GMsG03H7j8UOlzAw6dB4XEIwaGXECC+8oMYP/fOh5ZnpB0lRuvwCjKqL9vCtdSBt
6b7iHzlei2rCnQjiJz0k3soCUZHr/uWXkHVOCdnYljB0OH8NANrfWn+sA/mdWgN0XQwSWxzWfhZb
eiWEXBJs99omrkl293imy5VzOjACzSke3BkFaTERVpegZ6Vx0RguZ30juAf979C7ClJG/v7Ug/uR
EfiJ3nGjSht2Qno+577/dEiNUL1kVRAWgG0o4spjajSu9OYjy9BviFlCi48nUoEvmnzD/T5Rsan0
jZFXzg/RP88YOj/36H+lCfDqjus8NPDygDmVgcQknk1znr4SRaynncT/VyAaVvnz7d73C4ZVvIco
3y+Yl0QL98GmpJrSftVb8aufYrvNu9xLPGnMuX2la+XGt4FvuixWrsWRenZ9Bz13NP/iiBn38AX8
mkJLGjD3bX88aplW60/VcsXsvHkYhBvtxTqNct4QQKn6lBKNw81JEX301RUFCS05aFrOqiCvni00
R2UQgvLH6wOvlMCRqAkZKe6pYirVk1iYGOe3/3W8bbEcSOTGnDLL2ak16rIYTbvCBstS6INAoNln
x6UhG6p6u8O/lbF6HnHiMxckOKh0uCLXFACYAq2ip6FivFfySJZQFHDEJMMkWrGxBDuwsW8Mb4rq
TovHKYUK0qYgykPHDzMwTwqJ0TqSz60O5cO4iLI8aVBS2J2uNfz17ptI4cbsghFhKTdBKdCHgLXI
IGVX9XgKJFvFzgx4KMyyAtNEpBZ7RekOHTvHY24zzIP8ELe0JLcFuPAAkCusCI7hzrdaezTuW9o6
Hk1TCMjLC+H1ahTFrKFP/9/9BeVbEbrWEvEFsEwwMaj4nlpog7mtksYmGMK9c7eihwUKPiaOWbPc
hg7Nm8bDwLrvPODFG53r3NAwQ+/OXLe6MHyjpv/gf/rQi0QuZ04MpGr521thmz54Yp2iC1RODuEN
szb4TGBuLBMHQQWtd+rQwDmGfshF1nlz1DKH6bL5u3SgvRUSSzHziZxXfGGY5zAzRDj8j2dyiy9I
uAOY4GWCA1WLV43ylOe1cTPCGJVFaUVTtYWzrHGkQAn0rSyxJWbw/g4vQt+A9eN9lIpsyFG9NFto
VRUcA7+1BnAcqVrhh8uz7GIXm3mhnpx/AlpV0QlUz0pAR0pGPThHB3D6tc5Dim7CvCVsYkKRiTLG
dLYO/REoZfEcwiUTN7OqzeE+zGehu220mV3SInRnb9N+Z8WMtkS6dgsKatvmhPDG9aA6GqcQc4Ye
nXF000RdzvVVMBZrfsiii/+ld2f2ks4hrkZI9k8vgG2n/wNixc/NgByWQU2WJQjunKIgKCJvVbIL
3ui988ZGphabIsJ9a8BDPZlekjxPE8oh2TprUscOQM8w1SMqCP9HIKv+BnvFU/KWcOjgMg9GszHc
699cJjVwswDu6BS6EccnijURaINjpE/SylGW+u13XpdIWkjDrqtInJH952BzxVbInXIRgMICmEgx
jDiUWixH+MA1t/EhMmGe/jBl8EOMTHejqtfd5mWZ1kSkjVtDoTTlCUZcZS/CEX7d+DC6oPzeIqlT
yk8yQCM5dmtc/5RdrDxjEW2Z8p7OEvZnxvfhND0sJXVQg/h8k2Cl7RrfnPxmpAA/WGPg4nTdD90g
goKpEE0f2DWPxiui0C+aBWbnFaAUV2Y3SrfFslOU2xOAg2HOz5XT9YyBsyWxbnIcuO/baeOQGObV
vOCwDu1JnKYXYJ6Eu2dgnEW9kCzzNmvoFPg4D0emZ+gWwKZK/juPEDfWpIGmOhmFr9z4YlhdqmNZ
O0Z1A6vpDq1QgEu52C0Er3MbY53VQHYLK0J8PJ3fTCxTppi7j7GgEKnCifWTujkd9VplWZ3kLrL1
unJAmU7e0B8iMOQNguo+lG4haT6JcpldBhHyKNWvZGDF2dru38A8iOOz3cU16HvR16jjYW6k9wW8
bMyWyI4tmLNnY4HXTyXu4Wqse5BshmEAbr/+3+POBLyGxG+Uk36C92P6ANL+TIFWnlxAnQTim05z
nmaxEaYJIb1Jntxeomw0L3pS0M+wh5lonKxe259gDztzCZic/VkER7hVNMcC1VSQRIP65v/rStwy
hLOH+ce9EGJMZ4GMVXVZvt65b3ZEru+W1eOvP87/s4uFvv7+L/VaRLO0rYn14IsZVT8M7dcBBCGB
QEUijnDpyanP2P9q07ccw+NOMkPJHiY89bJ3+8YkWWLvPcaa1sJrAOlTHdxGKIVk3bRe1n1ziRO7
JJW0Df4FxQFH8vZ4hLTX6rax42HbXrFNH1NEIhbJ4OrZ9wTf7Mfw7bENa4KCme72YfCZM0SqCSC8
YdjidMiI7zrCbmeRTFqJLJ5obp5qsJY9BEc2ZeTOF8YWxzSYrCXcMS2hcIQLVDRGjXZ7mlhPBKMH
Dmw7xUQj0L3KBIg9p6YHpcugYHBZDlxmvXBQo3U80LgjTzS0XF08jnp+dOx9EshZnsCFo900JOML
xYfbCqnsqk6iqU5m1MIZIwUnhEaxntmDgYrTmLVYyNSzF1GQkDtYhXsPeN6gELB/2vdfndVlnQOh
RsuMxNrOjNSkhMJ87c7+Cn3xxPyz1vJ5/BcQtREw9FFaFhHqV7oYxtAF0FjdoqgcUfEFDmfStXcu
3PDlF4Jj8aV+LJ02mjJa3q5cUkBAQL8HKsJXSgmNi3L3KCO4rFU++rLFee2eju2jt3Bh3Ssn7NOk
vvbdbCDq8cEhhYXvNHheNXsTP6ARnC2uJmbn0MHqKVdq+B2mhPGN6JEtvR6r8y3QT4+ZT3DP8hf2
Vbs+7RFY3Yss9dE+w5V/GQxT4ES/lH1jw7fYLFfHTvrKFy78pBtOeSnpLqPapuC33wLdE63JGqeZ
SmlAheNb0XTsAl5alzIpxdTcSz2OHRy7ANmVpqhkyB54i0brigx5wd8OOHMyRwsgL99MqhsUUfEK
v6AwZeZeHI6xuPHrfz+Tu4CXjonmIl4UlfYAY9CIGLe0j/NdK4RqUKYWF1uxRvFReRJOQ9WoEZm7
ZHnYbRamXQHBv3V6kbZdlT/nUTRjIZnMmI9Y1iyPzcS7Q2V/gCn95geSsM22QUdg4fVQLJxUtTSk
k6mUS9G8QYtnPT152wmTkEQ3TL5BJwE0W1ESIjFzA+TXF/XM8+ffAxhgfyQ2G6x1t3iwBHHyZqbg
MnIWn2+4U47WH+TDy8VAbdd2fEpJYuX7Y3dftDVO7lsQhI7qdYrY7Fl4nu/mSMEiO6SDD5KC9NFj
sp2ZU7t6uV01Vxv5yRhZYvk0nkZUyPq7xc68yNFXUiQ+ULVt8wqLOj871I/APBrcr7CzvcQN1HAZ
PZz5r/WMSCDrKxfO+0bgTunFqpeKjkropG0GjXmQEHsABuf6SKwXvAmCK/mlp8Em0/UjEAqf4eLK
UlUQmCqSBBK2cXOLeCeTjS3VslkXPXwumklUx5xJKLe+4hOCCDDZrc0CiD3JfuKAUqaLZUKbB7JG
AbdTwKTT8/l368dDcKZ6w4Bmw2WwMz1stASpTMAakpJ/EmMfs4lMkW9WRIiG5uKPgNVMPT17mRNj
MDvVZDLWyT3MUheNW/EYg9IRDWuioKJ7uZ+4b6xmz+pRFrT9B92jBV3FZAostPEOBF599eb1L1Ol
W77Se0DEaop9ynIhHgkDOJDv0BcD5TzRJg6/dwVJVNKOVUgAUhft3y9zwNjtdrIUFkyXEWGOFMXj
ZtjU9VYZtI8bNqy2DJtKT7F05DXJUHoLIHdhMJ54zei0OXLCGnfQBWWDtFApJn264zDrGj7X3XaD
X65O3fp9wR2MCvTz6nPUpdUYqAr1Lj8vJ7+FSmoZcHQzTHXqoCqUo/ySpJqh1C2hqiAM9nHXWEyc
ibPzQD3DafwZowWLv22dZ02O4hZt6Ywad1KN/fhquaBhSt/IECdZn5kHEt/wnekWxfrzzNfz5gVz
+Ts7kOMdZazm6Bg/feEaqf0zVSLNxzW6zwRh9sYi/5rQE7lGG8xkYaNWeVTkZiLbveEwLMkMX3yp
5ymBYIqcZhrsA83/w+e6W6V2VG056OkCEGQ/P9bIuo492AeXauwmL9Jz/uWuHnLAAkX9FxAyTVrD
gkZBBtSh8fasU8klzG0wmb2QbU83himQ14GCleLQa0Ac+rMFDfZEB4JK6qGQDAjHM1pc1a6ib1XK
K3MQZeCD5fpTsVn8El1NHldCcpKpwU3LJ6ew4NHckTBoopciyl1UB9w74NTX5hFLOU7cfqUtQvWa
Iqiq/DV/Zm+gGIKwG+WEJU+hVf1L3pYxB1kHnR/ApM9qnitUsDe4QbLlxI0jrGwFU0M2vAcrtVCK
SlltxsmnZDPGwXpfIW5HoUvqQhRs30s46Cm4BRAPhYhmR4IOmHuEjeU4QZJBGixVICxqyQxOFLR6
inq0GIs5bL0o37JTqdZJ4kepLaYWlt2PpR9tqV+2TJghZ7iVyQBUS2Nei/yWHOR1Nz8lSYmOyQN0
V/1SZfqgD1GxSX3MqF//W3Zlv6W1GR6fy205sGf/EdysGBilHAB9ScnY0mxYkeAuT6BR/A6tSmni
HZQr4Z6XYvClGlm7j6ruwX+CJfsQqVhvsrpNMdLm1aTQL+UC/QUanttk/BwlyRAleOGu2iRjdKn0
sFL+PqTvi0+9gXovvoqeS6E5UAY+OpX0xQZRvaCp0VdMjI+CeGuZfCSSTN5+oTNVp7ZSaAEIKkSC
kd9rdHjKHuYpXuzaFdJO/Kg5F5eez9g+7So76Dk3V4f9bCNc/RmerFJlNkkWM1xDRwu2uT8duOki
IN9RRKDFfaS+M+HkKvPAqAiQC/3Ux3X3MQIbYKn4D3agzKEg/sFOEMF08Z8PYLMGo3foPzE9FGkb
SrGOIytELfh8SloW0evQzgiHjSvXgEx15NlPtm+s0UwrnPYPqgicd460S8qvqaDVaVSF29JLOmdp
7fk4kNScpsyztpe9CbC7gkYnQV9r7rW4tgMBQHJ2h1dCblCrtjc1ONXbYn45C4FKRsdRI8AgkjGE
VkCTuSqkt/s5R+45vJFRGI/DwUH0YCqXnYXgAcv/XzYhJV9OLmhgS63PzUiGVqrSBjqYbhxhf4Td
g2srmaKiFZlEAD5+7RmQ2zc5HAQv+wt4A9SN3zTrgubt0FXie5M0ZPKGx4c9YWCV04v/K0t3EJd0
haq1nCFyYTJaCYxDsrKwmG0N/GI/Vrnq0t23ryIa8HNs8ryn/9CScaQ/RQ/9zHsxH2xu3Yl8TOLG
N4BHnWDSVgRMNaQopLmJ2KkkQ4LBRY7I63OA/0hT4rbTtHNCBUrixgSGkdC0OYaxozKbqnrqy763
suWyR8LB4dykmV6j6GsgSjxcbxy0y3RiTwAKrvpecxJHsp3ObQogLTmI7HniVYQD6m9nRwCJbh8M
nCygaxlqGvU9+qWaYmrNazyPkWxR38gPHssDYS/AGXyfFzIPG5UK0S8h0xyHcvNze3Jmj9SNXGtT
ttGNYqVU8v4vQURiQpNrMFUmylGN26SjrNzSpz0+3n85s/fiD0/vK/x1p0BAPA2PQ/pENFPackRR
qeGdTyZjtzwAlpjOFttdHJHgi2fM4sv3NlqJnLG8Nmox8tsIT/nDKCbMuKlsktAiRJJEruhLWhRG
BBz3TUN7FcuJVO/dI39Gi3fUMfbOURj7QxFpjZ7YYlnMVblLstIGqpLNv92tWIVt/OPUSpe9UaIH
kErwO5+DiVvEndBK4/hIX8Xtd0mmx7B3/TQ8PJigr9l55SuGImceKMxI3IMEl4tEGP4lef+i3tzS
gYm3s5Dz8Dg4ODLXu8j6X7yTbbZ8ZsC4hghNSL0uSTKdZ+ftmQJRTXOtmUo7bvubdGucWs8jHCyt
sy1OBa77H7JYoiRqecBlsc/wRmi8sfC8T0RS0DH07EX9H8PBha9gkqa1RHFs/hXfqmoQbWUBIBOG
G9qWLDouWLKXZlTWghrj6h5DR9kOQEP/Xjkue6sro5zRUlDzJDPyNde9/ESS68rt/cJYO5pp2zn8
IByOAWvXsT4NmEZoNZHhjFQTUpUFB2TcX4v535kgfShoXeLBLQ8FPos1pVVcxo/1nESNWiICy/JO
QHkuzXVc41KY834SLFYPHVMCFAX/WRnN8CzNXlV0HrIpnLnCJFEVPCzj1+tUQTWCyJbLVoNnIld1
0lnt8WbAdyQ/BC1LTMDrRsvoMSNVej85QIAH0ZOvTrATsfY7rgr6bmCsklah6w+GJat6Qgxpxv+J
zS7hiD5HpuC8JxNv/XgeDnrRVUJZf1kgUkqB4gBfdrOPESottgs/PGZid8qG2c9yO6o+QLt3oVZN
9C8ufBmRgKJ5fsDk+nzaifZxG05rRzhy8200SRwKk77Td7w/+Ha/0/dXt0tpJ3bkD2QNcEjwZpeX
BI0VMWgCxGrdoGyt8/ff68hfeFN5M1LgHHI17L/G2LJDZq1PmJgDjB1uCbMj6uzS2Jc4ZkNiIQVr
r/EIn8vQvv8WLrdhVHqJ2ApJS25/GnMVj4w2CNF5YvLGE/DTQQG8f30SIKO808webNgpA12Ti76a
EHBMRfrJg6U8jRe5EaCpGQr7lk+WdRpDLglNoiDkG75GoAJVdxAf2hp8jaENmOs2eIy473dEgdwG
TRjKWs7VB4CGcLGOHe6CuhUtPJhPAthtuhdPe1ledyQci1/SbzUbZt7aFkfNnxvx27L2olxhFd18
YabEwJVXA8PLvShnOjBVWo9L9vwCT+Y6CWxHpfMnN3kybXjlJQioHtdUtwRdJB8A+ven5B1eecus
Ou/9E01s3p0UcUTyen0gFBW6nnho0h5ZNOVa1CYIT3r/djtsNMsLuMZgIHQGUKWzQ6l/crfIYhme
8aREiFPzoKMXaE1trvOIuBFs0F5bQG/rFvjbuFZ4+jpt/JrA7cCLDn2fi4yU6pKaP29e5c70EqMM
1C8ZC49lXnPX1n5jbBzXa0bseo8SncqBnYIMGAPJR1x1taSMuNSFf8J9lT0K/5Zem+SazUiO8DW9
PxXSmOkjKkLFjCyfkkCU64eooQh9sN5O68UUZa5Qkf54YGBT/W5T6Cp3NcPW6F/K+RM66FpqV6Zb
ZyC5F25j+BPex9XrMlltI7VQKWuspTLke6jejKhBDLC6wAvVShG6+gHj3ndkkskjldu7jiQ+WsXB
K0fEu5/dnXxKtZyBPc202GavdC/kb0NdhgEJj6/LO0HQ3nzyeKYxYuivORiB9kfhESmJePCtecQW
+MB6mCad5YDj+uLz19d4xkC/60aOtJ9fOxCdum28p6FYLEZsFgHKEftwsXZEb4cXkIFQc4DIsaVx
kNQHX7kX7+F0Pv1wote4K1ckz/HY5bsmYmp7aWGcWujDBF/YOBhhjeuQW7z2Ee6kP1rPmpuh0jIH
HPeht5uLGOwlNNfqbaDP7vv8AG+jT7x+V6haz2OAhaMx9bRTVffP/pcfRAldgcejB49bVMprkw24
LRljXSv/dIKVVnJ0S2PmmHKqojqh9fRQAra9R+uN8txu9t1L5fxVWtnGpZNfiSuCew0/OQrbtp4W
l1WT3DriqMM7fwQ1vlUgpRqaHEXjN0os9RydlyWxKtUnRUamtYP+2keKuIufi12g1GDdnvwfCFO0
mztKT5WoHmclVYN63C/JZObh16bHwWTgZUwsh90urqLXDIbMyWVS4f9sO+1wM5HwIdB4ZJjMd93z
jUHXD7BcMdCviiZaYsxgQJsMPr0RzEkZS18BJeXSoYhiJwub2U7gd5TxTyWZydtn/G4VMmA2HH/9
6seykuhabUnaZaHOjNMYfhpc0CcJPqE0+5emsTAM+ULI0UuYRSUpeBny4zP/kAOSABj0+wWSOQ+6
ntwECKUgbPQr58GzujvsCwUsX+ooMRQERAr23G+jkMnitSgvxmjrSzlttG5+jnWp3vPEJfc/J/Ge
Fg76AzDdymCs5Zmb5+LptE9LhJJ1lIqAirnQxFS9YsYTscEY0EKPsDg+bxXIvwWzbwd7kAbdTrHF
xRAyNRywILaJXEkod6jI/owEKujzycJ5OlG7K2kVMLb3S3zKBXfT1b4Zwip2UH4qqNqzJMmqFR7B
olPbsMX3Dw2TIpRHSgirqQW1z/kA6OhUkxsPdvFDmJi+HFlT2tYyVSrAMJyu0Wk2ZUt6YGNgxEri
wCp+bLoshCp6QY7KZGop9OkkaUD3FWP6G6aR+WtyxHKBp5hnQbYJbdXj5sCnP2Ti1kMKBDpfA3bG
4w5OoLoX3tK8fA9P/pJX0L+f9jvwPSYyBBBMBKmvN6pEfSRpj6cCdti9+Ldpw/pZ4mf++uiUk8id
bCezEW0whE1i6iB7XSVtu6Zhv1T8hwjBEw08T8Z6e8d+WlGcIi8uZBqIphWJoBKBo5LsLAdeCXIm
NN4SKiyCemdPDdJsFTHGALpkFYIU9zFx1f4vJ8fb3pVXMTD3FfLV4/XZm/1fGPYq3UUqdGBXjVMq
BAz58kkNAeiJeV5L2Nmdj5r+SdM/wg261sFQVH0Wi84ufsH2LqgBjLpTJHLJYhk5p5dPOGOq3x9O
6Z9TrZfVMveG/cc1HAWOOOgDerGjeo4lTBgfAiVzhyCP2k6ckTeRPxuyncCMmhyQkfZcGuWhwMtS
YCiPyvEisFSDpIamVtJhSuWtrryFQDDrcVBn4jgxX4sbnjFC80wwOYBjKFAp1uavncTAVltzBrt9
xwGAwBD9KyDFU5EEd5iUispgUP4W7oydf19SCHabbcPNCOV3kZY9IUguu0Wnwn2GkS8kkIc7mY4m
w9T8IGEwSEBE+qwYkFAMvryiV0AlcNXIqFRHJ4R/vxSHrPAXWFTCe3xq+vOoMaAtdZB/WSBzwhO6
NLbItMCyFcVBVN3H2HctoLM40/ydZ6acojP+YCV6/fH1V9Pj+swwtT3jwq4nsn5XaGiL25W9yhBw
yYkmezWVsJow5mjnJx/l8U6o5mama3GUVU4xdIo26zA/rpMKm0ob0gGIQk+xaZk3lf19aLntP5LW
NAh+gehxxZD7DlslQOPmwJlT2iZzsVkf7kjF5dq3v/umqNYvGcbYwhxKFuybKsq2gNX4Tm93Jjfk
YdsV6wybZJ6aKJvzO/jkSfxbIR6btBqL3oSfFiPGrouXhuzaHQGgY0c8W0vxY55omLoNoOUjgXTc
pPcc+TRjVGIifcvhVvoT1TAmYztWzggeu7Vvn6dLm8Rg8A6CCVpQGCe/vQxh4nEZIhvE8aI1K8l4
sP6ecq2yy2HgQBZDiiFNAfo3j82IavobDKjbPcvbbu2QbQSXS7Fm89epmOmTvKsawC9LzRrdHuLA
gcL9TY7Uet9HRyLWxgfjVUMMie/eAWkfPnL/232dNfvtz9cf8ecyptsT8w3Phltd3SvZCBjEtPft
adrh7j/5QkVHWwSa6DNieJgT04z9gqG5WBroIysSuJ7/0s/SFoTMkznPIwFLvuPti/RY/NqNq76K
rmcxYy6BWpoLiDUClNgQ6I7IOPtHO96z3sRcQ5xBEMzlEttd5XQAqVed9MdLmJdePHu3HTYAGl3K
wzDPs/rhpZ+PCgVPo0ahakO4lyk9svX+nicbYan2PhOf88kqXgJaWmYAx5AXmNwS+Q/ZjFWtpvOT
vVbUZfdIgAvqM6aPcgiZ/XDDZmqq7H28mQQVN85KTRZh2+qyFF6aQag7MhWXCMSi2aeQyrNqG1Tn
U16CFT/Gl5088f4TGuYlIWLRV1csU0fi4xNbNA3DfHjzdRQEB7MuzhSU163zSyY+hqelbNb+0TtD
2s5nNGRoABB+SWt6VBAGDXMlXwKCeMVnt7yVhk5nmFI1BlBLTE9UOlJgRim1eHFYtom7BG93iDwe
v6AjW7ngI8jHzl5hT2FEt310VQqRZ4Mzt/y2UMi0RGfryP8rClTVwMWbW9Fz9JxVBLfkFN2ee+oD
HfppGZij9sAa9RCqtZODHe/4cdfCZ7aI+Wo/hw8DzvcvWfzo2czymE6lXeZ4eBiKyijVzOKBOV64
wwEHQAULePwi/QjFhiCFsuHSTp10r+Mbcv6yiZWXRHc97NRpqgjQlUCR1yGkxnSCcHW1l5IQ3KrF
OFIFdjtYdCp5DeytHaFfJEndGfIhS3ODCXJDOwwvpR6MNc0//0M6Ln+Fgl+etNdjxjd45h3kTQpi
k7GL5YfieZ/A3UyyEaEBfTq7YjKpii34roEKLlAtsyzm9gbdfvhHTdOibAZOAwgpvxfZrbm9i1Yv
PCzEwSuP9E1Ey+5svw934tI7ss6AQ6F2spvuVjJs5XczVwJn4fch/DE4eQ8xeJrWQ7E1Mo3TZ48s
yKnAofIsYVemNAeK3T17yJVgtYMak2AZqFl4nyvoJd1ivmsx7maeLuE/BMDgF1datzQJTBL3uIl4
mHRA5teWzH78fLBxnPqYeifrh2vJinZoAGrBIbh+/z14z9E0gQ0/Vkxp942vddmOb1u6wycEQ1to
9zvT5NdSagWKfRKBLv/HgS6CPHlt+hg35UATDesZYyjfdWz7l8Xikv4fjFKrwxxwK06OQarsYti7
tjTB64ilNSpMEnfkcwgk/TKLcTrRXK7ZGDUZBtzWaNj4LIg0FDYNiIm0DvVhIicXoRlSS84JZpLW
/ePlL+LSVHXYHD/Zmvh1uGP7Z7qmNUwJlqwHMyZpLZBmygpXeFRScYHg168d7TZf8FoucOzUey//
NdQ4LXkBm7bQ/S1Y8LBy8B0+kmiANbgYUmv6BLX/FJiU2rJ+9dmoFdpwKcSBBhMMqLHB4f80QI6K
z5gYHsL+4Q21OwZ88ltErSdyZAmxFGmws+qm8wMdhRrrLR1mS5M74sTb10DdYGCBXAPlUAP6b4Nr
vKnDWrHwHQiahrD4aV2MhX/mJyNtnzuBqqG3c884j9SUOr7LvFy+Gt/KlTjnJQy7DvNCL5O/e3ur
Xf4TsRdPdO7IjsLMCQbTjjf/xzmhgz/osKxY5AJ17WBKqt7FKt3Qb4/GvtkefgxSlOHkfRLvO4jQ
Mnk7kU3nM7mncuWHYFmMlaHocTExH4rxVVgOMpvDpenMoI/5glHFvj+7j6LV8Dt7NWFZLZTsUWmJ
51988eZ4iPrNZD8A2AxTwYzs+bQcaxzKnSBv2VtvT9IV1F10jvxXehDGGQsTTdD6X1tHHfyuQTWg
j460AL+kWFdBSOD5bOrGHGRT/mVtPp/u9EHwd5FHvT7PMJRpcPayWE2C0edVmcSaxAHNgvDgM9LP
5Qtz83/A3WBlo8YNSXsIo7nj/d8+toghe3++3CrUGhASdGY5IT/WNxTKukXeXicRDUcmcAsGwCjE
ESCuW4Qb35T1ET//NvNaC/mVLUHAx9KNHyXiS+uNj9l4mPOfn9ppQ4C6+hmPmIEv0XDWsKB3hudI
Lp20yozclLy/9d5Yr2dGJBDSrNJg63M38dtCDNzRtrqSCFr5Xe5uVOc1VWDNdyti4KQwRg21/Aob
56m8oLCAUx5jJyEwmr+c8blEYC6p0y0BZOSBCTbyt8kX9gHZqmVTSQS54WLX1Q1tqM7gAUjEc+90
TtaroxruBV+cgsTGI6aiX2cYOFG3MiP2bNJ4+8k1oe1YpCNDUoZWuILqPQvHl6sVRpuAOXz/Cg6U
kw+auxEO+JdhAOA2yriQE7UD49SkMQla/MtojvF894ORNjOtUSJ0zP397hIZqDYqlJea9gSXx+qm
81FaG6qs9+fHRDGgBWsZ/Px0FuBuUx/W+TlmMHqCL+l78mk7HPDRNmzRiIkrnAadSP4bjjktxCd/
7KOLCsTb8RYVXKWOGSlhPrAHeBO3AjqJpZoHyIXq5b4OPutROl3ARUddDK3RDBffRoYzhCWYb2M/
1PONr91u2/JRLy8NPUY7LMoeMRD1cBsyFH/HxRbcqIAQvtQcl1WiLoy5Sj4luKJrfdVjkrcl2pvg
yTcdpCBHAD1cRmb3YhneBxJbl74MwYmNQEKEZDGoSO5NR7adll/GEu4aEQnPl8YUlLUPkZTShYIS
U1e/V+YcuSXAdmZU53e7IDTwEH5NSsQYYLN3rytd7YmvIfAB8H6uahCA8ghJa6RlUDgSql8SEUMi
geOMA0dcGsPFR2/g3a0zl6OrTwOAp55MRllWjxZ+LrcHm93/vOOLJLCdQd0pjtJG+064uZENoGB4
vnTI7oR7VBRE0CkvL2KeYrw/cTd3F0U1D3YhBL1CMbnLCFuHunKzPlhNxEyFXNkGk2qEwy3FV6WJ
zUksKTwdgq8nvzBrFag2EoQbQTtIAcvRONnGtiueTVOksyZx3mFHdr18nRUiQapYtCtl4ZwRrtta
uaKbj2o4hwhO15qISnP8K3vZNL913+/TM2UGT08ORZJqon/47+xgv7w8t1PLxNTj0ZuvVZxulzB/
a4VUgNnNcG5J7qgA61dinTktWxR8IzvlQYusaGIxd78Bc1WMyfDqxQ0gYC2Jx2ueKCoJL1vuGnSO
5T4Pp6VxMgTGoquWqs6Hg+11TYkDrCj8hdO2bPMz3KecCuKkrICTwXDDpVk/wO01siTeTwjf55OD
vN8pJYxpjaA4hT6cyxXZUo1OMl7Oyb60fYqv103WA6xYe+xkNnsPj0f4ud/qDKUEJvX6OA92gVKb
x+RqDzT3XIY/9dEHAoLydUP2ZXALjIDp2bfI+Z2PyOym0vQscgBRa+T3wvExA6qNqTQRDff4idBw
zvJ/pFuI+bqdM8YQFC7cNJUDVDcDeBIucfzPOJ+8VQy8JJ9WDxOD9dmLMmDK76CEuVDnQWuh3bcr
pjydQ80UZZjTv4yP2dw3o+kWuEqybK3J2WWpyiU7q99/5JDgLRIEsOK+Ey1XUTnwSvoVN5k/qnvL
Psz2jIg/LHxiIEQbC7BgD/H+AHx2l9M5VIKyt7jODct19ZMS2lPxfV7EcMUvBijAdYIUiZ9+SOtm
12Ke81KX5jXUg9h2B2tFDirsPoo3e3OrNbxAV3Bi9hp1e9mvs56getF/1VOSCAqu+HnR0gM34sSC
IHhi83OPH21z7FqiP6rWXXLeI97srvz8WzoOejVeXvtzl2Va5K4+i4goPQcUOB/45rgErYfAbauK
k+U5xnSEQWnYrHElWp9hgMNjoyvIplbH/3X4Y/kc1mByyGhJRCApnfFF6Nal2pBWnDOYdMb4u9Ol
DopFzdrkDoiuzxpDmgY/f9M+Bt6+jRbeRxSS7Si9ViZ1+DZx7aosQQ3zvvstg4qckpQPl1cF9DdN
QxV1H0g1wMoFLvkM9TfY96qsGLuWaxWQ8xNvQ6Z21/YRBG+Jv2vfvR8cr0lk7gDqY69J5waNw2Ct
T+DOeiOxb9oDIWSzN4Nm5Kk5XoBfrJ7AxAt/i7qBsmiPlfv6OMdDWuhwwiIcLA5Ox975y79Fd3au
LvC04NL2+KiAsvHLXbwGXXnnO4dNLHOofC02VGmAj1b/qJ8BVEmV7lc0kBQZklAHHZhPSAEzuY7h
GZ/QIDJzqaZtmUteVn2hzLDQ/KNu1Z/QbT3SiUE5PQ9NxYBt6ti08utQSVvm/JKcp1AQ3jSNpojT
8rZ+rIpN0f4x3Co3NVBBehwbSCZAHWG+SKzNIn7z6g3LKwLCX5/MEfff38QWAN7Uodb/n6SCg22E
x4AwkKuyYAZR1jTmayx8pX8mOy9knTwgEQb4/AC/qq3mnFNvezWkAX0mL4PYY+P76N5qpbOKAWdy
w+xD3+cXo4vF5XZYgX7WhQ4JLzwv0hAvcHj2zGIbS0ShJD1QWgXhl0942heBLQntz1mrV/KiyM82
AizNAlTTLutUZdEoxKppHBhLedPWSVX4BzZQewNj12+HkWu81blj6yFJYgkSy5tyn52nDOxiJL7h
VQz5B8xTlPbWcffv7nKGSkrb4M9QJX5H6hecZUps3Lwyun8bbM/LM6K8f9FOgE3a1O/0FoIYVXrp
Voc/uCtZfYZF2U76NQHxp3rhWQXkQ6S5kXxN2xzCJHjhpsqkpvgdJvosTs2Dy8uVrX0wU8s6oEuG
rmHklDeA+ZmN22CXcrbZdUE4UQDEz6tMdIZmkB7zCkT1DBwRFuGVxJLwwxNr8fg1U7xa3WSeLsIv
dk+/xO02FItEocdi2Raj+9PbeAEfrNFFIhGaLkH1uBSyeMo8c+B4bveWBiF2Hj3wpif1KKjI4bCe
fKcNbuhmRJAVykUSFf9oMzDSuHkeWCgnpG55pgndFIN8IYJE058ku06GHyN0CIorO2mzbCfSl3YF
v4QE2Uxm9I/YChtKSd3HSu1+AYfY/Q6IaeZ9YZFPlVnAi+8v/WsRIv0/86aWaISiMYI2s28+gxAA
GUDlSNTQtleocugAslEiba8TxsssdfNhei7iIi51F52szOg+NM7nelX2lGDrsIcT71OsLDMPf1Yi
Y1//BXJQ5SydHBBFh/Kuooa3GrvDQZ0+yJ2DrjZTJLyUJkB2UYEdjn2kUQSN3sHIsSiJd+fuZNb4
T1Mm1IALaUcMz22n4v9fS1P/9yXcACtd5bQa1BjLVrEfV3Zl2hHoodBFYYhtqB9NGQBAD6mFHrT4
HNrKBiPBCF1fgp3iFPzgr/8AEToCGjw0xXA23rKxf5ddsuWyPRCjeJ71hP54HBdbuHSx4eDmf10z
CDt6N6qQTEIQi235uD9yGZKPhYo4zx7poJjx7i2B0XRK1cu0onZW53t1VoORjFhRI1UP8OPvssWd
u9TiwGtGHqqgvcHtNjiDqBi17l4ZiNBYcSeWqXoGPbXimvBtD2wR1ff8X2KUTW34/LllDHg5sOrq
/cIsisjZ+SF3HOZ7s46gMBsFGYyKJK8Nj1JXYykTw3iLXHQdKLpt8iupKQd99wDfG/FB8H0oItDD
kSFFrBaDv/SUYd0dLZjoAG/XbK+E+ALjAMlg6pzD6iyTOX1JTyfffTIb9HQacY0ZqCgtzFHd2TNT
DgysuXo6TLtz41yojL4XHNAz+q4C1aJePOSep2tJSYEQJxCbCSWQ1gK2Vb3zpuZ8hzJ2dufsTnfe
FnPw++OHSV+Wy8Vhd9Pnd3zpIaCZReuKWj5ZUAWIAXHo4XC7eu0DiFGUgWXgW/tnloqDLKXzctV3
gHBUx3ttZTo/qIq+eZt9FSa7z0WWhSL605I8cTqwCLly4evPBs+7OqslfWaqOko+eH+Wm7H8D6DC
KptcER59iVdG8OytztbC/+s+0+H4a1D8c3vuCQMUQEz0b1AE3IPTEL6Ci//yvGombwCJguqnvF6P
KQL49W3MvUAGTxCUGFSx1ktaQXF+mG6t4rkWfd7QYlqGSG+9+MvOSZwbfNJeRc+yb5hHyLoMtmYp
5ai+MWBNnXrYgP//T1PTsKvtnK7QPszisrtVb5bWdSeL9YVBDcVO+qSgnBGf1b5k3vBm59aLB+ja
A6eCQ2YYXWYw+ItuDulwSP3MATis43y1O1GoLEcK8t+TatelK9cEkf7taj/xdT+4RkwdzqM2Jb7R
LEmDKnaJTNYgVWDnnd0ch0RkJK1U2Tqa6iL8x1NBbM0RnAJAENbTF1App8aH8HgCjbsK8ZZJEc8e
1W+sDCUlssCU1VOBYpQ/WnqoN71QlatsOZ6Z+DvzN3nYFzm2u8beosijgjsSmnSEDfW5yQSoETDC
BAqtXMd7c7goG59MZxEgLXWLqVyL/wmSPqUAz7Hp4Dd1tSgsUQmC19tPcdUZLE56X80vHTsmvBLi
qg5qfVAAI7PQy/UczGz4onDpibgA6DgcWtGYDq87sn2WIBnl6CGPcrXk5KmKVSzy2Y4evP5SBCiC
0ANKgeYHE+jJSekelDIhycNLZSgkvkJiy/bC8ocfODdIPcAnlrnnlZGtpDVRsUorZ0OAAUKkdbRx
yFmo9eiUYntMlDtDzvvQw3EdvQiGUBXNzhDRUaoqvLLsvJlstKA53q8XbLFNH4x6tkL0YdPUCcuO
E36XS0B+QVIZdb69Y5jbu7oJuPFlCeQb0X41oGuKv5pCY/4eKP1KvFDaDEprjTXLreFprRerd52Y
mg54GeZnxKGMFnNYG1vv2yx194VBRjToz6xWzg4oeGO7QxtYR+gj7F8d87BPdcLFCWSWBEPEmkn3
SaTJ4CZtDon8dfBNGaWfI2jPP8A1X72lHJ3SGIvsLTUZFgQnGR4FtZtzHoStAD+gUGC0ZtsqVhaO
+Tf6TDl56hIF26iNX4oFoUs4jSBldht9TiETjJh+Y2OVgKrfsN3kjUONmxh/+D2dXPRRC6Jr+jQv
k20SlKv9r1tyLQx2R/4XXLHPaQHLsclqPuAYBucId6shIkoPtsBKx4T0ySKggS4l++cvpGjzULYp
Zy+Q+upwMwfeH5y1lrugkvXalp1wrZ70MGbGcJO531yuKT3Zc89n8vAr3eYcvLVpe/De2RJmkXj4
A7DEU72Ea0wymMiVPstJ3u2gvlkzUYn8TyOHd1obYsxmjLjunmRkaG6hp/u6Fog8t2eI+myiE3JA
8UgFz2wC+JEakQKKFCmdlVhrnHhqj69Ojez3I2fXkanVvw8Oz9LW3/vZimBo9GJWHxMe1MuasyHr
ua5AdMwdpp7FaV18o2prXUZ/Br4c9Iq7PK8femGA4rk6rMNgiHf+SpXxxfABHJCAfzN+kbUW3qvc
+Ss06ax6S87Vgp+bF3OgzkwDWWnVso0KoVH5QYf8iR7yMCFi2d1ka+/X6mNouW2qTPlK85/LKTl9
Jy/6MvzGm7/GQ95iirrGI55KhIIPi+ZgiMSC4ZymmobQzco4pL0mH5G2xXduZVczF/Qg3//DNYrR
QjIPbJhrpkPVRQ3rTjERChJTgC5CZ7clQ1rSxw4hL3nxYXlKGInegx58UUjNqpeQuDuy0ryr4MhJ
YZuYKRIAAUqD5+hGowmsvP+f8GrbetGEVcGeqbKUXK3cDEQBl6M5fvgRaPN6elRWKctbUpt5mpGD
KBwa7CkW6OPSabf881LjMmZiszM3eOaQzsD6Y/7DzLpp+tYwo9YPKS06HezoU45/QRpvfASFpBSr
BUzkkqpTPudb0nTinaR/VZQyK4NO0DUEzgPz5xJkyKJzANXTEOA3XRajXiCh2b6qiHiWITQBu5b1
qqpiHzH/OgK5aEjRXSfp0swa/jtQU1nqT/8OuCBZTexgc80l09Z4D0/7pUofz3lU94mlkDZVKZCq
v3tKlhIvoIviOsp1guBdVrFxpTY9+mmSF4pipNQdSco9DpnvpodKbm/kvgsLUBKJKb7is3Qv8P6R
AwhxKmK0d3EkTF89DyypLAEyD+4XUAS/hZDIVP7b4WK6p7YtUpS6QfgNbf3wt9PSVH/1tvLNk365
UXIOZkA6eQkCaVPgkdvhkDHw9K75L4LaTfhrjONkyn0ngdFj9UL6g4FY5RAhlIa+Y1ZacGowmMOg
MivPcrJ/FM4ubyepsGeb/fVKHzOjGGaYANztAFdYtp+3bULBL502hXtPpeyrUE2qnBhm6POhbS0O
3p4b2Gna9FmsYsFwNZxuWNiAdfHsBrC54vpwUyiLmoivBfnsQinG2jIhuMmuKL1hPNLNRyolUyZ3
7IhiaPNkZBGWC8+TfoHEq9wBo3lkHJgws4MQtHeY+WwS0MaRb7JFfapmQwCeeMOZbnFBps82yDX+
8H6C9X8CRNt5rMiAJyB9tzLQmXdvA8nJt8Dx6W3mtmJGPzM6WjHiF7ZTmargKwTvnFNguKVUNQ6T
m7ZE5LjdIugBs8grwdrkMHftXaJsKuOiawUJpAQmAoirUsG6cot3QXIcPqC1bnx73ykxyBPlx0f6
manmn3G5ZJ+MrTNsCU0X6Qh1eDM6NZsd7xuF9suQ/BXjIDDou8x/Au7322pLJH+5y3fYAyccmIwJ
HcYjKas6VyEBecIiVOCcRxUBLUwQl6UShZseaLtWyfNYhs43gVZ9noaHic1MdeqqHF0Fx7H0rdi4
Mh94qVjQv0Ur39FwgXB+mksFraSefQJNl0+/kqBPrKwK+xIytjNtVnsw/iEKAfyUyNAR4Q1D6fk3
E7rWZ8HZo8BhaJfYuMS8FHF6aZ+KyuxcdEjBE/RMY+CNiof1bQi4k7s1qvx5THS4KX9ygvOCkIUH
KTHwC96ZFoil4+XmHoQCqQzfqID8SdaQHUyw0QM0k3Apq3BBuHvqui5ztEcRhKd3T8oOyaf2Z4pc
GZ6JNcnpn5AeVTYP+UdSxFDc5qNGJ8OVsc86VdcgVtIzYf0FAkoKjG0ZJ07TFPAo26HizGVRXhUc
QrnbezZ4Qfp7P1Q+tYYzhnv1YLcS8EvKdhL/i/IOyoLVOdjiJ34mfMZBEo8A4e/LRFVdhnCeBPcD
SLac2YXBSQi1NqNCxDW/ElBTZad7+Bz+0a9Nxa5W6mZGrC10DUubab2U4/0YHp3iGwZgprQVp1wj
rM1J41xTJS+ljn0WT9+pDezrYvykfdKA59eFuyRkE4KWEu4dbanR59vb8Em7k208dN0NmmkZhlTh
E2ESFCiDrUormLQIvO/mQbbHeZoTc287ee2F5LWMmZGpJMHrfCaF5gnNVoRSpY6EFBc73bEzmftm
V2cmsCqq9MbdA95j9X4jrdS73dBWqz70mwUf0xEJfIyBKQV1CUxL2nhTVi2B0cvb0yfbTF5H+UKB
gGiN+QUXgXSpKGwWqInpVjVpGD01pNZLmj81YLtlSuJjiMAUFWscwg8YAZ/N/rmxTFkmpAnMqBv0
8qd9PBy8jdMB7rWZ1r1Up6Bj0EB47hP7LXbiZl23mKIM5DWUfCCuv7GM3EuMBD0hWhVBT9JI2O3Y
YVC+3Y+GbyQJuSf5tLYpBYHdfe+CgOmUcSczvH+K9Q4KZ3X1UDkgJI9c1drHEmDhOeUZJ18UmOD5
NYcpR8Ob8pa54fgnlhoiTSrny0EhPsLvW2C77j8S03CtHQ+QyHehAixg35I88IwORoEZIPHbPr/b
7AkSIr3KfrYrvtEDrnJXrM5q8FFmj2/qRwaKcuinsC6NcYucQofjawjojuv8dIaL9D3hqoX4QZvr
pLm15wEOGWWd2QWRjWxW642cQiYp33geID7EJS4QcJPwx5fAmYUuKqw3kAn2s9acmAzqOXnR8CzU
BkKYnrem24CRI2ko7irZYXaEJmdP3vOTi1YtIwU9fAlV7DswffGELiJtfZeele6ZKKVkXJa9YzRU
NejRv2gNf0L0/jvtICbtDbErB8jY03y30q//CA9Tgs1oAYk7ozDQ3nzjqOx1a8k+XMy43XqvVtmt
RbL+1EMjOl/qUuenhbGWjrvLu2jHeDeVx3Cw/lw5d5vs1KjOr7ICzCxxuVHg+DbhWg/ZLEAXkuIs
S0nA5wHedmUB3QSe/A0rsxJnqAol0EHaSA+EBLwsVU2IH/2ugdCpdAIb5x7Pbpck2ge4p46ek2qI
Fsu7wloAVubFNOo5omJkI3m91ZqfLU14PxRBgBcO/lAWK9ujoj9YtY3GF0YlaPfjM5I2uke1PRsa
qVl0cW00loB4gqCi8T1Tst1+Rafd5uP7TY8DhNNBJFIRPopEUlznsqu+66egkF578T0RfLxtQGpi
I9C8COjcBM9euLCfgEO50wwI7SsiE2hfEG5brX91s+ZkW3K6rl4e0HGpZgZUAd/4nSsdaN+78ED5
f3Mfelk0Y3QawMdM0jXt7G6nulzr8q0h7e9UpyN4FFneVfBq1VFiZ1vCJheBoA3wVWZypFFZRGIz
R3yixjgeQ2A/j2MpPjfzo79oGlUO7ghYtr+T+9ap6R6DIDMmA4WWq9e3uU7rFet0wiikYCl/JEoB
NWuykc/ETRzovaUokF+ErnHFKrlhJwfOm59KUHwsCjobecLDsU3zbnHhML+9TXU5BLqgwymPfF9W
bDnESl0C+RHMP0e02XaA6/vYumKZZtCYiPFFw7s+HCvlFpQ6OzRSU6TmbLi9mpo+OVlchiaZdJfk
V+FIwwLMMU78Aqoy7p3ibWdRidFpPm82vpL3zfDroV0zGgChZ8AWq9GqvukbuljBYuPc2r5q3d+N
31F6k/vefIABK3PUygpTix3hNp//6T3t0YPnnwD762xDWoOk7WegRSUci8FvXgLoT0w6lQP9CRJH
OQkrlBqTxZfwz7q9ROFFJFmlN7VoVMzmq63Hyb+apoSLznuPmDZDRiCWQ+QEQW7/hss4L51cRvKt
XwBDa7XAZRwGQH56d28m/NgfHc5DdNCHQHRQ0A8hq+ctAy3c5hQ0X28yD6SS1Ns5Xv417c2+wGIv
QrcICOMPv7E/8UwietT0TEWsot4c/qEDgX2W3eLOhM7Av269JM0yfVWqPxdbjqoh78LTrkX5NA3p
EqUjdFUXvayw4B50aUkSJsbolsQZOR/na9Mq4Z16NriLFxg7EZeWnwTiY9lUCZ1Lrny/DIW0lS7c
uXK7mt7ea/Lh8AF5oKNROX/kjuZQK/FFjOULg78KUM9QnrubzNxLVXeKJBW969/YnmWLvPslr/KW
hyx2tFvxAwF5gjWv4/Y3D0vRFfIkqTVwJISb1J/VXxQ3aFcTUavgkpBYmKMFov/C5R+1azGrbKjH
b1q73YisK5iHV845ppqjPLJC9G2THI6H9xG/zJMA/fYpe+RNNscnhgRORb7UtA/78vrN7sHUenel
YLbJAzueKcgnWZwDq7QSFSk3wj8UzSkE2WVviktu+fjUPN3go8SYiF/W9Z49Bd8dtvyXG+EzNLa5
Kl56DnwnjDT/NBQppdIRcBG/t1Wpy94DEEqY3T/V/mZ//8oh+i5OEncxiP7/pe5LWIEhdV8YAC3B
rzghr1g86shktl7YQYzOV9p4QB8ytBKjGyV9/imrqwZ38rd73Rfb0Xk38JJpphsAuVnoLZsWVCKi
r2FOjTgdLnieaiBgS8rcV8xZ9yzvvDKvR7gRNpY1VJuuGQAuVkI6ESLmIvTSljDWAcjTj3XKuGyq
P3wpE6O40w9eiV6VYpXnJG81yQ9tK8rZr65XlHGcMD5PwOEFpAqNnugxnZd5RzeV6thdcfSGmlGs
k6or4JGLKm8730y5H3yENXg4dCA59AZmvLTxl9SPtmTWAKWSYd+KiEsAHex7AI5ElmZlZtBJWSK4
HRjR8YZsej9oxUGao6SIatMvWnIm8EkJjE1LfrfzOx6Gryh7NVwByv6pRbUvNBYZwv9oO+pIAGAl
Ua2D6U36d8QuiEJiEqZyOtd723vLfrPqocXYcZOj6HEZnr3ntP6vuvu4Pd7LISee9YNVEgZiGHvL
BOAerFT2a5M72eSXXokdNzuht5bCKYP027TYCAIygySNzaOnOuqPwiesd7g3eaD2sWxJW+9+BS6M
OQ4VcdWSvfVOVtaaoLQ1H0gHk27ehz61yaFQdcbo5cHC09kBs7vk66YTU0hkJoOxHDYpmm6rnPzc
tRXXmjQWnXTSE9K03HglNWNlqK5KdN8cM6njAI7BA+VGlZb4ScpC387ikUuzUz86q4jiR7zp2J0F
eT1HfDL/tGCcgJpw3bF/J0VSkVgFQYQQl7FhQm5LlKyh+hynrRupY40Y1yVvevQfypOYJaTH0Pl/
iZRxAFDoJyLiN1Bqu21T+MpRLkQDw84bqsJWZRGLexkHpmERhRYAjCrqFPnjbn3SRSsjO37bD0pc
jAg21MllYPmnp3HqLLY9r6+RIQ3S+OpL66FhECssHIQT1KZjGYyQUbFS6N5tXEYHHNUVO5EiP80n
/S7l2n+PB3NPy/nSj3fWcUxo4cpkzgJcJRe0UcrPkZFgR49fBRdsgfr9z2whgkFLjbtxBssSuCsy
coOOuVwPbbrSmIOmtjNKxruPLSyZawn+4qDyLFvMDYl+cNYJ7/aVABGiHMeU8/J6RPrXVxw/Ed87
DhmSNFtz8uHNDSS8vn+XRE1FJF2m2zQg8Bw3qigA6xCJg4SJfaCQEfi/J0tWKAW3111Qk+FNUtdF
plI9Shpe23uv8CDHCqnCs5yiuexlECtAN916ka06dAzGSNvFOWETtpVcjws274tTI04MjcmYx+Fc
JBuCUFvKQ/Gd6h561ZAH2oU3aq10Jkuf/g2sizoajlYk947M5FY43cZlNTSRtHC5aIl+L09kAXtQ
2BCcBgNYw1gYpt6a9uVvYb1RkcYgYaLWnXsA0Pz8qUuSboJsk6Zo/XdNFZeAHAWsUsoB/WyvzSV9
Fo04cevKRyZMSSfiloXnA3ix0+j4wkpeOPnZLSnX8zNkNnGL0NZBS9CBFb9NI/MB72KJBCcEj4ty
v9nrL6U3xYMXAKB3jqPg4SJ+mVyZTp8dYfsEbZUlWW7KIBGULFyteXQyTFqa6nhCyQyWlOP5eKze
TlV/EUwCqqOwta/ZFR+PPc9BzT3cydHkuV/XGvYkq+2xrHIpMJbZWK77ORYOhUzFVgG1nj2jLSfX
g7iFMBHKU7ByBR6RbYB6MXUwxkCCljsNlLb4JvnwGyqJkAlg2Jpl2E/NSHgL4qbkqgk8+UIhqWAo
ZXnbnSNOWB/QOgWVoETqdlPO7/DKNKpjaeRzlMK9CkDwUcsytcd2gdF+3R/YGjREtaXbOtseVP0w
h8Ad0hq2Odwz5kOQad8KB+UT7P8NkM7OoBMDRnWq+tVix371YrhVjTRaC1z6j+P2OH4+ElWkqjA9
GAF5HmbuKt2DzSAxLzWrDZODY9t4gVh5FAcv5YvnGckK0hEiwqzqZCnfNK3eilsfwVxCSVzfQJBR
V0W5v78M4OmW9PttELO28wIqkFt+Z+EA040heKgG9h5ciyH9acAx2Gl6+khybrWMVBgDQ2YrNlbW
/tAZLKkdKdXysJQOvP8btm4TJEsywhsvDIIQzu6TVcwen1coKV+VijqL4/7Mi7TQU3nG590WWfai
WJlurrqWkazkLeq9k/9Bld4AlVtfQtZaPHYETpIIJFeUY443NB99fU9rYYbaBNz5aEohv71nJkal
mSgpsnWnJbIRBJRK2WHqFcXc8H0nIIeb1y9b0JwDGyh45UIoQuxS3tYfWxXSs0EOi/QAcOvZejLg
94w8INU2sJTEkH5BNmI21VzjkZymAwkPD6n9GlXbCyD5BR6erUtN9rvaLSwBrEqxyy2H1Wn/nmsV
4vqSJsBd2gk8kfXOyFYT1at5/vOfZ/P+HAOW6l1Wiln1Czooubg52wdoEi6YTW7CnARvrB+hXf5p
/vchQnU72Y5aicYrOAHZeY0LnQ+DxhH7UD1DHbNMwNopkeo0Iqh7EC+PZmWQU3dbw7ATpItJM1dW
vdZhTy8LTzYxH+duoJeBMa+EVGS64yF9ISTk2wdpEM7xUXHw001TeiZGZwygfZFH/tanKID16Nuf
JlHVpdj4r8A1JHsUdZ2FJMz3puMuq9T/oPn02ohD4ULSiXqnbNoqO6KhupOhDPtF257AFSdoMncZ
FyI/8RpPqm9XKXyZChKzQH+heMbjAN4md4HFF/GWCcC0nn6cq/B658lrn1uvBH0Yw2E1M78cwahU
pJeQmCbMAl18o6zgP86WF89d64JmfhVz87OLPeSNPFRi9cTmDE3NmOAV3DQWpgExzU8gM6ts5UIm
6H/07iUqtYXaCPZNiM8Wvn3YxNnK1SII5nmC7FV1jLggBXFM95XiBYmCDV5MLe9EL6e0yiLri9//
sw6fR+FbL2Yr8ZCQ4y+ybFXyLWosiAyTQu4Kx/aXhCV71nOx8kN9+ekxyrbkoLV4W81Y8HBPJd65
A6O5DcPJiLqGIxQq8fVZga6pYD1zAdci5xn2NLWEshRJR/25Zuc6eenD43aAmzXro3JSjewYUvz4
c9nQeQ0e2VBcryN4jOKWN0n2CTF1dmb7kcya4/0LIQIosDQ0ZfI30DGGbY/fD1kySaPjtHCytNkx
mr3XwIvu0KIhjpVSv76aJfRqJuqNRf+dSQGhttpRRi0BVYYzU6AnXhiQDZYegDfJUQFOnEXBe5BC
pYvcnAl5oZG3whsm3DkJZy6HhU0V9/5M0XnfHncF9QKvkuPOTiKZZOyaKCdtsM2fUcbNlYlF5Jzq
gKHyvnLdvdlQfIou4Cy0MEEewlyeP0Nfoyby3LJhpwWvP7dsvsSlcMdnJBU4r7TjLKCy8hJQOdkW
EwYhqXwbIK5Nk6ZoQtOnuzfvYPyf2ArJjl/tSH3O7sJ9FIDK8Fs8+/wYUhf+nYZ0+C5DK2Qz5zlb
L6VOy2RadKMTGEnXG2XA7/Z0fxkeIpu2jhRTB84CRSgU7Qauu0pWeGqT8TSwXwZH5BSJxMMLQ8Or
Le0Chw0zdyzvqdNE5jh7xqG9hDXyisCfTByqF1IErPuQZpZ8IIOHUmffJSAhBS1IjkSku+o5Rr+7
0qsjxiw7m3CPk0p56PhpvAf5I9ZsFT068Gbl6H03PwoVb+hpfvIt8leX4Mx6fwHrh0/ZSxO1jFah
GiQTPj0Rzq1GEcEPbeQEkaO7CBYHpYa6uTW6rWvZQGI1LAW6pO9Oo9L6cNHOYiSHoVbanWpUI2K5
WKZgHe3E9/k8lUENgh6CDImmt3P6OhZ2+jYHtSJfWXw49mSFFxjGJ98YUKl4fk9h18LT+G3rXeoJ
Q0CadQ3i0i+g8olUQ/dqt+b9M8wEIK4ujWCk6SGjoJoQEacpW4CjXslLTq1vtldDSWtYxRra5Bu8
eUu9AoAB6CDGb5aRle9I94k1Hsavf3+0tcsxGTxlLiq9lK+Qqi6eppA9ZQtXlecu8Xk0icYiL2Iz
1x/ZV6JXy7JDjd1PhdRan4HJX4J3Ej+TWW8+nI1gYF3rVOm24+Q6pnRkI2OfJUObsEbnci01VB8G
w/3PtEr371Oa//9mYMwLgqw2MomnoOQjssCuSCnS7YH5T/yNRvNfDjc8t1vjk/3+xHnDbS8y3c7A
9FiVgtz3Hnq3Ll+Wo2LjvZNd/dRFwGsR4nwUOSG2WctDHdRvkFovJOMJDGL744Q7NkSoU3nUKk74
nQLFvS7KKB3fSd+Dr/KwI7rJk1/e4v8pXX92UnvFFhkOYnodrtXnnJyartU12Ve23aTTc/a1IhiV
ZClqvWi3qFiX4vtM71GGQU8yAB7PFpjunChmGiXJO6S6WpFeXcCkKC+ytdOuruXZ75aHKOf0i604
JTiIk5hfeffSM3yDNyPI82gkTiB1clyMD9ngfzKZHgBWM3phBXIBYWisJ9oAad5wwxUam4ZMIx7k
7cdghuYC1dO1sGXzJRTs+3byjivCUcUQtuQmpDRKVQcyVWwGD5rszRBfrHYJiS2mFwW0J+AGNhxz
0OJARVqHxlDZG9MXxpKCojPi/LdeLmZYPwlRgkKRtq8XxjkySqBvKw8oOt1cvaOnxWhN6fthRYed
8DcqcW2gq34VOg3jNhZ4FUOeXDrXfnHQfkiBC2Vme0yiaOP7rftXTNm6qHidk73lQG72cv/b1ucf
b96k/nxiFggzywRxUxAixn7f/1KeNexEMjmMiLPAOaAUVBtS/q3yzDjuRKQDFDW5ezZpfba2dsJl
btvviWVu+y5Ieox9Hhe34VmQftEpQZiwooHy3mm1ZEwp911vDeWwD4SaKFslV6HFvhT9zjztFQn9
iA5/uTDPDMhvlYFH5U9TsFxOkAU2YsN9j2LbLJu9n8yJw0dBn+sP6N55YzmiMJd6Fk+cPKnrdmJ6
uF3RpkZQ5Jqd1tAniPWDMtKcPTTO7cPRbg04nF0D5SjZa9ABkNQoVyUxRrsjAsAJt7Qt6QPVxFqF
7CUfsRiB4GEFIbsjj4/9M2rPE3f0YG96QIz9Et/OgOnXmsSgwEk64mV0Jpk0d4+9iuh9AfQ4biSf
qn6hTh/8AXiCj/VXLEbcBcHfvw9lYTrCjg6iBHkLs95HIgdZEVd58gOovCaqrCpOWTm93/2owdEQ
/W79UwZHD93C4dGh59xlRcfMhfLbl6J0CvD4TpozYb0uqwhsPiOLv9f8P4mxUtQTx04YKPvogjd4
Z1kSJNE2sqMFKYsuWXR0FotmNRNumreSukIbxkZOLLjzT65GixtI2tAHueK8ZqfDdBE85c77TErO
A34i3zRJQEm7L3F18OgixD0gWlXHz9++XudXGISw/mYQUL84xhbOj21vDpP+XrLzqYOogIX007in
vYvaPQILGs29MWRuevoHgODjea+ToBm3MzVKAyJjS3VQsWe/ayTgucOiumGqv3t9iXLdG0O+D6Ez
mQHP1TednBqgDZ/kRcj6JQMeppbkSW742TD2YTLVxyN4DjrxkOnCHAUJOrfAVeyNdYFv5tU4zxrZ
oRLS28ro7lbGSwmrz6QAjEIjIg1qUhs/OMq9jvxOK3eo2sUDZ+krAwwe9u6bI/Eoz9W9Ecin+b12
2E1ULVQqZ/ilFGfxcP7hoPOmlwxO/5IDw/9sfl8Yr3rmsh4IW/JLZyvLfUBxPNxPLKbq8eChXsgd
qVwu6YdAsIMQq/EwMDJkGslwqQ3Ewj7CUl8Lqz2SurHFs44Kc8DOGxbcFWhgnpXLOHM7JwFJbQkD
uhWf+lj+QXJKtVwWXIPbhBlI/Z/9ikIjn4xRL6Ohw5p0C0f1FdtbezZZ8oL3uslhAC1b2NW2lEL1
eNEisVsvVk31cOgfszBH/Zh0Lgpt2IQkkwQ2A+IdwrFleVoL4nbkJQhCNG4bYIvqsN8VqIUSE2gq
i3pkE6Hz9qqRVlA1o357sE5BMApp3s2nagok1H0wMZCeA8iiawfqNjNcyXbUhdlmPX4ZwnIeYeIH
hkJ5r5j1IscDu61fSI56h0KQr3UpckG9XRMh1JGB/yzoHcHAoJZF5XQuX4GrGmUOYM4kVgkZQbWK
E9M8qxwnkGRlXeUFSZaTr5o3/mbX72RKsFTV/VQ0CIsExQJ92eiy+XrFCllvxLuZl9iJfb9vG7va
4u0HbzfJccSckhEf/qUsj/mWLya5zJtfv9RYngjYkFOADlshK542YhjOC5CO0+fInxrQ4rm6t2VL
/W0/uBgOpRn8KxiMzyaa0u8gijFo6sbWhPNlphBxr39NEP3nzPDguD2HfxoafnDSB/9fcGICH1vo
zja5VdJGdavnE1NvECskNqENEPu33XexGtgTLLs3Z/9DVLIKq/OONzEqDNZ36BtQaRE2iZ5tc0Co
BrpDWUc2uTD8gssAVJE57kxQP91RMWUBbeIjRdzN21arLXsregq8jlGV2FcFDfIwMWabAPd8fyL7
26Mr6MtmyYPCZw9KQEnFgjyuqbkewnLG2NsD6t+TnkCdFwDdfjUQWs+5eT3pO2h1ZSCGS3SdKXiC
mWl4qmmMMpnubolZ1wJUsvSUcz5FxwNTxhJVRQf5OsSRMlz0/ZquYzBndP2zEpKlRWHmMwxt5CMs
GKSogj5NEcuW89X56O3Lh3JMrnHhYpPtOwbiene+kOuCANtkmqGZasyesRgtVQ1O0SLa2G3gSrmV
DUE0de+Xz9MYk2g8wn/jg4fA5NjE2/mvot2ZZpgkL+7l+SVA2hVCgrYar/fMHWLldAkAe2eZHIZC
Q61j41I9uZM2lnGw563s+Wdx2o/isY2vbxwwyFDDId6YAdTxWtVtQmAXJf+yLITWM4bfgfOwW15h
Zl4BUAdVsJNDdmCYo0/a9csDlGg8VWuDCFrwruq+VzUc8Dy4eYtD5rwo9hQ67HK7ZlYe4upQwq8w
NYNkGVfnKbF7/mNVGeyBLwTsKro+jcnXOYLGGzr5PE/iKtwvnga1Dcno0o5vG1eUUpce2/bw/4Pg
WO6ljgRgTzE4S8QGzPwIUeevm94C8om69V+WP20F71/IjDjWkDMm2jz9vIXQMfETjrFZ9KU3ooIz
eM4dfbpJ4DL58ova4zogmiP4a1nq9GjuF7+dDufxQ/0G042nRgy7tv8gjxKhDkBr1+HSfqIpvdJf
gxLIfkzM6I2mm/DI2Sa5uUzpcBN+Ej6d1MB7V0e99jbNTee6BkbPl9+5mFo/rZx5pzvcQXw/CuBi
/BBAbybSBDQ5nBIfNHuQrhOxvskuiZVWzVxm7+Sd2Jbe5w6Y037EH5mbgmsLfN16Ta3kOOmM3mth
7HAdlBR+QWcGl5gdzW2VNu+J637DHXd+Krdel72Xa2BRF4tBFqLQ4nnmIR2XBDxupp3aioT1M+p+
IUc56MLNHmuMdxFY4n6v0VrBA79A7MZhWXAXzhSSXPAx1akKCd49jA6R42YpToxSNKtOmq9kPHfq
tpq2evFJaTziqJ6IlGDs9fe3yYD8vTlU6B8CO2Ge8AvIpiPcrSA2mhmLeThsXGyu30XXUieXEbo+
t6/72sjH4fEeuJjCAv2V9Av8Z8bMwvhwHJKU9VGskMhALB/Fj92wStDAXPEBzvh6UrFyDJHC/00a
vkSyXcZRbCPpDUxcZ2T6DIQIv5+lDy0LK7AR15eBa/S28t0pfroSnD3aqe+leYRWMzYELgJbasU4
SRai75H8kFT0Z3RuAvfu5YgerHz+APeqWZBkOSFwwUhw64GqY9Y9YP7ZRylPc+hDhnBu9HJQsXhK
pBGnC9PBWO3moIfDw+FkLvUlO7DV16kp+I3s+SoyZ7WphEIynmdrFlGfAxAPbbSUwNfRWas4EsZI
WmJd+3HzTbbabYGt1KfBqBEdtSFZPTmfBKAhaeB2DrJ6PmgqI8eP01+u/cYv7Ho/We6SsKSHuM89
FG6nGA0zCaXVAzHpr9nYVU6YjFAIDBKAaN0dsdsSRbnX2gboj/EkaSgT3vRSkt4vidGwt2evjxSG
r30A2kDAh8skB9Ky5mjtu8y7HsGT4mSQ/lvG57oH8XZIWOOnUcOFHPlTZt1gxqZK7wEzhqbQgpgt
WXpkSaXotQH9+XOXOsKjZH2sc9ouM1L1prubX69tFVvKpDcX280hDEWx+HzUc7rlqLgLO00EpdGj
fUoKnbFexnFu1Ogti8a3zO0Su1ouP7dg9cIit/gwwYrXQtD3pXL7QQJPian1UGXyj20M0l4/XhpJ
g32PZmHut9S72/hD7cNZtGvx9j/+z7/x3QO6SaHdCQFXKoBslMeiSTccbfn7ObMJ3E9tltErZjwA
CE+APb+MkcA5aq9+5oFqfhnjAPJqx38p0LUAnqGWCgJ+dlICTwVpvg7fvd1Czm4Xa2NQNmOgPrPg
TO6Ryhci35UqymQHgoBGUEpY6pwtZakI1lhJC3Y9hgeMgfqAFkhGusTpRtNzkvz81HBIXHx1qdzq
9mYlXsLom+JAafV14jBNTdOe2AQELc+vmeZ7tP/SqyA6H4WmKf0Wh4CVim2qEUxBLHnYXQVffr29
asIsHGG7z6y4dMKJZ/3f30BH7v/n7nXRGaw8ZAqHBbB8sDPNaS5CmHb2qzqHlZG/0qTdwNulmWJi
cho1+hD47BuyX2XpfZXvdu9PKQakmmfrBqoDaObACzKQFz8v5gr0AujRwvWDHvwoZsSmJ1xEHcz4
6qesp8F4sN/gnZHyqLGqfsnTkCtgRtrtUaEIqSUSrbMiXK2w6iMunHZXRJpQcpRdTxrbSAuzfrAd
IswagSfrOKZvm73T2DYBTga/KgzulqS2uXPYJjjkMyY/8VEelVaVRs60nhSkiLMYr2pqwZaQNO5b
B0Efq/cYSZEQxuNpU/1S8IoY+UXyW3E5AsYsv3/gyQdW9ejchtfIWbcacTVFWVVk4r1bGdkOt8UV
q8tv1YwA2DAV/ptOlluiUfOK9m3hImqlf/ZkSNXJasGkNMMkSwG9w2aUul5rYDXamMpFw2O0uG4l
EcSmllo6Me1Wxke8TxtAUbUxcm+Ivwt6vfTrBnK0upGlzjT0kUiUPB6ktwMUyHhNgw7NasmPZkol
QE57LV+4kwqzCtdpz3dB3/wJYnf67J0gM0B8mSH5bPoVxXrTm8Tq9kyiW7vItnOwSGh/+w1TFVP2
hnCs+2zYi3ak/Er6Rz8Nts53mYXtmpPRISgQCiuR5Q/TG4Rxa7acYcT5DooiZz44lF9JaWQJ7MM7
fq33pfdNRdUC58v1V8FCl7X4Z6NRPtQLKbp9C0bQ376i9xqvFkqxrhQjSdRplqj2bnN1vSgz9Lhq
xGfN3QGnNzJV2GgVEEdEyCmdZnaCLx6h4IuY5q2piYNnJmQBHTk3Tr8JNRFFbdFzazTKQ+v+pyvN
a+HwwAiQYvyFm63KDuXqkFo03sIrl/XqjL+PMbdD5yVjJ8G8RelRrprLoIJEjAMh0xfeQxE1BkBE
vBZfFLn5Yq5yfX+15aqqh7lOOmA7hyazlmckz888Lob5DIYc7MQoZ+KAHLZxjAKu9+DUuUKDrlEq
jLLA7Ow0Uk4sj3eKBVE2N/V7TQmrvzkfR24Xhgp2BAZaIxLOQ+x2JdHQ3WC1sIbLHBKR2hySmB+H
cmTobe5kSj7moQr0mPyVOwVcijwxFw7/kl6QfsLjQcdlmZZ5MbG3FeHEBHnJ1yWP/s1AeehdSDM0
gnW46KsD8UOPgj9AzSFr7OJBpCZsTyHfgCjFLK4utHdZJnU4GFdfR2Axn49zvZvVlQ39q6jmnbSJ
4mx0fRHGmZkQ4SI4eENfQ6YOhaMR6Wl7tAB4V5zZUzfSGEOqp3+2TmP+ujEdMmNTm+nTybfVLojD
6z42sq7/mm+5qP8ZKm3+qUHJZtLTOLjuxJE9/jGUHA9DVa8euuz45pjCYCD8k1uZTNUEf2TcUeOt
AohoVtbVSocqNqWOzVSM5/Y5LDq9f0z1rIeUQ9LYEc8QMBPYMjLsI8AdTSy8/W2EcMHpx9gYPrhu
E8ZncN6xnd4E0Rvso2TljZsd9cKHdMIdqtVhXBzE+E72fcDn3KFkh36KsQpDB2eHyow0teSdnepy
82SmGFWpUnzh4g/LbROklnCTu4vmhWGKneXqSIVvIkLHURavAyM8N5D4E6kF/IXmUg3fhYtl4u/w
IADsAL4CBgQqoGhpAEXZcynDaGJ4HXY4QyhI1l8Qcd14o0KrshqY7HYdfSDeBKkr5K3P/s+x8uoC
CU+CftkML1DfShVw6P2fIs3Dj554d5cMJ11Vm8OESkcFQE6TcFGN5vU0wBzXIzof0SrkDrYsmlAi
I7roh2XCfFHedVlZhZ+xqnH7rvWxs19556gDbSVOc+FFYPNTJcQsjhAYLCzJ7V2/yLez+mAOza4k
j2E5Sl5JXtRGVHrTYsufamyRFVO4+NFdkSseIMx2B0dzo8GdKyuOoL1M/kXMuK8B7a1P/tpqvIPm
w3sus8+oyv+sHT3xLsWObfYSw2YUnyrFefrUJivy4vReduj4ZreRYPSKo3rcTZioEXQ9HXlRrq7o
VpM8usBLBpH97+Hv1OgRXpg7psZfQ/0+85v5nrXA0upKKNlz4AkcTox/0kXp94OkQOBCch0HH3Ik
Kdf4ji5h2ZfgiWJVEbyxbhyoa2kD+66Vf8JaVn3nUkOeJt/yd5JUTrhiPTD0UtpyXxe1d2W5X3Bc
pcTt/XU25m6vOmiQ4VcTFtVQJj2jKrxzxDHzTJoEwENUL3uRgPG7CzD7Y8V/EU6dekuNn7ql+nky
g1lKrQEMRFPaRP/EfB6f3kiAA0GFAdHZnkPdACRWP/F01s1PFqcchNG3Q2GpNbyrBpiWGRzFAf+1
LtsIfgzD4vGIltGCDMHdoeYg/2Iy/uTazH/JuTyOQDVKDolnPlSujHqQ4qkYBrCWHAXPGCu80j4b
6xbYwIjWzQBoESL+eG0tQFZtamPTz8aogid95h/67a9kdhoWSBbAfjiNErAqvJoVQSBrBDIhlX87
VSm73K/dli+JBRjNXc36y2PVnaI8GPdfDn4BMGHgwFf6KvHxtaXDO+PG41FxLlcrGKTDaLIx5sPY
0y3DQgq0qe/j+XFBI0VI4hgf7e6+0Ib8T/DQ//CTWsk/SK1uEXZzHWJiFjFFwRqzSGB1W21K9hy7
r5T362c+88YO0G2ZP0g9EJGbxoxfsrvlNNsZF9D7BaZbIIIzq0Xx+WLu9thZAUB5KBP7vkwPecga
amRrwOExhnMheDTwO95Go+Jt3hwMPFBPr5o2Bp4F3yJvjj5ch9KSPtdMy8E4xYZ7SlXgJUgmVm1p
aVJ62PuSpMayCTC+xwCW7h0QVdB6svFdkB2D7IGDaiP17Ue9ifvyAu4U5xhxGHkNqJNNkuO2hTJa
IbkhHgos0OOMntgTxV4FwXHaEHc46sQ7LBEo6HKdF0akX2NwQRrIxa2B/6+7bfd/jJg6iVkwH8Uj
dDTH1aAyyGalLEshWXdElDbpuFW/odlee7yjXXJSYe8FBjsTSFArZ7vdmxRhOlTIU4MyfPQKLnrL
m5jbbH0ceX3OmhoyXbzGbID3RzpkfO0hUkFfuWMQ22NiEGITYUD7hbt30nng6nc/DEatxccAP1K9
YksrMeh4X+HfICNHs8C9xpzdJDhovUIU+y/61958V6ruervOU4Yhev4A0PluiJreqK1q52KYcw6U
O6AfMRHYct/eBSx3gF5NZ8LUNbo7Ypz0YphGTpNSmYOpZOXh6PKl8m9QF4Hx2CXbUwoWnvMvaJCe
Ck3pnxYJFbgliJ0ymf8FOLMvI6ngQ1Ci0HRsMXFx8g1bnz32sKfPDmlsLp4wBrK3i7uthjwkczoV
PaITxg1DxLgqwyjBuB1306hLaNzXCzi+T8Amhf4TtEpVE2+RS9CD1SrrHaKXvqAyiBU7GPf4GOg1
oKBzljz9o2JQ5J0UeEzi3XKBS4FvGW0HKpdA13mu19UcD6OWYZiH1EwJ7trs8Xmgs2zlShQogX/y
Z7BqE5kO/H1rhzKsVvEvnNPS79vDrFyMKDkBc0Hc1h7lv+R3zH1w6xLHkSdi+mt4nTjJHtQT4fHl
6PpoKqlEUJnoAeoJFWrAhWAtf7mmdLB0wgczTxAQXxJJa1T6wHVk8/tJlqwABAZY4AwKTe6rgaC9
/Yrqzbijtae3VQoFhoUOas67kcBfm4JHL2Q3kBt2e58uwILy9D+zOX5aC6pvdI++JQxdLz/r8LjW
se25hW22M5yH5/fhFS55WBFtw63J3BZWPEVn51PXzNHVhc+dM4oD3dq3DKofQZRfXUW3whsQEAs7
DZbaPEIY0xLHooggJbKu9vg3XuhzSEW6W5pxfmahGDjAgezFXBFPSc5MDCcV8Rmk/DJCy3R2a1t2
SN3ed7N6agRGwfss1PucYPoVDBv/sWZY0fUF89Bb9sU6GrSmVeDDWj8YhSr61chrW+kmceBOd/C/
ZYkh61kdzjpDUepNl68rMGXHcj4x1ynRxCJ1HOMm8w1Cee7u+ns1fVVfrrRkfY3UWm7L5ewQpgwA
nHWIaaDV5MdN/bn3ECP/cEJm+UjPmfmxdISJCxeKuh16cYl8g9/4PQsVi9zRr+vlFA9Wcg4dB7Km
2c9t/M/9G9kHkEpyyUy0hSdTQxU9ypu2XKIUs/pYXRlu1DF1PFeWmLeC4fN5dOvG4p4euvw+WGkc
IM0WVKOuJHKhkbQpiWy6Jskr8ibI0cUTJElYpujqQywfai6+8GerPUgiSNRCqac1O6+Zwp/lSGUx
f7BMFtSDKZqLu9XkOU/32w3rX31gYGcO2fkF/0JfVRbdTKRMG2Pynst82N3V6mSyTcxNMzba9f3A
hA/9xhMyoVtHtdnS/enWO2WOZoCbRI1UAVdsSrmsHlepo5M5tV5ZKZKtBYeSNWRTV7gByupfPd5O
3YviGe/xS5keTm5Es2VRrgx3fe94fgv8Y0gS5d2uZwEIDGfaCYY/smhpw7kf7OHgpVjOVoBXiSho
mH8Fo1U5796UMKMK80UoZ2M1P3AzWEneusIGCWOSOsNnpRQ0+tS6majGiKmepScTB6V2PijygSYG
2j3NfHHH6vpoUDofn4hFE7AEXoyHIYJ4QrVDYlHuUDgMcoWW13xt2xhRBgOCsMjbnnd6Epi8lrHE
fHW7s9BMx91fYKOD1aM1QWjTe7O8RDwY6I8zaj2F0lmcRf1n3PvTQeFvPdYr+r3mRhKiVOU5/be7
2WZX/1sTzjr37YJA33R1xvjObXVSaUtRjYZvk+AIs8+6YGUdGah1lw1uecnOJyF5Mz5Lskjfw93D
VpwnbpXuXAipKTY8zHMNMUJfdvp12wkQNZq69yogxb5Xy+ULR+8GPLszKIOcJnbUkCjN4pkEHM5B
vQeUhAmfYQ2r9uKel9XfZcqUSkpG9n9VD4FMadMHDJ46IYUQYimzSssgnzz0bDUf9cFb8B/csRHt
0+HMXaVAW+nfJEjkKd1Cd0P75nu2K3rCgfeoW+6pTTRtJZZUlxsCXxbjKNROKCEtLXM8JeGTSEkW
bOJLDNQ2fz9H/gMi1+44JhRSAIIWY/xYCUp+K/7w8BP8onvBzZI3FddlGfcdO0LSQBGnsE5m1hFE
eG5rYIXLW2FsMpzbYfMq6Tys3E6XhOlcKQ6gHvxUdJeGtjti+Mp7wT2aTr1bF5M4AlSRXl/Ouf6j
ZhYOQjFikQb51NNzEpk4UUucAtgnPW5cmhvDX1i2ArKFbNMmEnwHL/PII/b5ncO/SVORY1hhxt8j
x0kGeNDrc7aNf9jvoqf521lgaw5KKubjcX5JeeOK3mNAdUSZYYphgHcuojVYEHqQS5dzpDwJ+eCu
RkKJzt7O6r8EOkdXqDGCA9tPGZUsYqGYNMp/ipgVcjLORqu02dFGyByU7lfvlUVPS8CIYrwI+3y/
NQiqBFfmi6ECE1HZMPUI60cnqY+Sv9XHdL1EGi++R1H6BQAQ+cwAhV0CfhcL0IkvVp+jRev82pkH
55jGfyU8XN3VgRySK0Suxm/k/JVj6N3uBF2kFdZTQFAN/33lMJOGBh+5codwJfPxvCN2nKZyrss2
+x3RP5cjSDKUP84bHbvAbY8n0PP5uFINZcGaOurXw18NMUOLuxCIwTEP7VQR8Yf4dmBRUf+Qh1MA
IhT1VezYWHJs7IaqcBtpLKXyzKsnD5RubRJ77GhG2aCHaz+y4OdwLUmlMZDjTMcPdJ3+oVLsC//4
Omvmvc21j0DIpUWLeRVvZJvF19g+XFFKAeb/MHBAjMjXeyxuR/oyrv9J+h06lVuCGM469jVVs59H
l6fF0eXF5mTzJ6H5G6EHBO9bsQvnaj1NhV8Bu0L6aPeOecNw8xbE5sqZGLkYqDE5WXD9JGGVCoSE
Iphf/gDafnawIjIJNUpjAIdNvuABUOiTLuYoN0PTqU/IbJ+jjqrsv8ymPFkQAlFc6d5fnEEgZVgG
2xKCWPPQcsv56SowUzTEP8QBGqefXReb6Xp+DY2lNB1ru2sb23J2AOd8Azl2oap70b14ZAYYVR6q
AgOjhEw7yMEdFRSKTqLe04sfPWuwA2OEIuyKqxP3cO28Fjmbl+rSTZRTiZurePsApQDgBGsc8QYx
5qCJVKZpx6GdxYEZIaGqXxDpbpVPJnCR6NdyzR6yDFdp8FiF9qnXg/rnn2nCrKylMTD/9d9iJE8P
4wFejMOZ66zTJCRvyhiC9VfiikvEos1IreF7YFXZwda3zA/Aka+SAoBgq8ui3WVitfmaw4FuONfg
oJq1PMbAnP+IAHtEocK3nFzQDdBbqigW1NfuWBZHtFKvvcCIrQzqQcD2Ndh3+IMw7z0Ml/vpdgxF
IMJiT4K3sD5P+UD2bFZ3EwzK5j6Jwp66z27KYzZnKjUgIpPTTK80e1By3Cah6yB8qNpZWliGSS8o
6Gw7AELa3xy5mWgNfe5sVkBFc/bo1Xyl8y9Vq9hhAxXp9IFIfb2sn7di1VP/QvnQdmfOtAlGCpzD
kbz8pPM/lUdi3o52UPJBmwwDaWFTEXGc5TpBCXqVTOxv26/zFoZCGa8DBZ0agQ9pobWqAt2pcXh+
21JI8NbFwYVGTfQcTAFe53YPsANZcrZhdltMSYTyOQYrS8+P8ZzjSxcoEQ7gXAB9Nl2MQr5MBuE4
6WiZDD8JI8Rw4fIXa8eBZVTm/o3nlC8J3rUvLsRpDJi5ZtLZHZxjt60/nxEWH+dgGa07ULfTj5ew
sGenLawe2jUfQMtajdKSxjdYZpwsqUO8aKelttzMyBIkDa27xm7nKOwCXs1dkN9W9HdKQOTN64ft
hkDzsEwhyDIqkPEY2MljNm0gShlq/Gdp2rTz96niRk2KUSYvAvqE+uJniGL7porC6s5ilDFjtIoy
tPhrfxZ5uQn+MwYN1gnbAD1Wy0yZNtNp2Fyarm3nH6bNIuVybXPIwdFOuBWhQFQY9UTY3h0NCuMh
y8SaAAfgOLkNJ7skiQq7vt1bkEEAs003Ylb3OIoR6FYvseRO8NMW/JVKbvZKK5EJhs23L9Nkit3I
9jKPpWzq1scqNKBnxhd06Vs73KMnu4vBsnlvF9KWZnwjBEH+ZXT2VMojPyr3zd4zztI2hI/15CKP
zoZ5IFbfbQaed0fe+YIiZehtwkqrpI+ttSrQyYcQr+dCM4OI/LerWHobGZNNNi3bIR5e/ungY8q3
R0twDKGvrKxDDYCcN9vIua3ByPS8/EPq/eUzI7K3DhTJgtWDo7hW10Jcy+AoLrkeplFJFnd85HVD
8b+8EcPLod+VYZik0gHFYjvO/RM6Fx98/kJBT9treokfAiebuvQPKyU9PkskIo6uwg4LcGA06I8p
p62ueyPFcJH7P7FEZVZey5Rl76EXIdivIVbwxaRc7pFRn0XWie3hnADj+gHWFIdDxxOH9u9dNwki
gmau9RliC19/Pdm1kUGpgE96VE4RzBuMAr+b9wleifYe1LumNvUvtCZLONDIiTU8eb5hY6aeADUs
n6QQJ51hzJPCXfPJYYB3lrvPU5R2ST7HycvWanrij+VNhXT5AZuNoFORJ1UchcVMtFUnGUdccsDt
9KevbPKPyWl/KWG5vlZjktXrxtSp0O/ZFPK9q870wYfqNFYThNNWftUcs8rjeIQNVjxLqcdXsb/v
CurT16VtgEqpD9HkL0euoPIm19sfX6pC7xpbiY45v0IVLxJ0Qey6Lf1Ko1VDqyyMfT6IkzQw0wHW
g3CuZ2WBkFJVFdqdWZb6UMYW+0p2rN4SVdRlCPp3/1z7DE7H4wSanKXVlWDQU52jaRgDxaG2f1Fb
wP0WuuxTg3oCWukqSZUxxvE+oCDcHpOULq1mHpKQAvioq0Rh3jqgS8T0ggvZ97f/yNQjNgarMTXk
puiBt13wF+Twc0zaIyOxkCDL70qPgebDtFa69/L/THV2C64BsVpAKuz8uW1Vot6XvKyPekowZoNh
C/vyWQO+m8hFT4lY0j5g6P83CPLhPZ+QNmADJ4Ey27mB82vIZPs/oQTVQMmZc4wZQHeBkHghLFwo
o5zznWIvAqvQWBRwaF2IjKYYg3TWcwNV04AJHUg0tXUOdyBj8EqP1aXEcHfFRrwvR5KgNZ7PbhEN
v5GhJZhZgOtOoFXGrXgD2WGvuGROIum6nMiENYdvNYWS1ojQ6Z7c6A0akZrmUSZILnZN1yJPmi8d
WKEl+cGQuUjocto+DSVMyVV0zIz4LYGu02wQdr0M3fBRf1c8JuY5nKIQKy45aBk1vHlvfQO5GTnz
Zvq2XUqrrooCbCNhm2KyG1nXFBDDyD+zOw3N/t5nPeaJ3lvwd8f0xN4tXnJvEFaEKWW7XA95wAu/
3cyZw1+koVAcvLOPmMtnC+b1U+02iTsrOVM0WF9QbserZrsuGoFN25CiFurn9sUWPtOLVpFg7vAS
MTWMs+pjoYUEkq9OXY8giMpA8feipVqU9TSBFv4N6SpxZ7WxFbXl1wmic3CKFbLH3Ug6yc8TOfIl
/6hvQX5pRZ/nt+g32+fW5EN6/7zkcrEbY5qUmuVOqftJVZ89QJXLbdNMrPXjqUx0z6te5CGygZ2y
y7rVW2uMNucAcAbR1dx/ZJlE6pnkIfB0zq8vdY90o7oEdB16jPiS1LSwk/4yv0F/paEvyyEIv1hk
XmHsKQUoDrwCI55/+0xCanv1VdjsH02sqavEuqtdyuS0sRTmDyo87Ss8jZnQNPysv/er6ONlynAy
Aa/5LeLmk/yfG+RwOyX9NRz+cTB+MCA7AQiNcntkXUGN9SEHgdnOY0tK5SbLIkoS0z1Vq19iOpSC
VWqRV+VlLbIkcBodxGwUx6SrvzWImTpiYRBfTlBBmxiKcxeLLOcLOo7AsNENsv9E/HNou3RSMGxA
mIgVn9cHS+6AzRZA2hZK9PeCGTev/+vZgVmVfXkm1LOw1ulFw0IJ8RHWo6clScCsNqDFAXclKAgM
KGjI3HmQR7PkTzU4gdB2hDUIjk0ndCDj91nZEUcUxhFAm98KRKdFr6Ag6Mk/mM+472Ud6LwWz2J6
j01LZdatsh777UqGj5xIJg4DjOlJChjb/BBnTf3boyxvGzjuZ8+XftETk4c7axJbktUSPoaTE2Pk
8dt4AIUM98Eek7fgWq7Xlhc+6pScMwpS5HEtRWJXtlaI5/hA+r/Jr7XUtugu5p06CDVb665YusED
YDAg27Y2mfZ/TABVSqCl7zHUmnI7LoNKtADiBtzsFPqLJ3iVhs4jgObRbVdPLfVtfvRB9w5K0ZR1
0N/B0a2r94Tm1UpLBOoNlXrLIH1egz6xnwz74NTupcgERRCIfrq0EF7IGnS5M3CJh9lIDbmEthU+
kfdx0djX7tAz4D7ySfhjiD8ahktRvqTtTF2CowxZKnwmWNEOBAzGI0BeKCaO3aGWOGF96G2tJ12B
lQd3039wkWIVqULZ0rpHUSYN5x2cqDpdH8xPdBO7qCAjADtRCr46JD659a5sCifIBKMGRuvy8gJz
/2Fz7AZHoIHpOiUhZD6LedVrfE9n8nP5FfU4fQThJoEBYq/JKyyjV6vrjhe106nBA9k9kOyP0tGb
uc7sEf6v/FvzUPV8c/KNVEVi+GSvRuikeil7jDtTelsNPwdovfwC/aqK8TEbA7TbtV3HoxS1LIwV
9WEIq7ofpShvqtvRM6WQa3EhzsoxqG/KFGySxWnumzF/VfYbYLclgCtCBRdDYFe1Bqmi4Phv31oZ
efK69rltAJ4Ficf+jNZm0EJPD/codIZQU49KXfwQ9GhbrQReOaMyzNYOVcBeEeFQY38cxJwsG+xB
22iiESo4oKv0f89GDj0sfLENeLxA2GelP+Xz1kpqkden/mefRn0+s0i51JPST4f0VSGOjO03LHKW
l5OFjTrLs7EH5AEZJzJb6gNAlwULm5cQIEx/J9lw7wdVE7pZRND7bd7jyZDA9jcVG694dQCSE9es
T1vWTYcC57d78juoBf54kcl3+wwiqeuRnM+WVBbztwGH+RkEcDfG+WXe9ba6q5mOdzp8Lzbbnaof
+pSUNX2oGnvReDBoQ6boCI979/yz/EP/3nit3wcu5UqmKsmmAiDLaLOWv7YnLBI7o3vvpddhi5vb
VWQTqCUBT2CTiSLDLA77pgpRWP8/ZkkFFoalhZMhfmh7MHjNaqvD+OfVWNUbsQ96Qed7dwMLFk5X
Y5sp6HcWQp3mbPv8kjqsZyP8Lbt8AFfgZh9xF6Z2kfJsoiuWk9EIz8FBdV6SGROEXZ8wr2ujJkhU
D6cxwJSx8TPc3iKKxz02IN9uzzbwKFUjQaBJTmwfE+yObpGKa6soZmf28+ibDZtUU7NT8iHEBUCT
JciJyqlBBLFJ8tLxxv3fxsypID9PPSBdq3DDKW46yMQS7zLDktSfZA0k7ZxjtmXw4Nfh/kh7bfFL
uW4xvlHJ8puU0suxtwWKSMwPydWJniMErirLXiXiqdb2oYoUAlR519l30yRosujQhmOm7rbjccfx
IdVtzw5E4m2cbuJr0+qvihhc7TGBxU0hqJXMlPURRxtXBDN7JwCdnximXabi12yuvJVogYqLEiqu
KHIQYXMuF1x/I1OYXiP7LMGbkP1oib52Q5IRE/lJ83O5SbBjIBTvvdND1aE7BDTDVgp8QTubuXfp
5jQfHzwQTExLvDmDeBvXh7u0oDeygTTJ1XP2QoB2sWfdQ/F0QfSi7ZtIhz9NS/m4jYLHjNkjM4hg
xyLYof7IW1PRGu1hNU4UYTv2rL/GHGnYYcEqBWQHt3HV32AEVpSFojZPeGKVOq5RO2yJBHZwGefd
NuAbWu0xRkyDq1kwRIDEeUlQJIqkB+k6TlqGRcjn1NoJvS7OwDAmKr7Iml5AQYCnNVUswthwpxtq
dMSTiJSO1IZ920hADhjVSiAH+rFt93b8nTPdc7ydJgu4sSxkwcrAXNqLG88O8tFiIgs05iDNt6uf
1cCS9FG1c871KbCiXaf17gGa++14jP5yO3se1wz1ahR6IE4N3Tai207n1yUZeT/UJ9X3gAh3POGX
lmiIbXoJU09VpMpP9KRC5nuclQZJYohWKm1RLQEHOI6kIIoMkC+3G949qyk9iJXfNfmzvLIcNbv5
nmDykCAnX03ow0I//k6jmXRY61j1rUODs5LHL2Q6owYd3qiDQQvwlsmr1sNgWOjMyoGaID+AmhuU
hkBD3KMr0s0Y2st7l62oz5Q984o6vZryU4tgkFzzCJdvwKQDmeXAPjCehj7zNAz03Rpx7MuAOijE
UuEDsWknft+MJiSQBCMXjOM4OefLMhr1hZ5Gv/KGPa+41IzZpxF0lGh80aV1vPLa2NoeUFbsOWBF
xJ2jWutwbv7qtI4zc5jdSrQP2rWh/OX5F9R1BqjviqT82i1GLbZahPUQ0UfyXF4qNI1rT6l0UROb
ZW6NP8hlogU8EuJfL6ng7QizbsquxBTqyJhcjzWWtr5WpSqHGR9K6rIXDFpwy8NrIqp21lRJJRWB
iCY7I4Q8WiVLugJXZjziXGBcvZ3yDKGFMFObbLpafkAptcN3WuMQfnEegBo7opz8Zk4tLmy5g1xB
D8U06tKG9GMT/XlHOqbUsA/UagggwVsy3JLbrmw2k9FqA5wPCBNloUPShXQCYJaWHkT1xNhg3O2E
33/aIHZ+Wqu6tchHkFbdvqII0ZszDq+SpVN3vYttleMAgmUuaW7qH/+mZAw7xRM9IiZAYCkgkitl
Ra0nr9AchtBeofSEbegkniWHd29+7qfZtNjjwFMq6W7PIDpALhwGJxEL0nm28x1F8Jb6SvptvBDI
PqaY0n6unyRXanezoPF9PeMMrs2wCL12SUSivxswPRnF6HU85YTHv6ezoHmXDZbFiPunftbmQB7H
9pIUuPtP4kksZajNmP7s7YbpjoCwekHJPBEyrXLV25lP6ak+CbotJaPTt9xvkPJsIFgFEgZ6B0Tp
gqSwiSF3lQQttqYoLZuj3f8hytG5tBdyKEe+TGbzL6hiO3kaRAR2gbfrC4mVHIHEklF9wrxg8UqC
xR+ntNZX4PbUo586TOqU9B3oCkjFKlPEyRrS1MBhuB6I+wAJ3DZP3J0UPhqkI2MvztNS/Huukmrz
GyFyrTLRbVbaqO+BxHQH/Ioivp9MJkRb8ph6Q/OcuwjA1io1xeCOFLcl+zYWBpATdtGzSCRZs1hz
R+S/hYo5xl33SmqEkRkytszlhxLpMIr1tij/FMYtAgpPo7yCUAZTVZmzG1QLC/B+okq/3SmZzrm7
yrNx9PmB3sBNYzCVhbA6s2JLk/55yuFfayFqPw7PeZToIxipuTf2dWBH3GLt5e0R2UZzq6ePklfV
v+1FfwSW3XyEg6dgQt1TLfy8OtMYIoQ/U90N47iw9Q1xRl/2df7kDq35IOpPFmh6xZchn9+fR6aN
CuIt0RZ6nMF2tTrVB5tsTF6VIEC466aVWkrBoXXvmE7JWvaavpMJeMeYcjLlxaMVr5feYJCEWP3L
CK0ea9HM1V7A6Hi0/3N0dbDHlFoIyyR9B2uRMCs8eTv446caXZ/t8qYN7B+6pmF2X4ST8yvqKTHt
VCKIi2sLsBoRdDEaguV84q1oAgyk08eNXhmCFZFOWWEWCwMaU/iCAdfEt+HF37HwCYFQTa/PBmEW
C6ErdSEEX20GouaNHwiXb+Q0D+e45rLiSEqqXUZ2kPvQiq1ZjdRHHA1VT7u+t3OpknmQLzMDw0Mw
3GP8Ow+rtKhjC1olCrtrsT3+ePcAvPZifH34vt2CDWGYXjgwKk5CH7ovPf1lifz0BytAnUNDgt5N
qJ8Gq5Go/DHHMGKOKJ4iCTz586Vq6ZxyuUOjPDQnDG8lqqUR5eCdqGGhYp4fakPjdHlBSf26fQX8
N/n+5mqlSQaWtJKef0JcRcMlAHhzqH5dYdWaBL89htKB8+1Xl5SUwtj/2DGYIxykYGrnN8BUSeuO
wr2HbvIoRljEV5iAzzfi8qqCqvRzyzheWUO2geWWeatGtcNhzPNfK+oEeAiSiWMkuJa0kyfvxV6A
HRT5+mn43Xb6vIwUCFrvkXlmxLwf7mz84Wrq4jY/v4JE3aDty42yz40S1hlQohnMvYz+l8wLdweA
L+XolhqEfceYHVBI51yyMPFUqrvCbuNd9+fOKCiulnBjgKZLTRJVojR69S9HeNf9zDvjk6aIpxDz
ChWa0yC4ZqMcce7QJ3OCI9pmxWax99foP5XuwTGLFot2Yd5SFsoS37wSH6O5a8s5ysistDhAVlpv
IIYCWwFN9YYE00aQevXDHEb99sSGLo67YlcHsaJWGmWZ0jJV6UmDN9qWrGtAeK6eIit5jQoKXobr
IV7Osd/gpzexoSfCcVQYs4UIg6HaKq2lmXjQaG269KkIbfRTyDJipfiw6meuJAhy9hiDG3CNlzgI
snQs2j3vnCRPvIU2hgT4pZMfEM+kc/8hXbiUTYrcfImKpJll8WJqBI+e+BWvashINHgAl0xrAjFZ
CnO6s6YIlRgHwNG00Uf/NXMLOPcmvJz+9Itj0rI2v0+lbI8WpruL33jZtSPtS4v2MHqQ/4R4vRil
GEYUxBVbBYSBtAYS0ZDNGVV15Be/7MH/9EM+FXnMmdoY/9Ym6ZNHJ9ZeYl74+4RZJnP5OMexeAlC
tTZ+Ss8e2mJ7/EuzOYj6L98i9llM0idKAXSvySfajIXnQc49H/GaxRBjjipRZsyz7Hd1eOcSTchY
yPKQ5wIePZzR0yjayPUIau3UDhhtufzqOt8jtsTILsv9BHSShUliLDFNAMHxtfF093nknwhqVHQg
4NSB6dmFezO0EFKVbPBXk+zl0B2sifeH6m9/XMNxF8IyQm+/BbCqB2t8BxubsVh+i+MRLtAvyKr/
3RKXb/Z+lx7LiJNfXhq41KAr5pA6/kEnmu9OGaHNxgc4E+HoA8W3Wf7bTwTqc2Nzj7GBH+NdOUIZ
NNNRXrCL72E3CUp/JrQoyt0XMQcy2YQQh4YN+3PMay87xz/SwgwpjiV7oSp9tZrwBxccnIQU0Euk
0ZyR3cMPsiIj6I01QSpJTuKmaHXLnj4cR5/1/nuG8xMhnQqo9m4AD4cObAs4oZZdet7RwGYtHkp4
+9RpF/JnoeLI/9ZCD7zJtCTMH09xELgJZJDTmDstcUYRWhrvxt/6RUTf5vAQI2wChjVmzVJyY87r
lpgDWOTJcKJDHGzZB9wc0+NhifCakHPLIEvcZov69TUiffOvO4ldHYW/4N/1H8eKXO1rNPln9y+f
G5FNa+c8jIi8CPzgY0W1MovK8r+h5D2wlsb4NBENbFel7/inZ8yNnA2agJy0NfuXxVnefbqHi48h
1DDZ0cvMASQ9QGSas6I3tF/b8GoevJlqrIKmvs5Hkn5bbX0RqaNrkln9aHLRNyFcoFZ37PpnlGY0
b/5BFNJOoBcXHO04H723lHKi2R3Af2/baO10NjlUFLw7Me0MQjPADU6jiRUm1jL2iTAANmGplstJ
yNSVqBFQ/V8L9o2AHO34F8gHrA3QG2VwJTWwh8iy8rfyFp/k4b5wVWxskMhuIBEGOVpodlToaztI
8HXShKIm0j7fhD4lP+Lel36ZRmZPPiPI3Mo7HZ/6SSExrqtC614x6qi7imQk1wyQ0Xa/n9lvFYG1
j4FS5EkB0ZSPSzpq1iPCMoTJklxyhE9tKEvhMDmvzT4iup6usKX14OBYRHjx5gvse8Kw/Ml2D4se
d+zk5cYtn42yTM9Vb/XWJxaZqLAcwAw3xylSUNZVfMlO/Gu/KW5IDZKp6G/y896M1rYUgpnjZJq/
p6PZChW82xRjPaHYBWq8IDqEFGzZSKhvvTZZXt7JqMUJJGQ8DSc0sMbvpkA25Mp9dY6NOPXtnymq
OACYkeHouyuyQq8fiNeHguWKdZS/OQR3whXBkWwbh3DMtFwip7o6HEYN1/AirPh/W7yTbuyP/Lk0
UTMcplAObQ4f52T1FijQ8JHXiuLprM4RqH7H8K5p3uF74E47Ci4cJBzoy18XIZvqoGVVDC2xHPZU
icwE2nm/M8u4geucGCu1l+3g/aWKc+qA4B70AMowRuXJwvdY17+R+Jo7GpoQWnpLFMKyA3Sio/GG
CDGEgq20/6ycqShcP5kKQCvE5EJctDvpu15coe+Fq0t5jPzqGgn9haL1WnpeO8kMyRxSvG84dH8b
G494PpsL3Tnzuz6GmnzclLKq87F66K59euKF9bo5zhvDSdZAZXxPqev6JjglQcVSDdKqjpDmpxwc
uXqhg11JgXgCSS0W4yXUfIfGcCYhsmaWWAY3ndNw5og6qpPs9i0gbWG2T9AXaFTURXlK3kqmrBrw
I0e39iJ5euES9mmSawR9bgAMoniSkg1eMlUnr2fMQIDAI4XaevLIwVfown7n7SwZIj9zwZxeavrQ
avcV+l7F8vM/EWmghed/GAbs+Y3DsHS5QFxb+ZKgUSSsPH7gH6cRcUU298fz6ULbXoPR52yR9klv
5MVm+lvbtm1nlEG0CbnA85TNLH+wNLBkQ2ZXy84rmNLGaGa2oQRjWROA7oD9K2BG2tWCfFqbtmK0
d0fkF6SspnrdwnOd4+Jx3ulGMPfgw9aDiBhD8egYfKg0ort4vuN2mewzuoaKrvEBsi+t8gy4+L3J
BdbaVMb9gUdj4oj87SmzqLkgQ/ZKE0s71svv3Tz3hzQEekWYd4jwKcCRAG3mIKiiItzc6Es+G+dx
MeLMFDoCUMsnyCsewJBgWOvGqIi7ej69yRkT2YgHkRkQdtJQop5iohSNdVLPEg63tsgIgg3VN5sl
DFtbtDhIJ62N5mzqlPSZVe1nELn/TnxFQGiVGsA8rwNuhEa4JOUIyxMLLRngu38N17IrgvElmCgI
N/myqYzf7tFciomGiVcOYbYjsZDRzxo+kwdAHKviwP2WUXhU7z94duj+PGlGyyr5y5jC7HkSND3L
g1Pv+vDBYz+R4sK5RkTvNtdSS/wSnLlw9qWbkrFUN1xLu9YusALT5AoYXPUjzYJljCqcFI93ZA4N
IX89lpFNOJb7ixZdffvPhNrrGpfqkDHO6FNrSTFibt717S5iTYT9pAyrj8kAprtJCkdilXxfKiJU
Z23864KsHcAMH+ND67ZcmkPZcU9nrb9Qzx9i7kAZRWePXJOuLyrNoUaGTekyAt3L7CNhlNvDLw/6
e9GsnA7HUc8YcCxJizP9aTcP9/8TH9HUQhmnSWuAdxuUo7+ix22+FveKrlCpRH6dvc5m2BEs0WsQ
DOTusdLO5Fv4fY5ag5EsmDqEPnWNno/m7Y6qhc2rFW5/ZrJH5NqrFHHE2ddaWqc3WTMl3DXfUlqO
NwzqWXWoMBA5TxKBbJze7BdeCKQTa9w94lZsECWAUOGrA9fnchNfudCzJMCyyr9D7P/6Ipt0MdLG
LQEp3ItDDyu5zV5iKFQmjxrhElGuYBfuMhER9BSsUZtjI8rthmOXaC9uP9Hqga9eChw0rKz13A2X
WkpZPjYOhIxfVM0pH9hJQBsXpd5/+6N14tSEQpczScHUKt0VNj1ddTh0p4q0BoxSyGraCD+EDLQh
QlUTj/bY/pjiV3B40BWcKTNQX4e8XEgay9XyOBVH6Asa9pWYAKEKjYIZUvs7iJKoj3nzvFDDKqKv
WleTBmco1yhDibzR8nYi/Hocx03Kgr/8+XR+O65v/Oox05yrLTkkcKqP/JvLOhQDzby3+b01a9ji
1SYxyQ+MnMVZ2ehYED/bJI7Pl5CICnUmeX0Y/mW1Ju1Di6dH2ulzrIG0BmRkw6I+vGVG9Ev6tZZ2
rdn+B/uJNqRsqur36CjzfR9yZIawUIQ7zg5OCOEdQq04Q6yghlcbM1ZbOP/CX1YCxtWLS7K8vOpx
Fvx4t1/ugi4ZHVmH0G0KBo+ZvvGqScuyg3CpawLlMAjBpkAsyxkZvBdZyn0pz81cs/kL1pQWC1iI
HjYKukWf7bjIa4hPTQ3Px/ur7tEelQqV1LATFd+0dKx5p3+nx0eJbZnEDhWMQVTm5v3XLTY12Vxq
tZncJtB+CoS8otYYkBXAkTWNEJr5S3awJBLnsuF7o0F1OKt1N8puyB326K7fPj0mB+UN83VxkuvQ
R+8YFwQjvEVitzsVO7mIdgZxaEBjpeOfHw6L6mTrPZ6FR7676EBsYydTgdKBPvrYJeSZg0vdctG2
ugZpsCUBhuYfq6OdTngn+0E9vQTGXOmX/2BLZL8J69eEdPyd2AqaopwnSZhE2HRtceoUKyh1mmDG
YlVOpr7uLwVGR7XkwJcgr182kUtjm8Fblfux2E8Mk/0XyoNsUVirqG4Nih2Elin0KhYUO6EvXxWx
6OJL9ieHSz9ML70VYxSb3CY+7xV7biEatuWgLMmRgCLbeamofxKCTYGHb9wXiOZ2ZGwUkqejAipV
GzMoH9qgvX4gmG9CUVQ9Znu2Fp03dbBVFNB7eKVFs6SftKp1JExDRydstrd0XCH/AqgAYZVUUsdf
b/3EuABjoLeMD9KesDUgfaldHrqdpIMLEor111mr237vVWlmPuYGWQlT6vqT2r7WN7e79DIDVd2y
Sy5dcUPvAw5070h6TXUcL39H3QNwrqKtuifDAHvH0nf88T4IcecpaTVEvxJQnoybfLR4aoMSp+kH
ts/td3MPqarn8oFDOeWFnJUEcf2xH0NeLTrSrDqXWGNoGwL0HKxcZa4XoYWdck/E+l6sbaTJBY94
L6r1UKwGi+/3XxLpIlLm1kgLrnKllcOhOXQYOWXhB6MKI6TlUbr1WHah/9NHsWatvi+mhCSAQpHU
OMsi32PQdvbD6WWYZLk3+OElPe8Z+lyQ3HnqAMdrLyv21ssqy9nyMFoOSbMQGSa7DfPok3Nij+Zc
GZPVitnJUEhb6iWy4u/fwK7wkuf8BteQ0Y1rLx1RMLZAXeaJUEYzOqol8KbRVbuOCq3IfSwAIJvd
dfguJVh8OOpy231PLsWn59kDk4+mjIkh9tbsGM6cT4HHR13Xqctfac1veLc2lIPGL1K7uoLQIcVU
9p7VTJIEwbgtOQ6XUGjqGzGlYJKIRhTp38KvKdeShAn7TjjDMpmWmKJVOvbX2WLoqZmDkG4XSWvb
rlFPrDuhXorpiff/Pc6AAUdmi5lfU7b+59oZG0uhbsowHbaTv4ASoGXOC3S6dCPlELZzHx5KRvs/
mY+WJjrOvMMVL4KX/SDYooJjcGmuL7tTZLf1kGY94TmYqRqTna5XRk3pcMyokHd8Ip3KWAwRd7qK
YOydyyNr3S8RX9P/lr/AHADtpMs2p/XnAQEmNTV0g80BQfqMJDgVcmyzg/dlS479gDUnpRTQreH4
cPdpopIEGkDLGndT7dMOP0ODx1eqyvfmGWGSx9HSUJLPLnHE665KqUsCRmRSgpD3cLOEJW/gh8wi
ZtUO5LUsNBI6ZwAFdUg0l5tHww3rs6aUEybQ1qBHOd7w0zviuasMjF4QKn3fVHLP5tDEoueJ0ecf
zn0aCzG+UCLJV7r9XSmb+e+gFM841MSXdl++77+5OX0XT99UiGrGwmev7M4IHSwzgB9IhUQXrI0E
rSMwCSyx9UyRQsILbMUB/3IiVYLara9fH9eqjYMtBvEu5Fv0zuKByN1WaNAk2a2bUBrIkXb8w6v0
oq3grbrLaWCjouFSlX9R2rCfOhzi6CDsU04wUXlWior6f+bbUjKNcltHXAH50HMrk7Wvv9qiQBDe
N+HPgMEDR2KPP5gyphiwl9A+sQAt14eZ2/DcuEy22JGjgBsYbfJFP4uz1ttr/PnBTMA9omLBwUra
6lLvvXh35tXbso131yFLLdpCHGn24/OGSwgSa64VKPXCID8CfdGYld97JuyDSNjMxjgDUW7/zi2E
IasXJX6zJMJ1+ROl9T4tLvH3Pmaymou+Cuh6GaYmEgyLaC5oukm415exZRavyzUT1y23sl6TpEXU
REDSacQdX33BsP9WSKFD2yPaumnqYv9vd6Q3OE2LgjzDzv/h59dUQ35KeXj6z+YzNZ/SLEBNJK2d
3nKYtU2Eo2R90ugZRusHDHS4neZdaMByKqNVX1uDggNO7N/dpC5yIQTQs2QOITJt1ezCJG3/kubr
+sFovcb9KlkkRhvMVsMm/fnU2FRyAH3QEXWwd2xNGCefGRNH5vxXCkKEZZZvZ+5ItDNsV3S6Qyq0
PPDHoMYuokwx7i4hgC38aqkSCVWnv3nVl9cs+8jcxbBJrlGofrjIktj9CsnPnOYk45NeN6IK9VbE
xG524liGHmW76ynhrm0Hkg2PsFI6GgqtLQfd9zT2rdww8Gbcp5YAHXoapLwEGUyx3kq8cHEIHDeT
UeYbSTb351NuMH7eQj4JX19MqReyU5320/H5z3o78cTBV7W/MA4PhsrR+J1LmBbAb21lcONfIh7F
ifd7yBbjXusFUyalHDMkTEItLsjSyaoW6NeG5qz1/J71l7zQCZvaQJmfFLD/JWwJCynkxmZhShp6
3JEG3p42ptWVRf1VDSTSk7lQTq8CIJgZwSkJlwA2mkxDppn9j2+SXfQKXAZL5Cfg/ykkoAItp4Xy
Y+Bf74PT61rG3tPnZkYvXDircaMnR/8g6dk5YrzLGiR6ivxYK6t+/3uiJbJGLHO62o9d7gObGFDK
1bA8IW+i3W0yKw8affByVXwETBgQABwK9Q52m6loFP18PS4hIrvTX0KVJgR8nR/2VweajVxRH9Ek
4uSADMVx+/WKubzBqftNqvFuHTA7yfxCp+BYhfLdfLsSM2Q6OX6S4YMNslyNyWoEyqm8MQNy911b
OYKzUAaU1jQJAS7XxewZZ+nRCHdJAhaUiJyrNiwwA28Qj1HVmK12zfyd25bY8OR4/ujERTB8vGUi
X21ehYY/R40h2tbM7h4DCP7YPAwTjLP8EYiutxe0jSF9mMaYiLZPckCQb6zohnY/KePdCVJQ9DrL
h33MfPdMbCTI0UAYOPor80ZwRrxxhzcUWoZzuETTHxq8jkuUwZ8dqX5AUsG+VKZ6Oj+pScqlud5R
934/mcFHCLRqhkN+h1dZ1BSwHVfJz0rFZNcDxwXRX2XVZ2v4s+9+reZKaVN8axm+lSNRSHtNJK/M
yb6X76J5NyNemb578+Vxf8Vqa0uVOdDYBIZXKgF/d7Fl5AbaV/tjzzpLgq4YaeS7tIWZ6qJZqiu0
cePr3VJ+OjMpgr2Vgmh+XoTrK2XkaKG+2Bq7ug9fc0w2ZrZARKsuX3BrQfa0U/OSSedB4VU8mevk
bU66XyUEUf6ENneZiXAcK4ZH42s9WDPjILABruAOXrhauoIcZTLewl9tAxSKVnLoAigT1LizQlDj
sIjfLiV0DWg1/LGzqxnz9pqog7YfVefN3gbQJrz87eRt48u3v1iMCIiQYTt5GBrknzJLluzwbg6w
8mWdvV1F2/YFxe04YlfcALpgrgxwYxdejXFYPPJsvkcMvPSSsJDaGwpFna5/+uqUXMdx+I7AlB/v
UiWIkHGUpUI64UxcCqBJnOP162LVp+MzgeWzQ7CE6zgDuABMfWwNYjSYiP9oKDv7QAi0F0TdPW5n
u1M1HJOWQEus7t5w9pIqijXVxAVdog+USiH2uTfwtPcSGFwbAi8HF7XKsPjZMWnNhKJwvu8uenNp
HQ2BFjVIMAnyk1KIfUfX+IB/1+p4TOV6lD3uq3i9oH47qaAHlLl42SLuC9sfBCQsl0OZ/RqR4p5h
CjBsoZj8GqJhTxe8UlpOOnCVFvLPFUOb6wIOaQhbqcCa7tUx/tLYAb9/cQbW/g1zXiwW9V8h8yYj
6+LIV40q4Ei1trwd/BoASHzYjWVGVd+1yIJl+O36BQVnXzrtWyLzXEtFJ0RJHP6rOfqyfHyUTkhA
/XvAo9f/3U36tqI4e5sJZHxkuotEApV/wpcNCxZ7L1/C9uVdanWKfX+5BIGRrKD0CuVK6OV4fwiE
xwHtwlh0VtVpDj5XOmka58F+yNSs//rl0bVHR9y5NORBfOMkUSHLq2vhAJcrhgewKS2uBI8g2xKo
lb8GIestoRhkVKbCif9GUpyJljHxs03cUOpR0/nty5E/8A7Imbth+wFFJTAVBt7KOP1Wc/PvxTYE
VvX2dGOlu81MBNGHUfvsmTsVT1ljSDHJwpFWFYOpMZmKjbmvXe1/mbFrWoBdAET+StZ08FuKhT1u
ZxDAuf/Drq2STwBk8pnIN3skXzKGc+wMfb570Ic7ykPREras0N7/D5svAJPSIK61/l4OXCIaOGFs
KQwF8ktGhAohhcVdfOpcyiYD3lr+LLwd3wG3MhTEwsTDGYt5aQZ9ONiRoS7FS4vMYAogiJxUlG6u
0fC9fP6kZI8i+SfD0lKbCzpJQWk8I5bS4RNMwvkeYSCfzQ8CRKMh8P1/L6WWQxpXUyzuL+JcLLvy
Y3bDNfwkBsbCfy7pyCEFeWzQUYL/tqTWQ6pMUlcqg9Um0XWEZDRjKJ9ehUezYjCuEUvkzsS9/fqE
5ODZw2x9K1EHv8nlCBByFyo7nha+9hgnk1e3H1ncrEGvUmE+sCqkeQWvgonhH/KjLRDXTWevZhqG
IWjuS4Ek6zNuOfrwAAklOiGV0Hw3ikiaLGitspg3zZo4g660LxpBIya6g1yKhkoHTu1A/idcuPy6
2UOUsxUxhNbdMLw4DffEtrvgw832yIo9ETEY7J05mhj6wo5O+u5+UOMu6arI+GZmx5K4nILqJsSP
BWMm1MOgkH3WcD8e9Ur1OCz86U+VUi0UVbbvzsXxozzh3is38vPr5ntalpkNsUBwsrGt/aEEPYdz
ZyOZ0HmDOQl8QunEcjp664b5wEI0ktkbQZboLAuVh3kzLnfFey0u8yFrI12aiuAf+VtoF5fa0UEN
2VP0C/40BDAHdICcrUYDnWB4xOn0OV85yS5GO+Zb7aEzX49yBfKpEnIFOa2GoZs2VctbY+Hu8GAC
jqQIa3KZruiA5jgT1gxe/J+Lf/Ue1cYBiYpl/eC5JmDTFwNbBHdxoyL8qRvaNNtgHCSGR/H41KkD
oM9rWqthQcIOMMUXWWVpOyvL0ok/ZXdEMcCLZVoboHTHJKUNaTD5P5hBReWfzPD7pzu7XDm4x2T7
jnAw356lY+Hyxyh33IMh+XQ+5V8QpkkAXB1aSwxZ+IAAL/DowHABdkWRhOqLZK03YZUHOktI8Dh/
DkRNa9SSZtVRNouav7rQ45jif3lr3c89Y9waT1fdAWG8qdyKuFbAxbHg8X3slr0vQDF10Ya5oZmV
T2DA25Qi55igiKZQjlbpfmX1zynIG4cxZjB/DTpZRt8FCDVZABJNhL/4H+mqa5AeIy854rRp2PsF
Jytq3MOhLVLnBshWEHdPPGwda1A/hY0aLTgN2DIEF0/FG2KIRUR/YpfeOSWWlFvQNFlFa3wrA8EO
vZPFBYtGiN1vXVovRnGH2/q34dsPvtpWIBbrQ7BXS8vwzjk+7IlFMaBHcBVcltaYkiz9TLddtz0W
rtxbdsoM9Il8SgPRNcR1qG1XOidZnGuab6405of8Un4rfCUy648SirOP5MALt/1v58SJgl6uPa32
DTU3l4T0HeotVLfXU01eJD2GwFdclsTPj2HQY20nEmI/R+0My+vYskg4UvKDax+axX9nkSDZxgom
WiSh5VCmJXT1a0SMbYP4GO+BkcKse9y91iAeA9gUxUGhjPXhTVVSpVmG+tb1LfgJIoDWQkhZkDuo
9ZgXIJQYVPA5tz+95wwZ2ryjWFHd+WDK5hz5GC/9fSeHcrxq8myc+PihjTXuHq7dJPZ7C/hdJTrM
ylrjiByhqkcqCbPf1q/IDVWW1D0eljxXEYDBmxUngt2JF1+z+Q9hSya+hFEOBwOqjrNdyS7BYh86
8JsvhTeFv7iScO2WQyuyRsJla0Ih+hqbwvbP21sOnxnREOX9t8j1wAYaG1jX82agFNrY+Bg/eUJj
IZZ8Hbtl7yT+BieAzdfESii93qhKaba5P0+uKV2b12rc4uqVdsp738cXCqHvWe0lSI05SrEIGjCr
N418pDELvGsQlkc6CMuGuGtV/Ksyb9dSamK6eas1TRq0u0j6x+5u96iJbQuDH6UMVVmdPEc3TuNW
XVTe4SaZ6fP4JXJEMh5aN0LjhpXj5uj+/Wr7aAD3aL6WexChOy/tfTBFe5OEbpGcXtHnT/7VKXrU
MDHIg/69oQBPpMKc+hLJ0mrlMjj5a1bqEzFAzYH3hAcqx52QFVW8mEMy6UELFIjiAWw+RQCx1bo6
JXTW8jEgNzP1axwIoVBfyy8aDvNGwxKE7Bo7Vb3YLEBPKtyuRuveVCw0z30d40ihCb65cI02x18k
g5EOVu48jE0gloXyBGXpXSpCNINFqf6EA6kD2XMpc9Y51F09qapjKsNwzPWYsTjzpuBXVrnFLPvA
tGRCt52y2ldFspBApI8phm/oD+l7j+6QUyQGAFKtw/6F0MSaBDppPCQH12C2tNDQwTrkyDhu+VTw
s3oqJQUyfpXZBCkuI3ftTTyWvNuNZQuw5RnhJF0Pvys/Oi1NLc9YN+7BZQXe5DLnMik26kxC89YD
nhVPCMcNzf7xq6zMYNgEnfFynJBtSqxQRe8JlfI0CxlDFnEbVAmm8JE16ATGAX+mGVAc5O+WC106
XeH24nqoDTJ9BVd2Ym5b5Jc2SgQblMgAreJhZzusIgxq5B3/g3uDlKAQqM2RyxNUuBOTF69ngOX6
wpSl92Whxxf0MnO3Ss2D+kwS+sNk/tszz63WNATwrczc5JK1C95oiOc5bWO4JU11dZ9FENz6eGz8
Wc5RQv7LzAJkK8mKgA5z4hUWYtOqbER4Aw5iiZp6fOXnmfHkRvykxrWdB4oHajBSrklhgrrPja0K
2vTstHwRzHhxgdGFGevfDzVMnh7Ul9k/lpklVwx266pvcy4+gs8RFgeVGimq6Fni1Sy1d9iKJnxj
lIDuMnYYtXbPz02Yv+n8A+erLoJQGEyvJBuPqNKnBAYHY01S/h9kDmyo8sGEef7vFxnTyCX9vByQ
YtNIKWfWcVs8Wm4jw9B31tu0gUm/3sj0b4YtVAFqhLCgdhtRMinvIrfp4S1z+thqSaO/QAP0ot6F
LznGR6qY+OOp7mVYCqy/ItvgfE0NmsWXFmpQtd5Rez7vuMK3tOg22IrfpaN2fBHcnE2Yj8VKfYY2
yHeW0EBCAOr4+nC0xUFIKOhNP4/ThLX/z02RSSAFgfdgCBaUR7YrBiIcuX6EcrpTKaruuM+jDwZP
nJWoy6yGGaHx6xyEUTvuwzqYrXTw6E2UjOJjjIqtGRkMB7k0goO5/Ay1qD6XfWGKbAebechlssaE
qrazJW2JHqvVYUH2zUca0ulETvnn4aNT3EHGeF/QiwRf9DvvwH0k33czpDiZMYCT44LK5Fwo4P9y
NhXLDkADUuO+ytn8Y/M6WhZcHIaQ1kjmt1BZIBftiRoqPsoYeeCn7eY0PmvOz651I+rGzfX54ClZ
ct3VmygGoTkSsiIOcUynCGLcavzeto+fF8sOiNQ7GUMk7IMZaFUG9/C4VUDtqczgRaMMBMVCeGR0
JVYjHP0p9Tof4Pg7aPSyjL2Zt+93gwwg2N+zlWGJ6jVpSxsAQYQITib1/+beSwuoUjwY/iUbCsKi
M0BiSTdUqdiWJFkPIaCV212K+IN4SilXBYht74GpKAAQpKRa8iBVt7cgSQptU2fOwwJ5HS2IJej5
am154Qn3yjxr7ifzLh/DJoWSUc+zGJYk1tPFcpdPDd+TXe0kfNNpPx+xWgK6wc8JFsDxQRe5F8kx
QHcDfgh6K9oh8cIFrTASlfyf2Q839oc1qP1aaMKPOus2IL+USDeORta/qTaj9R67pcE24lRfjtq4
9Q7sYZloMpnyDCh2gZk94UN+qmNjcAK2DptTJkWliFViYvOilJKonj86yhlvq1pgpy+3cT7SG4nF
R9Ai8/f0E3u1qqXsBWwmEWQt46D2+/hbs1gf/okZ/bbc/Ens+mlnBz8cwACfTlA3kzJTFQOaU1lQ
TbtnUCKgBRpn7u5YOItRBcKZZY2jpulZNOwXHPEPK7z1QP3Io7DCpbMvz1+S85y9dMm66FgaHwOV
SH3ZpNk9f+NOZRGV63PdASi1Y2K1wARy6u1z9aYglCAISAbknHNZxVcvZDu9kUYZEgIgvWwSJ8At
wCSo/KDGa+W9Dwb/MP0j2tmhE5JaOeUWpymyGz75meGxGk0khewosRmw8gcsgJAUGMYf/ECLInfD
HGTSNh6XP/Pe0mZ/8yX8KkTASsc4s+CRYC8270pC3JCSK9fw6PH7vD1W68/d2kWNEkVoDkqDvQ++
uFoNaZF8WHctw/toCALEOmvPOijgQC938IMSETgy2isp61Lx4y09NVjrbMo2KNah25FZkiI7l+iX
iMR5tcw6JDjvWmCuTSV0mfRXd4jZ+Vrrk8WRheJJWXsT2sZHUCFT/au/StpHbJWOGeSUTb7HkGYb
wqyjrZfWIboNtrFgcKm7H7YBFHMHornbs+QBc7etF7IveUtsLgwo0bmXI5gnRP4glXaZshxzI2Jd
XfQTxklzq9hjfjqqUR0RAtGzdt5Ef5K4GVtFaX9VIWlP9vzSJFKAMMaAqFO8bYHER2NUVw+nBiqk
7Ai/oJTmPzFttQ7Y0Evwdo+KrShrMVPwqwvC5tqzIArq/lOjY76WRj75w3wzcD2aIvf04O5bXhsS
+CpXyuwFIvVLKF+A/5Y3ZJMaE2oYfyaZdnZXsMDfELYWlEb5iMor52a0wgW4DG8vaUtJt1wn2Xc8
jK4nJpyi3cCtNGnx1w6LaiTHRvCqfhR+9LzDOinxDUUbtvnlKBzEBUylPIKlW5CAehGwH/Qt+D7d
yKSx2PzKdIgH24IXV3ilG6U+OOghF1B7jFnz6/mdc+bDRAJaynRUxtYKmDW2SGIJsEd54M4oHMJO
98EllVQSMLyu/w+348uUZG5ulMWoDsJkz5rkdRyX7sgoIiGdik7hqU9GCp5jCMR5WrYVjKkThve0
+MTtg9euYgM0egeHJ3H2I5yppHazt4tNZAiLR4dxtOzrGi8K2JDSvIo/mI5xBfB2ZeZ3EpzXnUDa
+eKFEjHWnS/9xvYpJwQdSzeGRcKFbaiAt7x5SSeZM4u/iHUJOZ1TaKzchV/cIg2N7c9L/FsnCDRu
rY9+rGzxFC5p8gk4WKDYMs7RyLs+X1k9PCfSPvvaMWbC4H3vfuZmtdBVrkdoemJ9hUp5efki34CH
5/BaiqliPQmGSE+Y7Jr1n2QM3VEpjEzTqFepWVOT6MlXNguspRYLBPUrRjLnPnlNAKjKfo8m0vbg
BvF+3VCq2BMt/P4NDbuAebZfvlE+CcVIyaLb+eBkQ/xrEeh/fQqRNcAD8UMOByRe9L9TPQPOtWw5
PoR9476G0zvP+KonXfI73ZGXgIY1aNdivVfn9vbxVa+ksz0hzfL2hhTx1m4ZVh9eim4hv1Kj8PSx
6qy+Rh5bRjn+kwpYBkhhWLV+L01QKGbaF5wHl4R6jJKmujUw9EaITGtth6bc+9J2FhR4vky3g0ww
EDCNVGsuTmTCcfO5s4WlgKeC0WdE0yUZgpXHQ6i9ZjkkqEHhRDGpXXE4q94xWNY1Saz1f54ASr4n
eADKkjNK9fJ/HG/PrMlM3aDkdtNHPcFmPM/Gd/i5NSTaCu+Vk054q5E2fUEamO/FRwp3aQizmIcS
fVFP03Q9jekPc4psfDUkqPpEMMXD/3HsTV/a+xeEV0kOZy11kAdvmsMSui5QTKmqanP4L0Jw0voh
TJcK04YQ4Z1pbHqbmypekkhILC7Dei3S9khk4kI+BMQZ2EiY/i3D1yWzITIGmhpOFKoo/aWsmJt/
/eLTuNOfTbRQHzCaQf588su49ZscJG7g9HZcwozjl06KfRyX7Lco2HTGc62EtHIsov2B1vRFa1p5
qe0L+L2ElrVZ796RFSApXnEIqz5eTsbVtSjTYX+w0sEW1HnMlDIxn1WVHydpIMMF2L9sz6sCOLhb
Sk65AWNQmWT+E8QuSL2y3JsvBfl4uSGLP3SldEkuJRMLwriGtZN0LBDt16DRqhr82SExUPJNw+Hj
8xHg4kvsExLJ1G7GKDZKcg4JQiLJnwKqmUZQtP7DmRFqSOusw72jPMTVZWoGAHdAvEbKtdHJAQ8m
ta1+n7xWUsLlHVbcjV+G3kkr1aXdESP3FruJYzXBdVRxSxh9VT9vv98bmcw5KfiR2y5JuE8REpW5
KdcOnyaq0+aMRMDs+QIQr7MBJqR8wXZNomG8f0XI8TzyzcU3SXDNNGq3FJvgyt7bWfyLpcKETY7p
K2MrtBWPHF8PpATRzngXTJXJ2f5lD0I6hLnr7IMDHqMd790rfaY1VlxQhOR1byOBJwtylh/RXIVF
kVrHofL1tX0dHV4wEapH9Qxc911Mtj5CPVQLKWcqrhbQTLdvUVtN6MMmzMOAYh3kytEyDTq9lOvh
OexbkR2bnufXj7YaHN9caH67xVr64gxIoIjM5YUbuMTkYySwxwmSM/SXcugQHi1UETV0cRNmRF38
ZeDxAYuA84cAYpnNcY06LjMgk6FbLW+t3aRqAJATVXJjm5B3jS7SMSg/PFAekLK+AISo+1ixix1z
z3m7Fsd9ZjCASoJdBXgcoo04tH9zDMDxUgLEeq2jw2kfPuFn6MsRlXLvXpeugAWcVQRDp7GoTxgA
MMyZRGUigzGSwFdC1feWKojI2RHJ9SwNu9QuX7Ksx+b3rMpY2AcV5HM3JH02I5DMSMdSQgLyKdlk
xhNy7eSe2ybs0qbYtZkvjdv//3bDdpe7axeFtvjXnRogwV8YJcEJ4fFeLJ8ADlNH8M9dEkk8pCHN
R27x5h/yymsDuvedPllnxVTPRkSPF3baMXai2q/b4WbGfUYp4wKxDow4tG4rlEMRlR0W9f0zbydL
P3d8nPNVpMWfK3g0ilFTStHnf5KphAPT8c/fSOLkMsWuYqd7WzJHvML3EfbaFaaMtbxqTnNIEPeS
FWwYVKCx7/5qwNrx/hw9Qp7Cb3kB/x+t18rP7eiZAnIVybXd+/6u/vVYAYXtHW12lwpC0epSQoc/
RQ2s++nNJYWmC4HoZ4GTucF0p8aRq+k85q+aLv7HRcrDRIxGWV4kuTLBjtcOT4bn4OD/A1xMAInM
yaUYbeNxswqAOg5GQCUTvWDc7U2VMz0F3Md9hx6S5SK+lp+WranvT2M4VqG01vofEnyw70PDkaYe
frzM7PaIMOPJSBLzYtfK3binz8muu6pX3aDDcT+LbF1cFjwBrAm5c8+Mkr1XiETcOd9PsiknNCiP
cBgI6/MOSlHghChroYwKjah0EiNEK3QUe+zMidf3Ov676vP2as2Kzur0ovoh5y+K38gzYT7Qgwx9
+HeChIZbzfHrxaSuo2j7w2Vb+7+t7qu5v4GaIxWXTTGdMxl/IAHZWyOZXalG3nw6Oc/D+c6ag6N7
+Ibg1crN1+oZE3OfxjPNB+azXBz/kvKt7ZCnSzxc1LyjaC+bqf6bmfOPxKHJZca7y/cW1st/uy2X
xt1+m3gqvBfd95QtW/i/RjE2++QC0FylDwjIybFkycGEkT8P86j+TkhE2WdL5+Lm17Rz3UUZDAte
A4/olTxES4XPoG6w77GR8rBbdTGrLz+26Q0jNB7unOLjAI/N825fUaBxzCOxLlGnQRXgbMHXogWI
Ibs9et6CgfWuoHOgBVGhHNY2GOtb6/9a4Exl0BvqhNaQVr6qpN2tuo5HpacHMSDfQJUvTJsDqZ7P
mrt+MzCkJzezFAQbCg10g/MPWZs+v4PCtfbft1OGu5T6+JTLMjdkaGmseNLudC10aKViPHCS2hFZ
MDECbQ7NAZqy6BwDImEgPkyqXY/34tdjc5wakKFtN7jgm9ve92dH/SsEykKWLIyxX8EL0Tf8gRak
vsSVVR41KbqPrWWV5g+62hjxJrMKWBJlYPirzvn4CMD1we06VJa6do58Fj4bgpkaS+lKNZqgApae
cIIqljBICHzVINwvtm3xDuoMOcJLZGuRIt9ApxQS/wY+jV4s8EDyit6TcewE5jgbyy7fWdjBysXJ
nOY4/fpUJssRFygbinsvqj5p6Ctp5inQu+HahIFQ1SCf7izMMCg6m5h6hSu3/YDGalOHQomSC4PF
Ce+7GkUl4tq2dvR2pmgNcBqshLEMXfiNw/gKlFCNwYXBIdoLrArORYoUcgTxY6xh9hhbWAs9/qC3
vBG+TmavipCkZlqrpTNgA6clU7m4Ce+VNPoy0b7Sjd055nXR8RcwV0UmUVbG8h6cFGsUPFNzQ9Dz
63vBoXT2ZpAddAUQYjUxgCgms7rfo25Nl8UZN9QPngXjSgGZTx5Wf1zFrd4CFkIUrs5IacpF6OYu
8WmjPTZv5pmg7VUfm5EJMNQ1kqFxz+BZ5rCjGGEcyeDFvZb2GTJMyHY8z85QvtwiOUUocNp0+pgP
j7ibVX6uTiFWmJpnnZo78jIcxVZa0paCcY0gK/0gtMxubElAWdWEmgwpKG+Ng0KvxMivqn1qoZNi
yZI4XzKucC2jbLZnIJzjPfFP4XYD9bsbPW9RQOQKd8Sns2D9mAEWJ1TzQMFW2Pizm2nNH7piXxiL
WeEyVitrHuGDj1WUiVZiV7ulZ9r8NQttXLbeq4APfp/DbM+eyuSJu0VyRuR9vNuMdRqe6LIL9mNB
A/KSjCpd9+WccAh0MhxsBqUmE2Y3XPemGL6GorFSVad1PIIsC2I4tRs7hDVZckX9Yqhc/oxTIZsZ
bz8N5A4lVIBj6ZK+/Fbvs61cKkWvddwrLRNS1E7QUhTPwFUYiKZ+J2lded5IBlptxiVcdWNwi/bf
dGfbqey/hAhmsGstgRENhLraM92k8F4ZfOh2m+e9UmMR1j3/6PypzSNDFqNckxqEMXXaohBG/wzN
i11ldnpMQ8mxHgmxwQqmodBbDUlmwhJiElStREJJAqX5xh+Fx0fVxA9m76uUw8ErCcoJMDjahi40
orwAS5WdBcC6pM+IqXW5gUTsvapwySVjJ6j2c72wtf8y+ISyt0QDIePXZNMuJ+Kai0GBkXSAgCkb
6pRG9fyoMg0ew1R8+ERn53camF/MZFe4bae4yzGLrDVtlUss6dJK24FVondJy7KGaeOAh+VPo8O3
6UlWrUWGv9Ml+IRjVAZvneX7tYzxsW9f6h6wkMnMLrs+2reziCSm5oGf7FQPdV3veyd23qkhExc/
rTXRAVlbXys5S6R+6xEJWa6lo9KDb6BXcf8BekpdoFng3cuN/fVJadB/cl4VSIHuxVQu9oU1BvGq
18UilnTcJTcFnrCUkk2+eYUMACLr1KgI/saGcicWpBbUSM1rYSITX9W2+q/FH6wXmYN7P6w3V/vj
hike1mPFKr1IL7ukC/E9bthcEyBRKQwML7E/SB+8v80/X9GmcoRGr2ErLSQ0d4TTM4WdgAGaRKGG
oEN1iCu9iS3R0/HotjDEwAssVf8MBw3oVoxwWe+Ig0Wl5BBXd6sdg4ZHAxmjbZVvCatacDkPGZFc
/jPYCm3wa+sDqaNGZv9quTXCaCqGCDzuI8z+MRKqv34j+eqNmC2GcwyDCbqx06D74H7Roe0quoIO
EPU5pyPIRiV/GfuMg6ak6GZmAQ8QN8MrXks8hCj+escKx3ud7aS2xWbleytP00kY8GcMb8PwGy6d
r8ttotJPoJfBpLzniERpBz2INf8ghCPZcWmaCbp4wXdjV0g/ybydL62Zw82JPCVeWMS0NWcUNbma
owjZCo1rMzIr3ejOOfbt4uAHm439sj1jrlz7t66x0VJOVAjQ9/21kKFRu4pq61ox3pw13p9Uh0kD
M2/+tQJJHAwmq70wv56yV/HdNV9tcSDt1ABMUq7kavW01w4nBy+NA9BeHbzNODN0NO/VzmfMoKQT
eF5zqO7FslUVINK++ijTES2gCG9xAsb4+RCepO5IduyoupzeKguu86mWEkzou/9SCW0aF+ng7OxK
PwPQ94Ea2jARpOBCFi3dWh/7iMlkjsDwdmI32yxNCBEJfcre718VsoX3Ik6GWuVAyBa2cJ/jIoVW
uBkHffi8YjQ5Zmnop9X1g6MAnkhWJVuZ1cQKgZ/LLjhCE1ZmtMBHaEktg1bhvce6GN4PnbtB0pdH
1qAFqEPfO7erCYdaO1bcUqgCLLnoWnPBC4FAcfqQkerqsG0De21wiApcjpfgkilPOGqWDOyL7fLT
0PhYp5yZq+KlWhqgShMrn744St9hRydoIuEuQTU9k3RKVKL4ThPlx7oHeRf5YMsY5blnR+7Z5eVt
ifAFy0J/1+HDTAWpvPniE5kgWodeDTuxbLLY9Y2V7PCoBx1A2qJbEzEeBRW2GkMw577I2toKdj9T
uiC7QlEexmbiCdTuIQBxMXrgrdguFYtoZyCzMYcugqT/4smQbujIuYMFnRpAhQHt/SytPt7YJDl0
p9Dqbd1O8aszfL6UQmJjgENmL9Oyc4mrtXNnwIOAaxU5j1mP7ZpdNuH9S+Bvpjp3sMAcnefY3ytv
V1N2x6XADqbxkJUX43dw5sIiTAhOfPyTFbMl4hEg6G7ymxpDsLt/IAg5N9HUq+BuqzZsmkoUH+LQ
mWTheW/ju0jtci2o/WT0IB2kV2pXW38XbTH1kmgmN3tnP8FXZs+mN4c33FNlwi9afSewOU84VowF
b5YOQa63TBqfstkW3pFNta4Dt1VWcwTU6TmrewLETKnLVJl1FwUzxJ81e+Q5Kj/mgcKKSj1w4Nn9
joRT/4P6ScESaG+lK2O+FqqOu8RIm7CiR3tXpUgu/fESLPASizgUHimaYFgIo+7zPNSBt+mOs+rw
Itoc6ELE6FIxJLf5uG7ljnourjf8QWaGPAgOqGYSPkipMAabBsE6nc8nsDraPyjUUB7AqvAxbzkP
wjpTH6AA+uu9qJnc30GwxymnUfcCief9cM/pccANkhAbhQeFtTYrDNKyay/qkXy+9B0NLIUB8Q5D
Ak03ICy7DZc2BRr01XxR0hz1/mqVcekLAcCbPsBqBcRSLYqpnRoGbCQG1UAfp2ueMURXSWkmL7Lj
sgsJ4wmIX9Wr8v+A/40auTAryDmnJ+Q3sO/jrhTEImazwa2JTPfpTw88JqgCJPvi+/lFZqVt1GhQ
8su69DpyBq5jjBdpoL7ToeR66QLcp2ijPlE8pielCjpfGSS8JryraDN3mLdMInynhcjxnfQMlkUJ
8eCSG/35+kwJtZqlK7HL55GilnmxrOzS3Irc8TxkFDrlBZWsPK2wte//DtWwy2k9MspSBBEmU2u3
jVa3PnBbhZODFRwX/tCpO9Wm0mOrTo6pQvi4rFuKm3tVNuOlsY2t8yPyqJPBawjMCYAIx2xOiuva
2ewVS6TBDTsiliPG7zYL+1E7dp4CjVnaF2DzIiAFrdYQz0RJh6Rstsyb2WUXmFjkI4kTSgg9kOTh
EoX+Hg6880loJby7CBDKFLpF2mmx4FLr+Li4xLmj/86Lf5FqDaiA7+/uKCQcYYOU4WxtP8MDwouu
Z4blqm3BhGws2UlNqiWRGuAemtzUbag4bLGPbOkXjqKun7ZeeHL5bra5jboMQmEnPNr4gHUnPjTp
3C/XBF+DR9N37NrGNPhWt8fy9Es+8BTVqn/q8aQ6QsQmjY/3kUBXVlTO7Y8lWKrbDE2Mmmn4cHzz
rhLfyYbvPftY9tNgIoz9u9pLrYRPpqetgDhMtrkYcv/9YhEzKArHWLHC49FPvibmJvqFhZQlgX0q
40un/ZKyvsoutFlNoiznPh69Br+o3AQunZvUWF5UgUNbrT87yOCm1ZZmVwwXtzG+tmhcmzDygKlj
neYy4XJqE8MhcmEdvEY0LFLyTiErm2o5RpAsCZm8J2X/ohndcNuAXbD6aqKErZaHky794iO7YLDI
6J+jDY6awFOPy8AsTxVVbOpx94zFh43QGOLqT3Dy/xXnxqaeXKVejAWDnXgfXFL5LFseCOkh57jt
klh59yfiJDl+lY3KY5yJOYFVktaZojIhsUe461OhqOCjSZDJwcJmnkQQ0rCbVGTbzw9iyiR1dhFU
sa2kkg4GEPwmFTpFRIKhHv/dnHuE1Isc3/WtlpETbY4jLzZ5QbBPDvOHyLKYxLzOdDv7VkQGrrzG
VfeCL22zI4DSLRpIIfEORwl2OPVxjdgawWZslFhkt+zxqXaibHtssBOjNT6hr1Nmb/BOPpzOxGyb
nTolZs/ZIi2JqDYhzzJJz9p/HWXqZfZMTSvHX5xIXpNjWnbvs30BwtemuPIHNEdITYnRDo2I3yIm
2fpArSqqsi06AwIgBS6i7zYiRx0Aa9mCu8KGVfwhtdsJlZvb3gffeFIDxWaNFMyaMH6gI1X0BvqG
jYscUUY47YZK5NDJJQ2mX0WYK4o+QleKZQWsHlGwfR0pEv/1+9/qeYgp/dV/GAHV4gkwLZR3OMPB
cDYJeFUKFfa30/V5oxkgM1Iwkxfi8OW2uDnmB1xK7OkZfDM/pg+pDQja29iMQ2Tcfgk0N/+Qj7E+
1zRA1n7lFjp4sIo39IaELAdCjYGHcadhdhOcE0NHDrj98dsiWcbgXP9qLUFZMtHOM1B5NBLiCb48
7gxTzndAYkfY23RWBHy0CeVVTSNK/ygf64QSEg96oqpp6XQcvrkk987RCxyXKGsU4ZAyC8Itjk9p
UUxRJ3WZwaO0Xq3VqHE7FRkKi06NkM51HKuB1474vHUlIjdmNLucFVvQV6f7LgcyqLqLHN+I6xDw
ufAMVDP2TYhcUj0cPlKkAyy56VY0JBPoX4VYmcoETZAkPf8HZ3xejpjgUs7MOWcsdG5Z5UYes6Fw
V4d0PaZukmF0U1PXh1U/OGbRPpVKv0RG3KdHKdkveefkfJ3DRM37mUBaya57kzjk8GOt+282Vouz
yBnUGm2eWWqQmxkPGf3ccAMh65Cicxy087C4BRpTIryYUFLVQh0dUY0LxQbG7foI3XCMuFdyWFgd
IMKvcH/yxILzZRFm1IQqfcv8wNjjeeca7xJxAArZTcrRK8PfnOld/V8v1D+3YlT/KJzjo0W5XIZ2
N6TP1QNYNl33bniUgAQxE5lR8K+5CB8iWsFVvG146aZOjtzOHBgz489Hb0Rz4gbtRvLfM670B0we
pe74jG0OXICjWNym5cqHXoD1TKhTHqxc4M/YTPU5L93xQYHU7ABG9X9pMXAJbzOiNnfskPYrAS19
iCj0Uj2d4G1M9Yx52bGoWjQe+kH0lveVSEGIQHGBQy3gwGMzRIFsLMK4fQosrLMuAOICji/GXAdt
1cNbbsZgtrxhg9gmdzKEqFRIDWK4dAe57sldgRZ/TKa75z1ZcX8/DiK4siqLoYHot+/9SEegFF+r
Djv32zXSUnzCE6WvgR38suhmrNbLKfD0aMvBbOXvPWznsm3sAeqtT2PWbiIuKOOYQX4aYeixdQqy
CQix/IRFT60GjfEQuKAVjj+yzyy74gYCq5fvErg0jTNooWV6tLvjlHLBcS4peokJ+RTzSsEq59Wr
b+slY9Fy/yTHhu+e+KeehE86/yRQHgW7ex1n8rZ1LWo8khMZZ3StGUCnvFW+bkQvld6760zskWNs
5Tp5bF0XCic/oUVvwuSMWos74LY6lP0c4k++ls65lIw6i/OaRyG3ENehm9/1X8m1Niq0uVzQSAQl
ryAI8vlrJDxBUmsYKe43dh/lYHgR7Z7E677eEk+Ewy0LulEVzqwNmFSTmrehd6mgCNQWJNuwSCD8
s7Lowp+kPPKceS8uGnL9BI3p0CdTik6eD8FMy4JCFLcRf9/n3bLVmfXFhUQYTNaRdSxASgQKocS6
BrgZ0K0YEHFML/E4J5sim1MSxhlC6PeoeOR2Tq5erbIE78OSMAFFsYMjl7hl8kbFvdJvzb+W3aN+
ujBmZQiLN1gJVO+Z4nsrLd0VuHloDzTkRShIS6lY+5OyFlKJUrRJvQXUzFdy6amUVGL95e8x2dAY
q2dTkOlAVF6Mulb1dveYYAWYLQqDrp7QSIF5U8Ut3s73aBiNeDbbLILibIj199Nt95k2opUicQ0j
LDu4tU8YlnbQvLoG/PF/NF7SG+tGTbW1VihRjk7zIEPeLOABY3eQEtFcb1nC3UTXsQO8iU4QjfeM
6VeZwy5D/xUjkGdQtGtpwVFuuI+YW9kFAZ4lthmX/hW1MKfih3rbhqnyGjrA/z8XM03uVXTWEEPK
v9X68n+/RbdhGqiq9bhwERZ4eUfCYML7YHVb1x+6L3AQstldl/Eu7tiwYKWzB1D4ylmh1c51KNBr
Xl75Ui5Y3Mea0Bt/EDJCIIAHWtYHwqo05DQG83b6MAukpuoXGdZAt1ZZGaVv4fAXo4J4y65j8883
m9Ia/G84z2a5b08rLSFfFDnVuYFQUkfXmie0BS1bDOjUDHum5bXhHEDGg91tEBem87wc4nBczsu6
tx6n2YMKtUALdeOKcDBp9KxxZWGRe3AYNSVIA7joPji2vX+WjgeSLp4K/VwRHEBbq6nv7Gn4wCTx
G4Ai8q3tn6YN47es4oy06/iFDN09GY3pvHSrmGg3M/AQv8xp33vgkf8dsLPNCeL7+qIMwiuyAuIl
bOajE9bmMLbc7zWJ0W/Z/BJ84t6dtMCL3s7YHLqMTbVohHZkbFvShs3xRT5LJCyZ1WffyheY/nah
xgxPtqsOcpINGh9B2dmEiWLuJg7zln/NchZ6jlw7W809n5D/KA0DrAXzCOFNyEKCTljSzRmnzBi9
UFhBNVbuS1i52VBSc2inX7jXdiyn2VE7WeJ/RepeW6i7XUcvtpO2OAcCZcdgFSrg4NMTpGuHP0eE
oGWUqK6InM14738p4R71lGq+kl1jsLNXAOZU5vruGL1D0PP8Q031ofBRUiHPmcI+06PVTGGc1zK3
TViale9BazRVhmSmPTlcygYno2haO57VZCkANuwezQj/H7jarXkHKtThQq9y8rqZoMPU8gTBQaD+
CLgLoPQE5qKQNM7w0hYGQs0+glbIpKzW23mDh6JC65ckga5bAprGycRo9D0y2n14k/UvlyIxyjdF
iGiCOKphup6CTYEN1sYSmLmQ4/EugG27gXj2ypT2BjeoKphbpxEHxAXI6TcO/j2EsxwiLaa3K2fR
8fEnQiTFvASwV8Bdfc0g9LV4VYurMZ8j7pZgX5Z0K/nLSS8QL0JUCJMpcnd0hd5cXTi8MjxqseqG
ob6nVoqAxkXj+NQ4r2+gufjmEoY64w87AIXJyE1WAr8e43sbeQ0Hx5hNLH1ghDrRKMG4NZwTjsXP
1uEfPhxRQzP3l3Lc4WrzG6n6U83wqMmF0EIeqY4nqop2kREoPzlMa7kiCoutYQuOZIjKO3D8Sr6A
I4Uw743lYOXxBNMoo00WjCcpRzKl1uQ4ujQcGkxh/2VL55vyMlISQBox4kVmzL7QKoJjcdXmZ4b0
imCj9MxxmB9Q1kWVQXcBn/dbFTp0J4EeF2Hq4jLYgwUlsV+6j3eu95tvLOX0FKrB7hMhUDF0rDyM
R9ehYclylVySiQ3lBWDWlsG32P6r6U5Ww13z0gvLblSJkC2mEs31yvz3g6BN56CLtV0D+yg+JJue
e20bRWs7Mv5gedJ8cr4YwZqH58l1GfThUc2Blbc8cYNSB+coUX1Kwbozni+XJD8xcDcGvs0534Ms
T4z1T3xij2FZLmkvoqxzUD4pkuFxJmfum+mnJOVXJ6OjLjYTWptvNEg4UWN4AdwDWMIiTSqNraxz
rXFJe4wXU5potWhNYHkn2O7GrBBMzsqSSVJwXFAjTGroGrVj5tjQtJFE0TMpREEtrhdvs0wMh53Y
13rNIWYJxyHK0l48jszcXJs32c84/T8t7x8t6ZmOox0opMrxyTq5snSWb6e8i971qHCPuZ1YhyBc
ZTNDTxG2G2O8IGwZViY8x5ziSFBqjQSmjktm1kb5DXgHkemC+Dsvv8H76/HolXVJfDTh9ueaCH1b
2YwMWcU80viRJ3cZbY2pEFfcyUQ/nQEBLNJQxUa/WrGu6oWLOjY28EmsLgQDGSCOzdAP9LQUtCMk
QkQN7jV5XIOzM2h6iNe5Dlh/Uqv3TWQX8K8CudFv4QDTqIh8G83oQNXS2IdeSX2VL1lo3WaC00hW
TEnsU1MUywiKQ7OHYcejljNnQCH7gzjulPohwJ2yeXUmylyiB/A+vpCmt+3gLT7YlTVuF4Rdic9+
Ud3nqjEQKD0qR6sFTHhIVEI7eZ2+dw6W0sx0kscpKBFPZaDxtWFGZrZI02HkXayUa/8Mm8lQF9Wy
Ogsdq4S2GUM82mYrOLjpruRXHExmZPqoG7XT3g0YyeFYhOmuJpWvr7aSESEYbm8da6n7PTST/YWK
XUrPd6xEqH/ESJz5v3WVkCN92KP1hFRGb9GRH1ir6mS36uw8hjP51nIjOlKA95+6cvNTjdvGcK2y
Q7gbyWBBTGLt53yC/6kVIBW7up8gZCnFVxo/GmKD1jVT2P0kown9Q7WX9pcFLLJY6g52poIbomgm
fbbVok9P2ynxy1fNsRrsvYVTFW1c4gZ8AzwpJuV3hcXyC45hiWmGOidgN3+2h24vZv38dXeeUlQ/
SOL7fugj/lgWqxRYGvZtK/dOkNOBejb/W7Y/bk57RQBN6ag6kjcJfwnqfgY+kaAEJHgd7Az2hlWl
8cZ502PIEr7z6NKuQJ2oTP1OoHCjPvxsOmaG0xXznSyibu+uKgsQlxvdYdgaqlr/WYhHUA06Vsfk
Lo/YvbxJRBwFTlIZbkSsyZct06CcVqyBejJKR9hvY4KaR62FaYJ+sMPgPnyJFXXeUJDDbSRGajBp
A+a/ziMvz0mASUlXo9jM6ISRv1ykKJgimJJPhERqlP2JyWE2BOiTDg+AYSWoOBfb0p0GNKSp9eGj
7+ds3C9navknSATpFnCiZqsTxdc0ZWvkOOnupHFp8/vT7f05d8g6UDA0UOchU5jqP2iBt9ygCBqo
ZhdwD1/YnMc5npuMR3P2DLroDMBWHMKH+yDXttJx7JoMVOOWRfF1JQZOfAnrq1PA1nQi7C55nXNu
RW6Y8VVrShYPMVOeriih3Esr33ICBasnbtUgdIQMHMU6yJsTYERpBIOibuqapvvkmiI/PSCzpTHp
b+gH+l8256YoVMM3S3oJZmTbT4zJF+HIWLblkwWSarAf8Aan9VF7gZZQVm7V9Kn9xciTCrvai1mm
Sp4YSuihWLKjYf9LGojxy0ymL43IULlb+foD/hstdwpyFkjvz5mSqo0noZTXQqIpPFkmYKbudK5H
BpxKLBBE8RYOWJVur1b8V0U3hQ/+OBEhbw3IkrpxUia6xw2XWebBpu5/EZWgI7fpay6eD8s+hJ2X
2m49i8kpdWMdu5YNK1y9vGF8g0VjYDVajBY5xn8IFFu/+pslr5rslnYNUw63VYYfIWBqn8jYmi7J
9TUKpo6XzHoVylaBfoN3yZ6c4R3HJ1BvAuVonk2PHQ2By1STEf3qB1DcWMO40r/prQ+Y3vdofHBF
w/CMHS1FdPAavWD1zeOQNz8fkty0KhnU8sONK53kPX/Ce5Z4Jmu/Txc/1feLcYBQJAgPPNTJYJcm
yRm2OK/bFLkXGpya3af8zjgqm3QZWVy0kPZrqJOcrQ14rPfX374isUmU1E5s8Hh84Hgu4mP1K701
YZ2XWsVSIieZWQpFsT//+tD/vq76ako0TXlwkp7QbyioP5nOaniBAWrY0wyHx1m/ZpaimnMzRW+G
E6Mo1b6R/5lyvrrHP3Bnor2KlnwOMLCWuJdwVZ5NTa1/IH8B8RXTvZ52otCxNXWPFHK3gvbA+5Bb
X6pO/eb+wjV5MalHYXqzzRj+PjEKu53CzuGkaKQsmeAE0Y1bZefqtscyolQszzu0V+c+JGaFbbXA
cO7ZxWGBpUjdOpBHA0rsfC/TFUD99UsmRsUkVSLWoFJ5KvZIq6UDOA5RV7gOH2wNVse9/3p80Kb8
9mS6fTHm4YryDPxvKAS2LT86wQTsrhhRTlHsiXe/bnIn4o4VhLt+byCh0CegxccLNakYqVikPk3u
tr07g0L0AAfpQn8GHL06Say211pYIXhWxwf0oHrKkPKXF+Lmmp+AUbqObmmBgOrQC4qfhwV7YVqD
RWvgIMdozWfN1kTVYUHWPpL5B2W8nUrMvDh5AXZ8LeqGcUtr4jaCQPsFxDWXx3knY3POxwnwdDbT
KVue3v1edPVx2V/j3CDWf5v7H64maFa73bXF6QUPyQtDqg85KNKEepxJnjgsMECrNj+X9M1tL5FL
loevVbyZO7f/+FLR9tflkE15KObgx7Hqbw30+C4g/HGHyfuSCO6t9Zg+y3YfMe/OBMKY/+ZuWZTm
HiBJ4y4zeJ2PFVxRnoHgaC2FeeZ8RZt/ICEf2NY+OyWz5pI5pLNXck/XNNnmGzknFTfmGOmxU8fL
gi6b8ldkpPvqhIhjag8ShVSsUF3E3mbxxQtRaJqBJeR4mPpyLeT0+TmD9oRVpfBHdbl2bPa7DbWz
xWhTtnNG207fjZAiZ6ZD1Vg0ToUpPj21yW/WQ+5HtnftJKoiqnTdN5UirJyoHmcKIX5RqL0Mq7a/
4fLfMy0NbWiTxhrbpV7ro4h4EX/mpPyE6QMZ/yI7SOTclSu9FL7S2C+LS40sdJZ88zBUbqFLKLLS
DwtNbldMQnXfXP463Ok94qj0aL7nRl5EfrBChgrElIhWFslG4vFLCGL4MGn5nQfSPxCXKVQpcEiT
gIj7aMVUevIeOgiesNb9mpHtsDRdfqmyp9mstHubYLSC8GxZYbK4EF0FTwqYHy/J6M4EKgCOe4Xh
OIu86GPIRap4FkrHWRKlhfgkiSrzGkZA7xIMURXrz+MinTE/uQSCKFFizvI9wjNzVg2sBrXpri3k
aS6GD5XnC7CBNS6r78h08AV44OrZjJx9GuHIb7K31uDBPACjLl56FfUaIR2osUOzLqY7CKkzwY28
i+moD6c5Jc7doezcKHp9tObWg9b6jJFB25Gn9AxULTJ25RX7mJiY022hqRwXTTexUiQ+ps5o3jlP
O4TXs0wqzuZYC2Z4fiVB/CMeDwH14BCPV+iF24DZG+I3ag6dqzHKJqAItOVicvHUgBgSaj9v5piK
f/9E+ScBh0bj7o31KoR+wbe6CvrXpXkCzCSsEJwbbEVYsgQVvog9T0Am5hybq9KLRjUETTElO9dh
oIoZ4rno4dAchD9Tn5YYOjyLnCe31JcYmqPx+ZUry1Snq1g9jLRDQE4XKpv7mdDHV7+cf2uHUICs
zzTPcxWdka4mbzaSxweRPhZgRfT94W7f8SgGXkrDmDFRZUTteBkPLSQvwvwJA3s8T4rvjFehOjVr
NnouIgH/SA8NP8/cSnwneKuEaXo9NIJKy+49kOzBgmppgPg4t/e+x0frrO6g3LQeAdvbVcGvwZrr
ARAZgKc3hRzFsCtrMIXDyoDZrbEH8Hcrc1q6H93m7lpUwSqISNsb9TOkInUX6oLfw+UsqBEGU20t
ifNPSI9NtskvcXmTjb7QxqZEsUIjAvlcSrHAk3qcgLaroPq/za/8d0AlcbIT+7H7De5tCS+mZzfe
ePvIzIpc2dd/AtjJLxDr7TA7jen8vE3mWJjXzRsItQBZweC/vIdK19vUXgNxLmfeaBmHbsZ7GwqK
0DHAbzNMrUgXxy8WgKiPcItBhHT4maJUTcopoBxpE2Z8AcVB18CPKrgyaZAoEQattDhIxoL/SRz2
a35VNGH28CURpLgLcP7JDxVC3B5ICYW2DBg+0gM9Gwddb9YGKDuSp4BGOdKKXMZYPqDR6CPl3Yb6
J+79U5Dd0fvM8pQiPtAAaPK8P5vQniFlKvdYMq1zGKmI549xhbDMJzd3G492rJWl/P6Hq8rkYCFO
sY5cNkN6aYIlT0viOzZ5Uefy3XyWEwrIOJXblOdGNMzCjybWVOohFS/PhGNpgFptda9lDPdED0fQ
llMtLOc+To3j3Wt/UKR8qK4GQMlotwasnufqhhZHwnWIt6LRO4ZtgR89ANxOcJ1v9uBHCvE6Yxlr
Bt5UwK6kSQOvDBsXHy5cWwWV6qSaLVyK6/7yv3Rtq7lYQ2XN9bT0Ejd5pyT6HQ2I9+Z5N0u+p3Dx
3RE2O0gxSRgGKnIuqmDoZNMeE+qfvW8/EkBFLKOZA3PM1/A0ZxTB3cAmhRjwT1YefL99SwqLLBJ+
ePztrYZsnlHhfJBaee2i1W7wfJeERrGlXrXO9id0ZpdUTjQg2L/NTg8sJWoxpygJAUX69DLqlG8x
OBmmwMHcH2sDa3tMVI8NRWcQcEnXTfdmWiPhyke2ms7GuTNqkxyjIHEA5SGJVjIYTOTdYvdzl54T
ottWY3fRqFUydJM4hndD6Ir/fYqOUhj+xjHpqRQ4vHCHkB5yz/6cp0Xc4Om7SiM1a2aRfrRSnvIo
0RxRxyhUrftU4J7oU2K2NomA92lieMqaw/wDQPDOyQbIcmLhJVmWvq4YrlVEpzJsytdNlwc4L1tt
x7EowMv06F6BkAZYLpYCEcqg6toN9I5GJq2SARmNSwtTbNgSM3Xfsonj6yN/HBYvwuZDyqrxo7is
AhBJQX7f5O0ZZ1a3Nn1Or8K6kMqu7Hjo6mmf4zJdH+94S0Ivid0k6jCV26V/OSPilF/xESytoaqe
2/0/wygD5cDfhSs/yW7blPeY0KxFo6f459Vv3UHF12b6HDsnzNrNgWp4KLpaUoQuHykExGlw7mZG
llYgIQvij2ITXXZv48OptzqVUR7mpOLjDcZvBPodHCLZBgliDD1/rTJggPQIKPoVhBtXZHB3anaX
ZPd1RNuH0jqT8t33mFPGXEbrX8GBmhPUn4uEkvumRUG2LNrIiV5+95UANGA0OZuK97d9M+8kybri
Za0m342nrL3dNu2Gy1K+QOCeasLnx6jjhuvp4fgIqMKpJbGNMI4tRCOjqHo/PegXybXMh2wiOLUy
2p4TPLnxDEmvhj2SchGCsl8CxuGNf71yNvTeUMdWzjLbHMbtS2maXUgVkIwCcm53AqsK7b25D95d
AbhPZGv9SbOo7OyjCN2NXtAYGeKiQ8C/KCo54yfbdP1KS4VlPw5dMW89j6e5o07TZ63+26UpUsRs
W7u9RtryDgPa71AFDS/pY4uS8bgixxBAEGxoq4depRs586Q17qsRH2/KMIo15G994UdBOFau1rjO
yE5svTCLoAFLFxiW+gl1FJSeUVHsljCS/Fi7bxVVHznZRyewCEps64eHczCTG2MaZJQCEdSaAGsG
fMwfAGhQnUOGGWAKyrCmNW+IvVaqchAmhWKDXW0Lo4COv6/IuLf2kef4hYCoIVvz3RV7D+ik7ICX
eYMHCnV8xpJqRX0Bq+5/1VO+5o8zDki8hcSGbfXoEPpbp5EhgnkYeSPk3KQ47XwVksfVK5nbswRz
rRinq2lsjSj8s1FR/wwlUKSJsv3LR7uvDL9oyEOLjBpIHeSVj9zdsE2U9pIDW4thluQNlmGsn27h
u7UnAaFwenWbLqC1QShjC4L3Pa5Y/bOB7YYibv6/BCRhre3zTBUlG92sG9rW4SLIhj/BFzHw3xVa
Y6HuFmLFMkS1SYVmscuZ1RaOrHKgzOteXkKCsukehdi14MC4nM879XiA1tksBSkG3VBiLaXMTzxc
3QtTipOaDB9M/kssWKuIp84GDacZsX+7t41TxO+CqFlZn+yVDwU3bX04QlDzb0LewLc/bbLELwaQ
m7u6TrclHE6Q91HUVoh/KjouMLLbENwO6nQoybgrgBFhTzJQfI2db3a0JXFLHLWVwxDCmqqWTeum
gdTpHn+wilIC0BEHZglw7CDIr3DQFJOubiFQ9N1NcbOSBlW84G202+GWViHJdiWPHfBIVFfbNGt5
9VEVcXLpRVxuYiWyuxwWGJlLs2Z3kmI8qnzue1hqd2MBe7aWx5xNMGyytgrSn/fXk9RK5yYq0RC5
T6Tq1wULp1moa2VpW2ypCwtfLYh+UGEf/keCDetR7gB2t9KxRv6bOOksq5s8g3jcFjBhXGTn+UBY
rGcniAbSWyNqhnu9hjPUQITG+8sNIl2LIsI9CQPOU+xRVTxDQmpdfcq89HLhHQSxkceDIlw0znug
Fb2YzXiNHkB4I9jYqWYFIHYXAiulXbrA1Fc+2Xw+acwGYJ8b0sNAeUcIbNVRtHydPl7xUmjUFlIt
assv9j6iSs3LPpJdV8vmX76ddLiB89k7Yb+/DsUrZ4V0WxtPpDxYTCX02/eVp+HlC+d0PighozlA
vUQmAPN+wJ5i3aK4lb2W0kKB1UN5/9Nh2GDjHsQKkwQhhIrDfnJhfbk+YfwI+j5zPekT+rnuBCwK
/0jd6iSGvIORYTPEUwrcXHrCIhadPSSQD41Dc6Geiv7M/VEPmNUTjLP6E0sQW0iVY4GNyMMmvEjj
oHL1DuNtk51Ex/gBi8tNLepng1PtQNkMy22Aqi7UYYWoDiroX3QpVG2iaL0ERAxLZAwiwmQFIwgR
pFak72pB1zXKSSLHRJ/E2QH+rELcOE0fJLAZkdT/IDfJr4qxWtUH/S9VGecTImQQWhU4ThvNi/fe
Ohm9F/C7+to982QYW152OE4KbTobKmza2f+qI1Vv5wMCZ0l/Pzo0dpSfoK9aM72QP/UBznAqZLIv
qYfQr+ubEc0tPVQUauPXBxMf4ftt/SwXWKpmK088kyp0tHkL9GHQRkTk9wkdCjOxxWIUq6f5SoCr
iz+zy2vMtieMtGc2aojRnSAjG6tpg4FHfCUplmRfaPJrk8/WumWpEGPA+1YcEq6n0vL3aZqcgA0O
TAx9p7hncJcHE9vicHixxLmoQMlXnKA+3UrUuAXxvI8Rsy9cyuuATKs7wbeCcKdPOpEMpus7J6OB
aGJ+nm/IL+IMeYOGJ/T4HvDAw/Q0nhzNMVNnCbLnSAvoj5KslL2+d2HP7ZLk7LUiS4ElSEQUCm6v
kWLuUtMEBDspD+n+YV5mECw1GrpwZOEU/2v6GpbKGcUVHPfuaIgyHxmFypw9w2MCju5X7pjJG9Dv
uVcU5cdKYaapBZgjaQTeISldU3TrOgtQxs8MERMF1/qzPGovHRGxyZlP4auGN2g+gF8+NW2rQUfm
nWXmiuZ+xVuaMdvSOH0F9TK48WpczKRpM2XB/wQr054cR3Gh0UIJnUicrqAdChj9/Vp0ZOWOep5s
c4XPnXWHu0ZiYqSPfB+rMH83D5AYPQKmV2gcj62yFCqRsCd6vjny0IS2HrthdbD3eRoki+N1pCZ4
nFD6sW1bVIYzC6PlaJ6mqH8rEsLjOgPjE2DnNWbTELyS7JlFIh9QgUvHP7Zv58rlQSzbuORIrVy3
8cRvPQmVs0taX2M63xxwgCgXzCHpSxuolzDkY2up09f4zUxBmil2JMpYTKulooP36chczOQwgnnH
XLcbXgO7Z9MadIijWIo/iwbP1gbPTgGPFvGUezjiuyDpNvA1u/uFAImSU7MM+2bff3Upfzacg2YT
QgwZv0aA9OUrURqwXsLKYpCK4FJAZFoFZueDABkDUl73KjXgdW/8P5BR2NGT0Pgx9OtlT+cUMqZ8
COvdbEL8itlF3hKFtzsHTszhycGCewqe4XJwbcuCn2BJb8NVzV7/i0p3cVN8Lyr3V/JsYCTxwSE2
RExWz5BVYtoRhd72qixd8utuMJr8EsYDr5r21u9y/RKCJ5jmMZ0srM2bLTHHeipmmD/cWcXYEi14
vvC+o7GXRvMHpl+smahF32ypXXaDYLLMwVxmPsKRQqPcT+cLtWY/FZsecnmaNhPMSNivXPxSeeDW
VmcqQv36cjMI8r1ntbfxotiUQdgi+9vspsktKY91p/C8KaQsT7yVJskTT0jsfWgSTOtI5lwskT/+
mS+Icnn6VTia4skJ1S5gXm2Lb++8UXJsQTl77tFxHlDKLyOrdYhcOZsHonAA5UPJ3JINT4N9onFr
z48BlULlwtpv3eKcdTTUuqfi1zejxmBU/HIolTYiZNXzaTN3c2SQgyIoTYj9Gz+G/7Ot61RA7ICH
Cp1/N0C3z2HOY9pJLMzyj74GRlrIAyx6Krk6U5Uon1pLPrqZGsZGl8z0jCLpYsWtG88KvTXfleN/
xgqd27fBBxhMCHreZdwT9eJUDnNBAnVvh9shSB44qoJb/F1+q+PFevL/J2Y0uHKNmrffbpojHl+y
R94+mtFF3EkqYdpzg6nLMhd+sx6TWmErxKog5qQKk67DZgbRptSffSB3tvv7jgCxJBTl5rgOk4uO
QMtXcVAn0OGtfOncC4KRxifY6xYTRrXNyW7NkyO8etpzlIai7mit5peSafDX/S9JKMYj5DEIp0Zu
o3fiP1sa1waKf0YAismI7dayKODuSz2W030H3gF3ZfjRCFk/wW8NWBGVYWatF/VHX9YWILlJPb2N
Lg2mgRwum8TKXnhc0H6qZWBWrN1lWxK5l4aOztFmjeeP0zFmNmyWxCcSJr1tR8f6ltqeG0h4pM/x
pZlKgTUnugjy2pPpSerPqXCNnW5BaOd1f3cGHKBuyaKQJNk6v1SW2jZ6CLwkWnX4UDi1E6SDJx2D
HSztCfVwV15lOENqisjVLTeCBl2XmS+/rgOSfrhfLbMWkc6XvCJ04duS1Tn9OqSMbBtHy/R+36F0
7kPHtCW49QS8FbYKJRVxswhLT53mzxk4MJL+kD0rwCxS1aNSrvXXXZc44WwRfh45TPQO49L5BIm7
2diDW0cPQV0XSlnLUKy4TGoiWydHnK9bbV/v50cJ/8Ll2jiCsg4Ut693L/NBHQ3bKk2QX/mdl2yU
blvQxSs7ocw9QCBGGExC4NRwdzS93z6e0mwRgEqE8nMO1RM6REA7GHJx3bhyLPbBHP9ETSXrL7q8
z8B5EGSQJue6wYJH0T4I81t6wBr/ZBZpxDGfRRzQh1r7teW08HKTJO2YyTxoh0MihBU+pH1nIheS
fivBUm6pj0AqicrDOHYfXGsT3pIxZEbQWuGcHQCbjfwhwlSYz8IZopES9cB3Ud7VSmshPqd4KeDu
EdavbAQ8jrfet+xwFjxE6GSie6FLgt5tMKpviUmHX5ZhNjAB2i3IZ+NrPB8HezrEPrAmsW2vi8C3
oAuROhZw47lIp6LO/viS3aeTAal4C3SbomwyC+Mo2v8CSIsIOBqWDEzRX8rg1DEe5GdyLfs/nNK1
O/8r7mVlk7TiYOWI1aCP6xlCXVkFEHG0L5d8DA/ofACnj2NXgUfVAf2FPWvHYA8iFQPAhE2pjV6x
e4RpTSaOQ1LqJi03lIvfK9wt3F7u8PO0FMcjOIakNojh5ITKgi0SZnOhE1pkR4mFWJcCEyOzsiJs
+zuqddTFVZP3RrBX38KN8mbyI8nc4u763hSs6bBNlEJt2PicKAN0OY23EY/h1vOrydTghxue73yh
xMwYBXwbdM9l1qNP5lJPq63gdrQgDyHgpFDc4ltnkaN6MZtCWei0Eba/bwkgwajBIsoZ0Y/XAVQE
/jeqsTN8/jptpJlo3wmxKeUzuNsP4Lg0+3miaumit7BpjopwlNwNptJXT6WZUNhkt+q3LtqvXwu0
HYe+AFh+hdjyyf23HKl1VXCUS9/MOKwOFsHOwATBxVDEzyzWfoOprtRqz/23Ayd3CBo0q2FLdf0k
qvuhz9PZFceSzHW9++wbZOWfXtDgClhc5dqgHpbvGLiktMqTd2eJ2xYwEuG+uh6HlVcokf+hOIDa
wBxh3++XJWoWuxN5OFJU0+oLrkFpI1qVcFvE1KSklbqOEXQC7/hscaF4v6hPol7LKCHMK+y9h+6q
pOeTV3bNhxicm9GKyzDifiWVrcmQ8Tcxs3mZYvsLLC/Tl+PS5PQQNm34+MACfrQeTBBbqKdkmpAv
DDzTA0Ez8AAd346Blf5GiX+RxJ1ftR1Qe3rgF6X4DeZg+sZwfGshFg5aMfl8uIWgA2fyHRfy2EJX
38on3DKFv8gsgsn0euvsAr215jMmnWPqDYk1zw/vYgmGikCfNQhavvaela/BfLwsguEgNLxfq7ho
YGAz+YfDN/rVIs7QjpmI4IRp7TcocKWqbAWDqYimWuzngXCH74YB0GWRr5lEDVMGl/ub2rEt8qlS
tB61/PjDXsTZLsuj7EipAaj28WULvIPaXLSO7woaLU37ebHcXoX0cT6g2i8Xl9gWcnENB1/1IKgw
xTM2P/PFtQ5fyShevCuMUwkLBMkovQWnYS/6OA4xvss4cLcOneDj1rY5UZMSsAaFo21XJWN8eV20
Z1nEQY2oSVWlcOH1UowAPV99Kw09k+F45icWuo48YMtWAmNpxvAwzHIyKTyOiT2Xa+H4YJUGXnM2
nlckfjvLSO1ck1iJ4O//cTb5Ha0qqd8zgN8riRUWtw8K3Zwd9StMvse4NTdweZuLkn8wiWEzsnVK
7FU+Onj0rB+blq5nfIOXPENifuOZoEDf8EqCn8aobWT3eqb231NrsO+sqbDjcZUeYeTXTStr4cDT
pIypm50L1XhV/FNeXX0777w8ofTWOvRUmteOc+W3rMoMTyYBb7CWX5CoC8vS2cepDS6x8MMMCpRR
fZXMMfNoMQLbG1Yc56wXPsLXGy8cYQIEkH4/W8q2LjB56ZhOOs+oPio6UL6JZcbQTm5NCrbcjfXF
pnB5eLNx8tcHYS3HHbJ4C/TA+lbWAqcpLpmaFeXwxpg7Qo7nzbjCLd1vOusImMxbV0YwSaeFiZ/w
C4RQ7R062tC5LGNglVn0piy/lnl4/PXbcNp4mrTq7PmF9cMb7ZVLi7WzEoW63YLQBz5dX+fNV2SL
418hcI4ajY+IDUMXMOTe1JwAA/VblEcgzoLAfl3Rgjg7C/864gZYbjJx+N99JdjCfZ73ihpx0gKn
uZ0v4A9P/FF8R9YYvsHhVlkDxKdkNCqTY4scJ/CoGpbTWxL5PiJFV6w4W3MyIe86bVLM2PbTS/3V
qQ54jpZcG/5aZCT15b2zefWWGX9NpE/tbvQsJJoj7ujcFE5VjUCU5f03bXs6MprHPgcSztA6C5ZU
c0LILoVoAPI1fc7Bnd8qWkCJ1FMvfKXn0mdljiofSsDq/X9qFkvarU/2gVeolmiB39P0fX8zS6aK
/76gxl31RY8A7c0NWqqM41pnkkJLHCrw6BlL7O7/ibuTB4AynnC6tXgKMyyxt+7yo9bRNub2UVrz
zcjFtHKDLccryAgbevDC/knNKd11gFc+HTSncsuNvTPOtau/LEPZIWZaZaA3CRgJ5sjml+Kbfron
b0dhrbAMQ5u788Xu0mlTCqlLmxpZCMb/5DXLwLCwEfZD7uhfAqJRsy7eMpUUIlw7j/yhla4+0RXs
gt6gPM8jAl7/MB4KY+F5yT90xEEmDiyj5i7qtKgww7XKhRonPdBQvx0LDtTx8aviwRbdI/Yfgyoj
JJl+/YXgHSHa7K5FtI00+F/KsDJ5w9EC4sva5u3F1VqYWLQLAz8tngPEkGFsO6QpSp0qRZIDWnS7
oTO90r/PkmBG1kjC2poc4YBuFbMaf8Zek8RBum1AZAA9wUZfBxwv8AME0ZYsERQWONnevNrzydyI
vJoYrmUbo6Iw7MrAwjxSwYRGQDNHbRP+nqlGHLunjgUON/u4ud297+hXdBOHDxwsUQMjdawAA+RV
kLoBJopwAdVvTE3LD+j9wOh5uejnwQ8yr6NwCbjsjSvKCfj5pJcwEl2ACD3dzd2dzdsA8V1GlZCb
r/Cd1fBVIZLboVrX4m8n9p92vyEA96gCnCOskHz0p5TiMKE0AecBpQrN/ozhbFLPXk0n37lbayp9
fOolAD6pAJ6r2UueZiJ/LcgJiSqcfATV0otMCyasKgJJ9GQOhRbWHSjx/8LUoAbOmADDfnzc0Hn9
iigGYJ521ilhpEn8yRNoSQrMSmnp6hCP2cDvnKXCWhFjVWm1L754VbLwUCWWLNcdU5bHMyu0hhiD
AcFKzwbN5Q4e2lWeAIf+opEz0g/FdknbLsFqGRbgVEJNBPSjXPEI2HPfyxncOgPmhbJgPn046WBM
0d9y8RBdDJ8BUy+A1a7DwIhmXRUZQgL1ejI1Y+LvV6s73ZlO+li3VZAjoUYDe87GRYWavP/vedhP
3IJ09iMs4enxVIb2N+5UHUoF86dzuwgg8myjZfq1gllE6o/G5LaXeAdDHwwfB1qG9SDsxWL06ACZ
JWYAfbe+YiNWh+2k7cFQow76egr1IyaVsBdk5Yr3fcHgMKOgladVpqy60S4N7dYaagR+lwDRtTSP
hnvw2fV2tYo3VgZLu7Umvpkdb4KdhRW3RDbRpZ2YjJNSSISGbjI6DagYkbGRB01wFcY38RFdHc3A
+PBpkdQ7pMDEPN3+6oYbyNcMxNPy9JA5Or+XMHnAVFlMQ2Wg9MBNzu6VaQL5xIjJYP2o/WoKEuZK
r1890VF6O1RNUWz/3k2e8TZSO7DoX9xiHdN9bC/dv1qhAXMqDTBIdhZ9MYy4MgnrEs67Gjh55T69
PI/RXfymOT+tQxtShjSJ1a1SNImIgULkIN5u4O1xLIF9GcYYR8k0Ls0qaQ/mharEqcthIitsExPC
GO2eoUkI11U5uaar20FhRzuYJ7RHLb0zKCK8oRjUENh9B69Xb/94jnQvAYSbLSn50/mR65P9BxOZ
irZI4LiR627lItkXBmMC+tr4WSEQl9YHOX+8etFBazh0Cyxe+ubXkruY+Ma08Mv5WfEU956qrzEo
PPqz0EuLkRWz9lJO+qR1YErbFmcCwUT3Psn+Sc9OJzJix0pwDiTsMG9Vx8OueMBYP5FCKvLSm4Gh
A932JN/Uva08S2iEcF5zlOKqy5euE6WWy8G1pE1OL7RfMgA0wbLQqnAomBhIc8v/GGALQ6BICwPr
WciEr0Wisx+DEqXSqlokFNdpOHayMAIcJCcYqNcaqh1kiMCQDABRwzbvhsy7eFilwrin0tst28Uc
hWhnqy+Y3Q3FLtUga9IcMuekxwj8MzWDgjGJUxdBXYR27TIxYwxij15/ae+9s9H3IxdhIyoKqlBQ
kCTdpWoioUzJAS+I68DaM1ilYnTug1mO7RiOdN7+msrywkbQxVGGBWGvhuQQIIT31xLr82LYQR0W
cD9YCZcPVOs0PvqT6VvBBR0k8uaBoMZ9u4IxC5c/aSw1QSd47gF/H9yiRB+4Qn8M1bDZHtuL2ypw
w3Tuq5/dxMdTPGUmpvDJJT05+IIAtHHUb4msemlSyNmYd3avqhk8KBwW8GyZwFgMqsK4r/gfjsQX
CNT0hf/sQ+QIGixdpgza7E0aM+PJSRDJf07+D9CvLTlLGP/YGEHNR9q6Jnvj6v3HipHmoSA/7cSx
f1kj64TpYG9FdbeyUH60HnsXwaBRUNs4vyV5DvM/rVNydHYQuEgbqce/iAbewkbpsJ1TnFHCsCK5
pC9m85BPBwSY9enoXsewnh5cMJD41tf8JgTm3ldIgDNwgdsC4bdsm0kX7IlVobTcGWSnnR2MTG1S
/w0rYQcLO2kJwXO3BtmMfLeWsSQ8cU8+s8ez4RBRouZBv6utQmyiFVKVDLBmMwhN8weiDhWrDX8W
WrPrJG1YUm2Pl+WN5HgZipDqi3HOy57TbiprlFRQdDAPDGQZL+RrBiChRjBN1NeCOQKL2xiM80gg
J2kqA0tqKRHvDpjBh1UWFXwOLh35HyJuXo77/TNKCnuyWTlxJUKJf0He57/T450uMm3G03TMf58B
qoXeov+ItbZqYH3Mo0nbaefgiGyDDQXN81AWzEyo/I23m2Gos5IppFea+iDPjA7BVUlA65zMAtnl
3yw84vz77FxMPhXQP51dHJIqayio5P5rZTPC8jcjD5KCyBBwSLrlOflpkc9dukLY62Tew5BcQwAE
QsgasJxO+HBq/UaPKpw1msZ8zOFuEWAyQ7IRs3lW74uJdnArFrZxT7rXFhyCMkjqGayPn3Mj2qJ7
6CxIqbk8YsGZXrXs7+QdqFmhQIDG7dQ1ENYBNJ24Gcg8HqhIJma7qqLdmYPZHkXG4lOwUEJlAiCk
ghnuHiQw2aM1jcVajKB8fuPbScoNBrN5zM/tpUu1BMT0Spjg0Ah3maXb9i+epRNKAURomxgrr3h5
QVhDlDtdcwEjrIJz+hm6hFJuxNxj9F52ZpT6o5mbyVHbTbRIA+cdBtr72GPKw6xBs29V6GxR8u1j
jFfdikIVC1dRXwPW9Z5lzWU5vMR2J4ae5p2hZ97enD/rnZEFXyLbhC/a0lgoaIahzVjAR876tbb8
3573GtAscO8xyVjbfCRhkP0AvZhUGpdo+oQ45jRUFnOz94qef0GFsa19Ugu4ZeqXAyE4DsBJ3ZO4
n8DApDsckPJPr9FA6nTKytDn9AC3ydjv8CLQNKXArMI+TR9GTS76aEDH6hI37hFfkvTBGFExaFDQ
ZJYR+tO8C7GBQyAht+ORBpiBZ7cdOGZ5pXoK0iN5nx8io6vM67yzNL5nRqOAo8n11TaD+9ve1fuc
yh1UNJZoKvU7sPoW9xrFLnKfDEFzw3UgC3ikOs13XD7zHCvGUilQ48f/DAvGm5dasgF0d0N20PFR
Z6HWuWoCnme4c3CP74+mrmeqsBOLKu4qG8ef0m2IQ07G27SQLoCSbUbBc08lXKSSOv0FJvjwITza
mav8Miq2VAUPMgLhO4plCQgHmEatKfIu2VMD4U7JKPwD4uT0lGBAmFnwl7h5J5KsXphaUwRepiSI
J+KxvwNK8lNFaJixlB65WRevaPdp1UVpYXPk0RA/KCngs6v289jqgpxV9PCrc3GKXiWk/b7KXFRE
9Y0azEYg9cIenZYp6S2iCl/qBN3hlYYbfG6bRCoHbWeCCr/Io24VYYqEVKtnrSvSHhpMuoXYYXNp
RFEYOVrE31V7Eg+4hSLue64ZIY50k0v09ixSIViC4ia1pz6dfffonc1+0od8A8YVTbP5Wt7NpiyU
c3LpxOfJMb4+UkiltP6fxIOjQ2BNfCdzGAbiY9eNhbgdZbL8zdXxOEg3j1PBkf6uCopnBj7nijkl
8xhCbYqI6nyt8n9awLQc8J1JAJKVUUkGDgtfASmEh5wHssI+0CF/99Fem7hgGzWCVHUrfbQ5rUUQ
DqaZEaXE8Fmz37ay+VbkGC1nNgrrjn/a90f8fDmPBYk8oewz6mh9XotGEfHMS9Zxv4BlEzv3I6m9
oHLe1/9PRhEJCsFHY8OwPRUybxq/kvKPITbbSySKrd2tWUeUsCyCiKs3vy/adcH4EqBU/dy3wRMq
Zhzj1NhGzHhGs+Tq7g/J2N1vQL4XStmek9RYmPJ0WFfkirzxDxST0rWFVp9CKUgb56ruAGffhli6
7+llr9X1Ww2FJlMs2Ai5kM30EsW7zNw/Eakk/Coocg7vRQIkSsoFbRs+aDqoNwQpJWGtezhW7Dar
PjXB6AQWVEwhdC0YmSuQfc5XucICHW5C9SKLwDiQI0EloYe/ZDI6stAWdifY6ee23BhD0BSoaMSc
ShGEDoQXMIAU4xwXU0VQLaBdu17+Sl/0+wUaBOQiGNjymbj6JWi/783uiGp7XBb9hinaczVLKfY3
KBfAq/1vdmiVtC+GhjyDw4jhSf/n3geeWmAWzsNnfMuz/m2plEK+mx1SYt4z0KoGGFJKo2wLtZqI
K9TerxnvEJm4kCH8ru6J8YsVG8vmeN2h17+3YGzBLlwoeVvnUCIdKeiSf6DbEafE6d4rnj8fuZvr
nb9ySu/WxFuGXMFYB/9/yaU0zI2OnHaJKRCepZMoE797uRIaJHrPVzFFFOO0xHkwNg8Wa43dsqXH
ZbjIlOzMky8CkxMhRAyUTpsivk/z8yD1/Lx/zK8A+GK0HrPAB2axG0oOHA9dwxTLWHcJApy1KtLn
AK+zKFBt76Va0d4IqSN+VYZokIW3cbZBk+RUs2qfjNPlDP/UiHhwloPJAIZoJpgR5C3NdxnBlTJB
i56piAc5pvM2EJt4nAfEPSmRzB3ROjRGk4GTTRvNCfSE3xvQIL5F/t6hicKgCLG09Gcf/MQKQjxd
uCKQnWruDNQkPmPPq5Oeed5d1lBR4pFWOvGNlA60EQVsfMjaO+QuW91gUOP77gkFLvdULQL20ez3
lM7meOV8TbbkktSdQeJjYssI9AUymWwurnPHrEfshI8n9K8BAgLwdIg4TJibTD6Ci88AulVNmTOY
3iQUSKKte8gB62v2YGLATfbpdXUd1FhtXuEIWXgOd14YZdCmqNXQZGtX2RmG/4UBI0TrhvRP48+3
OIvQHSZAYKuUBrz+FmOTUDxEekMjJ+kRKhDPkRu/cncT3q1rOVzWOSL0MsN0ntDGwAQg/s4WR0t+
3euL7vrM+XWSMzfMhrHuAXx35Y5G5FriODKYaiGjdQJFp41P+jAEQbvkU9QZq4lUL9jF1MiZQHKc
7OflfjBHM1oJrUXMkIEXv1t5HFIgSkuPOzTNdYd/kkGLbfZDk1nET5xogYauIWB+uYLwojcnwfuN
S0VGja+D64twBug3S6wwpciJTAXdT9GXUarhcgIIfhd4UYa68K9Gu3Wb7L+IyaWNUqQQwI8Mi1zm
YpnY0EMme1HKRq9X4LtT4ZHBrdrG4tKo3JtPei+Z7EMTEEbJc9I4JR7eFZewh7WIO8oP0Gerdebq
1rFUCVptLX6RZhrnpZGdgLX3o+BrQxBySIFqkGqjsXZq/fbRSRtadVKvtm9kT4ck1RI9GOBpjdkJ
t+rW6gP/rVtrM4uzQHSjjCJVswXMyIdy/dRVwjFd1yDPOvsDxee0WfzAvnI5MkBihorKNvQ0+Znz
xIN0/U8rzajaWRk/RGpnKFuveaeUDtaSBhUuSx6qOMe1Ej0GfWUqR6eWM13kggykIcdl1WtuFaW5
FpSDGfYU55ezmjxQLmnJJvwD8+hM31qNY7b9R98Q0EKbu6us26VMPmxUgJprRKNWPgbVqdcTTCL4
MAclVYeTYM5qo0KfjjwA5sRuuNEe88paFP9o5hwVHVyXbFaAWerdo98X/fG+D2xR+QIZCDOHM6eI
yweAKZMEDN4qG/gAU6Bx1HeIuRkWpIChgYC7G0MzieWdg9tvPUt5KEPUqTXpNM1Z6F4WvyZtN+I8
3koRVd30/96R2vnj7nWITHzTHcUgXdClHORluGOorpG3nLL844lfjczc34K7qpa3W/2uaYGtktMm
GI8VUxxa9QNfdAViKSYtSBxGbVnSUyAL+mseLIDJzH4Qq5cB+qNmBCh+NjcPtc9KLNprCDhwgYLF
Rxx1QmeuywIY6sxElSIyFY1Yse0QfcAE97AaXRt7Dk0Fve+H+fJtbjn4K5FRvXAJ6P7av2vWwnH/
s/RqbB2e7+olGXtcKlt0jH+bbi4HwJpPwFMtQadHsYGGKZnnoeHtut50ShvmXE2ZBLB9fctKG7dr
WHozOdAT4xT3GYL32U+GoyTaofKI0xhc2+zz4pYPThBwBvtl94lfudd9XokJNDFIoHkPqjEm2Ivw
EU6hPikj8PF0dobX+yuzWiTrPnS90BXO+5XxLEXj0x2pHmItdt6pRnM7oRVUz40xG9QHCXpIkcKc
FxNBMxd4vIvXkxMGAzUXgbVlefbwihQs7Bi6h/+H/myXge4t6pqtkdPnYCrxJLKU1F0lXzWnIjoB
uOsQ4Daw326O89geDNp7TXWQCdEj2IfmfilE8Mk3iyhofdtHzFUYqav25Pjs3hiCZUs46UDD6otI
C6wzQJTQrqJRlJVCtvxqqGrxol8pIubXGTB0+L7mh5vhQOzRl94mcUMCN1VYz1zpslLXPU9h9fuU
mwAdzUamugu9cQMOw1DZPP9Ozxm8R/OCCpp32YALbA7uEcgLfy5I6LDtfLnvo2kqvtHnKtsXRnsv
+ljOlLZGMKmoFAdES8Dzrn1cZ1uDCJ8DfM1BUgu21HOqA2ZEkaNUe2wzG+r02zpxiLCetPylLoAf
vTJdEo1xEkcJWWn5759se0+YImrDXGd/kEwNkOzbHHvlAbzCsolzmah2hNLdiTQwCI5aF1EmpS0m
3pSfiE/VdxNR0gbg7qLzSEHXSBsfZo+a7cbqJPvq0PHr4UgVVUhe/EbNuf9Ahj7mDnaLtQrgPf3t
gaTQ2bU8iUJQHX7E7aNNdjE1UAPkmFl93GA0mjMTrCl/cSAzR6zRNILzBA6qusrZE0qZAFJMvtNv
HIwbyou+RRKBK+7cO7K4PWvQ33NJouWSCEGhazn9za/ySZ+JBr5YVYf/5gOL+SjiVkEvS0Y01Wo7
j2OFsc5f+5DgkeuZNXZc4l236/+jhIeMlSKroCmxjv7s1h8pBWO3BqEX1IQ2Rl1NH3E7dWGGJrvQ
dG0Y0u/VmJv/akyEdYXhEk16h/QkWuDHjpEmbgntmXQV0dMXnE2/bQp9ayLg/W85NtnzdCGNVAkr
fdxVmTQ8/w/qIsr/c+BtGzrjKmEugQTlXjp9NDsIxYcEh4ZTB9mWqiIoG6bONdjVv0P+dPZ2oEPJ
rYV0kg0GtEK0oEPw/SMrkKwt+zVp7xWSPmiT4OSthj5sFcHNombaTTHpOThWXnPNy+HmIFKBEWS9
bBgrg4dBo+E3JMZ5OwMQcgDEtFMHLmjr1g7ALJAreBRIpANkvA7XbBbGL0hLI3J2b4L2SpRrcNdQ
JUTE+qsni2wSRcrlcLXvlEUvD5SRBC5+jiqK6fd7Tztfu/t4ttN8RfoV3vTUPQBDBlcruzmENyTn
VHxGlcXpCBmtK3yMTPxOvFyFNld0EThEGLCyMRPUZwGBZpuULAZx96DHzr7VbcY3MerRoprcXC3U
dZeP6uoeIJIxfgb7BfuZkivCKcHMguHqH/GyiBOhTyGwH3ppXJZN/ow12ywaXsINTjozKKkQm56b
oIfD5U02Nk9irmegEYvHJh043zCEt8g6P3Q28ZQfru0zanooJLE6sBi1alz5WNOd4lF7ExYeyd2A
EoO9m5MCVDzRiabM5SUzVQdW66g5zwKehA5j9AlRZy9MkPw/59irJBpb/GgdZH7t5FQMfN34etTr
zLIU3k8nf8lzzZz/sLrO02R1YxFGDqDi8HzFSBi9EnzVnnuXdRbv8Ene2iwhCJ8X2Rv6Pvz4SYi9
9tfUOMSXVHLSY/OchGaUF5MkYAWdmOLexWKt/3SyBWoGw01ei9Orew2KlDIw+RqsmA47vb7rKYGz
8osMMxC39Pe9iIjk+PNtHOGDi7JcUVMa+kZPUGQIdugBmk1F1HrdU7wq1gINbU7RyY4gboD0okkg
RJ+dIBVBF1nT+8lCWo0IFc088ZLGil+4cEldjhJCmkJBVUIu7CLljiaPACVIWtYpSoOqDBAljK0W
A/q7EkaA88alkVBj3p7rsDzC4JSEDT4TflMQl0b4AIF3phj+jlAN/fFU5i9OBMYIC2jBeoC71+U6
29RTzVWQQIpvF4NRmpGDFz7tZqPlKdosBcEffb3KV0nrSoOqUBrVtlezuChhXJBchPZRI+YdOEzQ
LQlmzoCWfrhBWXhvGqOk0Lt8p7yRBCspEOEfjBiWt5sQPBY5wU+/xald+8NmAWkyZN8CwGAswT4W
OmQeMCMwOxP8EffOApMQvjbQ9eLNqgPXMOwcay4U4PguGZ3QhKKvhYp7SwM+R8U2jpBHLqDRh9rC
D6Lr1ap5r/dR04BQlGPJgmYpF65qcWGPZQHIsR5iW8t9YPBVHJyRxYrOObV/WGWj3KPtjblq0unl
gNJE0WcmvK8hxIrR/vWTX67slaLIPnWHwrK9osk0fyHBqlg+NXj/6Hrfvdm5KdVhdsF9dtFxhi5M
iCVUXh80OVl05xMvjggU6yN1q8LPCPpKFkZXMb/LiOdfQZMw1E5O3BDw1lW+aHJY0R5hDuvO4Fxb
mU1duFfefMtgFsw5VjjHlOXFuwIBwqYL7S7d+1lY7Pbftd9oh+Ioo7gLt4G+HMBdkiZ6w7RAFbTm
rJfVbQIVA7LnYFvPjDgX/eSlP0lkyFitjaOauoaBhBY2eCFXxnpU17rQI9kAbJr5483j3L1zGvQI
QcwrH22Wm3WOrdqXObpTsOdjPwgtwNqqQfFt86AZV/cx7ki7QLI7EvhHfLqxP1qjwkIqcogmbbEo
rKCQ59FE63dfDecD3XZkYJwbSuBeya9IpMRxUJBKwPhzewnyx7HgX+GWgkbXXe0qXGP58LdxtIEd
Op+D8RPnw52BW7jIXvosFrXGskRpnnmWj3gy33jfHU70spHSgv5QTcRpxcTJWK0flXR4aAk5b2ut
8kfO6Rp9bWda2ojpn3hZDap9xu5rrcGJTEOMOpB78Jac+pfQFwDGIfrdLROaFZB4NHxwV1ePaQDv
qzxhHRWaUOjrINfu1WzlvHnmTixHpJOZiuvE5bdEiFQtDqHAUE4cBwO7ihNK1o9jq7aP3Pni4JP5
22QHNzKlavLC7kloZO2KR1WhwGrq5zYgHlVAwbgs+FMsrTqhIMyr9ScGPglLDPUH2Nbn/FKLXkTi
bOFyGbTWK0++7BMRZeWs5ltVf8jnkDW+hF714nwAEwF8wHCg75wXVJ6HiPjrX+U8UZ59gq+1fDZr
6RzJRvvWSPQrXaJ3XDcvsVIKbJ+1whfW4m4MJpvkLFXND1JdamQRySoOIGLuW+kDVnRwuW/8Eu8F
FxjguAmG7RoP/7Y3/iiTjXnva1S0rJu0meDOLc4SwgjhQu6sIn0z5MyiRzcaiNatRq1HIu/EneFg
pGGh/d6F9NvB0pAQluLpHVyZevhpt3/Syj4AlIVCl45VfjWHdaQJNKjpYQZfpCKSevPxZQ/j09aN
qxeaeHJttY+tZoTipx+9wQo5ydAfG+RlqS47+cpouPhKyD/hUSfBD7opHbNLuOWir2O1vp4/wDvZ
qOgXr8uskorwm5lSI024zl+HrEbx/0yVqj6R8clNKVJKzW8L5TFMIph/GvWKX3S6p8FKdoisEnSg
G44V3r3/Enttk/6Z+IPmRX5PyQCxpLdJk/tRb1OSHfDgMGS+MUuiH7qlRimzh5avMp4zlcC8Kvcz
GtG/A5NoXLVROieltBkE1nANBFrG+x+5fMg85B+Fkw0fYGoNKcLGjzdm7vxRRTvepQNV1y0ny/tw
pBhWmgdtVdbABNp2Deb3bp6UeLDvE9geaGuElkI8TdGcbpDA2Eb3kA6ank0ydnA+p+OZIlCUFSwk
5YWGD5blGVLWMNDFRoUIPTcdZn8NesZ99MzLaIAQ401oheUQWMVzQ6rzulffiLGLXpD/XfwQsTre
Ff7m3E+xlA5LoWZakjU9BiM9/rbTGykcGhXJWBGkBM766vDPdFwgZmCZJvjAe4Qy2QPd/iOFS7Uc
Mbk34epvWbPsrf4b/ZNOSWECedSHkNy7vyGAbB5QtShQGpHDDdYqcpKnr+9jij6wKJfpJcdgB7oT
9sYwgCKJqHPig4e5UXZKSseF7xA65sJjox4AO0xnuNrYryP4noq6B0gkeXQ82pTqyR+Uv3rWvPrW
Wc3Oi/Vnk1uhZ9UsvlxjZjsBmuR4eC6a9C8TWFsAtBgyoHt59Bx/IocYSwIULSjJzo6FjEdrNuAJ
ccqX4Oo/NwP6yBVkvi5SgHkyH1f5hiIzitwtv4RgsArYVBCTOD7c7bjfCe9Zbzjsoxhkuuu7Hcl3
TQ/bTlrlRma/tTPKgQ02wbrHlYlQsNZWoX5plQmerpXaz7LpEF2V4ILrbmJXyC2QoeCsz+LrX16J
sl7VUub2pX5pqWxnky+VpF91CE/dzgytPYWZ39X4laBLt1L4PenZQsXqbYQuUGdT/LYczjcamWxJ
ytkpfkVbtTCCh2FoModjB84kUfwyjAOdzwBN3SWU5am8i1RlstKezLQAV+iPGEddZpiOuliiBPb9
uSvZdxY75/XTvq4q5jKhJEyEkuDLqiZQYVUVj8pt1sEl9XysZcH9UVejqtTGZrwAT7nQDx1nrcla
1h6vmuFpg/xc66xe8qBpViiqtMMHu5qLm+rgRhIHNMuThVHdbeeEprW5Knmic+X66mExOnwP1hts
BOfU9e59VCYJixrY++Dfnl2QUUPeOY2gSg+2tFBpNIdXo/afQkU5OjGlhDt1FNicA1Zs7OLIqt2o
cbUVGpBo4DDW+ELwL4LqjSjlb8+CavIvT3m//+jeor+fddGRPWcRdeGaOwwEsGXDLdtTGXg5BmKV
cPjiyqcv27RyIv87xSvNZ/G0XMkN0i+F5CAyvpFAb0QBJdoGpk3dYdreM3lGAGjnDSHYSaXxyYDF
dP5aadnQ+mvVL3pQOhkAyZbTgYNqrBORrwcH0q2XHeC+PDYcFVrkVyYnROBDx9KMjd+4T60EXCIB
qipDuoBF8wZdvHUeGVd5DPhe7hfJT9r+gkHK2tw+AwphJRSlbykYlB+GfKrgHr78T/iuXBM16a8G
76+1Jea8qj+jLm3oU3cPDHWB4YJKAAHOKqv6eqmpzh63d6tp7Ol9HszH4QpOeGu85AWydNxQCYyU
LL0U++Z8sDczCwHR1O3wwXeSJd0j68PvZGcVJNtAGBwLOhwrXPF6qe0g6I7cvgmA07bAk2FrNy7g
Tt+uQ4b/nZs6wrvkksrhfTUPiAXP/cfw4oxGHT0hooPZFBL86VpjxViIg8dYC4ELMyVSMIoKsw1z
uDQXPDJqFAmqXY0gmZ0ZP7EHjr4YXaTv4AWJUJ4EItd4lZ+hE2m3HJf760ZkyEfXNFrXfzRk1/MN
atLCA2H1mEJo+1VijCdLSL3ZFCg/3M6LHdkmacvj281bfF3quF57BS2QILgDHPR3aJnrTeQ7Iugi
rbdD+M8o9vBgpiC8BugdS170KQW3wFlGICk69SyEpScFbmZ1svUZfJVI50xl6Od7B+OO9N6S1FFe
BtZHODGUsbgj0FOuvpUDx4bKSZkqoJqWi7KUojetyy6s6oBBQIm60S/dp8b999rJfcHOKV+0KjS0
UX52D7Bj4ccj3CF6xWIK32FRWzxAbYwU8J2aNjsKMWjCBIz3mGdRKte3vkAHDb8uJTWYw8dL+7jY
CzVW5sEERSRslTB5JigVoOicqG3N+LctSpH+7J7dF05dv2AaINE7dQXe64FGX9L9bTRnQ7vI8XM9
+ok8wFlv6e5V5G6ZNSzs+mGuNlZFBXO69mY0WjyrIDWsR3fAdewP0AwBZUfgjm1yP2xZHmDytdww
PebV7plcreSGdIz2A3QQSNtNWEed1ovVOz9gqq6HhOYeyCbqbGHcHtz9+gHg7SgZMlUZ3A7XB29w
4QjHe9Vn2HEbAzgMjM7l4f71yGPac8T6pdM4K4c+PRz1LGI6L4/Lj3exV+6Xx/xOxSIenpEVKL3N
LRnHtsbj33DZqt/3k3nEfHYwgivbmCzlXfXlsbpZ0hneL7t5Tvo6GyuabwlnLQ2znCPYj9wqdzCZ
9AxeKCNjm2fq3DYn7k3boRsm+tA589E6Xh+5bYxoSPexU55E+DlZoy17iYkjS6LxuaA1R+1INn60
b3mmiXzHtIOf+Rb/p/pkVKh+DuGakOPvqeHkOf8B620UD0fHP1QO6wEWWcBrpC0f6F2Y+tmo3Tro
en7EW6xy+kroNIUPRQGfQk/0PLN4owAx+X/Lmkp0o0Re7L0Tz45rnxHxrxKS+kjIMdy6gYgUDg/O
UUfJDRmWcwKFxTQAxd4HHZqpnpDT0keqK4brn1EifQQ4TelDmlXCzC7epbd3BZUGp/quntf0/zmu
Ga5v8quD1HDRI1NWlnvz3xdY+p8wdj9yuxLQ6J/BAL7OXVnv09bOAh8AA1R+1vMUKdxgiuQocFWn
kS6bfhYt3shbdFNy6xKyf4swDA/PdpOoEbrVrtsNGT0/9yPVnBEN2dQlvjjDG3Dk3rd43yccKCY2
jRNm3qAXLH5KRMs5VwLEv99WNW945Z312xKj9MxhdZN84IdfcV9h2Cl4komL2J2AG6Wv/Q5gh9b5
9dU96oL1V+OFEpjv/Q3xxbsLgNu+QJeDly5qeSPTHBOnPYtLMK+cQ77eM/84y91/5OGrEmqHoBO2
iKr2MiiwMWzcKhrCZDDOM1qwnWiONuqkAk4Mdorcv32g3byxFaF6zp6iG6jQqIHg4ONUNowQ7zD/
8j+G1cugGqpgeIlb3ADbNqa8mIa9VDWksFJVJsk6I/ZklRlfzLm55tId03nXq0MePgsRPlIamVbd
0/flGmxNKlSrNAvwEuW362doIjmMjPqoL63ytGlD2IbSx6/GDjqAWcwxtWiTSv58U/a96liLkIU+
+hCcwtCw0AXj4x70hNzX9tcD/1V+3kgFFxU/iG4Z7aNEpk0crYjUyNbXued1/yN2wdxQAtijl9cz
aiz+gOOffHzs5EK9Y09p2uO0ZhYVKZeJSi1rNZvH5iGyeVDUiQPFsHTtshsGrfUk0SzXNLqGzO2O
LfxKFmlr5IUblCTqCl19NMXiHkIJjGkZN0yyQfRocwoFzIyLok7BtB1oI5dwHZErtciHtfOYT6EF
4s/8FSKbMARe6H3ib0RBOY08g9NVujf0/DSZnO6wpO782yBYN0sqt8JsRjLFQP5DPCDBu08U1Bm9
qDz1Y+7C5f/NwNhKqH0C0BmJ7AjxatgOJNmlfJWAy9hQNo39XcmJmmdDB7PGTyGcDOgIwPEpsmcU
WQlAOCtK/RO4seLiTfjHKHv5RIsu7opFNyaTARzbQPOhhD2WecSCKAPcFmXc3s+28tyBAD686Cuh
UgnmiEteRL2Pg91gxrOlfdK2yjBWqM0bLjlvrcnrOrNUOLV8mCWNu21RiLz96QePkunvxISBVl+g
fLdYNmc3aTjxQQxEygnFZJ3kOvUmrq2xxoJBSK+eGaKl/P6jL7ikZGPS4CW1fD3B/jR7SsflgAT1
797w1dCRpFVP+DNW47X6P/QaO6Rlv+/i4vWbP6JAmwO2mdsWtkt4/dw1Ef/phC2xTgShl1m2WNc9
t0IyzAGmZ03iLMeV+6DRkiQDRx36tkR48PnkJi7layuLrJtAzbrJttKbvT5arXc7QgAu47d1Nc2t
bEiWgsoYq86S0C4C/OW0hppUYeRvKfryya76KMlHJox1zuYPxvwvZrW5vRtsL00nvnQfGkhzPX46
E5kfqgX5d+8PDLPkElHbNas15s3tES2FrIRW9c2cGwopYIMAGYY3iLNGiRi89JKeG167phcu6hSA
EsdXsV0k994jjGoGOP1q26qpeLG0XwnPbamXbsQp5FgAqkyIueEHHa4TgECorqXCBTT+8uYLlqWx
4XZp22RBhmASn3p+C6lma5zfPMsAj3VuEeqTD2P/8gfTYTErH8fTBjsYYzyAHcT+XDacMGqG5QpM
R+zfx6dD/jNWAjzYe2lEWeiDHHqd+BW4fKIDb184LHQ4l88sEBk13HS+D0cOiJoFs+6QZxe07cLq
PphBVVEFBMWvp16TDcQ7TL8JXTfId712DVEr+5hBMojySEIVw/ouoRmjFz3twqDcdWZc0yTUECrd
WZjWjzXxngM4xbKDAtBhGNM/SV14rn9wztNNzbDRidcK2OVxd6kQjXlSYT6ZZEZpZGBxIaLEebVE
/4bohFh5jBfwUFLqI1sa9lyfzhqz80ms+eYRFJqerg9vfSPHdzhgGsznbgXdmKNlwBLz0UwSn5dB
mxDDXGUPs3lSoCV+UsSWCdBikWOM0idEIx4ycaJgtsqzjctiZpQ6otDL83roWygtOn96Zhx03c3Y
KrENK29g03nU0g0oUk/J5DlQhlzctHdGVhl3Ok0T44QJIWloydhotJjSyf1BoLnb1eFzjjWhVM84
rTSYSAci+2yZ/I7FK38RkpDSutN+6dWIezvJPENUwmQKIcRwFe0ORNplOceJgN/uE2Js0dUhy2g9
0YaJDo8SgqnMLEF0ajksXI0c8widfcRIGtDUGOwtplxdxbNEhIsntPT9x92qJfrWomblTbDD5UxA
rYPcayVsv+dt43G227bTvKFQrrZ5Eoe5lnNesrKYzIGxMWoH6IVGlYq76XvWs1oAEvbUhTv4zKn8
OpbrrKPuGpv2h7Cqy19h0heevFPWKcQwMDubvKYKQb7uPuknpjJ8QgdwjcV7bSMcd7a4mlJXx1Zc
/T2mQuPrEUCeU4+CWIhtBoAOFLsOx0TMybi5LOLp5FKZCkR20yHDbKZf9DXb9L9HKjSTr7UZkMLF
1zCs10gkUf4COfFyt6KMN19ma8Yb/cNmKIviA32jCHEM97ZkrHwhydUR/X0SbtxagHpVKX0HQMSY
X6XW4pDPnYvXEfIGm26Br/eo+cmX11pFsmQPngqUsV+gpbFWjuBJ7A6vSPEoh0zlRvrJQwE30heC
P5okXyozxnw2zwQmrbzVL5cFjP9kVoSKBkYA8conB6zzCnuc0Oud9annnujeHvYrAYLYQfpgxD2x
C+rdDebOxqeHg68f6zNmK7HTxWxDP9fZYMANKKctELWCdALoKLlYTZm+/ZltzXtovJYH8WoceaBb
1lR6Y1SopUHUclYF3Z/IKkQMdohGoI4jSW2V+PyfvirMy8nqOn4sY/Vs46aXzaLlXvQhUboLKnSy
p12EeOaAJ8dReST1KZRtp33PGj0qvK+AdXEC42GRZ0LXdvao49Znq0Gt94M/1uMWlpsW/vEhIx4T
3Fcn8nCay2qpRal2dQKZ1XzgpfFz7346hqGPRhFqy1/vgEG90p/nWR3Wxf5SKXRDmTk2rWPQyAQv
ik8etT7XLMdWTa8ld/hW+sgHHIDQjcNVzIrB9r09gwGhtd8cb8yjz3nrUi1UcVc2yPaMvSc8O24y
WRIlXPk8Mw1lrrh+e6m4/BYokzk+/BkVYX3wOt+sT5cZLadnRRWyX29VMWVt7ojT7Hpe9kA/PpD/
+RsAD+ul79k9hFoyw4hiyMsEwLSV0xejUat3SbffPM3w1nK7//AxqDtgNOnHdGd3Y97fro7+rntC
g5rlh9iNxEte+p52CFSKp+xCq01/YrvodJnZmR5TShzz4Egwr2mpbdXlssCAwFQvpGf78FB/ykKZ
lvYbP6j84xT8iMzQiRRgB+QXZIOr8Mps//asbmUn1+Qh3v2bkpg7NNv6AuGxSLZh84bKZ/2cBXfJ
tFb90SxPZSUUtlVTdt9JpoJitaI+hQ35M4CfaoGSG0TgTjVwRguCFPWTupUwueJtffjQstnz9EXE
a4RZKCO3Xkqvho5wFucS/ybFQ30HZUBvhLTBLV8IXVWO40jSbAicqNk+kL1sKgd4PigN2B1YVI01
u0zQRv25kALopzGCt/HcX5+JxJsAYM3LLcUDkRRmflRQ5OZ6TcSspNuqdSHTr5CICxpYBXjskA2P
baqYrkN1QM2dpmPcmX9BXJl/N2z/xm7xaCeWj1+KpGamIIRgW7s802gFR2vr56BSt/KLH0fVc/p+
j9HM+mgY2CcSYUXCRiNlpGSg8NEzvVtdQ9L0BSP8SR7ZGyLC/suijgOwbOM4y4ZjdmXEhuWsr93D
ilkaWMmW2rrejKUtsyfetalusKt4cAgwWAC9qJWtPiWGjn/8oRblQnFXbbvwHzdW4ooF8GMxpRmM
IaAnBUBG+UKHcWYxC0lNKSaJUnOW91gDgnJ5wkZRLVM3OtYaypf4YPN7WcnPehE0yDtnvvNrrPvg
ftt04O1t5qCcajeLqV3afRD+nCit7NIyVd823+0gQROct8PdDcr8Nr5JKaRFm2nrXDm1C9C8pnEV
wcRBIjGFj8XPouXXQp1StrPAK+gYaJe0shxETQ1a/5+DBnkFCcGLlWHrFiVT+TJZyHQ+DN+kIuc+
jVITyFxz0ziZ6VfUK4lZK6K8IMhwKwClUCZvJQWqhMyKSAKOqmLAhTO5CEWl3CDll71jvLmOcUdH
Febv90ZnAWI1VpSb4c8yR8TuY3UpeQeYSh0Sq9ENfSmsSV/PQ+DExiry9GfPQwE6ZRcSNsw6gtYE
rf5zkr+2A+7DWW3Z4XnXPnYa6tv9P+nC6+R/sp2TFg5doy/2h2PriWds7GdZKia9AP/es1HL8kpo
IY6m8aVRoRBCl/M0CLLz/WshJt/mJ9yb1ddcRF/ohZEdX7LVNblZwySZyaJo6tE5N1YiwaFz6CqT
fyyDf1vvfzLJ5ie6oUJujKiFiwvvylqSXJU0UnunHYw8lHirv25D4I7FrA2NkMG8O/uVlyEKBoSN
PACcwdXNnOv6t1E8fb8roX+aidGJfeysgRHScSIOqBBAv1kj6rA8WLChuXJarXzAr4x4V8VjGjrS
5sBO0SevyXt5tojiDICUql6Qu0bB9SMXcvaa5elMR+oH36mITHUfajIkxPLS5xM3+4+pt0nB0Hfw
JUbnGbnzgOW3xFJJGKJA9vhXsr+cG7vGVpsdoUWr75SjlLitgNboYEjdU6xM8VFkyK80Vb/BhIS5
Xw0KnJOJtWGcK3cPNmstprDgZ+lVYvp2I0KQBIyZlc4mkLcstMrX81PGwjMOwNruDzehvC70zxzw
pQNSCFBUpO7NWfI6cdiMlsFJLSNsrCJAHj/ylisnU8Crf9KmOKDPVedsgNXxDQVf6en9Qi8pgQzc
0PECYYJlHju6yBTcg+v3A7KuA8KIfZBa1g6Hq+6tRxwSpHiknyYUMvHdy8ejVMmHgPTnX+2qOwKj
yihf31EEDOS+LpSEzjdU4ZIlDQgHIrSjyF5TRD/+GfniJfueU42SEUiP4L1iHrJk2tJaofxV1O9F
mbBl/FrEQmWFlZDkGXtLkj+J4uyszqiYbIunU8CjENDZ8WXK/jmGesWyQgto1/LzZZ/MpWgXLf2E
nacfDZe6D7UhZdlLQJspi9WE0sDqoHG73inMyJCPx+QqeAeEa5DQcTnPfG7OXgI6L2nPndm8Oke6
/dFTqLCfwz+IsquAHTGlz12YrCm3ZXP6G4+1TIu2LFtWPsgV+EYtXHjOm8vcCCkt3xWbYuDvslxM
n0xAXaKR8X28HPR3Tmh94P0U9rf4OLQ9iGFqjcw+tsnyHZqaA0KK3Uo1GlHFnwL8ToEvWNpc9+fO
0P4bqrngNzmV5y5vDapP+hPY8NxN135faIWrqobcx4p9nGr8Ef1DfZ0rpiYJe0Q7yHfy01VM6hHR
4OVY+du4ub4FxmuDz/J0UZg0QKAFt3kef2jAGLzx4Vp4bvzrjdnL2dIexnomFYD3aR17e73PBLj/
wIrQj1X+mp51vualNlsxKhzw9cKeLNd3jfO6pvZZxtwsArNstNE5jfA/6YkrdVJJ+m24fkPwkw6B
7kYg5sxFwIAXBy3aVxJTTKWud/ooFRaQmsHmuP9eaIVBMtWe1ynXtf4yXiHG7BNaT6dIuVk1zUzs
UcFbW8qnV70OwKSZPJtw+9MylT/r5YutlMfuo1QAVP2oSWDgPTowOQkKPCHFAd1UgkMzw4VPVXPP
cD0HrxQ1J3JeSolNd/sFl1TEZ7FfDcOEuBelHPkgtSomRD6DVfUi7yHaIgNM7OZh3WT2KbUE49Px
7mchnssXb5tcDLX6an6QPctMo8YyVeSPtp8VJGGbjvt4uUDUp9v78TH8ezfFQRfCs7ggjhtM476Q
PLKDjnfuHMj+PVMgQe6lKhpXbgg6lJ/lKc0KIc+w9vu/rP5qsRLKHOXv+CRtPnQ+BoRWd5HObhBh
maeMIkSCIcDWV/46nXWlKFPkwKBiIs2tefzPb7CHIfzQWEg4UgTp5hcpXlm6iLssKUssTHKBPfwj
3RoKmmC2HlHMZGaLo6yadWF7SKJzGEj9s/rEzJ+vGgwGE8Dq4EL6wGBrY+QmKJiU7Eu3gAJVJCLj
FED2+P3BZQnLcauqcVT53zvE10TdnZ0S/WpxPYBIRrm6eJamsdSHHz7L86yskCc2M/Gfgfnm29Fp
Cj+wlrtFqa/NzioJk70biS8H/iGP4FU0JIBvS8BKzWaDwWXdoOU5iishsAtiYEWpP5ZgrVkml7LE
cciZrxkry9/L2nZKQU9MGz8bcuh8gPBpToJZxaYI35adnouF1EFkFPAqNZnskZJHG/eLZrN0Aoa6
Aejrg1pQp2csbNh5WjVzDnQj7Lws5HNaVEdKI8+VTdUI0l5bHEZ1VJ+RGFvH4CTOjNHn3le0+EpO
GCmcA1yk3jm8u4uqNrGArbqeBQKtfc9DKK60cX3k+boPTFtjPQdmOqReOtC47yIspJK5+zAkAoe0
W4SU5ByZUo4A2CQDTOKIRPMh3hrdeSqkGJfHwqBCAwKpW5q0mn+V0mo5jWxaExKirRIuUy2Ex+1r
8EULumDl4sjXCm75rDq8Cq7SxHaNc+TjexRNa29aIvQB9GilshW25f0Ty2KGy5aHakFLzyBKJ1t6
6Ol37Dw9dRz2kqSxOats1ewr5tnndXHZVyu4bD0NjGiBgKYsZAwvkPLd8ffd91C8caX3BA8oI87O
Rc/JbSKqF8a3azdkp7G9K2vWaNkWX1k11eMPZx90uE7tzSYSx9yRI9RWHmVvlzbJ7kA9JJtZiJhW
Jjl2DdSYhrIKr8DBI0E8e3Go7jCPkQPZ/yGAkvVkxq4DVtxo2554EENssJKeyB+mGbEa/JCYxCzs
U6t2O4lMGpyO40DSplo/MG+hoYzZD5D2wsFM3ZdcaNYw23B2Xjgem3v/dvF5ZOBWk+2gKx48AWf/
6qBrGQi/epKBY2b7tLDGoIGnRgnTWilDPNY2zM9Cpm/GUOm3PjS/2KU9Wx+vjcILUbSEIFLifZ40
z0ir7IEwuwA3zPReE4UnwGb128VwMMPqUf5sRZ6ozF6WzYEzWK3MhV1qSgP1UdQr3KeITTxSInyg
0NykZFVb0Wmt1XnZccQFO+U9F1LNRpVeNRK9hhuSgrr42thGu496Ho6I2w93OqhdMNH78dWakd/5
D1ylFlrYuZY5nH89OYAovNuq/f0iDivUH++5FstwmHHAsx812k9oMrigryGamNk8ZNp77eEegr5J
8EB7tNTxI48x3kSDvz0UFM1+/VM+37aeZjpIjzRw/yK0WdeduklRHSoqF8o7l/czyz7+v4SjAtXx
g44dJCCHc7Qh+XzINF5YG/IoD19olvW3a2o6Z9WKjBRvA5KcYd+JKNWnKu1xu2PaBEdp+Gfpu/gg
oCTrT0E1SmqiYNbHWhF3x6sFwVwqMrxKzFG0T8r8Byct99+z5dP7jta5079A9LlSW3KqK9y+2ZiY
AOY4Cgc+sg/poCQF8KbyQSvRW+zqAtbFGh+uYfdgS3NZZQpIHwBIPf3Qs5Prx5iuhbrjC5AGiJ1C
3Bi/o+C0Do1H6C15IkVdlrPupA54zvLBpC7PwuFAhrycJGXesZXoR714e/hr8L5e7FsN5P/D4jgY
+G/Bv2N9Dz69Ihwb9Y7YC/pD+geoscRPFIJfWUKZ6rxyKhecEM5Igrsha2WhXqpSXl0uuAPWJZyv
x07u1Jzd1KtPMqJrB1Rp8nR/Q6URRK1tP6c/Loc4yHxDhOtkamLv7IoVHvsXKOzYXnBZuueorPR4
DP8E2j8aY6C8/8x2wWDOusyKa705AGiZjX6DgBVUXPBjCrbd9raYPrsLTeAyny3ywk1clY3CShje
f2B+HpMEac7aEqij62A4RV2iV/aN0vkJywTXGNgJj2Mp8xstYCpPFhV77fZF3skM67w8zBNpnQa9
1hiNn/TTvCRYoCXf4ykvgOvWM2bxmfi6yQzsEYhbTQay6GWVFZYL1OiXNoScA3XFN4o8u1S0ntfj
K8RySZtL442hRIkHufcWr6cZtuBsPi2BRARe3jUDL1DID9l9pG4XUiYg7L9WZd8R5DZN1Z7OE8vx
O+4HfKcY4fMXIaUa74MeZmEI9rfiVRGyh8BUZLJi65akOuI5Ui+9c01BKqLkYZiO1KlQNJMGE7i1
ni6x9h+EdtfWD3QyCVNcIb46ALceRpBt10khCBmUiO2tuZtpXeuccN5NwvKdnoyamG99dyiK1spZ
00ZyqSNYHjR2zQJiJZgwJ97FgZeghYceQrfJecsjnkRUk68VtFLsgFHv42y+da2d8hBE6B1KHKZ7
6ccDWbbaTZgVpGEw3H/7vWKAKhihYjpZ48BRCgutkoga3qiNWqQG2frA2v/6bjrLr7E6VTfZndep
Obyf+91Qu0u8FE+UwgYzyVo4RGMWAVrAwiztYZ8khT3T8JFvGLhkkFFYai8FSooNclJWGIQorHVu
PFIBXzzE5K4JC/lxsW12pQPgAisdTkPp4KqIy76MQ8DUHMJd1EFDicQeRE1s9KprCxHhiXpmetTd
B3EmbA8AamGq6jFTD2SIaK8Fn56pwrq5xqclMzEMwmTL11BoHjn59HXP+i/6r79qcMR7NTYOTpLZ
z0dkbTMns0hqrcLRHKVD/C2PyZFCBdB8PnJgpBeXc3pIUSp0ROe3JXrSkbGD6+ASAiQw1bosIwen
G84BpM/j+Ps/bHAYkMZOIx7T+HHMcUdUVdxGeBQiRLCXLg1+lEnJkjLUdTxq0wnGnsvFuryg4O9t
Joc88SeqcW0N8CRUzXoEM+SeuSveHQz7UwDBEyBXAIaHzpFBa9xNszCzi7/QChEK0wckmaOpNc6k
BrUnTgAdnlUFU3A+z2QHWKOg8ayUpmdNnLNMkh/zZ9XW2uFi1vnSQTvPbhgBy1TBJqHRjXifGAJv
5Rs7u1eTk9DQlRq9oVqwh9Mivt99lU/Ux7zdT6Yz57/v3ibC3sAhmLre9C2I8OVT8ILmqTjb3Aty
qd4JdhT4RFSYrkeBVSt0w9xEtT7axl5o0xPOpblmHhx5v5BT1iuJwzu1VQmwI8PUXa6X3MEBWSio
C0HZumQpyL37eeksVcobGrwFggF9my+T1UZijg9Hf+V1ZNRMNjXt4igXUH4D9bJmgMoT8eZ2oKcB
+i1JXEJakM5i4fueqZ7ets+ZTYKYOTU33uoA27WnaayffJA2YaYMSFpgmS2LJMZRWBdVDKre1Qf9
tLo5dSSEg/Q+0UedX9vtHy2DlrxP37I319sW7vijL8rihCjz4KqMK5cmBJmk+UFMAtopIoF44DAT
ikqQ2Y+7tTKgKop6FsdaCSdAuJVZuCGOpeWsHDQuH1pznlfH+QqCAah2P6Tw8o02sNDtRRdJQE4L
w5o+rDaSJ9wF85TfjWt16d1+ttrhL0BgIiOcCBNpNjNbwE5CTL7Osyrv0KkrYBUbvKM9BQXTOh58
Y3EMhcM+mpoav7m1eIg/LSvrbzFVl6zZzn/+ilBoYA8Vs5OMiU/1IYqZkfXvi/ChnT//elqq+7fy
XSECsm0cuzf58XyNz7Meyz9NK/u08g988++N6btQTdByCJPc0h8X+15DtvK4uxvB0zdNpvAsSITQ
mrEM9pobUpQcwHkDL2r94CotMBln+oKcb8cIWaclqplmJd4EGxx9+BGue3PCL4awYj6r0FF8AD+e
KLp3/AEKQn1bF2kNjzylp7ud4Uk9qn3VjHk28Rzv+lGQc+POEQTfoDeAjqsZyvQ6eoevoeu/7Rlp
KsGUx0vJDdk5gQq+cTr9NUXRQQ1WSXIhiguiYjXCC3sBpFrDve9AS++OU+grQsmyBbtpNzsAx/Iy
hyBHW1f7M1dqUDcndokpFcpUX5w9J7K+tXz+sfJNXqVBwdEixqGgZm6YIl8JppMGdJegjYr0pXhX
DSj9dhlWVx9GFKQSuTjl4y/oNp2ebO0gdZewx+4Tx6EJGjFFk9DxCXR9oZ4Sh3s9A/VU+Zx4Z0Wb
K6TJbINPwioijPruS6fxgBYNCoWRYaLiboIsdG+rsXlTCCNxzkICTj2RbLEnQIgX70xUFFAhdG2v
wOFTH5h/rGvqUkLII8T3c8kjwxmVcAMhV0ab2/Jyd6Hz4FdZyx5aphEB0G0qmVyV/W/YxwmA2Xwi
4RSNYsqEHF+ClUYsrDyxUJUayUxpp7Dy5V3DdzhFVBztDhBFqL324oA/PKaW/gA58JSO+YRkOxVy
Lt0460FTFe9KZkFj4u7Iwg23vdU0/Zlz2C5smsQblhYHBMeM1++kQd5K8+vi2hx1er1JkFAKAu2R
QO0E9SgbvlR3XuzClp1dj2WrDt6sMxLDx4/oMKiCPMa9vWhEEz9pHpWeuBHnrS6kkzW5GxLR3INS
+cjVwZX/jldVBdgUmm1hqXFcX6cC7n2yRs3KPChMbZ/KaZzRQbiPWBIcWXq++WYvyREsuCRjOtac
7dKTsNtpwKiwcg+ylp7IQcEtn3/ciKa47EzZESrMDV/o7FKvr4p0V0X8V0sOuxnFR5hOJ6jn/+Ey
SLXv/fgT+39yTvqiR8899CAz3PPzWUWnjgemLIWbA6HP2WYupz4GMIgtcChkiSyk9tb2iIw8/Cgh
ExB+n1e4J4cwkctUINjJDmrOs0PmUH4garSPCKYMqoFZSY+PRTtPfqycPqyhloFGklYjncvpyUsj
7oDo6b2qcPAYXizExqczQo2B/tQvWvwM+piDnscdyZ7bljNSJuVb1hjOj6XbW25Tqs2sqTvDto1G
nPbiQaquUnLNBvjAyZKbA3lbqNu0EiLd1E6qJfaM9v+wa86PTfXTgvimh75aVdXizOW3B++2Yd5Q
fMJTHYLHEOX/+muRZApTs/urnOk3xAWH6Ijp2sSn+/iCzos/EwLq9VG8yVb9Ex7bgQMzmeLVb7IK
OEUG90slgknxhTEKnlFUjstX5834W5wou36JateTn2Z53FQjF9zvQmGcGPMiVuy8ZZPN5gICXGC9
AT6HdgYIYbfuxRxV+fe/nVHq+aRlOlHme6Ufu49u0qz8mfuU5Td423czYaWe4ttGoB4Lti5y6+Sh
I4C+4mjmWc/WAazuHahW8uo0wopMO9s6DtlS/r/8dCVq1DqEq0H7Aa+SiCjs4Et0TM23X66CsPGh
tQCn33ZBZxniv+fG1b6tR6vdQfj6ejoVPj7ZlJJticLesbum1/gQf5UUGHhd+O3rJ8YcRj6LVH8Z
76KjRdYQD9KEe3BWYCwZ09zTyVL+KKeVPy4wNFrhCZApoTUkXNEv+gARihQvQsJXHY2YT+NUysuB
py4z49ATthI/uFMRM8LzFQB5pJamVqm3R+v2/mDKu0MS4S2vc9+Es4x8Hyom5aToukhoZ5sQi+B4
pm37fnyxuhuBBLl5a0ngDUcMxYtkzqZ1TVOraV70VDOzNGb0kyog+KzfvP1vicFjWeMV6zIkpZM1
rFeWvlSTyelHYTuaNqtP+0UUSd0Y5xUf3jfaXABStTL5EqHSFisi0xP+f341K7V7T/7BNMN0WMcs
+B47ibuuTKWCwLHCoaLtN19BNk0mTdIS8LtpvlFEcaDa1eCdl9srglKGdGVxWrh9FkWFh91Jpbn/
fGANRAb7R+L92MsM03252ymUIdUMy/BrLZnbutu2tD/q7QpDeo1rVtoy53R80wya1CEat+m1pFY/
FMIoX8UGyLQ9oMcRPjL/l573H67JJKiLqRvPzNxVZSygCkua6FV88cGcKZH8ZiCki9U/rsrHVo9U
o8GvzQbFwvONqmw4swgtmyr6TjY+NWWcRvgecfMZs4nBvVWaTV06H7tEv2aSnP+g6S4tgl7TixDK
o0VoFRYUMYOkkVV8+jcHK5oeBoookrnWX5l9IcLt5H2ckc52DpYo3qaTQV1HUlS4xW+z1f7ng2zc
+zGedSlZsUg9+jyYsxYokajhgB20wQGU+ZAM292JxCkWdOvlrRYBfsrVSaNznfihVr6vF4v9XrUU
exCnJ53n2vZqn6ohUZI4GW2aAbMvTIu0dSJG88JFZd9P7FfRGkTj0FFtgbzJChihsVO/6SzbLwOJ
C0JnHprd/WB6bL+1wjqNb+OlumsMAc2FjP8u1+18aqGe5+ZavUcputZ6wEjEMd872D39qhpM40YR
RyUl26Xa39rcdiKmrefmkJ2d1uJaxBuUxhu8QghjptVxD1ZZzAdt8zA2ISu89yKwYePooTChxAOZ
pcl/Ayvd05i2wMob8K1r1m85rkDd5Pk20IeXTSPiDnSZlfZR5FpSD6WRXfxq0tnu1n18kowsiQ3n
3IDVX0o42TibLtfFa1C0r8OI1MXDpZvaoUpQDyxFiuf1b3oF0XDul+e0F3Zujg++g+4SzLzDriLg
8DT5/SVCyQfkJu3wYM11ckbaAxRgK7oE5vsFwG2Wie1zvjsJzCPAh8nlcIl+ntkxWrsCCdc/j23F
pK558AgHCrifiiC1noG51GYrd03+wgd1/Ik/XxzBjAq0/Ja48ZBOPpbVtSMJKSB0hMvGY43CsK1V
1+mQaf+lOXR83U2nWOEnp5T3lBrPWbm2+iw/Dj/vq/k8O9f8r+H41Zp+jaB2q4RVu8kTUkzxIREp
iRyz03Rsb86r2V+SDgzBp+Mgkj8M/PA+6nFZnho1Pe1PnRBpJ+m4hfPq1iyKqhgf6QaZCH2+qjf8
3vXgEtGI93FuCEQLd25nfI9Gs5MrNpyq5BPU0r1f61bYoegpccEgNk9LJNp4Dydg9PATF45Awyip
BMnOdn1kdnMpqGGxrP5ALjAqTKVkkRDKn4tG7OMcneHfTIUVGYVf6TAYvBAQnssaJtV1BYHN1cYk
sQWFgR8GfhBpjMEQEod/iAGoVjIbz2UtvhyqV0uqBTc7b/DVUI/EyXLEpIuokn5a+Rs2AcwPfivi
T0CTJnUJLbme5H9bAb73357Ze8++vjyatXY0eYbqqKmXdxhIeNyzlhlCHZkdVMyD4nhNlD6YlMjh
m5JLoPUfclQr9T3sAsMcvTvv61q+tqI6fXv+vwIJaLPSMFmoyKDWNd6KlnQGdSZHuFrKu/XcNSoS
tmcRBvh/qz4dc2lhyl0RR1X4VYXulyYkPqhdv3jFP3de+lW7bdCNV5JihF4AMY5zTggw/qTAX5rk
fA5F61/p1gnIDI158Pn+1QFXJ/0zmQfxbVI6PInfgidFS2E3eQ1J1Hl9s86IxCIWUvOPcMDcVKri
gQUlpKOxapA7kzVzmEyFN6PU97ILRv+UFc76zPT+dSczDlyD8+lS0ClAMve8IN58FxgHRvDYdbob
gCOfoJ5ITleoBpYiUESNRzIipuutCFHDzeHBVluuDYMpmGJ+MSLcOtQWY+JBPqZOfvvmDrEMqYB9
8QWdfwQ8Tp6v9XiDJKDwoUtG34kyl4OQKb6uRRlkxEiWIgxeQA6PyRFfqNrCMVRq6i8AjasakqCM
3eX6PgOx36NaY/1ml82rfQRbOlVxf4sa6Do/xzWL6d736mJLJlRM5O9XQ0xziZnR6QhylD03G64C
kXxI30B1azqSEg0jtXHR4VPA5DfB9OHxo3ZZMK/uETg/cNDs4S9obzI4/Cqc/R5B0ckH4R3J2PWK
EUGGkKo/TuqzsWpUovpwLU1g2r6sj8ONcqNUQdqp0mod/IMt6BngEQRHTjxhm0eUVeVNEc9evFQX
OcM9c+cIc9TQ9aQmP3aXO4paLdE7RC1oBfG3Lz5dye35Pb45Yg9nVeQjmy2yYbPnuUBikwuBuIV+
jbkIvEmsZXglDpQCXsaQly8bOz1SR+E9OcbDeZLT/Vrns5WqKzi9gQprGDBFsPfih9XDvpa5Z/Ii
2oEQQQpB7m98DNi1YAodneNlk6CiQEzl7AULaeIxVSApuyePfzXiG+xrphX0C2AGpy6ri9WFcETa
8qyphGH3OPUi76/9siakxeh6kOLUTcZjFr2chr+82B+XJc39MAPZL0axOHbdig6C/DCrKK1R2Gx2
5P/GZj31GKP6W+2G4BjBGIgPW70jGfqlxe4rLeYHMFhz9Z/B7QffVKbqdci9WF1hlP/Orl0Eqgb2
an1RBnE3jO3hZqdAGY4CNQ7+MvvRR7/Ur7gn0cGp25MD2WV+9COpTgUMSL+V1jkMFqxOKeQ4aKQs
KbFquUkQizUK28T5U6i6Eu/83lqw0e1bVtVS84aGPhDPXaENCDyf2tczu57CS4feUN2W/U1utzcm
AHK6Y8qp//L4pqlffLwlsBK23kzH7+mlbkcJ7kh8teuIu3H7YDsDyDA1uyHE9C8syTDas7hugT83
D/5VtbpIAAZa6Q/hJNAbFlE4C3M+I2X+j6ALXlQHrkoFHedulbXEUfnMSOT+fEjOQXmF/e2FgLF6
Tpl8t7NjiRxAB6CBzJKWM08BCYx1EJv4h+LR8nt59xZ6zQMjalpWos7bigXiia7tmXtxQZ1UOj3h
dbR4+O8I5aptDh+271LsjErmjWn15Xp8JK1Jfd0OnC8dVV4BfC4TSkg9tQ79woLmOz9aXsGF7Ppy
nWSwGJXrh5yd/TMDQSfAnThGy7KQJo9DkfqeGjQQrBJRgTZUU7VtDhH6F64BOUQQrc5j82zZIAS/
U+ypzpCbQNK5Ab0Ny58wA5kq4sW2gOBYSh6j+8vTPt5Ic3hgInLlx5tJcRGP1QyfroV2jSwwRGHY
pQ0E/brZcePfwzF1EeSakhwnF0kEtlbVuUcOI78H5fHYqTUxaSwMAQgdC4BoMS8DxSgERePBQGxm
x7ZkIjw1SJIlhjZ3dtXWg5K705PlCcqPEuk1OMc5vQGScHU4yU9AmYP3U75MFKyCJCBwr9f5EiVk
FUBSdh+qLSBXDV8GlpZ7K7wWknaTLEb8s5fj3pmb58UsUf/glYrak+z/E+sMOUz39YoG/R46z2Ho
cbDLh+mSR4Ki8l3x1gtdUXmqvI9TqQLCp3Tr8Wu00Vf/qRc+7M0mR0Fm3GKBIcHZXJ7Fol39pT7W
Yc/P/8eQPhuzGsyCjJAIvbDAO03/YbZPQ0NBaMfTJ20A/j9qfT3AYg/mxBk/n1/JGquMhwnpyPFf
X0yvMk4TPYzhckL+BtNWWjUEpkpE8Rbs2E1qHjc1A04ZTNF89KJtxs6DNAPZPKLQB3BTfY2g68uU
V6oXfyC1XeaJje1v/imhZTSjyruL0q/+lbRmA/d2K9oPG2O0ALQWWdHonn+B/oZi909s5bRM11Sk
fj/XeEdiVzagu4rARcDz02BKOIJeDhXCW6OVJKJArv/9FEXRWn3midE3MmRUKZ1EvigD7K/scaxN
WVoFJbRmEUl2CgVP9pDGpyDTE9/2D3xKILopU5rxtXfCysX8NBtZ/WCc5lZiN0fNl79ybLqHiS5u
XaCq3UaUSWww9db4NWqjrsjx/r8ndCEyHVLGNr41V09pmEACX8ZKFu2iE2iRD8yctn2dHnEqpHXS
I3VvkMlg23s5xZ7PJmKGyYnDg6GP5pxCmtrlChtwM97XOo8alUWiA+l3e44+QMAjveIfWxTMgiJc
WvMeMEGgQa9Y22uDKMXYfhoNvXaN05IRkx6y8xgw17yb8qjlRcGAVvQm1dx3qR9KXXh/A8ytx/pw
nFtCPaFUIob4ohhHaaYCwz2KFfm6lh9n1DJFraXefIH3BgWgGXLaP2btUTOkx9fBfJWbutUhme13
6nIS78Hhtr4wofRjimgxZIKuQq5umjMJkhw0xwdf6vmvQRfS3xzx4inHB/WASYkQ8uJP4mRJL9GT
gpANWf0uSPqQIECfWYYapA/+kPuhCa9Dej2TnZWvBu2ODX2aZj1o9PuM4r9s40eYJE/vuMQSzPXO
+VNb8ZS2PgQmBRT820p673gmQHM3I5z+xrqetD4G+b/9nhx2SIQqtLBZzEwsBMv2H5uyAy/Fx0Ah
5paC2j5VOWjW94TU9ugH6HPrvOv9yC+IXn7fQF9fuKnkXnASy27inGQUyL+foorPoEtbrQVQNaNw
vAclB9uhKIm+8i8iyA07iN6o9OphWEQEob5l9qtCWH5Jsd3cHW/cWpYdOajHzqdEae2Ivw30eBsc
jz5VNxgunmWViwH4O1pYeaUxrBgtu6aPtOJg41mjHUFzrR6tRSNkYB9yjsuu89YmPs/2l2eIXDD0
R4mq1H53/+o4hMN3YpRo0z5sfLPCPq/Q2/obQO6gQrIhBWudHexeTAcz5rOG6C0RbmDY+sKEsBF+
7QRVoK6H0BWq4rNtEOj/hPpddFRurEoTN41jEw3cHNWg9w1WwBj8dUOChGzi/pythMj/z92GIsUT
LAX8f3Lhvf3e8qyZrBurYk/MzaqBoT6Qxco4QxsA9VdfopiHAesAwm8sixclAUiaTOWKSQ3YQg7l
OTYv04i7LaaXsdpqDfE3GlzqP1o+FFZ+Sqe+ec4TfoOxTIvzWZi5R5dQPxXILKOfoaPOQ4B889lS
9Gn4MGbZkqteS3KY6eEicujSE4QZJxVAqeoDmQxnnOolK+pL4WNabPA5PbBseDyY3cmW3yiKg4iw
bLEHHsLMvSMvdra7Pq196gvc1Cbg2MyU6a/B9y3bpQi+h7nYI0Mt4pzk4LYIwusL1ydv+YmmTwvl
uHIGmCWs+4Za0VjzvS36+lJc5FYZYpQ8f8i7wAu5DKz5K6gw6BxoNSvNunqvjbcfdyp2pxMxZPDF
GGq451oWkMVpOnc+dfCr+nEDrlOsKE3rZ59VehDDf1yy9EaYvrxVNTgB2RzWPsPXCGLevUaRxygS
IyxWbq4lU2tl4cwfeknwjkIiY6efZ5m47bdYKgRf2yOtd8p9Wqa8axhrjmpatfn/vQgB+QwM42h/
QimIkCcMvrxtnenU2JWeng3+F21AnZxwPKFW+iIm9PCFv/ewZKB/Gj+dE2ef/bm10LceFHoUUTBV
WWq2SEdIlaG58skWiABCqVN4pZF4Kk5raMw4mTbr76/VZ2nFvdPapI4unzAaAyY6j7kJmVmnhQLi
NIVGzezKwPBaxYwic7Bq9qgyma7/spaov5Ao0hVS6gVdH6reBU2ObewEgt6p510Ec2ViADj2lvQo
sKyrRDxoxANmXe4vuDOCi/nkfZchJzlzdpDWT8G/RjYpI+FPH+49JRIQdBktIvgkAVapUn/1FZmj
vc/w6l+FXGZzsbvyoOtm4XLcURfqx77+IUb9iwZC5xiytlKUL0rGqo0jLY5sbmK8kVfcVE4N/NCn
CQ+oKSmMv1SvIR/sbMqQsWAFahNF7Be23pzhVWGcWUT6MawNsRu89KfSynw62dQMKW7Wcspt9sgi
dm59+CJL43TdGJyCL6+VRWq5G3CatGEt6BpakcuCXkcIGmYKE+QEhAokBn1VNxbHS4MHOhM/UIOz
ZnRkbedjwHbPM0kiStJfppTKx1/1R2+0jldQI4whFz86k8rWAQ+/wqPmELqFwEItNz1NpX7mBRu5
FazqE24xQUghizVkQG0W37gAGBliAU8ct0RG02bdAUDbbmOk95BaC+Ms6qFkQc+fCvqJQ1GeHtE7
Oyrg6v1i0ca4Ugh17MSruULdcNTIh8s6zeqCUqviXABBFPKnxY9cdRc0gxrXu2Bw4G9gJFnCkpXL
nBefZgGQVZFle89Su0mlYR2GV0mvfVpm3+rFN9WpKTgkBUed3mapoqPEnNRidK7Kqf7Dkzm/17rw
pTO809AIzSHVBB2Qk7iAUF04e7673y4GMr4fjhQBpuMQr1iRDyIMXWrFWYfZU/e9WC8TtnVQW7vr
m1OkBqmm4Wzi/LmmawLmF9TOhOUlXiOiBL29ASdSEiNXmaUytvnaKBY9Ppn+kiOB+ctdqoF5NfcC
UaX0MYjU8KiV1dbPzP7wPhU6P9xJ5G8/aakxRHKnt1vHbMGsewdqRFbkvupNJ+sFfv7v/m+6RnNM
6ru0i6H0fsNxIRqeATrQ/TNdKAftsj/3V8ya13nmGmxaZm+A7Ree9OqkA1E2NkGy6bd3vz6Eopxu
OlfBj+g92QVQnyAAI4xy+kgNdim0GbXOo1GwBPD55I+Pjuyt2hjkjlxut2gjVkS6mcy02MjtxE43
QA7O+M09cKcIol/vbO6k9gMn2X4kTRrn3nm7KW5RdpqeGf43+4OErqWqaXD9hxm5rLtWt/5mN3v6
gCaevTyRIday+N69ISHF9FgmTKqZVxvUznpJ6dYffN7zE5aBwXRj2ZKNWPNCgio6JKoIba9xhifA
ojbY3kxOQgg9g08CiT+L5hOn92cDvuA/JPgsn/h0qLavVjPAf6l93c8KGOutMkxVjrQuIlxHNlBE
3lq1yz5+/EpwF5TG3zXuv/Iz69v0sZcvL592lDCTFw3M7O7WvXXoECe0i6azLKsLubF6ZVpm/YxF
JAYitt+MTgZxNLUcjwhaWfNvGHZFOwmtKWWUOAG52BAav/C3ymYQCbGtGuM7rdF4Ypxdmgq8ZfYp
TOwcr3YKE1sgdTznN68k8e5Tq4ltFbTN6EZd0tAwb9FYtwnhpEjr1FgCiIJ4NBKMsXNIChAwF3x8
02kStVaDKVDRVHi3byTpJReS9eB3kAcI01EsFOulKhMl3Mg1GXd/GTV6j6NdtQZSa5n9mJHqUjLi
71767mgNL64nURh9I24fnn6/MUO/6Y2L+falxySbhfVGL3jT1pUTQfI4p7+qXeiKcihGsivRRbC9
WZjlI+/RkYQGzjT9CS7QM1FuqFzCU6sIfP4cQwsQ06crHTqmFAFPG1CbKP2wwplwiL5o3eGrxBiG
ZcF3jFiM9IdUwfI5wZnOCd+Bctm+IR5VFupSeJTZKLSRZuB3SqyKQOlsGzw+t0FdlROMOogJb0v7
HKFeu4dwc3kzRcU1G5STxv4yT5kKEkmF+MEXBEMLIp19Y1TbL89Nfsf7m2OfkvJDSWU47B8t+4e4
lORR7KbMvd5P5TOteGHfpoOVLm7S+xile7ueFcQaPONJv6cCuI5hwkTvLhIUIOrQwJj7jTwNc3N+
OvZGi5QE8A8BUFqYyq+TZ9RiVj28oKWct6+zcvrDAS4lGh7m3MBy7q6igJIFAMWLRUVR2n5YEn2F
eiHR3zkvHC5F0KT4UvR0qWWuYHzONbAArXdgXXMEV5l72+1pg3HaJY4sCatwKop1fGaEaXupZIrx
/UfUSckerDEGmRIb8d+MASrkinKYEqAKNbgr70IVYA9YrHx/oSllq7S4GEQE8H/B3cj4T+SOAE4w
zsMVwGQFmMdUAJIL3VYRe4Jpr3Qew8ct0aTB1WLEwUgoZEOa+yxfE5+WTqToDJ+ZV2wwcQd/6571
3mlv2DD/GW1PWTXUjeEhHPrbUsB0cdLOpJmYzY8McMy4CQwukXHRoU6XQhU0H1bd+cD/qVkmOTqC
p62Hl0oUFgSDdzRPm/Tz+m8qhep9uCGyIxfnQ9s5hT1h4cgkvv0TesfuqD2LsoTCs8ubzHGgnH36
16dpegOlJi+ULFMA2jHCuQ7dgBy/Qb/rqqnmr7LMGrVs4yE+OCk2LhUE3SRpX32FF6pHPh1beUfk
MGBmvKeZAxQEOqLheNDSOu+9i/F16BELmK9J7KoyFKsG9gmV8XrgASyUTYOMpOp6O/XDM4Cs+eRq
RaFoiJzOkdH4ddZrSUCakBO//TBIwbmC5mwvm8a4XGSF+Depy+UM6KBDCn1xYSRYtH3CT4IFQW1a
CAF8GMYTdi0kf1JWTW58/7VWoMWsJ7bWrxDkxsdGa9sLUMNlJfSfIKVOrB3apKaLyIkSw81Yw8Gp
zgnRa2m6ik5odM1985U4pJFft7qTnvDY5+w9bGBe1sDVb8I8Yn8Mv6egjBbwNtI5s0SipxDUJD7W
Y0yw4TgHMs4vA8YMQEfjWVHKoKGmYuBhJL1gVvKG/pDwJ6257pgaYNIM4vSKXJJzdjt7l2GQAFRR
t82o3dMh1MDlSeVNZRw3FFgBbS6ijuIKdES4Zw/r9lf3eh9ZNY//b4pQcKPzRf5gq6MnYmDjdcG6
GQyUVx8T6sSmnILGk7tQa/bqUCC1XSEE/eA4Eb5fdfiWgvQK5S2rGOdXT1C/nZbTBgsJFyD5YklK
Nm1psjsluL8j4boAF1KPea502BJf8I6yb4PK61bmP6hkzXo3+wjxuaQR5tnbzysnQh31CHpWTwij
jOiaUjOwQO/EF2G96LvW9Dl3bUqVLm2oQ6YV/MjEhoMY26kCgQoOc2KhG+fDmuvOS6cvsMIkt+i9
Bgy/9W3WFK/CpKGCVYaXjlxpz7welFJGrlUZg7c8arsYccF5s7ALJGw5PXlbuEaf9luuOvT7WFto
peOWt9IqhfqcIMjtmZfFeghbakhNBtXg0K8aOQSaUT/WG9oLzSpYP0im2Hc61FqrRuXqZBFX9+AR
2dwSgnao3JVJq3O5nKmtQQwL9847/fqHRe+3MRDL8uCoLB04B8s/HDA4f8NOjjiJxhizlH8sT4DM
8Wbr3LYYH7LvHAzzJwqPnUEFwFtpRhaV97PzgCVkQstrWF41dPABbFbsbDyyj/L1xybeD9i2dgiz
VFQYlucfW4jZCJKfU9dfZIgDHIX5lGGH7brq0IDNZHMHXFk8GmOp5TIxsbZVwRQlfBdcb2EOseIQ
tBd11xTOu5RFGC/zhgi8bXtPY8ag2GQ5cbUFdseJIlK7J5PhPCujSMNw1rRXR8dE218eyaZMzWN4
Y0zh9gj60S1qduvJGj3UqmcbZSk/xgLpaZYPFUKFfT/Dk7VX8e1bYUUTEr4qV+bAs2ChkT8a3+Ov
XJ2GzZLBdOjq5FOvOhxIZFPhKVtXiyM0cjkw5ddOXIlsTW6jXyIet3ozYj37yYEdMDkWl2e36wp1
VE0uyl48OcwIXOqxXRNPT4+QtS6LtbddxMqVUadqG5znvtB2UCnkLnorH7ejJZ6a9Bl8av/VTc9Z
6VaKOxclmSMYunmC2XlPVAFTQJQkiX7x+CUDbjnJsE7Uorvl9nli+jFiW/xs6scDLsHdcpCufRYP
OOxlWHAEh5CIRx/8VB+dUsr/ooBVVdlm3fDKU3Cln/t9h9xmjF9x52VpAGklajmCj3CpL43aEjso
diY/4vEwyIO6io+3H6U6P/wGhruK++45HeCZDAX0MZKf80E/ClOYLAV8ZbjVZhF8bxqLu9pIuknK
RWmVar2uRg8uHdpxcO21LqibYZKRsEl3zZGFMboznynkBVM4rDyYDzFh7A84L3ixCxlhSariY2QO
O4MzXLspwsqPQBfPgotJzGpD6rlfzNMuqMaNhMwkh56/kr1Gp1VULvK64+UT+8SHYxNq3MbpkIjG
O2HRtL+V/cfn1RBn8Mr9167ICRbNiVid1A3wZ7ebtwSF2VemdfS68VJ5uktbKBE8THl/7ViStxb7
f2xypQId4ki0m5WpU6+D5RGxYw3d6GBaiwW5cC+UM+fA5wPYQftKpWu8tf/q6nRbaLqo7MeYav0C
UPUNKq4OTGXWrfP4RvH6Jbr53y04etPUB9omtl0UufvXBLbd+PQ21QvZW2qK0aRSL3KHNDI8P+Ag
OJkUjMB2V+1SBS+0Q/S1UYtAnKi0dTiioDFf/YA3YMt+C04lqJbAQoZN2FCofeViDxHMEp1VOzJm
NuoGQ6Qq/KVs7jMiL9+icvDfSQEL3lNKSlbk1VVzCvRt8sjToBMbF0+m1fHY5sQmLZ3frKU/Uxif
bOx/Izt6iYpvll/sDV5DncoRQgRWHJxbc5TSNVHjNqz7mtTBS2z/x0KSMSHIdC0AB80Ev6woAOsg
VX3Gk7MQdtzTIOL1zLo0UZfuZIAMMZh1LHKdj255dsXkecBX7Us7KYitWz4eEWggOyv+ufgNV4Ho
VYW3T+R36TOZ3Qu9tmz+O/0ex6cJted5Zi+mOXYAP+ZXsMuoL0QYT1mV76gKTWMe1ZZhwm40/oC6
qP7dP3fNdJ8Nh6xx2CflAM3mxZiMIUKIP3fQTTE9uelSOB942xFTzjhJxpynSJorlCOtyg29e5qx
ijgPhIkTtuovvEo4s1pdL/aWLEHR6QmpoFs4QFt7KluEJpQKHbr69VfHndQsEOPVlRhXyHon0SJy
8udW3O12YTPW6anDNddWE25M5qB7EpnnJ+9crJmue/pcFwn3179+Blb2+a6vJT7ij6nf6FKZ8uxx
LdHoqCqXQKy1OzrIq+h4LeBTbMsvthoOPdqzdEZLXxWYXC78gbsxVL8QWXWsA21Yh/YfLTzZlagW
DxcwyO3Uw4IoLPK0ukNKtVJ2chVAthYXt0UiWb0w2qB3iXKCaGcKRMxe46nrtXE7El18un5TuNGk
YK20BotNf97bcCEIG+xWT52o6XY5AxRkRHj86PJ1sssq8dm/pWN3Ij/DoLDLrxSdMJjZFmcFUmCn
d6f++pKfYE/h4204z2Vh+LAMeG8Q22raOBRrBtQ2LkzMo0EEX8bsryiVNKbRObNMX8luv3UrVmqi
lJzrfKHVFZE52BsSuZ9ZYtoFGjC2CdiPaYb8GKb7Sw255cetrY4F1ivMtdspRaOXflHsmlaYASDf
ku5Umdk2nkvzMBrGg8D8t/OFiArwQiNF/nC1qOjNqkuLDIPFQMjsENncGJmgZaEpLd7Gs+74YTMz
/Be/TBrsnXsN80MP8Czyr7ouzkn8H+6/L+FWJewIAr3u5KLC5jcbzLxlkYAKWaRLFY6b0ET9ARAf
Dhb1/BAogPhgMUaHD2xNkL/I2hgybqPIx7inVWx/Pil4kPjz6lLRtDqPU0WpnMo7WyVB4mv7hpvK
S4IooiD1PGljBDUxXH5aKmVrScGJFThoKpbuJ0HhFQ85B8qnVgxxb1arPdwryskTOTSoiwsYF6aH
Zo+zDVS4vLh0YRkFNgShvydjZoNTxP7K51TciNr+nPv88OFE/vRze1OTL+9FUJi6xiwDXp5YM6FF
QnECedPNumqBinMAQYlLXABfjsoNN2KACxWUlnXyXvHHECW2fWrryki87YcdnyHmtlKUjMR8E1uE
XPsirldPq3elc7vOixnxYLVhSApH+mMRlJs77jJgJDerTX4m0JHNou0MOqXIMe+042uGVjMaGeN1
QqugGOrh+Cjl+aS8fTBLeZcjkzkmCx1DnsU50/0bp9SItEEDIQHHtVApWEm/YUURkViF1ZdUpPS5
gzJxGc7vQ08xh83kQ+I8qs0LHfkJaMJVQjhv9nOyr6T+ypwujqx5JHsXuKC+r7GS7uoNCw2GxctY
IDEsmx3CMB4fzUUnUEX38u6U+6k938icxqvnvFA++P0+mK4u14i4xX1KmAFcrRIxCBIFu0QHg035
OwSbkvqC7ZJ+NRuNsaHX6oTghTqpppq5YmD0+F1PdmZHfImZkCUiR+WOmUF/HNgGsZp3Zo187QD1
lbXTGkYGtaSBanhqugXr46M1bfVA32c290a+icwgc1YdcMhC+a3dD/4H1nLyQ2IQFHIVS9uaPoDI
aOyznMo4185NuDVZVyvz16gm5a0b6rbh1Q18Wdk+irnWUbXJRPC8XNRsZkOlt43v1QejpNZSNqGj
Lt2zx9kmERNmyqzehlbqE12QlgmqQImPWTlzKaQuzS7U6RWR+0SDk7pXgCUCQsseCFuD6ALcTqFf
YGL3n+d5EkISuElY8+h8Ga07MvS19wv9iQu0Sd0R0DN6dTSDGcWrIxTFYGqMoofrF9PjEMLfIK7W
UbavtsYSQnKmO7IQJu4u+sK0f1OKVmBRkby/StHn0atZVdupDLIRgJ3/n44seKXsTtyYh+P6B4OA
3utT2xNOFo27AVAyx/w+o1SzK7xHLfxkMaWyIJ2TPzB3cPYGqb3B0fthALv2CGGoHMgwvP8tvHEW
iaIpCJmlF0Bst5whxiosgIDLXqTlOQkvpmH8EdzWIhY8voamU4hLLQSxBaoOD1tFuMl+rmsGdtZB
2kPnT8Pya7E87EbWuwekOHZkZVQU+YBiDDq0AfOqZHq23cU++E7Ob4NDq+06qAEMS6sShEL7Fqay
8FoZxU0YbrQnRcAwXU2liMm2vBadGfUcLI6k9V4QG+7BX88hDSY11FulDsvHTfj3y0yfPX3WBnM8
yMN82QEqXaB2aHSM99m1SiB2l/CWaGhWYoGy6dv8Vq+Q1N+HEIM7FdrHpZ9QEjg8jWhBjtoLNCwW
o3BJj/6yedd2UAKPYKb00M4keVBUTvWB/ySrupn8sq9eg7JgrJgFcgm6D2rTZxePIlWcgpiwwEN7
xDInVTGcVZioY0ph3Xuucc2v94QOAEhFJo0CO/4hvShUeCMscLNWb4FYliNFT+aOsHXjlwv0M/iC
vJcHlE0xCssNB4NYtKBoG/VzGH6q+FEueeoi+12DtS+XqVySthqcqlW3CMnd+UaPt0PkOXjrQT/h
EWNHmtJt7us3t78qh9Ftyh5t/Ai2DrOrjYnLappjtnrhxwkajoPG33n2WFVG/RlnbxvvSTMNETwg
MR8Kf0jZgFJqzaWbwol6XjLa2iMG6o7T5pQ0cRN/xlW8tXIF36Sjm9NE1roiu0v/ALm3eHEJA7Ts
gueD35KWdvBrziE9CEaKIuH2RtCTHaOD9XL5PoTqsu20dbd5Tq7PA40uNncr/sjxFNO2s4eqLyZQ
QYeaIs+QP+kz4ikiNTGPo8O13xbUoMGKo5M/PnBxpKQOgphCqeHtO9+PQ80EmYYIvpRdPmb2C/P1
KrKEgSUjchKbksol9FaQgc6KNO2TiQoms/B9FjF3730JHjTjqlXUDxnWA/1o1CcriLhN0JbEaydz
hPDOzoiFMeFOrXwRlCHtUMpQ1uvxoBRj0gck8pcFuVcSP8ULJlERZ0LQ7AZk2Jv8Y4qSI6msQplU
Ma9/E8+H0StcsfsmnRBzaokK9E9Rr7YdDwmF/6Um4fNwSh9DdiD9RqSnu3SkvKLEvFNP4IOf9HIK
CrMOfyq0pa0d/xI/3slStKSKDxhBU9/Z/WtHIWm9E1vKakO19IhIT2yGfMeal3+n7s9vLrGA7TiS
PZAycUAlwbuEjFyZjiSwuQ2NegmvW4jBcFTlQj2I38VdF9AxzkG5iqAh8xYrAvFHgU7w1VmCciqk
Y8m/kxEyex5RRtW2GWESnEX7l4ymE+d/ecJJmyBu05SEghTJb3aG+/anOwLfb3yHCYG1TSWznk94
P0XpZlYS+iNjnLK5FvhmzuHcePxoLDdlfwCu9Npi4DS7rYOVr259fmCo0f1oJ3hTqkVGAj8dgTBc
uufA6tHe1fAUQ47YGAcnyD4yPFk3OmvKWx5+imWJIZfEnKjMFaEtBIO0+YApGUOd9WSTfPdoijDU
5WX+nq3pGoxX4+syw/o3/2PEeaxpN7ENPCMA8DevIl5rkcM9D4JH/dfwaN4FmRqW23GZWmufI+O0
PgZoGuPeyAIZ0Zcu4x8whdUKvTFgoMeE9iLOqru79Bb059Lrkq7bkHh76dq8oIYeVWteWCFPl2od
bVOvh92t8qH7s2z1CtuexldlxYFSBzHeOlQ7ryh3oa80RFOf4Ned4/n/M1C/Q56ByQ6gN/YMEAVY
OorQIMpyMebRtw0gleFX5e/7wmj8CRNYF4VOmqeXGjBYPYyO8GsVvozR2VZvbb+xYluTt/FXvP34
4hqs5FpeKagf+9QlI6BBHEMfFJDOpYL456PDW+FawZtlhpcfxpQOjPW4I9vL5z0KvS7cZi2bwNVy
QZlHIKEULJ2k2yORdjniQIRf1n2DcuCZ4q9f4wbo5sITS2IoUpXlGOtHf+HcjTquSuhCPfEEsRLB
pW95Hp/c7hHoghSNmWJi0+9+zdl26kY4a3x8uzAHeMcCaHdxzQLLTDoRFbUYTWjx7kqd+xT5Uo3h
6Sy9QKDxKaSJaATD63NyqlO+2pEh3KhS04TaOif85G3cKlVxkh+ECOAPeypUIi7e/r+On6ofxBZS
abok2iillgN/NNL1WweOSKVsxn5RAjwgTaRoc9FJcaTsZSk3gg0DwO5fDcEMcIgu6KPC6hFMMpDL
i4eRigOr4PV13j2x+cSvQIyksaG1Qjyp+aar0u56X66KhgCI6sOuFv8c8BmJbkEvCg3fLFi/R3dh
Ky0A/AUCep8DfD3DQeZQDkIUIgM96boSvV4gdxVVYv9iHN+vFwsKVE62Tf0aERYDanNs+eehobMx
B9FVd4h5knoqiHqn7+KXEm4WyHaZ6l5UPBHl+1Iqj0o0sMamvhntikNJR4gKxUDXbBULxr8TC0hm
wF1itbVwYTcR+QK2eVd7ExOLjrmq8QuIs8qvITud3FHATIb0A39IuvMYseRzNRwI37gfV0NiPyJz
yLlJReJBsKmUEhCvFAncYJfRR0Rnz0uuTLCsSExoTBcd/f+D5fZ/1sCXl+uPpRK73QIgGj4mqrIK
HHDrgaawYDiRw3CkiwbjsStdJCXdT9HjyMGpFNv2J9sqm5FEV5YkxXXkFKEcip4Li8fPHMBZ05Qw
sFZutubKuny7kkusxdfK/evz+LhUodQjcCmd/vOdfc1Hsy5HivRdr6qROAFtOeV/LjGgIyiFrCT/
fWtaoFn3NBA60KYzhRMe1lwwCcBHrp+7/NqWIPLvM6sjLzD4SEDpvXjK/ic3+PSP7HU8etL9+IC6
Y4nMDpyVJWhXnnWnDw9AHlg0lZvHXR5Cn61Mdg4YefNsC65kR4ye0ftvZq+qr1bgprixnrRKluMH
7ZoBJ+FcaKzsH4jnAoGxHjZq976+RSC0ApbYYOGFFIsC2EDvrf7501CNKUk5rZX5VNsYIyAe6MkM
P/gYiJ0IDqcKz54rrFLgO62vgUBLUiyca4so/cx7IqaAiUXpYo9lQFLHHKWoRgdVmWQc7e+fIQvS
/6oN2NjDkNug04KfiYmmA7VpbsSL6YPgRNRVT4+7Hx/RKwkbb7IjC2FyQJxCOc7xtgbbLnDb94KR
SDJ0rq2BsWWaTWUuLZlxlM3amXjJxNRPoDqagOPRAhxEd0zGnYyn/r7MgeIEgadU8AGyy1nL28b6
agS2Rx+uCZS9zwMenqujAJR29GO2/roBoseondFOCBBkGpTRlql6tq3C+W5nwu3RIW0RtHQ4CMHq
908Q0AQtFJCQ3QE/K13EDfD3lRgspl+0INPesdeWwQZQLKgSCD/Ra3xgCFKDBXgV2k13hVjGYPh3
sm9j/oEd6cCBss/6v44ew7QEdOsGeEzOnzmp3V76ujRNUGGcUJR1FNQW8USwyaqP+Q3Eyu6Et1CD
oHftteGZcTonoHeoRWr0GiQ4Q+ZfYDLX7yZ9FzdqhK9JD0kLkp9GI9gfL5EyY3ZpsSuq5OVur2lE
nbFYl0NakhvOzDEoTBpscnEM7MpKQF3gN81NEVSo5dKih5YUfXqbvoQCgmdLmDBzQ/rBjO26568r
0q8k9hyZGRaPaDKsVQavFvIK02FYN/f5jp9UdFpPZF87PYqTk3bwoDV8AdIrZOwe0AdDeJtdihpq
bnBwav/t9u0Mz20Q9OkJ7H4BEcgguJ0pyApbHjjc5Yzz6MB9ELDfnIDVM8sO0mQ3EF/SNoqBnQgU
i7m/cfQePXKShYtKgkjvxkquUDl/Ja5tSSBSctrQ8tEqtdyT0HD3F27F1r1djW1k0Hz+jbJuPYIp
BEZptHxDfvMSsKzBi0axg3BUNdEzqQRDVv3qfO3fyNegZdGFdOpupNl127eP1fnr14MXhNNt1wY4
ScYIR0jHbEYzVg00cis3iRKxZgZznxK7jxKqyHkm+pzz7KLvUu88eqigIsvn9j3OCQyl7J2fQrWf
WMhJfM8u8haQPBCI77JzSZI795dfXwaBBTdBSdlFJCPzBeov4ORNGD5COvSx3Y2LM6TDiWQS0DSA
aM1Bxsfy0bXl54t3cnSriTl2p7/8Xqr1xaOzawz95AXYd970u2ioYvRPMu0m/bxYYVzHkdPD60/2
63LMq98/RbtoFS8ZfZ0Z/qXieVL/fDrpvMJluaPCnrmZWYfXMvRtMKCfi/fLw3OeKjzsSWxFwIJV
B/H11g8MyH7Es1pyjasknQ9Mk5UmjXqmveS3ssRiXJsXe0IxIJ1gvcV85tC+j9yU5/V/QPlh269w
YAWOnhrcbSUynEe2sRyxJ4g9HLKqNWvVjMyWhKUafrgmH8nwR8MOyCGda8QMAyLLrbIiYXHivzwQ
aFSvJayhmgGRlaQAATUHYt2qxFxm9kEFrrbY0ngVayIZXokGXlTFyeU/7mLAjpwCBZNIN4Z8btMN
33YvzqGWZcszxA76S/lveIeEuQ782Rk+n/BBB8o/p23Wb1bb3PAB0zpjNRnEKRoYmbZ3PamdxAoH
9Yb3p6BlXhN6Q1cN427e0BWWBk7vYy1y2iXTuXN6BNxVHBidhf74RnRGYcDNfZQ36fK8LYW/1qet
kT+I0Nj86MEJcv4ZXsz2f2bLYXjUX2YX2xFzihiTDkjCC2/cQAc/+F45A0xQAwVww91bM7hkNojA
Lb2tPp3QobArqTTXmGbGLmiFbO3mP5vlDAibEBJJotTAZ9KTyXyuGLSKXPpc2XBE1eL2vBAybSpx
ojzCCjo8JzkSArFDg1lpBrnjaRsjKuZHZhO5eq6xPKWkwM4yo+arIej21eFQiS+/g6mFxcKhacE5
fiu/lpH9P43lzUtphRT2y40+kn9YXFCGEgUqCWW9RG8RzisxECH6525VKZebC52cXRJL8h2b6eMh
PmGxIGXtZwKceyB3mGMBGPgmDqnZCcLgrsI+5CeFJihWwnO7W79BGDOCqNEtBPPyk2CftvL0q/9+
poHRzOI3KTTnmWgIWfcBLLGpur/TnSI0KeiMFyWQJUSH3hUDMzsfW47Kwv9YpFMFFtjgk2Po3cVC
DLMqd4XnY81ACkVH3Pqt9DKm6ai4gCIbH4Z8fv1UFLbWGTyRTCw4lHpDyuNpxbuAbBErv78cgsxW
Y0HJqEOizvG8VLylUS5oPt3jBL+GgbBWn+JmcTHW4j1dBm/nbMhjIQToUu5nioxiS8wMXW20nEPJ
uXAq9e4RuU0pEJD/bgEwg95I2msLdno2ggxHuOOJeypsQUy7ZULWsENjJqLBsUig+Mesq0UURMCk
CA0fxvuU3gnslEkmTHANzxu/HXuYsZ4rlYzd4nVGY37Q/JYaiuHD/BttAbmyC6yVk1lQl9fBMeLQ
cw6BffaptLzOgZLuFultveNeidvcw4/TS2ygmA0UvGJDz0v7ZWmES8gZZMOy5IGBbFbW5EzdbE36
t4xBD9Z/rH9mknN/kOtI2ORaDAD2JskEoJgHrVEWEfb1S04VjB14FB4dTw5PHBWQD2EiRvXRYsvS
cI1JcEdnwlmzBvffdsA4OXKN38wHZnRExKYc8E2oafwBi1eHPV102yFsnK2nF3ndEFSufpSgRw46
oZYz8lFubNR6DbN+tZz6qpYbeV4CWa9CaQelFtBj0tnntF8DHwTvZLKPDPAcWmGmMMIy3/V8C2cT
Wi8QrX7rv84sgqEn6yTzqq0XC5vWfaSJOdCOK8cM5ZydpPjSz4Xwr7xMk1mqQGqSHfQJwcY8tUEW
VEj/1XuJQlDdaQjs7usVETlrlmrIaYkhJMvC3A6Vol5Iyldwc/csqmNsaiBish7XkIRcOQxBf8PC
EYtgWzb7GuIwJGz+ovofOtRo3i3uXAw06VpV8CqjsTx9BlFyHFIOUJ7lyuLUFpLiVx69eKQFKmV9
RGgXUYVEEFDYMQboZwFDH+Q0BY4tjfbNTg0ToWgZ7YLc54YNs1nlLF906sWHYCCxNq7PKqlFxk+5
xi1Oz1SVwUuuNIafZT+sUrr+z+vOvYydSIb0HLdMY13bDmU4wZV2ZAMpqerNh4mXF9VbsNfSSeVw
mjC2U9EfMLXvBSmkF6FMlcyUQdXU/69bcWOKbtOHrLADTmjGiwZ7DYlKrOiXLNFWvD2pB+TPU9QW
19HAkiw4eQwQayiZLsL+P7gPRwkrclL9A2VYpmPXnOwkf38DHYp0PpZf3Bj9fodgBAMX8tOBzRJN
6xvuzWbx4go2y76yTRYhT2H3d5KylMR5mt2+MVXSSVNGyij8X1xKLp31Ro3lZ9oY5cxk8kmjYpat
SwrN7YpwFhW+QsU01ByBJuBNtXSPmlHX3yydQv3xdUWTDW16aTB5cHQ8dr/AHtk2nQYwwkcBJ8Wb
fOKKpmzyK4R/Do7XOKl5HtwFfTWsm4NOCAQgABnbUldow+ChIoKbYfqknneLBzcxxDrGJAEdXjUD
m3q0GVFrdfeG80GEIF9N6psWecI0JJgfNWAM2ZpSXMeV7qgyNfGqe7ozzCTgcqEBnEmdqEiFRUVK
ElXxruvYLE4Qh0ZxJTKm9HjP+WnMmzoT0GBEJa13thsYnY4IpggEI7Tq88nsy49odfHWQ1/n4f8g
tBJaqkWQDz2O/KCijev1cDPtMzuf0Sl+95sVOicQjBX/AjTbYqwCu2e1AONHrHkbtG6/eyid8lKw
1WzefAFL7diiOfNrc+PICKyJYMvr9H5ohYnDsOGX0VjvRRh1//jifJUEsXxAIhxx2vbbfBf6tNBB
HDjUqTgYTQelmFUk19LML/z7kj49mV4/v6EhAdmKksVNBp8YFQRZdzs7JLME1/+gV56kHpn/tfM+
oPkjt0vBvfn0iWJ87uPf/7WBjAfayeiuCwUbgiJ4YeBPGmF0iIH0yLL+OxVRoorKNuzQn1QLUuJv
YYG7+nE+f1GpozL3WaCBQaUZUokrouUnbAL0UJXoWjCB/2qAt51tReBiTHK88SkxRu3xa36ZkqGR
xLynf9ECQEayySnbRUgqD1kLKlhKxwi3Y3ctccE1+cAZ1tgnmrkfQ2Of3iXWwLzSoDdKO3BYRLqQ
SJrGbFrCbZcaBBqwDuAL2JIQVqPwTuFL8+ARh1W4J+AkeTUQZ0+8ZRFVBpSbL/Y3c6TRmMdV8hCz
wO8MjzZejKWRPd8Rn6/RFs2vWz7ddAcLWsL+MeZObGAMOGPIhkfCdwj60PJyQjCDFx5ED4laPmme
VjxeC5IHS69PU+Lstad6prmUqNY5UrpSH18AiUFr4iqyeHQ+HQ+DJsUOmybhsF8h0k732V0iH0D6
FzRY+FyfKnMHOcRdFc5RI7omhX3weoUISSfcLVMUGO9w17gkR4s/x/ORbgTR544slIyBIY5C3R7a
GkuydGDhsiGzPlaKpSnrWmwvPSrTzpG5/CoKMaXmM0e4a/JqBisg5o+f2+6UekVkqz8do4DKHHi/
6QPO2BTOGY8Lez50pqFJjw6Y/IiJ7/vSovEhKaCwGcXvAwxHW/2xkjMpE0HkVbLq+z3YzDRJJmSi
ijk1BiPi4Ph/iYW7V1bQQAWHIZ+Y77loUlvHOuH2iFb9JMbiAQx/qDDsQ5dmedDCCt0IFoX201AX
UwVKGobGOw59UN+kci37yLmwNYEcju3jp9whYyBVtaTZGPXTcCiVdKFQSYOjpSCBJCmV0joYXwTS
Be4JVZiXcsoDZVTwgZ7dgJH6b2peU4PVMtDzwf40gev3YdfhMLZn+OL6e9Q6AamfQUWlW6TjzmDn
yWs7yb+q17TBxLnoFpg6QAXG/EAYPTwTZUC9O3skJPPbTXa1A6DwLNSVrncyEiGExu7FapqojkXy
l3bxvj+oI22dIAiArnuN0CBmUu1r5f5cAxqcLQOQ0XubWwHiUOvIlMxNm/hiRtvu4xxBpIQwRj0E
m4PoCWeHbZCMiDywZNxOBheYj6WQ/qYv6XEXb8xwILilWPD/gqZL4FHWyyg2pazOTU9fRIhjc+KE
0OOHOc4egcRadu1xIf7hjirCwQ5eqInCknUmYLiJ5lxJUDWNWuRQszn8bu11EGRlTo4PutzE0zwq
XD03xae6u2WRTbwMqeC0Li2OmGs7KNVZEtNn9+iuUyryYiPdqhP4RiYmz3pW+rAmxo2rRDru88KJ
meXrElEBhRLBK8tEAS1H4BSnHvFFPkgXKUJXALAruo4YSmWpW3ZU8XAU4GJrMqqlXgN5I18yjbBZ
/3NrgUA519rwOsoCifHbeJJFUQS/bQYDq3FqRsayluP9+FuOMhxK+McnbsLr+bj4HU2+yplxDJRU
tawxsJCl6XMSWiiFk8Ze3acarD6PK8GxJYMh8DW7yld71qmYYJ/CcYlOuYrAH6UPkHx6KKDWxoB/
pdpfDnfbWa6sPcHYEz5uRad8RU9j8xO5GsCyQmCVw+Bg8ivxOdWAum7VqiuoWj+YVQuBRk+6u1mP
7hLSdp8jjLw1xLUhyLwbsfi0PjhjVelm+FTWHg63uKBi6RbZM6p1k3HiBJFqlUmlenMBbe1tQA2m
fgR5hp5OpDETPPr2vVQj/9bpSsqpvjFeZZHVABo1KsV33HMuHqljntmy7wk24ylOkarB/+fN2kL9
5F/V9hixV4wq7TzcD7yxVWko1GXiW8ACTLkPoUzT3OF6jIcWycak7yXQ1/zEkM/SJS3aJVyiZP+V
I/O9Z2+ZEE3gWrYHMYUXGClwifQg7LtJz3ffdAah4H8+BacpQjmvDP+7ZB3CvulXgvUXjgykm+fc
9UG2xTi/vbLz8n/Hjof7ZT1dQPgrwIWKKcl7sY6uilds+bRsMURVmcB+jqhNEIIEdmN0xNByyQUp
QyOKH/qCw3D3AXhcggVJDc0KECpuh8oXxPEOW7nycOBN3YA35o+idzejSNurCEnmYJPWOAiLFaqA
+ZQy90+68A5QuGTSyAO7MG+Bea1+cLyY6dMXng8+OtzsMylzhTuwRjE7e6YpcdJz0MyJTggdXmVH
VUaz5YfGWhCCYxn3RSi/baUkBlHzHUI7bw0OzL27JpGReCcIKnvBJUyLsBNCSN15uENuCJQKeedZ
RmsdcQQy3uegPAW6Qef0ayW5WBoF2urINK8+GSyYEaAY7Ajbe8387AIeVN6gZjKRTVQCXzGNI0rr
Wd55v4vXBKsTWzBeU9KhV26NROK4SsAXTzXzkYrJDeIAjD9SkmLPWfHU7CCOg2vv359cbasdzM05
J69zoXdyvYlxNFeJ5rGpwjy4PlOkbPWRxhl6tGRZ8jnXuL2OeuqtTvqivZnZQczEJB1VslzET2xg
hYbXb8ehINLr6U+p74OjvkK1ZIN2Jco0/xgdYj8Uc9bYP0qBFiBEEAdIp5n2D4PUEoq6F+f58Mqt
K08vo/efp2cf1UeMAy3/5tJfZ5nPw71dbMt0XJHwJ+/0dbQ63CNQcGVXDBSOmtr4C5W4L7DMWruS
797/OXnJ5gz4IU3HI7Q+jAplpgWNtpaThHiwCw6zH7207b7x19CL6BNHkCx5UaKdjA8/BJ8pM+sY
kVpCtY03slU+9osfhCwtBHvyVslKH8h7uH6BvLlhgIRlpLyihhv2fxR/6p0bfpwAu19ftauhqTKz
3NfmexhvqCTi33HNuJJV3Kdg4Mw5NAAcu8VzCHgrNrAQ3e/pKVGpx7zQdFx7gxyhugoVFBoCBxDv
mYXoOIqAr0//MRxlA620xadMDM2UOBwh1vsSQ+Do9rEKn7wAMSqhPhznnDN+tp5JH2Fx28WxtVx9
EQgOog6EOaauOQzkna5ttpewBtZ6UXdsMITic1dJLub6x97G1YRaEdrdwLN9Wku4OXj1hcvSqJes
Si7XedhsuSWSuagtJ05qWMfRoxiNMfpiapkhoKdGHkVepgh+LDFXaoMeDzRm0zqPc9VGPbiSYjAS
tfD6DojRHpXQpCJ2+qg0QNj1x/SoSbHCaIKipMNGgr4/g6kEW+/cM+sOoPTndq1HJ9nl7wYsvVGG
qkVgyXWXPfRCtHGhUESk0vEjucVpIMiR1HDnnMUxlGYz65gfiatYUg3IRZbtNpz0YINHFkqZ8B7u
iU94V2f/6OXuYJ67ygF29Wkkh2vOzTJT3rF+6V9QPd04/BFPUbhFoJgcjtL+BoGZ+FW+7WPmL5rn
yxTiEjt3yEjd1Gg+KDPEMek+nwi7sjYC78rNdY29sK496I6G7tTEyjShAwabImL5xa8U3UJgTecx
kFR35f8iBIgT82elW5RClI4umqUqkm+qRcksNvGAhUf3KxEwjNbi2S5LY2Y/2dU6qUJ/YkFdJMsz
9SRhg1R6fZGTuptxqVviK1MdOTfw+0+Z8FtHM2XM3IPUWBfeAl6OLEbCOysT37MmsugH/fGIGAD9
wyOGE+KXOg8F0L+79y03AhyXwjHi9GL2cnmMrLBlTMqID0tmQT8dODpx9E7iYGcY21RTo4GmnGMs
PHa7+E1mibvPC7fjwBz1XWAEZJXa50dqpZ6kmDxQXm/MQmKDoNPzRBGJzPrD8LVwiGpl1nbO9adV
e83ZCfmoRUNrlB87dJmOdIqSZQpSE+z9qIB0jJf2Rr8HldOLPUiMnc6sKcJz+TbM7FNBCA3G6SXJ
JasGPadCslRdiDHq4FsQHv5jafK5G256NhIwriJKdvIIkM57pfJtJwGFg6DrbG1/dtibrsfIjXY2
9ZLpiznaaZhIpjzcaTM55NNVKA6jAY4cCgYG8lrj1PRqXbB/IUYv3r/IegjIK3Ykwxbq0m7Wvdvc
IuLjrzVZXh8jghxCShvW8/nNzxbSzGfbwewwzE4qUJAq4PyYtjjoxpdZoTBunsz7fW5EoxZwHleF
4ckoa4tW9I2cBnpzZCbFKiy9sn/inE40cS3UmtHEIUCugg5HsoIek33eQF0fe+9Khf3NWRVa8Y3u
zm+ksAT74aukvTNK7Mq4LsvF2wNS6mrRMD9NtAEVTSgNRMJgFSPh8c9LMhrpvXlGJ5SPgDv133NS
iqQm2UlBuHT/vRf9bbpdvZloQ12U3mgH1lplBx49bHMs7E+dYFmker5Vw0zrWVCYOZp00FXwkiNb
29okROc9iR+mxSNV7vZwR15Nt+f1YfgIedyNi2zQ1/nheZkUcWZlIcLu9+pK7+7P4YUwCq2ll6eF
Z83Y9gOm0wYlriFbSRYClePzYbLZrrE34Fm7DZA/fN3hucI6c8AMclZRZw0u6ku2O4wBtZCUDe4r
EEb6XCoREWFhDyQNL0X3RucjzvkVy4WsOtTsMHMtqt7JywOlZlexTKfGr0Mmj3OZuJJLe6FToxtZ
KNkaI1gLnLUbUOGw4WbqRiRtOOzT08z6DvLq58qrHOykLk9NqnyGGvVTDcP6BXJk9gy55dWpQTt7
mdxjbh4cS2qucngJoUhAFs8HXTiJC5+7u0OQch6u1IRTzSoM4q9+Y8lAjYd5FLL66UdKOxp2f4gI
TtWHw/PqarVbZKuAHt3kN7hjXEaslcpqUSSxj5Y2hKWgG9ucxWsg199g8vPnG8oTWKD55x/VkdCe
yi+kgz8hG07fG9+JcEEhewANHYfIQeG1TJdiYw7DDsWUVe2iwf/Z3peJEAEnep/LHIZdA3L4CPPk
eXwL+Ktc0AEqcC4WRpcvjJqtx/67aBja1qh3Ek7hEmty7Fbhvt5TKokN2JTq3NDcJ+urQEY3glQ3
HM2jXnuyD/Z4KLOnLHVTZWB1wrH+KPjsigMOjO+ZMNP21hHgt/aDPpo3njLn2551OqA6rPwYTZcN
nwD14If1w7cyfnMW3RfSTX2I6iRqh+23+cjfaOjurVMtqinglwVauZr95DP4U78jwfBNB2zm0mH9
wvh6fQBtAg6AfLvoE0NgCRIysN8QiAzU57o3Igh09HsFxwSOuoaV2UbjaHRgTDifg8ZqIH2IE63c
kW1B/YJI4Y+6IMeB7mmambrG8gYsQ1ZrFD0XqMx5LkSkqRqExVGZ6qzrcctprM8MGPw7L6OmYAnD
Qhu79sOM5EXZsO/jg+dcjDjcspkEiQfhosZKHHF2Z+FZ9ymmndsXr8y9zliNUWjxSS7VLR7eu0He
S6fVn+jtbAdHj+R0SqfLyj+p1w3Lr2Ld2SOPQu7ErLVw24RsRQKhrWyZwybYD0XwYnJUZjRFasgH
590DmMXPKmwU1A7d95aLpl1+QhCCSZEGhBzG7liJMEC022JOmO+bIEwVZJ+61KNSrMv1oTPr0ntC
FxA5lF9Oj5BWvBGXki63NEqDzCBZcqxL+gze9qcBgcv9Rr+8UA8K89ne77alkJ/eaHt/Eu7eLSpM
qYEBSSua4chhMMu+hiHvBTrLJ72SOQSc5P45/bBBjY0bjN1lTvumaYy5XuLs9DNsahhBZHPHQv+U
Kz8BgXbFX4EoX+RJ6englAA6VsLUm03QsHv/Ar2djlRQPs/s5rTSaV+vMbcSinQ0y1vs/pscdzPw
VaamfVsWbF3Q1RioYNp0Lzvfu/zsOKHqUHQfGJhA/iMk7rrS/77T0ZFViAF0ZeecQee7tiXILtoX
VsJi2Nw9gujdnt1BS4c7tgj2l8vdB7UDS8knJIaz/Bn2R9dey8Drgg346yfnop6j9ChGJA2Efsqt
Xgd4xrzvYx2vUTwsCX7WZ3UqVXPRqhPZEkd9na9Z4XicBVVagVcTuTp+glfSXjpvK7Mc2IP4xjGr
8/fM1wljlbXG7rkDFM710jsk/Le3v1+/Tq0RebQfJj6yQ+BDu7jGwl99gfmPajhM4t1+BYVp4/9Y
Asct0D36XIR5TERmj7DMZF1Buovl/QZihkP3Gk5cj+9TXHVxRFTU31Uu7JkHubDGKkr7I7Mewjqq
rJ1ZISuycHQXgXiUPgOMw5oh23DdcwrD89NBQ0n0sovHwmQgaJzr7O4wmQl9DWxVe0BgNJhh+OON
xq/cwZg/wDBpfmfxrJrWbKojJI2Zv+cEL5JIvMLOJNg+9jPZBnBzEc9UsQAOtE6V92/mRNIWCw5c
oQyQIJrtKuoGMmtmyimXxZARHaW6MaP3Vk74yWbrECtRqeANdy5k9ET+7FxUIu2ngcFQKGoUhB4P
xxKXKT+O6H+sDrYqFVXDbYOtNQMKuFSG7N2k9C9WATebKkedxBoZL8epTw9nuc/fVcek+adRG9Xe
JZ92x+JDALE8Z9a6CFi91RxFjWyCLSl1N846qVDs0hIB+1hk37zQtV2iiedhOiUOGaALNsW6/WhO
OJLg7eNSng1W4eK02XAYrGFlJqTS34TovvvxChfXnzy3j8JQky7En3/dzy+3daOYVjzytGvTH6K6
7/GFHI/oVma3g2437BXhWGpiO0dBqtkrsxHquFFcVU/JyeaP2mFg8B9wBCpARuNdqrGWEXL8JPSl
HkB7QqrrWpNxVgANpedzrCTRWwAhZVn5n++xuv3qdmRs0AZfptoS9O3yfTbkQshEZfSkTC3FCXP/
4mOeMAPE2VXTxkI6+Bd5aFA3H/4iHVofedNPPxZU6daBO9qpOk0rXXtbE7zkuhPTVyS9ONLkeqPf
5qlsEe0IDSdYgMYCXrEVxug/3IGiHxjyQiLsZfu3isNosASTWqlDLmvhMXFTZqwkBVwqdCGnqFVn
/nxJhW1IYkdfndYEHp1wl9aMIAvyAdEDxg3zhJwC9r5pc1ynybc0pgfoOWFRTC5dW5kQZ/kim//u
5ux1vuoGu8sfTzmBB9pbYIPD9tf6//wFgQNgqq5gKazcAjQRVF/HF/ALennGSaLFQYzSkow1vQ06
pfz6xD3QsxWaOGLKsFmedEp4cbQ3C68zgpXr9DAPNVLQovFJqj3/UH5Jg5gaW4UMomUP9wuSOxee
V7bmG8EoJ/FSLd5oWrQBwYCG+rpS9ufGzXzdD+YyCzfLdqC+4GwjRe26B3UpxbZhfzSqzLCRgg+h
dQb2PBrn6TeL8zqFSxPkc98Syi5jbR9GFXyt2r9C37JP0SfR0ysV4xeneC1VOIYODqAaqk8mPSZQ
uJCzWNIKmvi2Rl2yxOD533TuhkkjqGtlS7Sj1wA2BBz+uKN8PSQsKDmqNW0XzEOCqU+i9OflUiey
u2xMsjauj0A7CuHh+CM2EyGHj8kbahByY3SlmZmTp/G6Vl9IZt1k6YLQ9GaTM0MkFHJ5GewKRk+8
fOHb+MUFPn98490Cr65p1Lg89TKZtXsPZIj+iFzPPlmhO9Dyp5w72bHLekqfTHCy5fyQeG3sSrSE
nQ/veXhg7onJx5O+QUgts+io+NmwfJdNWCmSMpUNa/o2SzrLogexMdzDSZdUnI8znFrXPhGYyf1Z
S+y+XywSFlb065jmBaNwDYhyS3HR9Y2CYLc5YhkdT2rj1YGTrfqivNSmEQvWCjM7uU83ra8GXsjj
mJXuJI+Q1oiYeUE/xULMa/VY88mtDC6Go81A2O+7o+Mii3LxmbTnNoJWEDlNEVD3Ep9NU1spdAyv
oQMoLgQGZz0N7adrMGBNUp0P3CnwBnKygJMPoHFFze/NjDyMxi+futKtjTOpU6rPx+33qEZQPsER
fB9naCKg7x/3eqSsAoJAQW7c122DvjNdOAg5ajkw/CpMx6Kb0kWHOqx3dxdm4bO2h7XfE+jqMA+c
OX1kMZjnKsv8vZOb4PewLdJpGAbdo/jAVMLSmL8LdkD7USzhEvAi1Ujvt1sHAFf6cSxS7QkKaYDt
FGHwPTJ0zYZ05Akf+ah2v2gKCUZ5oNqkcMVAyYDN+jbZ3azlSCBW/ZEQZh8Lfb/qxpcxSyfvsblr
W8yp7vmrQF1HQlcrKMovHrxJUf83nt/cSBne9uo1JfRdRkcUFHlPDPNKGW/FM18LXXwudynUQkDb
2QcjiaF6pmOMTGa/fF8yT3BqKDNBQajV1rgweo4HwMh1QGoBlMQBB/o5MYjY2YQdaRcckGucIjFc
vBjQSkxkf0wm80fECkhT54xCW149KhKAknOobwRjo21JjDu/TjLez9TN0mqlU/D5Bx0M5fowE7Mm
8bmovuuxireVn/rnagkyPH5o9dNNUhoEseSosiKVjQrmekmbyqBWa120ukchN+SuXLjxZUnWu9qR
LOGPpS6ZsoyZd71EGFRXIsuGm649A3qzLINNf2rwvdWly0NoCcRl4ij1PB9A1DcXvjQkm5dR1IBM
N2wd4MjXuL1LaMiWtug5osweXkdTO/PVxTWUukZzAQp28fkG/4sc1063uTcowye0Ga4YjozPpSh3
f5QL4dp8dajhdbA3/t6jXwaXUtGXkA7mkvc6DZ4Kn6J2xnUVoVAxD8Goe0wkYWitHWf37rxLauM1
0PkY1S2/FkhoEE6gCD+fiXhw3zZ9b6ugWaqJL5tGBgzijiT4u+Djvc23hPoBnaKi39Iga9Wm61xX
4M4xzkVqjozIHpRRGmPBhC1ChlFvzKcR+EeZRk9gdFykHmn4F084IybniWNIdQ33MaqU4XfyY6Ai
Sy3umg9ZQ27h1IjYAKORrFHnEcuNNHnXl9hAy68XIsIl1lqsPB/ivr/xDbmCt8zL65HN0T92ml1A
u5lOzsJhGOX+a+x9B5cXKzTEHiahFV0VCJeomIcm44fknKOfLZJDJlUiOc67fKCvHn/rUYgwiGSu
hlZA7TMxwQ9RMyZwy/6BLwXG+gxDwigB4k0NDCZGMLCXWX2sK9KEXh5zJoIAV5khGJwGJjbUjJNS
v/nV+YtPPnRb4wzL9avHBiaM7lT0BWzWlmynMtXFJF/81A4ut8mALvU4ln14EzJ9+V+VysJeI3ca
z2nzDWsZPUuOG7R+HlP1Gw5OvTEEDWcmErdMfANxfMX7Ei6SRXZ2hCje9pSojhinHMvayP2tPQVX
mZIuLlG7lEOrfR2EjfPFy/L7o8D8m3RUavBMXB3LfZIoIMbNmePVJKT7tDkVtdUMlqPYgnDMIfCk
ynEofTPnFe0zm7vIE83YolnvNVTrWhjiB4duLqc+UEmkZupaUxk6s54TUMmbPIjtwarn/aVE4w1V
OgK/F6VbNvCgW7emH/l5jm9hxQ1aLAPOibxNOg4s+J3oXoBZNZ6v5VbI8U7m0t3geKmFVMlGLi02
DR1GN5FUD/gRFN2Jrk+/pbH/jdyONOv4ATeFZgy1/xoN+/NS4VwlLqRiS/IUORhcOslpa/BoZZGK
fSga268+sasEivmVbAQGWP+JWYWHZkVOCHOPNqp2vtAcGp3eoNnuZkQTcvOKakfG4LT3bvTa7vHo
+sDDtO1LTP+D4+S+nfu60ojzbrj4Ic5YR+LIbJLqmJc8UOrEiOfjWGa9rvGKvG2JyZHaEQ5Iz511
yPFe61flZCGf74obEb10JuFIKY1nA28iehA9CtySt4+heU+UI9VPK9F9iR3eg5TI0Kx4g1udJhYW
aKYZa1mgh5hHNFNNd6nhnPsHmxLZgGmx8DzS0VEaabXBh4M4Z2GgjBlQySi9kJlh/Dz3GRenKDxx
nHTbopso75WMyB6y/rTBBm+HJuGq+3dI99jFoKRRx0UOt6kqcaR3l7r39n0G+NgoTlg2tbqZtUVz
DnhAI5deaZFJqkOLVQzh5vHPfuZgXCcj/st9rxhj9A7Tr/py9aGyUeJmkLq78WJ6r803jKma+C0j
fqQFjanEkLL/lD/GHrSRWCbNLX+0iQNJiD+AG55DfubHo3ECWDmiEDPSsNyORSyro4i0trU/p3cq
yVckWPvojm4707tAZnB4A9DF4d7OAnekqmnZRDf5RgeHoremx0mD4RBrKrtSt8G8vHrliZjH60cH
D9a+jY2yb1QWYyI7i79cSMOEIxjlm8b7l2kss0oxS73vaxhSN5IMQMd08OaS8O282v1/uNPDQg6l
8QD7cWS/L5gJxRt2r5mS8+IuKHXvd0KSl4QmalXcMdokzvo4zVM2qd8YZIec0K95sKGsfP0gKP4c
5c9L1VpmqJhabPzgqZfUA70kRd4HzaelenbLN3R5dUvriyKk9zeYULsATIqiUHr4DVW70sP/VfVx
RAhvIeqT2uD7AEonBVxFf+NtCP/aCUPA2lU5QVlFbQZ8yM/yS6EXh/1SSO7m/vB4naPrRxg1z5CW
BEgoVJmZ289OLDpbUNmySMYhWFJ+SD3YxH4+R2kVRGhttA6QFVWZLl5y0LyJRLaIagJ/uMomgrug
EaWqQ4BOp3SY8XMewVloV4bB6ft/6QhaFVFUij+CQ0/mwklMEr3zx9zzPhzckqQdDsZrsF9M1k/q
D5o1xp/GFlZiWy51sAjlUJqNNctJfTY8peh7zW1QS99TMItV6mH8l+Zm5bYLFRr7zNxzwaUXNR/d
44olBPdAS/GMCV4oYJjUvfDIriGfH+V1DwzHvpL24NCXaN9ydpm2+ppB05wXmdKFcvtpDujmmDmj
VFQvt3Yrp5C5lhkixiJ4SNXHJyyJn/8MZw21Qn20UK3udXwnBXa10nuWoAbLHRyF8zj280wGxplD
pQ8+jMIIOqiOmLlmIQWV3aLL8aGnG+YHNHzUhveW70QnYfBfQCJI1w8do3b2Zcbo1GCU5COKLUDu
qebjh2PXu/2QMDuStjtd3xd9b+8VXV1qfru/uV1Bz8qGgQ4x2uSvhs3Lku4Oi6YZnel6xco9gyFu
xTqMYI8NPoWovJjzKbvY9rinxYOAJYnhXDCs3dseEalSbnQXQAWpjhj/QQdl15Sf2fMF1IW7/Gh2
n77VebYz8JMMfjXWokRZIHrkjuD8kXgm7ssL5plde4xHwKKwvGNuc2Nuki4O/YIYnbO9NdtD9ylL
6RviyI4H5jLWSIIcqla8spTOHmRDuppuu62s5kGnzWarwsa9NIWoO7GlUqVcGuXkiDcrfmd019nE
MfTtYpVGtmLHXRL0l5n7M//cAf/gQptiYlKqezKEbE+T4HMG8NI42JW/CarLZN2yuHv5uXjSUu4P
Z6YlunBAuTqtoxu2Fh70/XSdrGTMVQLXWRZtpwYZRJr1oz4vMQjYfd+Rqv46Rm71bVblL57n14+c
I1xz9l8bugKw7wDA9QOzvMhON2B1ZSmcjpXiw4kinSyMhVAkYq4+zJADGiPFBaeboWsqusZDbLAK
ayQEBmNKM90Vhlp1xI0275e9YwOa/bCdf21rUK3w+pV11RRKDRACcb6d2p9cEv7Brzrxd13olXIU
OFD/eZ1Go8KVf8v+k9vfFsJ99J4PZI4jTR7KHso9Cf+CGu/vGtT9QDe+VEL2EWmD5a41cxJR0diP
wZKUslOlHQe9cdr6Pcfevq8FUYcnubWnJCW8DxX3nwPm5gNmACmRgoNiYuVbgY7UM3mKpKsZErfe
hwVFsT0LCmJswyMFOonrOuTfosCCZpsySY0y0bhZPFoueqiT6ZQybdRHkVN9c/80aoWyh3G/mzEJ
6yho3ZGJFF85GurPOCHWdNfg57BbyxZsLCtHgm/Cl1wfTWqgC6lh3jA7cp14sXiwK7rko12pwDvK
0LTKP0rMX+T+A0JdcsFPDrTgGPfhAFg3wgnLhnh0acE+dx2ocSY356MseBpSO4f2j5/l4mW1V9D/
sYF9zs7g8ranW52MSitJis0UuHqOu9a+8aWY7Rn+gquyURo7/xJvsrsU2TlBeCZxkJGoDAvzdlbC
v90adyavmHf26B1sG719MlN9WBnPzp2LkoxWGxjST8fFv5LxmtVPaQCqnQnLcMckjOc3HqSVk4kk
WrksC/VSmP1gPuf5+4hlUkcBp/Ed6LMLqtW4Y0yjokAieM+AHTv1ymJMyJqm/abm3F23wkY9iIsn
/S6am0+cyw1LLD2o3O46rDCqM9VAuAHBpeVNaDK+s54PPpJYInisywQPVrm4Oj0XOrGWGWLq+qRJ
KxFVfzMIjF40P36RnD/+m7lnPH/oySzQHNxhPU8OrG7hDsvvOjF3KnuRSN3cQaAvq65cO0mydOEt
vgNbP+o4msXZ+jy2fyhfg6Ohnp1N4+e7EH8yRflsS5XVxCrsRRl5ychQG9ZEw6q4K26BmNg/H3ZH
v2D3beTQmZOX1WHAghsuFAtF0Tob0JEDfWyxb4G0vUd/Scaf89SiAmtt2qbMPxS25UCBW4Jcn10q
BrAIbzzyFgfGzsyRrR9stsTYR9cVpSnvb8B9gPk3L+gY15xNoo+ZxgrEeVlVFJ4dRt9bGD0WrP0r
dmVaCzrBGnE+A5gKkyGNK2e/wUQvEPUgsl5eeBTkvfmV5xaBUEpDLudUyqD4lZG56MFikR/NSW3q
jo0sD6W2wbzgGJFzdsWL26FQUlAIp/oH/4Q80e6MQPmweUORO3JwuCAg9mf25pKlWTr6UmdTsLfh
NnmLkU/hB/x958LjFToN4QTI2KMqmgP6VHq6/COe5hbtOs8I4qYkMkzG8SMV4tQs3CRgj/9Uop8A
IqQia6ve+wotbYkeGoHcYW/wFKtQBdE/1us3JAXSBXiOlCfSbaZLrTEsQkBV1873WOKTOgcjFPFD
qLHgTofk5V19P03oUPxidiQcWQGhwj6YntolLoZmNQoe65a1LFwRfADiKWCxXNenB8Ipn5DZtNen
NKKE0oyyDDztYJgkCgomNX61W4039CG+aAOpp95UwodPAz2zvMsFKL5+9qybBrelAB5yHWoLjv3T
KL/jr+yzen+8SGBFYVAADTY3af2fs5/7nikiqdKT2b4cJslMAlIjoilqFiorZrDxf2jISjjPDvir
4gjBoL5G7Wk3bhRo2tpWACa73W6Ml1VZ3Ym1g/UONaLwByBoDYx7cch0+jPyHRtWjwSqK4LqN5B9
yhX6JZzLvEDqxnq1qOBErDgQ+op3vPu9h4uGO67OSWtK64yDCbTKNYNyNTa9PJhvo6kdj/V1+ckv
q6+YsVJrAaTs6qZGQ5sheJp9Gx8n1nJGAnygqSGn/l7Sde4DgAJi3IBzv4k+ykNDvYlBJHpoX73G
HTems7dtpmgg76oOCJtYq68BYX00dt4TIsH1AJZ5Jr2U+1Rx7yCvjZoGa26kzKGWv2x5rlnf1QaG
7PIuEtWYgXd60Z/OVCvb/5XGesYX6G1EAlZ73ZeY0nxHf3o6A1ihzjvT/D3Pg6s+Q8UY7l3UjD5N
Wxc3+Hk5THSngU96vukhmWpXiW6+hzEgbMmXQbSxBhRoqVvhlhIsVugqETweT4mlSSOJYh+3JKC/
oZrQI5bUM8+dwpebjz5e72QmeyNRYxbnt02jl5mmogrTsE4mtcAekqNwT7mGrxqHYTAg9jcopfqp
THZay8ZLD3GDN/LIbdBTVqXDp26NN66VCpmDk3Chv1XrYuLXLdbQS0C+5KMr0ijfxvso5T69sur/
wygZpYABdG+pevO/mo0LoZ8NPPm+VpI5dOmIlPV/WRK6wX1AXx+iFHgOzHLFvdi14qxW8V27FYOj
8blIK1l8L4P+0BorfJvaQ8+kdewQ3Jn0rX2pc7mE0EcpyZ+6akvhAKodxZa9AOK6bWeRFurwtsto
WqFaPijac1ECvzSEzTnDA+HTJ2YGEeqP4mwHPPitXhRLb1MeDX2PZ2Pp7RL+R32DJw2hp6QbKdIx
WoJxQ+1GJ5mH+zRcTxtwX0BeUFXzNOFJmBqwOAZX3s7rPxn7HP8VttgO+uJmdzb5kiFLpv04yBC/
FZG+6UIKB7mIxMijFrMyPcC2tMnkgYngTMinncqWtHOESVAjMXyDYzDFvIqVbEPUePHguJexFLOh
bQtfTxoyZhvWlA0gWZPo/MCqVPHonPPmsmVxYBrBzlIHKc5rrqDGtHyyiVqe3ekLPyT06R7qya2U
DsWoc8xxlD6I2qH+ZJlcm8D234CgLcvp1mz3ad1allLKGYdkMnETjsA1qFfxINT4Y7RsT2DdMNSX
8l8H3wQf4swtl+fzLEgVdTscCWcYfsgl2hNYox+Bb0ZdvfGscGkgX5OWCh67mgJLoJZeeoZU8il3
jxARhpz35woWHIMYMQpXinzmagSYKul5oiXw8tqZN6U3UIsAQQFdQWPNkyZ5C7bRwIiJhwKrXCF7
M1OBxz1sfnd4hf5JIp1Dgi0o/zBcQMb4o6V4qJ0sevtYa0G6zt3zPmOshYHafZKKOKLIQNWhOmhD
IpWan6/U50H7+k7SeiliWQFniB5BCEDj2RET6pi3nx2mRwSY9+q/teNiDd6Yx4OxshxAopKzLoKO
kl2RF9iyrP02PFFi6gpeGbyXR9f34BWBPQjjj+RFp49GdXz3GcMSWlTMrNSjkvg/CdJ/uiNN97W2
9ZLepbD6DhPesEYxPMC5aELCMirai3B72VOQ7axXsbIL9q08t/qPfxCIHYlxquvpVlQ15KMzjyKt
pGWo6/gNy4uPOCP9Hjh7FAZKEdXJpBdLo01dV/By53c5OY56JDFuHwbk5ieSvBAdnI1dZeuP65xK
cgndxBdiWtB3SAyE+XEwRgYJfYKS9Me5280XSaHtLVKwxlFhM68BjczHKmlB3rdRIdbqbjAdxNIC
Vthi5fg91lXnrXN8eYXlQXAbEK2qUjjzcd6v3pTeVLENAOGS+PbTB4Fv2yuEbP3Yty97buOw1jWE
IWsmlonFKvi74D9uaqhEBGi0xU/JOSW7+oqwRTn5ydsEEdgjnNYoE1MXBwg01tgRN1p29bSJZz2Q
Z+rETXNJ7wb5PgjqpabCseiocIiRtMlXyV3fQKh926sZQ/xTDG/Qj+BL4b8ScPnyfyD/MglKA6yC
eLlZpm4X1nFAKuG0+sNb9Inarj1QJGCfm0jYXGssQnvppoySpJPUkLZFqAe73RB0+9kvtPt/tllV
8cfuJ4V2PlqgqmP5JUBWZ4sS3kegpCKZbWRsTnSkn0uZTuGwxhSU2VVlAPeWE5GQlslKL6SptQBo
oeKtq6rP6GPi08vpdTzg5Z/JHRzG3OK3ViHtJV227qGMPobdfvvokj5pIhjnf4SluKG8SgJuQot4
Schk5TX6hN/TowSDyhstl27W9inhouUTBy4MC9iPVxReqxvKwFROeuSn2Pbf9eXLVC2YDBoUF8LQ
zqXBl3oLOiB1J0ZKIQZswTwXwN+DH3Gu8PSvfyQILjZ6h77lXyp2A8hYNVgQZ1wUU8eMZmRRFg9s
yXClnH9FvkfDdP9jgd3/AYEs8lgGIJfWai8k0amSahYaLElu7NptdbBfVNhr1Q06YYAIA1Jfu7Rh
ThzvWDWd4xbT6o11iL5+QM55b6McpiX1R1xVB6YhOjyr+i8GyXnLTwUW2GMnliI63thNVhzTLqcy
o5DkfLAkAPpdqw7G2fTGQJC5sLpEzLOC61DJx/oguDo79GoyZj7Oc+OfP01OS8wgI1t01Q18ps9C
1bvouWYonE0WZ7sQognj4AVhU0rh7kEiD61jAq6yp8hyDHRAh+Zp2+aoXeGY8EPRx1e8rJs3fSDf
89K5Fmi/fNRQBEjed4H4+YooAFXKG/2FzsWm+eSdrdKzd2zw15o3rORzoNtf0jcvOWrigOwOa7TT
Jkh7D/EhQ9nIba683REoepvX1nfwHWQEInBpY0+Kusdk6V7T0Dmfgshywbc6IM2eNOLVXvLYo0lr
h26z6rgTGKK39tzPVX/16RdEpQCCpoalyvZ0OrXkAlT6LscUA4BC4SnGBf2GEJEtmOR3xQkLEHvK
J/6jUtpbB686/cFfKCYfVLeaRRahCy9TnwPv+nSIjoANEaCWwN4txQ8Nt9jPXOZAIjsRV7YTZ8is
hsSKy2mLMRVfH6Y/dfTCXDJwqLFKtcCqzJnMvIu/u2sRsj75hfpQ+5vfuMTGxr7fvj/9G2fma687
Lo6EoSKhuqWbZiSM0KNXSr74Q/wW0EIMpIUCNgDFrZeiJfKYHZjSP9TaVWxg/RKLA63IfnifFPIX
2cWfpbHTNLi55OpcPAfMaqMOCzmOfBw/LnjwFGtqu3YKaUHrVGXDzzhgVYQ0OQ9ffzH1SN9aVqJK
xPjEEfn8svlXDNMthweNU5/etViuFz3Un8cqaIgIgmTwN0mwfdb7eVOd4OFnPkOE2SYoyHatHGOV
EJlqVRapsVI54QY2HJgrhX6f25Auw8FRFR+oGc7g858pLvtgMfHCLEMDxqGyZlKS53sopElkhY44
uHxfaRix1vlMMWHsjgL9IkGL+3dMHi1OSlJv5PD29Y27H8erNVDLRrXwq7PQYt5TR3pfq/nH+8i/
exqiW24OE7r4WA8sV4mveCTTq2jNqN/9JHWq393No8kX/tPVlJn2f9J7n28GO1N1Xlkdb4MtYaX1
Cm6sn2owaA00WskESYIUkxaPIhsNv34YWJcsOwcREyVYfdCvshhHpMya2qPfbE1k3RXHQZgpOZWh
kZcZraG/VRcmucOYZtg6oaGAvKScRzu4W9xUEYzhP4OGJLYvBl9RAKor+C7fxVn3hhkhRlSjGtMK
bleNrlz0iT3P/lAVmf6/6+WmWfLt5lH0JGWzR+F9o6qsNx1CNjjRI9ETnoAL5UXJMPvxSvx5YNC5
bAUhN5JUsHAZMndW7se/XpNuZAaGEyRPVp6ybcfvA5ZR58Rqwc+XTC/uDxaYDYqCgsmzKRaaoZ+8
6wa7B7mZhxn1TaZTwZwkXeaGedG7Y6eraJVFfYchFiKTpd0m/Heokujj4IDPePMADvOE+3VendrG
3Px9cLLD8wwqV8BzUguPNYtshF7xDtd9xTqb4NxZK6ZkBSrpQ7Wet2z6nsuxW168ygb/YQAwVVeD
JR+qCraTxLxkti4WL7Eju6fh23toO9ks414OOrmYNSpfjkXTNJXmPw5/ON7wUQKVLnswjqhtop8m
f6CCPIqgXGEvzgNL750XCZPxPcxnjvQiIfC457CcfJkcVip40R/niT+JXJ5PoB6JrAZRFKJ5mby+
Sv00QJUO/McWKQF+58s6hws7XZZtQhfpIW/MFf7sVKuDEnCtwG9MN5M1pShQzkt/HZR9XaDCEntc
CMrsPywH88SiOeE4wIobSSDkWT6+rE8Vz7F7Z6Gv9ZW6zYPQryzJetoUPcnKjB0Vsuta7Kyzpk7z
vFmpGlqv5cEab1cCUxorE0FLcZZSA6NFEWuSQpzoV4eRdz7dEvWazLcZx8HjEOV7Rvv4KlExUd3o
Xa2tu7oD18Qu2b/MMsX8pxNeMpqL9T6kveCVd7B6kd/50RD3hy7vr52ErZatkAnGUR3iT2JKGfuc
x/IG+j9KmpADRExdkLw/IWqOnOchK7X0abvxWO/z+8RmBeTzJYMc/8nQiavRwvS/bVl+hAsFtIX2
sXENZjHQqTGnGGksbB4gzS7JccPTdOPLfjRfMYUQBh8YoSRDcFOFaJzxdrucYZ2cqnfhKolzjPc+
DfSv7RMsAYsiq4t1ShG/cXoCVf1aUwoMILUy+jVVg0wqKaDSqi7ug8SvasxNA8TFS8WslpklNYZU
36HCsqSSUbXjyfPAxP2ER7aB+sO5yE5cAqrEImjtlsD1eqoeIUpsWofN9JC90Rs/bFLyEGzdO58t
Y8IwVGYTpBFW/L4PMBaoon+5RbDHWkA94FAuoRPKIv7fLnV9APZZePIWXaBTUknQSuSSCunz/3AG
yQWnRSBRtdowkz/BJ0kRyFRqp50QvfhsSmiG9YsRnZhkPADZeGLOrPPM+IO0qxAcqC3fFKdB8pXa
aDInlfbyDcPRKkGrPZuNgwNJ25hKVYqnCPSXYytTBo/Y/YONtOsySAznMaana2n3tpj4/TCo59XQ
aWqXNXXq77GrpxSoOS/lnG+8GqAucfbo5t5cH9N0CkPXI5J0ReotNv2CCCjXEUcgHEyD2Tlkdiv2
+uDKbS2p7HPklecQpIGdX1SvI0+vHvWf217RdMTjto5wSAwGrW7qVJENNDygMELs8mz+KfOU9mGw
Bo0HaL5CnCP5+q510WwrGE49MAbkSUBJCdTTeve67/FVmgl3s7eMKnxoR5x09n6FJ2BzAvt/Z4Mq
Oau7bffpZPOR6KTO2qxKAlVxl6zKzoio7NTG5X3VUIOK+kQhO+PvTGFGhThNhq/FmylM27oTCn03
pka7R6FFQIcxZjN90WSiFBJ3srOHzH4K02Hlbb55u2WAVd8C/4m8kHKVkkzJ0jm7hMPkQKxhb+AX
fe9F6l0r56z0JT81jfKVy7BNHI35Rmlmn8xHCSb45brMO7uUvXKDCTF8EkOfY61k5gKxCnOePM4Z
YiaTWztrSJ5SXB1D6nNhq+DhMz0GpPEsK1OcHdTHGagcKYUI+Nq0enaCtE6N4wkE4/S6GaRb3PnW
jnVrROsbCXeQIOaI2oKG4QYxzR5Rq/cWSULkln0faOyGkb6yGLzF/wpzvYgDL0wp66hOy28mOyJh
OZdc7IV2FkCzA+awsGhqEgyKUc4imDe1Rg0iW//9LEd07TyMidchaTAWfsE1avGK0cyNduUZrqP5
u3gU3fldtwCvuhUYzipnpnIO37pMWYyrjVNZxrBs12fx0rldURXgzAZI8b/VGPZGzoODR7Nl33MO
HL7ZwSua30qhWolWCG+4PAWwfAYTRyuFvC66sY2/O/BJ40FnYQLPjv11Rv6iMHTMg4FaVa4b5duC
rlReIKZ7Bf9jhjrwPTWlguymP7B2JYB0Znut2ytz3xKFbZW7jvsO4oW17AiVEzaX97U6UwyrbXdF
BWepxv/sjjJYuWPf63NjrqTNDZ2Wq6lFej2jfPS3g3mCfIcFqW4356AfT0naB2Wz2T3w8DRzxwXs
/yOgHaz680Swm9WQB+48MC/V2rnAlVq23StyD9ucGsn/mrr32tGlnhevLom3T2qEo8E4GE0hTl7y
gDH4myhCNhL3ewgHx2Mh9NyE7ANnY4qHxoyjpaPKdkYhf0IYtMHi+oraVoc1tEmWyzIhp3MLBJoD
8e+RfiWq8Z56Vianirih6qg5nmiR1olJ1CJbueGFnFozChsLMp9ZK9EGut9jEtLRdC+R2HZNEAfa
ZM9hcM2W01Hxzw5OPTQFt8kWZrQSe0TvdAjgxDrY1W4YLGmZac7P92XCDp6Y++TbIqIudBzgX1TP
2A60F8AX/55mT0oJtQGPZe0/guJf8NP6h7fdYx7Ke5VKW5WAGg1HlfgcrQAl2FsFqWBToYP0xGlQ
99ksgBFtO+OVwD7LTPEn/STolWKWkGqpdnNB8q8fOdS+usWvRdlMZdUfo9mVZPg2If/AnavlqfW5
PRRD7TweOLUb4AAkuHrGjuRCGBR4dXP0xMdw1pUq4RzT9MSndwaYfIj5xrB0lSSFWF99b43l4Xha
pr3wwF6oCEMeS4SOFX4WweAgxYs2E060swo74GcGgJ6Bdq/S2ud6zKzCqpyqiwr2H0V/Se17QCNo
6KEAS1B/b2DmbsACYR+0MS9Mr3SJTzC9PgZrd8/7p/VZA2c/JTcVzAkcUYd8zlVAp7hqphJdpwEC
6lI1a4ngy1cNQq70DBO/mapUOdLtDN/pQ2n0AfNBUKvjzvThnBfVJd7fk3q81hk5tnBn7YBeZ7KM
cgrGw3SXSt3eFpxe+6egIMTNOLGXMZJkF1NZ/yl/IMAvF9epcAe91wqohn9q4E1O7mauHCAZz1Nf
NpHrwo+zKEvth/rQH0kC0yzZYhoLMGkotmGGBTCjratvCYaGcU7F35Z2CEaOkSenbw/66PVfXb6c
ttxVj+Ahm7MuYBS4SSCCRDkXEFmq1jyoyFt2+fOf3uJ+BivM/80O5rji8P16imYm8zwIxBXgS57s
6/qLyKz6n789j2TQjc89sOw7WtWB21sL/JwVsabNeG6HKtukP+B3YvOmf0QsyOoj4OmLqZbuuGfc
lCpIt0OkXaa2IAYxG7Env3EGUtl6IvynmgLXKw28/Hn8HrtI6s8APq6q/rtUac8lk0oZ4oNmk3lw
hvlXtndnagZYPjpxRErJ7OTmZJEiP1nvJJUJiq4b0F+RHsHGIoJt37r/DA/XCrcxSrwP7Ckm3IKb
IexGESskc5HG7w8EXw8+HRQ1S4xG5NPjAg7EtgJyLuyfERYE79lNJRWxdUQVjOrLkHwJqtnWa6Yo
g8syGjUT8j/kF//diCRt0enI2QOCB7HpOs3hd8htD2IJ+GdvwyEwjFsl0tkOE/ndvXqWY7DlYEwY
n77Ue/i8N5f72eI9eVZfp7+u1F5olMkrDGSec3NEW4z47zuaRZvNhxfP6lIpTNLskoXYHWKFCewp
O1fEbRuO4wHuXYFENIMr93G6teH22NlFjVTU/tAqhD4UBAgKS0MpvIi7acHKr9YU+ImrdoaxN2G/
/Wbq4at8jVe5MWCiXc/tmGsgatpig0eBL2I8e+QMb483YlcpsdFaufg6ML4EvkVyVo7wehsKFpFI
/eES7Mh0frzHWx42nz8nJLLvP1j6LWbSYjB/GqEB7J6oVDVkBaA8rn5VFNxYH/qHxpFlruUFAbcv
QtT8+NTomcZUzGCAvEwhfwccz0Lko/CTwPBuSnsYoieFiPrhUSANedmmod/wVFzuYsoteD/WRhzY
IKB3QskGjE7y3Ty/V6a4d542s+FczaKvDn7FQdZFn3XiqjgZPCXRwJ7FGhFuE2m6+fms8wMQCYY9
DiKkWA9FEHjnrXff2HzjfkTaxe5OldTJoOwEE1Tz7MgSD8lGrqRN42BLLN8yhG8W6KiNXcHyXpEu
jaJz5slhGbhBX1zeKSFav9SOwuVRbXJ5d/9vKutTGd0rciJYH6sHbFk7ZRcj71gFFqSlZtK3YmA6
mms/vGMf/INANuvuoHM6gK7GRF3gBZBjotK7kNZ4YyyS0gL+VVJRcP3MQoTlxaxCmyGNr2wDO2zE
eDPUfQ7PS0igP3Vsn3o0CV8DgxabFtCINmqFrDacySmIp2wwe68NDqcMIQpoMkmUd1VF4zGhM+uV
qeoR9IjcRXT5/xQwmPNNpfF/Wj1/9EbBP9N9ukwbPxswrv22C0rnIJXXZyLjaz0JXMQPcRIPxC9V
/db2RORHAMBjoayjP2KJQ7cBxdCgrDOeNzdEMFw9ROVcnED/6ifjlMI7/LQIqT3prUmvE6VdyB0m
p/WSealWcJMA9rLqofoadQAH90CzHB/oY2NxW29vL3wTltMHl4FH2NH4W7+C1jklBYhVisMbqI6K
jMm6DQtUN8aE9wEIzKYh0PKSJREcMK3sf6FshuiIpH/qAJi9hJlQhAbWBAXcqplBYrQSS7HFvI3l
iS9hxPOalTXreR8K4UrtliX6VteAnWpuP3OUKxCPc9y3cbDeN8MyGJdE4u95gf6mOLU68e2zbp7a
Dlt/7XA89nySOG+Arr9EWFvbcaLaslNwv0sWTXYidvVtZHMMPe3vmpG2J9J+wEYU6Cys4MakJZnV
DOKv/4+99Vy9d/gr7XL8UJoppPwF8R7lI6G+FuYgjzP3FxgPh17dP1JXfY9lcW0KHnNV3zjp4Lui
iRxkHMHxS3Q88bbMe78y+oZ22AN6LSSKOQeleqSJJuzhbnEE98CFtUOjO4r7Za8tnxy8zwvpS8PG
fEk1KR8Zs5EU3EfWQuT68oEmbH2+YNU1Y+6fHHL8X27N90MUZz41bRtSRRiAaljgmyzv7ZTo01u8
2wyOAohvzLWdcSj24IZWOYxVKc5jB9vRJKGrulHwf0WXf0foV3vCq51Z/v54U/HlP3oaQJUzKLnQ
/69/gGCEh1bMAf07hzbtuRt8Oswgsp6LJhfuX44QXHFB1H/f9xJ2bbcy17FukUUWpcFB69mWxoe7
1asy7nC+7I76dMyxfDO7RbR9p2d+zCSWgBUL5Ay/8Bm1Y1Lo6KFi9iRzKGzi6lNtYNmLNsB76g0m
SAwh7Y3/84HHtMiB6oc1RtPMQ25h6gcJJHn5GaHLh+9RRdM8kjja0nDGONZEFlIUBuf0+Op+DG3C
Yh6WLWleOjvJZizN1MFUNHhC5vd9TYUN86HUVr+209pIxIrKoBCfFbN75waQIJ8NR5O6Y7BWT4mq
b7lPKvQy7M6kkzzW+UW5hmHOFHZbe3wGFc79Mu6LVAWYsnScvXDu1w0dIuXEL9NyIAN3astsGOUg
LGi120IaSUugodicXqkEFiya2kwfxuGYwy8i0Uw8u5/Ow0HJf0GKPHuL4fp7oks/unKxpXFU1ghJ
YYW3D6lhHrCJEC3rz578QkP6/62m/8kKr9v/h0kqEvSzi30uNAf01HNzuflIwBSwy3qLrlOLIejb
rFGxF4DIuWP9Yu4rrgTi2yjzUEYQnqDNCfImYUA7M0/0wdxrCLdNbKly4URgDKxbmycev1otEVRh
h75TZGVAj2kDAQOB4Ia40LwMwK9H/euNn00T0+UP7qAe59tJlUPMEEDzFgma4K9cHWmmhmL/vy14
JY0X8YC7QAEMqsCJQx69064nTM7euUI4nRGjbeibpw1pedL3u34Hnx9KCjy/1zhd7Tz1dd9Hw5dN
WhTFSsNPJwr22ZEcrvazqplDz579B+Bc9lTG0+D/xAq68CuwsfzU7rlDHfEwAKCib2YDHBk+Imex
C9+zu7jJFKBDqodl07BwnsdG2DbGWkxFKnKTkE/KEgmbhqgoN8FhmXFNmW5BR6NPErZ1TsrXIZ3S
r7e4RJgTzrxaQtuEVaMkdJDBq3w0XXhLKrsyz2lxXq2lql7xZQqBkNyzGWiy/D2/P/QkZU/DResK
x8ifyFj3UfYOeoxQXBJ5RlrMoqAKFq2plOFbTLok3dmDFT/Z2ubYQqLDrH3pm9/usr9gvuSumRBz
cbtRz339zBwCBnNN7UAW466xrX3inlNcyDm1ZsgpBcLf2qj4uPXcst3NdZPEB6T6Pnps6uC1MiM3
b4IW4r15eG1NdTWiCPrspLbNCvWUaUgaqUS8/VxhQSKuX4Ue045QSG7+OaadVclWpzCZWMMgnavx
kS9X4QwStEP9Mor2nBbSi5pcpEXRbxeJC+ZkPl+YxMQArRSWRO+18xn6W/CwVTA1immi+bgn8NBj
5fAFukn6Mtu+Rkiqn9YdyozFx1RF+lBTYFaTZYwiXo9ymeQpAKD5zKMhwH0xXrukaxQB13WDCeAG
6PIaqDkbZZGAsjaonsUn3iPQdO1qrJBcfFjR6RdNj6y/rmsWV5Ds/ORuAGCMAYIO59lf8zcTuUci
30ByB1VY0xTNWdQZKMLQoLZGrj/yzKE19d824xg4cmKz1NWV0NLk2TFF2rI5aWjdGctR2VCyLmOM
ojwk0yoTlEz8fIyrkTUww5lDjn5F2gWSBUjxz4N9DFPr7vG9+jQhlq79ZT0OkSvI8mTbIO9akRe/
X07QxQA1YiWD2hzGBwtfYGaM07bAx6XVbGPU7QFOjiWywMEy2QunaWzIhbMDkxVOTP5+sWTbwKvj
AkbaXmtRoTQRVUJo8MjVH7AMPf+EWvpx1agyW7sb8bsNVAb0Mw363oPO5KMOk3BJ8v82dMWLx6Fd
wKD4oHoodPuTcwG2I6iRJSjInY6JJiGF6Anhf2nmEARft7u2IVtUgbPCv5M/7dPG5ZZe5kVOJxpD
Ih1DNdtb6xVLDMrQkzEP0ibph+Mm49kt2TnyE6PqYFvd2HcNOGjs6bhCs+KhHPevitOL71hTjjHT
DRAWKqK7Kyq/CM1Y6HPAOQZrFkCaM+VXy8qaPVH/2GnfnSnJM+aQjhRwUqAfM4p08YaDDqD8xCwY
a1vZm0FgeHxZsB6NKXLlX8zMbzKXuRruKUMwe9441i4PglGZAt+RM7CWBi09vPAGW+DSJ7h+3are
m85cQustpRJOC2Md7kRDSVsLPEYo4Ob7S/8MaLtwNf+8UStRkveUk9hzYBUXyEwqnmNqGlEAfa67
fs/4psaeBgHBwGuVo5qK2d0o1oR7QMUhk2t11adX3nGdkkLrmUBEs2++jg9t014I98haIQTGfXJX
kC0D+6yZ96JtfFC/A3iQicJxAtpWb7YfZOYhCLT1tLinvMxXq2Z4kBtFUtmXTakUmeY7Gv9QAeOj
lOKILq1dVFk6gBK+iELKywtgGH0PNxPzVSmhd0PMmCK5cM3lMwqP2na1jIhsc+PSRJu/tKnV8ryq
PqxrI46mlIG0nkZkoVTnk9Z5n1Mm31UcexM/ZziGpLvKrsiQ6xwSxRohPBOlSc26ToO6y80EZlv8
FbC2BIznykHi7QyEVSQqr3gMwHQmsoPF+NV2oGz14J+hvgmyVmW88d8VBJUGtQd98ziNWPsEYw1P
bQyNeBwJC4qSbZjU0HHpPnfVHmj5nNj3hdgYsq4PVaKustSCwXaerqrvQzkdDCIV5r4yuYEXX5KE
8pKUC2tA9StYNZnax0LexVwQuNnQvYT4QNPDlOPy8YdRJ0WfypielRGiWTo8UmJaxZaCeXSJWNPV
Tqf3zcq/2uW/cv2cJtBAkOA1pxWCge3KCA5HBGYb2fWXdp9/Hj1HYWcA7tRRIdZptf7NGhug9Ejg
FcB0mNdEOYSTi74FytsR/8UzWwxrjmSzesUEFeIS7pOJMFxLISbWAHHIfpF+dlVFPf2pGyTTy1wU
ney8Sf3lktriUIR3cwl1sgBypbAP6h1lZi79+uuI3EoWnDtZc4AOuQhelkYwt6BqL3c1pK++IQpP
OLY9IoNZwWt/ZILcoQlC65D3KKXR4T19Nm1H2Zkto9zhUbn2SxFtwvm13qq4mZjTFFDDJU+VB+Nk
w8BCTpnY50/kWhjrDcyV7j77reR02w0UA4PxmJ+fIOYPq/05oODSD4HVWhxyAG25goAPrLC/qirm
fLAZNOOL8DksPPZFe5dpQOSKF34TNjrIw6Nxa3xemTxvjWc4MEV6bT7EKl7usQ5DSGgVI2zZEf1n
zEJnDRI0AsmUC364GSw6aqX2AF1Icmp1bPL6Dn6hzrDQM+I2bWXWaiGLJHcxWTkr8EJV1uI3qoFH
qS/V0y+l1yZa1DWrX3n+NQt1uviv3sV6MMBRRFZnorMzFSFDcQOmdH44HH/M2HwyReBTQUT1jhef
u1c8jqSu89gIn5WkgEv7DMxTT6gOlSFFDe5zRqCPn5g6nA70QlY4Xw4M5NFPX1TQGmxzlJuYhTcs
6vRijqfCsw284bjhMtUzTFVHXs/FgHqFEIX50e4nL8EDBs91jiHPGNYCzyY5XN/xX6pCmyLTaU+g
Y+d4RSR0k6skpQocaCI8Ora2D0ySTfihGXd82AwEcFcRmB0J/d7v8ckheFgqf+6Caat/MzcfIFXX
CgUs7Rxx5ihF2jns+XALSpYrIvBlULyMJW2X9zMnVJFH8cE+U1w02iHwUMYdj4AJHAvPOcTM+rqW
89nY8YvJDbEKSnc8vXb//egTzUgtcIn/IIZH6D6I0013xG2lioryZxLi6nd+33NbZ+rPePuj67tc
A4h8a62wgrKzb1Hraz2jW2kB3m2abPgbvLgJMLh3suoJbOhwFnphWAgn5irRVeabYHHOiWKpGTiH
Pllt+n9E4nxO/Vo5z/KVcK/xuBkl4OmVDhPkDSuduhAB0qHFbLeHEgQ8Ivn4dM9H7OwHspqDtmHj
waK/gkPGPj8vqcaOo+WT/1ck30iLjVteGwvykJi4TuC8PUrq8x295kPAir4uhoxJ8/fus+cdHu/t
ujktz2garSyP1OFViTRx9k/WSIK9ZlOGbp6GV31hBu6JJYYaiMK3iczMIpAgdht2AdgW5ET2Paj5
lLYEhK7/AuQtZbIPvqzn3JKt4fbjZ4a3THssKIQ8S8SjP7VUhA3XaH/GePRzdA3WDMXz7SGte6Zi
vLLVq0RsFB1YlqTTS66gXbyDHfD/IyTmC/dgXiqnBzqriBhCCWZzoPOODMpQPr1Z/585Kef7qnp+
RVr2qwdp2YFqa585pVmpSVKsx6crl40QVU8wK3iUTJO7sg7ZqUynR/oaRhAW+sLUNkDLV5VHdVlU
1eg8XsGgmFhA0sYiFS0TBtV64CGDaS8QFXrFbw8pi8FlFEvrqYlDZYdD4SWantOAEuFejjn5l5b/
HUzDoWhq0z2eXNyetF8Yyx8/2tJ/e2twYN7kW/QH6lIpwt7YPTYzRMumlLdPFg398NEj9hjJC57N
ePHqHIB1IeHL7BDScEKefxTHLHK1yGZtghHqoRNikKDivIJeIhJGfLmueseV4QHTZ4svcfWu21dN
FBiHTsLDJZumej0kfzz7LnPYSQyY+g/h6SAZxlWDXKDEywPgiur+h2D6J5GzquJBGxPO/9wOc3Ke
+Ezu7r/x0wSVT6zAxXzPZGAgzC8NCkA24GeuRfmsR2QeuAmOK4zGqhTXnp+n4xPbYtcyOlWhODIa
QCX4kHp6Zfl9ShXLZDTMdo3mxY78u5uf9f0fn0YwZF99bPmIkhTW6zD+4c5CNBsQN18yFg/SwVXP
eH4V8pFL3NtgS3i4SiykrQeNOts7AJYZxJcYIC5sr9a3KDidK7uvOw5xcbpVw2AuK5qS/xQCeWVV
eDoasjtgCphlW3tgZj4J+Xp2dvU/aQC7sgSsl8jEY6GuMkua3bS7gqBeqpvVcCg0rnOsMyF2arsa
qxayQXTOn6Gf3JKeuAR3ZrncR7zmQxMFE1LhrwlaKLL1o/6zf+QHesxEptwQv7pGpoAmFEgTv8kD
m0iv+TtlVXyJ53DobHSt4APETr961neY/+XTdTQPw64uRR4PDedGgm5kgMtGNyudaCEmgoW74p05
+tx3/jZbM95+puP1/SvMN2EY9DoQHRfm6oFjligFAkt4EOFm279Xqc53bF6VlLnQ8aelNLasW/iP
zn9+PaL8yJf4jnTi0Rl3CGf/+LGcyMb8rchK9rW/nsgeZgOFNiGG55vu222rxCKRmkAs0FqNAaxM
TyvfzuqwkyNHMj0l8D5pM1kzhYHBsjwaF0bLzb+fGfu1qb8Hs1shhT/XGmWWFL8TVcCSsiHqkU6k
KxL7rZJb9wmEX9Hma0itM0ooLM8BG6pHbpiHGBVKk8mUhZKG+EIm/swpLIj8K5uOL6LqOUSBdVNV
T+BpBvhGFVoTOC+hY9XmiOH9i5jifN83scBmNd6tP284ZD0Rv+ujciCuDmtyzZR5vaTajAhxgXsW
jgQ0fg83CsEBsnCJJNBQGh5FxYlE0tTKTihcaUX/SvpDzGNdz85vKK/mvhgnSnKeyiu9lTUiokVl
gLobtC5pZIQsuonSGt9hgbXdxEdweFE/uPua5wgzJLEE3DN7H9EIxhzWAX/TH0tmyqXkMK4AjFL0
RUgD8MRutaeHRhnr7oQ/lfwBVylKiGBdFuCSYlE2BrDIvenhgVyiW+JjajbpvlAa9u4NLOCjToJr
qIKTUNfz818Q1/juixGl4sXe/5m4m3hIlN2dwvqwmxDFOCT6j0UFMxLrOzeyMfJt/pVYKYWdKzc9
8NrvoGGTI53vXNc3A8PvNx1EW46LBEiBlu3AvCvVz4ChX23x+sWFUXcVTEwE4gsj2n5/iE8FNZ8q
dFwCqXSETXmkP/M00Qs77a8xIrkLDnIrJvA8ToHlUbMsuhuWkMxNZvSSYCiu1NiKqnYCSwLpHtsh
BUWK4jO7b1Fhg+yjm5nE7PKmwZI1Im7kHJH4GI2xJAIQ8lR5aA9M0MTKiqgK0biQGB9x9aOf+4vK
KeNyeHVmultAtiDlzHHLW0n6o2ukoeZwOGr5jnFTucAbyg/yyAL4jpFJ6TlvT/5GYDD5hFn/E3gl
zmEGiDSQK3c+BKGTSLmYEnHri1CjlYFJ8GdxpQ91L6vJ1fFKC7ns9lzw0JMQOAehkAu1hs3qGNax
lFFd3/saLQNbJ0aKoRgF/6AMdj3/07jzcvHFzwS8raCpcVwuStH+RYrmGsGnLDBjm353NFJkiHND
G27T11ZG6JDpUOIhPnwgqCg2kpofimGVp1XPeM+bZucuE+4FwTr3coP4SG/U/CieEqRXoJl4bz6R
5nYdrL5Wou5gwUAIm6bb3Qu7vGDNOAyL2GNWThNvwy4W4Sqo/rEdBf9iSJLbe1HSgQhJ9i6BURk5
mJ4ypeDYkQJB+pSU3UHazmUNE6wDP4/2Gr3ked359qPaBAywEA5JxvqK8jYRZzHYEtuJQkTvZF5a
rmThEn4GQ5qZavOYBsSQsLpFkT33J2PWempXM3D9JCDX4FPaKOpPiMrqTBCpabZSkPjU2kQrrXXm
1ySgqj3zKX7bC5jOcrkAKUbYR1yPAe+j4fQMjfzF9aKNJWIRAt3Ujso4htpLdIY2QjwP50RyHoHL
GlgIor0ZcPuF2r18URVDNISyIvkWMVEtLsenp4ZKMkzDFGBIfkypiZNQ7o7UrBxJ7Ps53XAU5qD4
nRNBvYv86JP+xf/r6YwKxu/zKA7AQHQlax1pzqL1pbB6uTnElvwqicWcA0pAI2sZcjaFObK8Zya6
VFPlWsOYy7V6X9ZimnsP1O//8Pj6x3PguUg0hCaGcJFmO417bXcIeiLSEBJqwVsAJdmWxwKgkmDC
mkZeV+HDU3QEvQ5s/HgUA3pBq8Xe9Be3FGTyWRhZvY4a3a5VyRq69+1HYbVHgAoRawq5ERKNgjXp
PCpQsORKDgSrPNcuPu+v/5RHpPa2ka8r0/8aRdxDqoNf5eiugJ0VOW9ibfScD95f4Ql+DolOIVDg
9yMLE0lXgPkqwlDPCAzX7modQtAcQgQfsbkCmAAWwut2qGecLdxJ1akhVXWtgozfqKM+dxTMCwS8
TDKxFqUx8Z16gdp8YmaZrS9Ii8DgRfVTHBgpteQM1dkko8S7Doc6lNSRlZohhBSVUiStbNL3KLXl
fIbmk/ftY+VQKQo0cTRcPWsWpLsN0jkt6j3LDzd9XhpUQhMX8RXoIqcpoAyRv4398ieFg5kjHixw
wi/15uKDzKI6Iu2Pccvnv1JIRtCKgZ51R/UcXI9IZJgNiWiFc2s7AVXarePSO+aQa1tQvXNA+gdn
k9K6D4DmDdRlrg/mP9sJhr7cus1gLQG7esCkmr5G9oVX0y7ryeQxpPpX1kDZsLg+A5yI/u5Mft81
D+7Me3pfU391VDy5AibKNQEKUnRVnOE/xBdamxIB1ozli94GDKxvVYvSzffa7ncnB0h82JmWnXkX
qRXL3fUzqLB8gLrLu7ZeQ/h2XGj9KOgEd0FgCboNJP97fKQNBVDyzxKcoQEMzLSCoiHKyXirawF7
4CHquYKp2WxghaBaeVWHUsAgpHOQdaI911UqaopL6jwY+ThovO6mbOaS5yMOeJq9JB+17pUk+kB5
pxPqjrVEIJXmXc3aWsCbrIA0XkrfFfhg33MyngeCR57HxaWMVILkTU3fg1i89PwdsZBYQct17hAg
n87G+Rk42Bd35I4w92MyYlkNd+jpObldFyKObcGnXAKkpRddaHtNvc1wq4mndAzBFJvVzVIu5klk
ju03CUcDO1fcJ6Ay3Pw+aC62s/fnAaoEXbx6aKTCT2QP9p0remkKocCCyZRMNDKEfy7lFZqslQwE
8GUjPjiqLTq9nf3PGA0je5q4O+97IyjDs9dDV0cLIlh2uYnWsEqUBPVhlagO6ZNouNr380lA/zC3
ekQke+AEjYVMMw5QCd21sQkZyMpqLQXs9R8skRnUna93zf9e/dt803XbHGKjcVQA468plfi2QpdF
FsHCNgJEjdvZzu+LjY0T/DrHoHI58qelw6CU0kpVN9oNz1rHAQLiXoTbDASGX0Xt/57/nrPjiwHe
+ZOks4RfmLyCQg9+WvN9f9btXcDl5AuZlMsLFqkUZv9WnqDP7C2ptQunZQp+YGxPD9CPeil/OibV
m+qCp0KUo+sjbm9A/NU1lOg6FqD6M9UoTr6f/TOXXB/ccUOHMjM/wFAdiAM5JCcpJq6TbGjtTsaY
1jOdYHbbXx2kF/zXiBctrlSmW8WqwN/yVGS+9NT6ei90ERTeq6tt+g2zL59MOfDrCD7tw0HnJ+1M
ZirFTVof2ZVgRj43ASs9QgIYkwrK2Z3CSqmgY6kIFpek8d1fEDY4xxub9b4diVkw399UaLD635T7
n7HvRUB87crm9Pe0YX6UgY9SbBCWmPBtCcT+cc1yoY3zc8fFMP6cEaqdm9qgnXf/8ApI7pFDo162
dV+xjgKCgMCUx/eliWpg9UplNwYkiv8uvmpwVRjQdpBLASFHVeQc9hd3/pcMWKs+BVd5kxTYWJ6q
NhCum3Icg1oN6AdgJ56B2mKYBP53xMcNdnZtOoZoBJZdx/k0OMqyaqHM+ZA64YkO1+1x5h/pcYDT
ZSH9++2RRsNQaUPuWZeT+NCHH4wtCzRGCfNmkDNkX2NUeuBR7kENixB+6UVeyv/X3ROX5sB5lnnY
ujEy86B8XqGuX+hFmWVkY1Px6iloZDCKI5JxFbR8RaDcnCQpIKnNtUMxpRSOo8+X26ezFELrelbR
/gsub7F5jSdrjsFHIiB+a21u03+s6jVJVtkncD3PEbITIx232OWqLoMGBDLuy1iuX2lKJ35YOAD6
ReIS9kmooiexH+6w64jxpceoVQ+WjYNXjt5UUXCRaXPtnUpVo0BvuL648uGZGU6wu5TSjpltlzzf
R6eb4jz3xR6XoucdhfwAWVeT3bi+K0mUTUZtPJo42PuBop2cqHBrfWvBdxVdGh6FmTRjNZrx+sG/
y0P2r+gAygmstnNCiQH0XHln8Bv/jyBqKENyg0BjuWiuUJG+avfT9hNJec7VDCturretGM4vfD5U
wsiqgtBBfSpKHLTa5XtK+07CY0BMXvZulEOk0DSx0kKT9SWfWvoVlSrDudEmbnzTvHR3f+vWm2zf
vfpU8EnkqWgEoxjL/uoFCXcOaa2aY0Qxo8xY0T1OLaRk4rACRuMtkk0WV3brUwPjsHjIze6hB2gN
waC4qiRvH8RFTtuAbqFl1Ay2bV2AWhsKIFxNckDn5o/TU73+ExWr9bMbL390Pkj04otGQPkbg/d+
CKGzLVavYTxXy581kPy6mnYmbdIzg2og8Ax1mPGYNqscUiHd8k1VU35LMzzOJwZIXjy1MzosnGDU
z6vzH3eSpmnkX6kJksRvrtQkwhgZwx5KMgOlw4UBxGRO6WWM/iwQM6SHtShP1i2TGElyEhANs6RQ
LQi0c7k9Bzvwq43HHnWeWEgCfmrKM5EfGJF4j2syB3PEDCUAn6XDfgUaLC4nVkOjLt4u23EuMvFZ
AtXeaSinLjUziMPtNfNZ2+s3l2p5DwfL1Yy1Axoj0tmceMaSrRVwqPsccG4hPX+U9WfxN/IhmGn2
9l0J4EKEWxHyW68RiTdSNulPMp6tfIVmqnP1mVee0uJ/WjqMthg6610AGm/Rb148yLVOgs1Yklbt
RpqtJl2CcA7gFEBlOQCMQ2Z6z4aIpj1qO7y4jjauvQ2gjOfUCE1QVnhV5TXVkOpM3QyiZ0p3ZBcs
rH2mkPA+/Yy7KuYMw0m5bXUyamtnfiA0g1tR1QDsozUxN/rFXssDLNIA9E2eBDSlclCnXGU5CVk4
bN3TaLDhDy+lwxCkBf4NYDbi1uW0tdQSNE9UkZqmK9bba2B+8J3NTuVJUgIPpPaZ4vSKbhh07nIH
gfqsfdtg/3IkA/2NiHTTOoH3r9YLt2ImihE9UtVYtOqBh2CDKwtYWTgxeSfPVavtOy33z7k4ZN1M
FgXfisQLZliWHumTh47wZC3dPKg2Dxt24zb2bRxKfdPxos9ypX6KOiFI2dFLowumFi7pP7b0H+Op
yuS/REodSQKkMNM5l1NL+QQkcsEX3RmW+fugcyVBuDrjrjWWE8Nje1iXe9ozcVC5ghTQlHqX+Awe
/aNYylXwLodu/nAMeLdZtLl6qDKrVTurxYxCvEL5dRslGxdf0X8UN2xqvs6kiLrT+MAUCep7mjXO
0UTh4S8WYJ12+rOMGV+1mL9KnP7AEctG7VcP+tfqucwOPSjWE2BTQsi+By1LAxI1iMiCCJ0SOdxX
T2Psb7FPbBarPXvwmSTV+h08T33BUfD3umKOM32XjbmIo7U4iciwSRU9Zk3Bk7U3TS7QwjJshvUW
i0MnxOlTV1iohFFyUCb6qsbNS0JShLHw3pAOEqxH0KaG75zokwpNkCLv6b5O9K4+MKEGJEVd8LxV
WLLi2eQwB7WhdfuNH1atE/G2shU4cAKZYv/e9mCFa+h65nHnDjY4ZWenk/GmIeQaJRObXTSZaSLw
ITHMXQ8nKwHP8dJI3EinayhX7tiyZWUZM5EBIOItRDa08WfQbynlJCziJL2ZxTci3S/XuDYwafQw
uCGPHHfcx1omO5jLVE/Pu6DuedPctTwRSldJrZu1JneOrk+5f6bCMm4IHRcIcY/B18gGQyq5Dykz
7q7A+oQMAJkq39KzYC1AfXGTj0XBKvW273sSZy5CNjNBsJLCEawfUJtfM9mDGpsMcaPpKD5sI5CU
S0Pm9MuQQHftJnsCENBZJcJGbC1PqC+rWthWDmxDwAp3efntMmV58KxE4Yqs7yhhWp5xdIR0yddl
R1LufHAtNM1hflE3RQz+UH+UA2GfqCp4vAdRLS2KkSStX2xihBEGtlqYt+ewN5SsP0VsAZ122/Xz
Sqhghq1G3UWVFqG4IkcwvVK9GayqCH8bD3Qhh2AppiBD4CHzpAppFmi60QztUpLb5+6w9gDg8mfT
daQKJnqoyNuCKfRc2JAcSXuU+sLtANt+KWnuaeoTszYFqZnVbtwUPp7jhLjkLYrpJGwBwmaf7gEx
7baUBC/JjpvYeDEfcqekQOUdisGKsvvsn5tyeha8cKT6TV26Ym8EVWUSD1l8qAPTiNAf8dAEXT/6
SteaBdE9lJ0onRcwIpcqSmSuQUHV83FDKODGdknKLInHb2NaQnjePQ2fka8qL+P5loQIXhoa5FJI
eTJ6B5J/9gnn0VFLQFxVLvJWC0PozZ2LeOy9CmHWWyCLS3yhBEVcL8B1CtKWtFTBhQ2l1A1le/oW
Z9ecZ0VXP0EDbC5XSJmr+1RAwA/mrC0d3GLyl3XtZX7BnhsZx3MfPJREnlHmImsiaHs/V0yEYry3
jCKEqhP7XvljGwr8vozwDmL9a9hdbRGNlEoEzo7YKixk9jAzRFOOMTuR3UORAoXeL+3vl76bUgV8
7fR33UeYyR/1Yg0tXpE+eWxLRfWY1BZn7a7C6LCPSCKrluVzzCDcq+KwJKCshn2Ugq6ugUvwihGa
WUryVGOVNLJgxx1z9GrlUsvPGfxjE91TOxSPCkeIEl4A6YVQj68OfceFeoFlBVzOX0+lBN9KI0v4
esburgYd5wtxUbAwloCXsg9rDy/I3V2emtekfCixy5yvSa+rxDqWxcloxk5WSd6n7SqH9dpCxW70
ZJmXUwS7mfA9s2t/L5Hf8xkzb7T8UVTjC/WvWOGzADoDBD/4I7RGVdkhcEv5ThDldX7jIvfunDDc
yvp6ySniGOQ23b9ZGcqIBNdAT8YDTafv8fcRXdHZvHFTS+u61WUcPIMD8bGhkaRMD0Zp8tO/iXFk
Tq1cl4TnTAzlgVQBRlmWsQ6eLTOQCw2FCY7rTn5DfajtpsFt04fzOwCCB4XcrYuz8TshcbOAmsGG
1YH3nWcdHa0eZPQCjIDCjV7FqKqRXBMUsp9Oo/Nc97WXvZQ6sUFN4ypYy29RmqEeIAIxgnfgo5I3
HEGu9hwMUxEgrlr3WwV+4ameyt58sm9XNOVN3OwjLgHY8Jj1/C/aO+8i0IFdzI0fcUNqZ/S/HPik
IYxsz6x5rEpvo7cvb8P+DK0rkagwJb5f1qF1lKQWUm/yzkJZo8aDPU6+s6kdpNFpAN5JkBy0Dcnr
bRKa7m8xP66M9JHdlORaP8xA0n5gpUnUZd/KFwqbeD3/hAnPknP+Qm40yHEZrimqqvdMN3zgmjBK
fK/o9PL4HpCKAIAGrxNu1j6LqyULUsAsSrWOF7rzPUIDxHWsncFWvmvQj8Zi0jJVlWEbrblF+9Nf
etVSfZ9orQeyoMUuMdtc4vY40f0dj/IxmoqujcfI5ogTEg1ziqDgyrQ1Dj+/4V9QxkjDDp7rUyEY
WSvCpNoXEwQT2URTRTlRLKsiYD6COv1eD6zgAdIJs2wT/ILYsb4uKB2sV91Sf+TbrDV96vI/S/mX
aU647d0rZRbLqR9oXcw4ZVahUaq7TMkdbReo7EkwnVxGq9By9i1twnVCcGtBSbZU1EH5m5shHPMW
Fu65QSUH4PUf5rVHRlprUQ8GDHrIbI/WdQdaIih6BTXUDgiqPuy820D2gCc4XO1nb4LrdpFjUrvp
+w6U65ubu6m4yAxYEP9+f6QWT+qLZ9ZsGAO3HITjq5Pxl0r///3eGwQo3C/QcDfCoL+UemfLZPGo
6JOBcPWYhIen/74vr8XCyFuApYJBgNSbtMka2UOEqlICFKqlNFKWuTi/KZOrREcyGOwRxkmKZuco
0Ui1rkkDVYvt+FxDllua3TaHFbZWW/usk3tUy7PsP2pdFAtQnE1HrRPDZLOs4h4OYkmAqtw50Lep
0iIcNK5hjY5FNVnEAAzfSA1OBMO3RPipLoM+z1+Ci/xNOe4ePR4fxkZcJ+pdSh4B6D5GADS5JanZ
N/uNc1Wbj5cevWse1AlV3tKzn5EYJfnU6meqbHnoFK1jWSHBZYgDEnV1k0vuXFiwfPvXn7IoecJa
vKozQAEcFd2oIvnMEgD/OhV357rB7BUTXImmYqrEQPnGJ94bEbRDpKgNPQuLYUQUIWUIfoR+2ICE
mQqQ0V7lNx4CxvdR9MLW0nYpbO0j8t6cMIwIFWEYUkMzEeu7o1WNrtphU4Ye3bqq8KwzuE/aPdMa
9aBlEoUTuXp49Kq70e3v0ibONfF2e8vcDIO2Y3iu3SofPVKKWT8+y+xieAs9JpDyd6yzcv1kzMhW
8ihcOn8CC9tVBkJrDmhq2O9m9uZCafxMOXj5lUpp3wKCOyfoX06f5sAeqO3ArMHBzShSoJhKhogT
8YputSJELCQBNm49JQG6ltqgSxjXEeXZ3Yux7AHqnAIb1lXu6FH1nE4/PmlnumibZxrA9+nJPcZx
YShd6qd94laOoI5pXCvPiYiHc/LDwQj9f02g2IKIP7/Youw8Cj40lDzb2HGKelPGv1YcjgRSatx6
6tzJn5KoiRrr8YPVP+zaReqdiXGD8HEytSJqASWhI2rlO4i+ABlT94bwFGFZHuAaz1yaarYtPfoa
vL6yA25r6q90B+KKXa8B1H/1FAyyx94IIi4Y+hv2cYpK9xVr+ECeeExM36+3WGhqVzBN9Ko0uZ9e
eg3kCgPCx/4qs8z2R0j7Kf+XalPAuO41F+t3o/4pW7adj4qW4juV77uFxnyYScbKau20euIN3y7d
IGURMJBmTaELsXr85ivUkmbFopy6tqYguJQNl4DYOyAmjyL9Uxye5KWYa8woQqnpxbA/MUOPQv7W
kEO/lnZ8fkc06i6N7BpjbcebDu+c4si06SzMBMq2nf3ldIhO8I39oRTCRPDbgfTHckm1uiPFOOvf
9EDCY8iLyzoR3OqzI470bGR8yv2NvSXNAk1CMAwJwJdBgj2/JCaAp4bKYUOkyBMoRK5DT9PWWKm2
JqGf1yQq6U1jvdspd1Bncipz491Ik6uQQLTrfEqxQoe4brYug53EXOgra1cFVM2uR9lAEGykzS90
PxPd8vVVkNXcjmhIbKrm3kudREen32Tv/8xYpdu+b9ecL1aA0m9HM3YManj49A48+DhqMnvfsYG2
UzcH6kByRNhR+2f5TsJf8vOshVy/JcF9nrpySCZdMVZC2ZJVT7QFUmC6Q7ecXY41wmn8vB4Jn3se
bg9CM5dR4KIVXSCIW5IiZ7/dLm69QukgSYnz6lSO9yEqBeQUJBC+5U0V5/2za4V5FLu5SDZ5CNz6
pF5KKPmofAFz7iY/9m/PtIEgumYt58V48SM7JSaOvC2CAgItcnnl0+f4zqPkADvUWLwz/c65xgph
qfKWEkRb/EW9niYfMXn2+Lloz3Nozpnjxk9ZgLo70AU2AyZirsZFbiySjbKSe3iia9sMAp4WMkfD
yfvtKwU6Dwe3SEXfq/YQC3JryX/hs/K2dWjNtIHxzgV+1oHMpxw13jOFbmIJF7OqwDfCySnWn38a
Lu3R2ig8YdaKmpZSSG8Gezgt7zTEezofn+DTFGPcECBJBF5P4vT1lpFj7I8f/r3TpQJr31QUMcOw
TUSfgCJj7m58yBGa4RRVdNOybjWUoQcQJok0YMvVSZbLmfdwYjZU4P01U4biDZU37KTUJiSd8Opx
ligRz4R4rmBHqF0yRq8Qnfsx1oDccv6WnuQrgtYKP7A2tQsMXQN+dIuXnZs6tEK3B5cjmpqjY1LB
2lFfi8jUhsU6ScwLyqwdIrJJuMpwFRPmzD8MXGls/E8/rE5aqy3FoWNChvyrBCSxMZP0/U7cQM8L
0Ui4Y9JfZJOc3SE8OSmkywtF2Ho3DNxef8Jqx+ERrTGD30KVHKwdcsNgDWzA6OhbbNY5jLKAXhDA
iHx6gTBc2mMx3wlO7yfutllizH82G4W+5qMoJ++IcxWN7fhvyX6JEfhxE7aIDc63Pg0xltB47pMR
LsAnvc29IDvJ+58+QW3UhWecBww7F2wi4cI6FiGY3CjU/tZhr5ITUd+vsHxR9QSGfAJG+OV9wE3O
FfF2NwA0GDrd1h38NrrstR1KuCIymARkJic5IXNve9eEXZrUrhTo3/XQu8j6tFuDlbNTdCXoedp3
gPnTAy6mCxUcE8a1G7eqWItRCP7bnnR5JT+qnJDRvxMpD/huWmRNfnxhaWfzgQ+yJVvRDCfmP6Xo
Qb4trlkloBzbj5C8qIGZwHQNFLQs9CKCpiUFs7eb4sK/xIc6b3fTZFl4N7YL/s+rG4G0H4Kt18qa
3bFTnSsHeOnJ05VTNzj/FDV1d7fRXF2raWL7X6VSau6NId9gitahE0ZH+5DISm9lPAMEC696LnR+
Gz9ZdGQ/l1EXdsGOjxn8eoaTvIEZeyhPFz9I03X2fJ2qoThNchJuLvYyOC3R+3PNGMS2WLH+SNpB
JEY1ZRFXJuwMppoSOvZpymyREeBI84Vu3+x+9t4wYH03elCJwmBKDmKJpSLeBfTuPviGXyigpTti
ooKesPOMxEwpSy+I5l+v1d7gqsyDZKiG90C4PxcJIK1jscxX96TBQBPbXrLuWPlipLA+/ypCbei7
tI5qwhdL73efZ46cW4MfKmlTlYbgI5jBKiGjrDonZECLxVdMv06kbFfN/84FWW8UGn5ftXY2pqJT
woKxnnO3jstCjKgbi5QRXaVS575+ZtojFV2D5AHaJBd6K/aU5cni50zH/xfhj+w6Jp7DmDg9GvO+
a8X0rKtWX5vvauakEoJB92ety94KGRXKTk9sC/Ydivk0ut0BqNaMtOlArZYhhIeb0i2DX37zXHUF
om0UU65+2JXfiuSIW4g5YZpoEedofXRWGQz46/AeosOEIE3rMtP1+cs4Dnc8p+FRaPg24GmP5lDl
SPAHI/jVGdrozYh8wF32B+Jrc6q5aYgC3O9ROUdo9cV4URpWnIRisnehkG2TTzMVW1CoiOHVwq82
yH23i5C3+JgjrxG/rKSnlbRVgughPyi4Qxr4cNEG+EtZUB3OumEsjakwIPz6lQPVf/bkRXYtkwJE
ISukyyFnRecSzYOE70ilGvPmCiGU4SpRodO8LrSuZW6tjMQamv+dlrBEVQEWwoRQtOkEPiLpSgpf
jrc10qKKQpjj1ONlncqBqjtqFBc6T/G//H33Uqu7MugNwif/o3HpUN/BAayJxKIwhlzGVpmpNpGF
DglW3qrBbS/+uvX7ouSUXIJeBPcBFgCAUTWf31GLF8DZJ64hqHb96Vd4HgJqXDYPOJkt4DptmyQA
csk38Za687CoZhGfNrs15LOBA5udJM5OHI4fG0S/EXbqsuSQN5t0tlZWr9VJZ9Hewdqi+gDy5xQZ
8tCpj7zkJ2PXGfOrUrfqfDYLFnZAC3W2gG2VWuxjd4tI+T6Vr9fCbAcgua9yjYv37B1fV0sqZhoN
eiOISwBfvvY8WHyZzalmcrHS/BW9oyyoL40UZpKe1pzaj1DcZ7daIaoRtHJDklfCfy3c5o1fiSoO
H3waXdG99VkNo5h1nZemgrMY77XGNGP88wv9DOkXaE/3xD+OVtyjQgs17VnkXLVJwIHMlJ1OUvYK
FBktFP8F3dEFC9jxpJYI0j5RsUWib2qzOZFhtwTwZ/JeYuN3a62s1EKm27g56ZHMshuupeBjgqsH
WqSMXA+fcDLHaBn8rAerTBPQXeQ0fCtpBzcLhYgp1YYq1svFRCB2e89UWTSdzie/rsj4Gk6Y6aLC
09WiTwMX3sVxyipN3MEOOU+fn1baToN2kPKrjaeOKXqhMR9bP0fIbsP3l2e4d12W0L1RpWQV1x1R
Kw4NoWkr8NlalK9JLvk5ns6dvQHazd1Jf17ch+gCTJbMhF1FCGHMwmZqZKnKkfkYXPqb0u1ftOqh
WBNXAafMOLpTaeBI3lZZvY6+ztri5/i8vKLGBg797grztUCiMOx4kPiYL2S28NOcp6rzTiP3/xqX
hrzHZsC7CCjnfCIubg4VeqoG7C3Xg41dLzf/IlHcA2U/o6KJJkWMvNBUBlLwOCdjkfJbZKsrhtXJ
1V7Vni7dq7k+kA3z+THBhMXt3wrazSxy0VlM9ISaiAT7OGgA7z5y8NvDXambYXLyNjpLvydbE1po
ttfJmG5P2HpjhvHY7PnzmhgkiwPA4GBMSEhFTTtRxpwtRTfOIxvtJ3NfeVId8RstXT48MOjhC6kf
a5OL1VtfrdCITDaLsZVYfpc62yhgfv1Sk7JsUqmK7dDHdYTQ266h6NyNggFyiXk0Kn+1MHjjPyq5
FxooBYB2usUNLFlIUvadRUYnHZ9vnFS5ujgKluzoDQEU1lUZxAuxUvmh4A3gRgggBhxO5ljYncuu
05+z4lZFbYnz+UXhRqOdR3aOVPS6JOl1biGhflT6t6zebC62wr+m/DzoQ5DkvGwvfY5JldQZm/zK
7IFK5Plful/4L4RX4EsWFSW9f/2ecohFJ+MSP5IQB+mPv9w1WP2ZfOUYC9Wm2qXOJDEiRcgvt2Ut
B4K+BJ7XhOM8iHiPHcQ1xgpsrHx4A2oRwuetIGz3W1xDs9c5J2Luds9x7nRrqNqavueQgKkXo+DT
3e/2+SqyAOXXyLRe59IXLhuLoNQmDbRTbAemMHwQP45nXrUXq5WTE/ONJFyLvVUwyu2VuxgjlPIj
y8WDksr5thf9oI6wUqb+uQ3vdvNs7wB95vfCrumJm7W2FNic0ifxwq9WfLW1N5BcfZlj/7zeLnQu
DiLJeGROESPTN8IQ+NgdJCCfUTrBhvSftuUVKDYpFOXU3dHxGUAMTbhcj9sgJLxYnGsa0RPyC1Ls
YO2cZ8+VkJb/wajS8AaTW03QSKnnOMiXzFB6BCKwsxVd7hxt6iRP/2orn5f1IZMGfgZhMibmacH3
+xNH7D0vZHCQh40z7+x9GEg9v5Y6+33a6MAts/JwdwhtTMoX/jWTSgFtgGc+kLojzDrdp/SCFCHM
Nb75G1iuPBsMcXFeuW3cKnFFvkClsXMJdrFsSgSeg5cM/opi2t3ZfEEMTO9VcDsISPszCHDd8e8Q
p+eHWZ4ZhiLU9OnTGm5zS6XHFejDFicOPpHBYIKNLWIYuHQrHJnPYrzySWZzbqgZqQNzPld5XeHH
A1n4/arNX220OrIVv6B621YJER7t2HCNn9MFH1JENnEdeKynBPzIwZhn/UHRnqIp1IyVEjJkIZF4
Dn6ZsYQSspk2RhypU85pgE0WVXv9Zj7TKJjCY6hTDwvzBnf3/Y0dda8ZTCDb3NtRwlqf03pDBdMA
+5AKCtrvfZZbWwNUpa2t+SGoZVomdWLlWIbf0an7/suefQvXw+y855bKmDX7jK2QmuDISVknW4TH
8ERx9rQ70WBMi4LnFYO24mGwitcfXD77zOoqa1E9zvQKPI2IRUPvWch3UVqY8eTKZ6VJCbJfm06V
1OhUsyGzBXdU3CihHxwnTRBP2hys4qt1xRWU8qq0Pi862fBEz7c+mxBon8hYn8OuRO32IIBbUPmL
rAsTtSVgtc2ZcefOvPLWbp0x+M2ZtMyANMYRNszMNRTXTdo5TbInapIvuSi4/mgBdQLXWOCJ9YQv
0mm5bPclpmNVkqZ+HIEmPNN8eJQzG7LdpH8q1A7ZNRBn04GGlZZIPxFLH+ZegZFbz73ka5M4d2wE
8g2ROW3m/MyTbLdKFjFi9Ii/R3gBvWM1OwNeEZbCroi7ZN+EmJnab4IAmPgA/NAawTR55Rd4t4U8
RztGBD6n5xintqUfVLpB2BJiSvvFdVcF8EHwZIzXaeZDCojBRYfBQ0hhnQNP5QcVM2RmSokR30DC
ZAsUYSqbI1lGwmbmh+Ukv0pZH4ODKXSAO7HoLFOCAlwC0PI/oeio3KZ/TKD9Zr2wKcq1O5LQxvMS
0No1x6xTGrBeSNUD5t5KhF4Tzfj4tjxqYKMIaSdz2atWROFqHe0d3wOZXZ5IdubiF2IiEpAQcY9a
SZg0es7N4vIXNz9UhqVC6+lYxwUy8Jzor/2WWuLw+E9Z8R9IOWpmOf7FUaj0cRyzEEJJmMh2uzm/
TYGEpflvJEOtNYVme8+EgFHDcvMFeCIM4Opc7qlFAYenYsFu8HbKahntMOuQOlJb55F67FocSYVy
8xMCSKD1L63L07154FFN6XgyaqaP1uZu8m08wBPCnCY5EKyyBDEquqVNuoJKz3G1F9EtPuu7CXv/
Kf03sR0coxNxxq7mz4egXWaDeiD5ZzR6VJaNwovZfEjsFKjYERcjDqZSge9f8jdcikVaypZ5XD3i
JX1UNIIuNMgK9YU8q26w0+vuXBAmS/7CIKU8EfklrhD+KuJqbMEYCtcpDiSxiT6aotq04TxQJseQ
B8SvyPhqHBx2W+DK8BclRQ3xig6QN6iGbKsLI8j5yl7kIzMDwy/MO54rSSFikUzhCuHZLOOyehEy
vqLrYdd3mrCBfwU7qjW8kg8rBybiw6t3cOYAlP9utdJl3D1mqeLndol0aRFdhRT7574xbl7br/ZP
AjCzRE94BOV5WmLTy8Q+Zn3hVEtE5NwoPXnlEY1Cj0zjreJIzLR+JgMy8E3UitmiJ5zP4VahyjkF
hJfwUNjrzq/tZ18D8gJNrfy7YwV2yTUjWGjaMtHtQc9TCoLaR4uCVhuL3HrdpASFRRVrWz+zhfPN
JAw/IXuGkHi+lRvtzVRNdC6Q0tCH5WKpk5Earwrl7Bv0trV4X3nSWViCpyf/hBF5B/ISP9ZdZWFt
qvQVyn0grHclcQOHz0b/jtjVC2T5cmmQ5W0ytAWXazlB4qg6yMvikS4tkq5Cu6E1DK6d4Bbuu1vV
n6qEb/sEfLnGlCe8Av6VjIggsAqRLrREs2b5LBtGc3mKFMhXvfn+Jg/+ErpMKz1UTb557ardHrlF
F9dg1rSbe2Chsd88KIttDZbCxE1H6pHtd13cmES7hpfDo0IDXS4fUJmScESiG3hfAVTyCC3snMNr
JtWNQYlkyng8DKLG4N9SVoLyBEANOc5sjJfUB8DoLIOtwe5Y9eooYPMY9WBNYivQH5ITOJfdJIUC
9K/B/GSohz+d0Zm0V/7GDnfdtO8fbzk8gw/K6vVLg7uCJsxFuMkwZK3SJUL4L1gLhQcK3B19p5yI
gJiAjGGODRrJnURKs6T2KiytBJmNnFk0+0pcHXPD+G/0UJd9OnKvybQWKDBFOdtXw/GjPdvojz+S
BdF24no0nKSeBLo7QdsHCp4JrAIMT6J0ZbVFbwihiGLwJ/an+n8JLIRCdvESj83KlQ5m26sfgwOZ
Xor6nz4YUWWTOPdh9y/+B3w/CnxdhrKnUsXmePFtVo41E5Eak7/dwE8/Ojlho3cHqprroJTpjBKR
RgcxhcYaUtaCCf9gMwWBgv3wEEKQ7E74UpyIV88C1cKKxrlzQlVBGMP20lRguwK283rrZ+I6rX67
n+VaSkFsBN8ouQMu4T8UrY/lwpJvbPBai0sqh/XhRgapl3AcxLsKf0OlPPe2cPaUIb6kidAmuFPK
HgbfYoXQlqYuRTBaHqsRgL7PEo6KCWuNqZPogJUGNFfO8D222qG14fQ4i3fzBCIJa+enaF5DKRX0
SoiSEL+koGjnqSSyAiIJTAaHcVmhUtfFeF4H7Q/8KGhOQLmhnx6kmmpcKUWyGdz0VyRB5M5odT5G
Vc8DEWSYLcuwZ1EqVewlAkwtlSjoTGE1/1oDpHVPCJB4OgZpTYXY3V+08tFwbItof/HKtB1amUt9
QFMXk2jj6d2+xlSt5948ew5bWYe1gKP66NNmfrfWU7HnoYxCYgadooJdiODhAntb0OtuXe8aNOVe
0i7M9liJKS8JSayVj8In5mbwZJK3vBXYAE1NvEp7MNrRdG2wirlYOx5bbUGzJkhrpGp3loTBEmDw
okqSfgpwzUUjJUiZvofowE78ElQbYZZxPLgE4gJwcdTNW8BrLD5EP5Ue1jCfS7WuIFYz97+A+KnS
pU4Uf6JW05M8FqyQZvhm54YxMHhYr+2nxiQUVXe3TsDTvfzt1e9ac+gWlE4hfMIr08Skm7BFaymK
HIlGwVlKWz290ViPyzMR0iWk+psSjbbi90jnibHne7Brb9yh3vsEIcz4Ib4F+3ttETqIKgjM9uUh
XuHVbK0RYMGzQrINbaC8PAMvlcUn4oaFYYsZKGaemF2WrtLVGuEoa7+bUX5rW4uphx+1SxjSbUK1
+2Ajt7rO9FcbqYR803aBqcOALzqTkW8wYr6uZNmb/n9Lr2h3K8PcIBtXthQ5gQ/T9VWwK0a+sdB0
tMdGxYgVIaVpCV6N7OgGIjk4iffOgjGF8fuoYtzIacY1/brTZquXzb8lvexw3Q0Dsz8189Xu9Z9m
Q7Viu5fDF+n7Pc1skgflgtZuaJyAD6OD6KrnHzEgtXb3ouNUmvNvqIZoIdXFvA3VhqYfF9EWKrzK
J4aNnoFOzq/MV3dPyGckKLZTbmSguNk0XGhQYed67gjZL2WuNfcAg19/Dqwxim5ZiG0lLgpKQLyJ
eBPP6dpdwJNUq+U+GCg5ZlPligbSEIXjdUo/Z2z69zfiOznHrjYC1TFMRKOsdlRyC4HflkCjRG70
HbRTTlxesKnj4dA35AS+4XYMwkfHuu7q0fhRUar9GCTO+Tsaxeph0rJmwB468/4f2/0qzjp86q/b
e3d1mHY/S/Bb+Fra/Wmx55BIiBAbbrLQ56F4UAsxY8Yq4Ewdg9hafTTysau1w5K2JQKEOJvEImd2
mFeJpsZeYV+vzbVefojUmGJ9526vJDVVgvaVcnfyhq0EYKi+Byh69wJ2YHH9qpUSSepmn0U//VaR
NOw6GCorVu2o1vnhYuKZJ+1CG6G9uyRTzN6SUmaCAn4If2B7vAvAguSdDGaoSawG4P0tck6XlhsA
bOT+RU47x/2z60+5xRW1A1mbrFWkXuzM1fnT4P7+11SXhgcmEKRPDcK1NvGSqj5C9YEMTPIb+8QD
C09FJlE5YOHKoumuRYfnlJ9tY3jraEO4Kwxp67GSml1a+O1xRRhbmZs7L8O0pCnTT+AQXkdqgvj+
+jdj7NwmgKjatsZavzaOsULI6bLvLsCJJwGS9FhR2On6pRDolCvHO8mRkXIIpCmtc3LeLUkJZjUy
w2gRLTtk67+Pj6FHwVU+ExoE+aadPZ2KMqxMdVYpC53vwyx3wslkMTb8PlaXQT/oBRUEWLspQhN5
kv4YRVWYlKhmXsOjYrSzot6IIOCGeVMnOIThv3J7DnIDqzx598F2bc2auViWbMstQVFjF7NLG09v
THUTAhO4UGY2iXZvLq1VTSFP0lohlz/CV0luFMxjazSlUqEnOVPx26eKQhxEGincOCo5ZAr9P1On
Ao6sZdapMQj11NCvgBK8c3SAdNzwfANKyFB7OWMcCKj87Gz0bZY8R0v65tUN3mKiJ/JA6xks/8qk
zphbd1Zu98BTCTm3AYgcVkg0JQ7aU4SJP+nKL64+z8HDrnpXQknddvFA4Eqr1FhbtdtqwdR3YR6v
Tm/Apr1BbG2KbK7lKCQof2cp2wf2OKMJxbzPP+N93oxVR5s2KXiYVspkzBH0zk9EU3d0GVhQIGa/
AW3Yzxjty9tgL/Zji98EUgeYZn0k4bA6xJkgab0BopYaUzc4Mwwk5p0FVGIZE5wS8T5IxyjILQCd
w8YMAxpOqcA0SradTVWgnO/p2sLfUMvNGmX7EiU76lpRBNx7xCLRjIovmIkLO6OOa+Ugh955kG55
GkLYXEQrtZhAdvXgconh5ZHzSoI5b9sVzScr3GJUTSiPDbNmu5j2tGk5vYfWf8tAP0lI5WYxtfFO
qbI9DLrVcv8p4GZumD3SsD2aSd2kkoc+uSF2NsCIm39cBMxsAw6L4omvDdtWz4pV0CT9+qx/+usF
U8Qlu4qk9kg3h2erCmP2ym6/w57Bb3suP1sX1KBdL7TELX8czQ85//ahseD3WvASfRTn/DiSvffX
3qHElSZ2jYfkN1K19+OJg3RkaEdmUxaY+EXiIih6MOhWxGuLAfIcr4ECPT85cbXbjopnHzZZgIiF
9xNmmmX77KMDm8BxovKU4H1L+p4ozkoxAsuYJpUtuzeNvnfNaJEyoRE/XFiGfxoAuuuMtkZNj72/
JJ86ldI7pAbeHZMKuNo7P7Qe5kOstModVRFlbPI4J0vIAweQ6Ac/+7pPitP6tW5cu5dEkU9esMuD
JRX2tQx6iGlvThqwAXODn5giw0hFVOBup4WvP73iFevTu1VDsWqU7NYSsO2eHt3NPpYbJs+XJhHA
RKXXPvbBWtIrCESSCvbs7J7kTrQPQ3HV7t7Fev8OwYhL8ZrllXxs78rpbK3qLeQA5thVDEL/FUwE
FpIKErP+VXleFjo0TVKmC3BVqkPuc1l5o5sA6HF8X8BnwDLnQtkQGR5r4OPu9FHZjECsTqMeDOKz
S/zR+z1O8ZVSy3z1iAwSl5mnBeVoo2U0TEZmAhKb4U8Mjxf9/RdLvRoP42avIbdU3Fn+1u6vy0jE
MAyfFFN+rxzKydf6Ma1dlutxf78EoEUSgpzaf3P+mteGR3ngYY0AhXH0i4n1y0PAem4hvlJLwNnb
gOd3xiAVc2VnSx+sxVgc9k3E1bqYCcznx4+mEjs5ZXdIw7Vu/l1du1vuHtuV5a1XpwKnoHz9h0ms
Z+hkTz+XzqLLa0HAS1+lJzhRQWMGabX0y/whBDQYSChTVGqKrgXgjuhUd+opUjbBBlroBxLT1xQr
bbKU5nVraJc7m+XHBnExvzjnMvQXnUWLPSe0W+IzJQ5oSOySaS0zS3/a+fPNKkXQj0hNRB9tvV46
y8djh4fjMKVi2q/+PIIT8yyhMGIpAcWTO2d+8+gF/Ot1PGRLEe/8KVkBukbj3KcYS3mCvjrtMhrq
pRSeJFUOWwQ4P5mNuAY3OV2isEdZ05CDwZX1TidA9MTW2B7koLUqIknvnQ/xWBqdUqAYPpjku6vp
T4XhKqeNxch9h4gK4yfd8XhTFICmxuzkvs0JCLheIKU40+KnUl7XZnzHvGxKSlPBxCKKuAT05HNK
yB8//NqUF8qLcGbhNSYlQvbbGYpHKnAt2tAdBd9CjhDVs5fAHsPvWGcEiL8BP6sDEkvjXFicqjgF
BPLvhlIsI2DctnB58R2GqX2K2cR95Mj2R+vQ6TLox6TkGzMyMldftpkuejCa2K7c8oRKyC3t9TSA
+iu55xedn5oMaEGQpWZIwwgUTSqlyXXVYzmzyoy/3JwTrM7GvHbscmG8uC7AzcAjj2/rNYNmlAaT
iS4wNesV6qdCC+et2dFB+QD0lBdJp3Hl4jrO2FZ81W1JUy4GS4ndEST0XSBH59F/N1dEzGh33dN9
9wvu8v5cFDLLgRH27TI6QI205YdGULLzDzMW3qOBTwdL7H+W2i5AOB+aodi8fQaCMl+0sVU/GTXY
fkspMVKneAeiUjyedx2Emstjm2WtzUYaLzVNMzBhQyNv3BJDC72ghZxOKrbC0ZlcE90b0jVTfX7H
QpK/zFtfgCgWuXAkl0LeY2f2LA9qIp611MuKymjofgK29ygx6TpbQw9nSPv1a6jIr/p2VmKR+wEj
Q/nGRwUFKAb09+sfFFGmrX5VEDWJ31ksBwV+J+vuW1lCjrexNr8pEwdby651790INNdYQdkQ3XeA
ev4UgJgitu9vHgDy8Xfc4KLOd5GzWU7cns+xvKEsH4yffupAr0bIVog5m49orllwcn3xJOS9JbMs
kIOb3ymSS3/rMus/rWcsxegZm2GUvrC7lP7bE/zNcOj2F5pBNV5dDcif9mnwTmArR49vYnGws2rD
7snmygzKnMpWfNdCZV0+7T1zvR+TNFdP6yGPFq/hrEHZQHTBFh5h6WTIFWRM+nk5XaWXjXBy5rc5
Prgbe8UpzUlguTrmXzbeO1FRTEzUHFUGt6yDjnZvo/uybeoI52OzMekGIcft0ia97xFkHwW0Nhod
/ty816zhCrdRh3mEN8BtxJbImOVxwJ8FXDG6p5pPxWid9o2B954HBHqzLDdx1v59XS7VcwRt4sRB
Z1Y+1s2VJAXomk6D2WXiDxSezlGnuxkvpG0aVh0PD3X8ryLfmaa7pAGcaHj72geUJ2jh03WaCOYS
0EtOuYhx054NB8g5+vKA3R1B7QftcxYng76CQVOoUiK+JE6fNK9sSBwjsNT8qVv5e3pxu2MMd/hW
cXfcGwdmCL3psE/yKvtnTD5dAge5JkYsTNDbRlPF3kYgI+foX3RULPc/MM1x4+OxgEN+ucI3PHP6
FaW9vtMcX4v/k6xt5PggZ0CVH+HnFVqodyk2YxaOsikoQIIj64dBht0h4TUhOzhxH6Tm5pCO7a3R
E3nwDnYBn5bN98m7RE5oD/a7vCQ0B7B5MFDv1WtSbmmFbCv7rJ+WtZUDREVfQ534TzFxpJVpLtyO
xmbDNz56aPpVKNH43/RnsELmclFBrfJRVoQuk/9oQ+tQJg+CbvwxBcndiqIbN1YyQaSEWdaes+NL
A5vER2vJSMiVnropAudINIQYLOCX482xAeBGdTl195tvEcuq6p7nUUTNIcqzWJ4HfzrovVgA+ajM
dVR+Y4QKCNRyNfRi81ZZKHAc89evnVycVCGDR1OcV5d375AQV8B1UfPNxscjBbuj7+nP0ptA09Ep
HQ7lw+bXWzZbVnKACxByFisDgncxP6davfAgoi9/S5wcRz4lSUyvEfvoQDT6SXImZGlLsuujmWJ2
Lap0P1uNEmaXoi9zXxsun/MlvTohlmOgEyO2ZV39xM5N40DUWKR97u61oStQEOa4TeojWeClCfbE
VRgnkFfe1t2xlpz9kFxDVEzwVDUQnnvIAMBmVI0BcFUhS+SkGKb4DPMBZxJM4K/Jcl+7DAuh6ZWN
7USQfe0rrNzjABDWZ2M0kssH/7oDu5n2114MC5GwJUHust34cyBCM0yxc9vhy5oaIbwMxTwW/+SX
t/Tfv7aoE1aDUZ8xHMEGpR2Ai7tcOUm45swzLKVNNAa36AQiLWSCOC05PJojCsCOX7DmgrXrztZy
X1h1xK46MkLnkAVGG9+J/Bg8u+nkSL1l7YB3ZmVwfhqK29IhLIPhUhoTR3jBkd6H7eYMUI+eOV3x
WIxjFPYSDgnh5CrFKk09WjZNmKe5c1W7S1+VKj+e/yXOaaOpUVy13HHuhz42ztLHqq+1EfqWFcAt
oL/hkh6ZUnR5SGUokbSz5mrX80QzpGvXMcxhtpH2JqZ4KrOFIDMdyuUZuB9kuKVwDuxGYHmbcHxs
0KxzWuLfZryc6Y/LUnHrzcdKhrBlXJCluZYpL/45fwhXobckt33dSVmbhu7sXagsVGR3c63jilRt
Q9ruK9ehe1cU3N3iQe15SVZSq/X61Hp0DoY5fAaqHcYyPndNvqiyz07II02EG/E7zc6vyVF9uiod
AweRVVfgfhn0Hdz78E5BK0b/wlvP3Dinh45rMG4AIp+nlvtkdMxf8g7VNTQ2se2bRA2L02apkzV4
WSSPvipcLjbydumCsW4qIqElsz4Q3erJjV0tzODV7BXmDf0ZUt4iyR81WykSTxmM5XH1g9rSQbOU
kLYUVSNkfpp10cQmHs31N3fZPfFIGDUSb7Gas8RtzLOi0J+4oPsXAevtXi79xka7EwHNf5ZlTPT1
097mDrJmhUebUMlyIW8SRflTADH0MGhjAbHQ3WtZdAHwQZGnsDE8oGobmY80HIqW4XgJmmknYLcR
eY6Evha39mdPeInSYS/VgxI+iNRPlwuIg3ni0FkndHjlZlAQmNPY47OnGeMHFBGuhW3FfwjLxtpF
ExDK7HKqkWR58r8vNwWryIZPgP4RW0KTLzlS+cGMv1MZEHzNMYp3pGE+uy3Cv0+ZdTKsW+g6rV82
Z2ld2t53href1ZBxi6nmhMmHyiYVr7ttbBw5sTaS6C5ykxeetr74d3z7uuZXCBzGhxyhZ77ismdW
6ue8IzaOPgAx/cSzPmqs4rkXDL1fE4NNGozzsnXsE7/MFpK5DAakxOW8nSTckCBQNBo+uOjHe9ea
S7hRB4R7LY61zgBhBvn+KMEAS4qYAA0KX8AHiT1SBqJDthaNCPg+1X6mEcPbqaJShOTYAiGlnAYY
q7KDwrBy+x79KFGpx+dpeV485BDcMJUMku4AB3MHtjkt6lW/gIHQjx3lMsSjA7eUEtGgKEU6bjtc
h6tpKd5yNtRJuYA7AyhFA6j62jH7jJHj8PA5PRU5Zx7b703m9vyOIT9YI5PIVOIXK9UtVi4CfoKk
oVI/2W9HFjj2R738jOAklHbrq6zjeaiR0dIUaTbm2Q8CossR2ViuvjR24i7EBpCPL9bBO0ot7yry
45xPmySDSwrsqr6xisEdyMuV2BRumaIVcxBO1AlZIPiAoFMRe9Aik0fQlf7gy6QioTKVxW40f+Ju
iRmwwVH/rOXnCBSd+2nrz3pkKg/DLjCSpLkr8s6rq0MUqM/TECaXf64wT1kK4s4t3cMNSn9/SAXC
6Rh4YfQM8LfPdZmPoHWqIcmRbXwP16XUY4If3iaZgX0JqwozVIn3eGKliomuaIAPQa5o0/3x0fuQ
XLpm6ueeBNYEFdHhleH1ST/OEWE6M2OROso8Tg0X8jSEH8W4r68xSmiWTw6tIMYGCZs55oMXFw5Y
DR/LYghC8nZPFzWTrwawkRyHzmKNT5T1RwP1B3uMJBYTX/kxTv0sMEr4vhMqtCfKqzdgAuyq0LKJ
wFf/ogfuW/GP+M+5FBdgqxKv9eeDRY+rIvl9TN/jnTv36o2PZNk/35c8+l7DJMDgt8uIGx016Unx
/UgJLNcWG2rEFXvxnC3KLosSj6WeIsJ0BdNDgUAk+8UzL56OqycY0KmA0wM6U9WQXypVNPteCOL3
k3Dze4knrxoU1xjLwDdVnalw2GG/rmH+jkW6L4wOOh4c7WB2m2DfxbYFPVSrR6mGrYBdcwYAt7w6
xskEAoOq1PU2HR/vgKif9ek19fm09Csdj+/LQnjYQZOfM5OfiItsdhE5a8FWGIt98YZVkNKa3HhT
VnHrhNwU9kxiCQXTfXR5SLZpcz38UK59la16XkxHrDmIF72hO+JOoum2NztLOvc+PV9w9VrsNSsl
b9Desiu+iqxb22Vgy5qkrFOIxkaSb3O+2C56WhLDYEiz7R8IviDLrVERxdAWUzQI92zrXk9aemEw
LAJ/ovXhuUI1GqzFxSmLKwvuPUI95oZJzMM4Td0crRUpm5y0K15DpKAuR0maBc7/WWXtFLLwDJ8H
wRUrLMIvBu29rSf7RDHw7Yr8wecbgDh4gv0e8DxEchdVxPiJE3mk3BMpUE8dSDcRR8WlXUskchHd
FRelMik5ML6IRuC1ILKDsnVKOoL5tbHLy0gDjW5nxUJ95OE1Yemeh4wH/qzi3wT54ux727brLTBv
Crb8nGirhCBJ2VmYvSvE6W15+Vld4Z0Z8bJI6hMvNzvXJxbyytBHcXSY4osrYqmlV0O1dxLYGiNa
q4QQwifYl/uTR3g01wprnHdHT7qUEEhDmrNYLqG4BU1o9ZaSYSfyanlMfIN2qCJ5CH5c7aVH1E7L
3GNml608gKEGNE+j8MyhSyR3SVy8prkgDJgt/cDagKyABmbnSiCXFoEXL1KW+ZOaS6yoHcno5M1R
ZByxPEDdJhzSV1nHTCfyRe+YaEPiL6Qp+OdNIH8fLnPaKL7Vsfp3ZKtN6hi6yd3sAB/yZGt2ApNN
7YyVh/rhIvctaR9vZmK/SXOKy3q38xeuzb3uc4KWOhU+rl12MDlAibpFIil2chpaw9saqmGNpUbu
1hyfsSOXabbY5dy0UkJFhzBveVvnk+xJjigxIhdr9C42fl2hw5ZX7EEncHhKNYcn2C3wH9pbyDmQ
PWRgcqR3qVPHzUJaWRMdqZp4DnzTNrolOUMS8/j25jBS9MNY/Lv3+3WUg465swZ8VqvEYApfoXf4
6WHnn4Mi6voDmwBMKX0H4Bftk0voNnv0bpv9Ce+uSQB57Ax72fJFS8KGuOAC6nS0Ie/5NCaBEQQj
P0NtVgwT179U/VRedySV8HccE8nwhGUatYj5w46rzF5dQ8TEjj2Gp0uxmavIBl/djW9uYAU4UstR
WeT78uHJd8dVQAJ4FKi/A19Qd8wxupt4amBKTumd9hZVa5aAKtobv166U97nKnF3jfABIAxxcTzO
KEGKKfE1oP5Id0ByfQxJcDkDRPqPeaWHDFKmItYu+VAqzsPab2QQcng4PJxvM5+cvMtnAYHDOKk0
vskwIKI3DZ9HFbRmS/4gyXwQCdCRCo/y+mIYUTfis8EFwzbo2kg0HRwZ4QcMwtHadDNXCPIVyT1y
6Pp1osLCQgXTexBYhbG/Pj+lwBWR/pLhzXqRV5uxKYXp9HDa5x0bzrGNWhvjRl2m6GmILF176ohR
wssnPjOohPP4r4cHtCX5yZbEn1ArFdw3vW9Guws6UssJ4XNnremaMtf49ELgvnIGrt6qquqYoqCJ
5zINOkq7KbWF0PfwC2snXQjx/P8AuixLEKaLS06RKMCKc0zW+98b27iN/iYbcbn2OxMhPyBudtvp
fM45B4jVMT40HM6MiSqfZGe7BzGVLDdlu+2lIeVCu55XIxmDS8JIhM5/SAthdikAzyKNL4usvha4
RJn98x5wdif7UWZ+vqDlLXkFgD5fhalosTcnDBcrEaBj7oqD5cObezLxabM/r6RpOz/cQ6ERtxCS
WPys6T/171QCd64GkpOhhoJq86UPMBB9OSZm8mb48vVDqBeRvhfEHK/7Tvz1kF444w3qU6dbywmB
KVdJA4uJCV8UmcdtbsD19+3/H7SLM9Y4h97mbvDSTLsa0bIqjcr15RbkKBq55yqjhPxwms+toJIp
e8iisDhU2A276XwlZMH7KWqMbTomoeonvfAxjSuyrvjTPsJYw4Frjxb0aphlWVn57yuCF2tbiTjO
OSarvBZQAl9PKweu1OGofClqJD5ZkcYZQP+PyrK++ORf+sRsuFas3nTLYUcWXMy/7KoBIoNEDxCA
+jDF9Z+inmv4+1NGtj+ghpDnta+Crxmwi2ePGeYpuZtx4d/EUHa75lBAlj7yb0tS3N4/2CQPPjtV
1QuZFYfSJnrcjMfCCCpp1efSmVmc5gsU/ais+wSZMOi6BMJKAdyYkXB1jD79OHP7rUSix6VS7Agp
FyrG9MOMJo/2IyIHajwaV1H3yJ8pNv+0xKtXr2v98fe+RpZ0eIlaz1CTffoTSC1DmrkzP6YwDmZJ
M6u5fYYLV9XwLxgtazKcbtYVhXoDcbmix00px5kBm9WZT3lpkHDcLnx3xkTUuXSc6qw3YCUC8ajC
pkmCVEIj9F2zDz6rqDsO0/vf9ysp7rvVEhswPv2QQa844XxzaLzj0zRmfQT8w5byCMe+bzb7+rqV
Ay3ZqM8rVZtKEJLCv6tl3QCM+Xc171WdkY0Ab8rxbF66Z4B9tsKVagr6z4KJgs6A0mIUquf5MCSV
z3cnlGB6+v3a0J2sXNnf5T0Gyx2vYNXDeM7e++7B+3f0o8pqu5JuW+KJlevAEPJXaiDIf2mMWRjN
a23ARdXvfGJhd4mOQSQq8rr1CcwNAaUkqH8RPeqVpJ+WnyNFkE7Okt/wFpfuE64/9srEwg4glaNF
PR5FwmnYPPsZu2NFRT21geFFFXG+d3OIL2TbLIkgvr8leIakIK9V3VMa1rSc/VAdfV1KB7Ci87aj
Yiu4ZxMI0epi6lrKjpeXWH1OCnonTE136taSzhvdssGiQB6aNF5Fa+UryI842HUMlIXaHlXkeZZG
EGTASgISabOadJR312I+BiB/RrL1s3UXIBWSijvNvXC+Z+Pff5yabrh37AE1R0OoiV/EYIIazWYf
C/R7yIf/+gnz8WGm+1Ize2V6Tebk/l+xC6buDR9UW7g6hVDiqiWGOi/VfWo7zIxhkyAqV9pcpd09
0j7pWoQtRM7yidcC03BeLgi2VVA1TCqgjDoepKNwL2mpSwvu+9ggEBY7ZNvrBJp4ffmKw/njJaNB
OrHxYSXVg72AHv8k/9vQuC6mlgXumNOMOZWfW4xxVUxTRZoptzh9eY8Edhe0oBEg0WTvnDAgBEb1
IjM4zV+SFPO9OHIseIkMKIeDH0ExzTyw+pyLgTGDaQzb78RFr3kLMSjL1sm+C0v7xAeGlUraCidY
n59/IEvDNra8pblqH+R5z6cVw+9jnVifNt8rLnrGNkHrbQo8z3qO3TTvhvBfbCgc5vY3Inl02SeL
eCmC2Ffc4XYVYcE3rmBbsQWIY1nc8TExcIRbYSg5XGCYpHAv0nEquxDRJ5h9VBZFQA6UqW4JJxgg
uRd/m+Ldbfe/w/lpjDa8wKeBHDqaTD+YeDm6RGsQfablyTq7tleOBqh4ppGQP2YqGHlT8/CxhOvW
wWm7NQIh4aeurJl1edF9HqGHpiug5zVOOHuYA5EYqCv0aDH7GvEHlLDotuuAoAias8NeFjSPnKAu
SDwxrCqGqsnljACvzLbiv8X0iAju9TRYSYTdUbpZVQY0NFHjl1WfE+64TchOP5PWzi2aG/TTzJ+0
UenRPovXU5L9L7kxeEVsUb9MdgrkK7u+ucGgSkYYG7McLPhsRGYkTS7pPzSxxbwK/Eyj5y0cMu0V
jXjbrk+qMhlC/MikmOHzbRq1DChTlHruMLX8I5rPqrH71dMjfDywThzrLpc6YE4T/vr85pUvq6AL
u9/itsKbSRgMPlP18CGJvVziiMj09b3T+/Yf2sk1J71UI2nM2EObjkmi0AdNRkhIo1yDRE6FBt+T
laAm53p/ZqkxH+bILIwcrvpWsw7b0z/3/5loQazR+YLdCQv8fgW9Jjv9PGMLNdkcdErHNng0NgXq
pzBgvaExXrqmOTguvvm29WLwh8G8A4PQqcSFF6KcDwl3Xv0T2wotOroHOdQIAvbmW4bGB6e3EHrj
PU9bJkjX9KUOYHfiH1SeFtZSqTHHp1e6ebzDrxFuNAN0qZP3GPqSZO2mcCytZSjJYBdytsMDjddY
aA3zDuhruFgFHc9EC4Xs3Bz+2CB3Nqg1BQcTe9IZFIELoP0huOf563IlKcVYNlR2xBGqOwv//UoM
oEo+9YdsVvzrD6+YHYdTHayFgfDvYDNXCuH29JBbgLNlxIzvFNMdVOv6kWuFRirJNEBS7YyHZVOn
eF2tEBKXf40uLkG7MfzIsqTHFG+ZJYIk00z3mFYEZY9qjWUrONa4j32CwzVvG6e5FhM8HRJAlWVd
un1PKVkPQyZp8P5UepV4m1jRGPD4dNwe4hrktrLr26GB8ZZN/HLgjzPHsHj73aT+7TCSgW3EE9Cf
LhRlLo++oozkLAaZ0AJwxiQNJsmmi+lj4MkAsERnlfS0YT4qkpRuS3mcR+f+Ig1yiMuacu6FneKG
+3WEVakIHhug8GydRtS64hp20uJ7mAix3367vPvhqPZyt61P3SEQAUI85Sy5vhVyEHcwBVNi5emk
RA3+b6YfpPAf74giVR7DWX+04hYtjer8kOTwhM1CJblzjfNw4MO4tOt8jegxZLHmWmhh8u/SgXWD
3t7pDwUAJ5zfRUzIlbetMQOi7Q3MJCEv7Pw9vXIEt3AT84qADcvy/uan0ThoTdfOnE/7R5EHZU/N
EW/2QuTW+CgdNhDyhezpUEnR8z+jrbjCzpQDWDHE0jFIH1Dno7ILjYNX48bCZpkjBY8etgUyL4KK
cTOpyBvqbla6Y5QjZzPGz8//jUTMlEs6bg1R3kQ+CFPDjokDdyF97aZN/TX5DFnTTsLct/BevK2/
JMEBzBgMf1h30pbzBIlGkfs6CUHlAaC0UjogNxisZSfVSKKzwMlfIXkOBmhw2151NAEx0+4MAMWO
hawSAendpyiJMa5bDpulBzlbnQHu1Dc68x4KpcuKWSeRMnQUbGVDJ1+N6HGa8QcPN1I6dGKGmUfd
tPe653w8nMKCAf+j0nTPUvJC1TMDFxYVTk2tRUbRMU5uHv8Nwj7IjHZogfTlS5W2O3kBINVyIRfk
PuTNOARtGY7accwwuk9XVfqjz97asNVM5Ze39Zb4QGaEV47+IM4a1GNI0mSHDal8c0G02ZowmMic
3EahZ6bg+ngXajYq3S7GYqA5+d3NqWXPexb2tYnuYkIho+PLI3k2OESxoB+9BuUkK8oAfCW4vIOj
UYyVSIiVITxSbWjZzyrZbLAZwmDpVd0jNrqP0VgiyiR8dEZQEzy+fYHnJlCBLKQccHBzTMpEwDwQ
fVE6QqKvDWmFYIVPJ1rpgS+qEpNzFDQ6MmpuM/GxBxMasnfH0V4PVst3xu2EoYdKlgVXdJ7e+FbT
VNMvSyDKi/r6lkYi35wLRdoKQmAL8GOheE1wnvCPFVaQpJFpnrb9ejawbN5RJMFlf+OGscmchIPc
x9VrrFR4PWQ3Ut7F/QMpJAfFf/RXEbNARAxhA8RFfVjQivVZiV30345MyUWKPS73HL0v8Vv2vS4V
sizsziIMEel8/A7t5IRzCAROzjsASVEFeMy0zl2USs96BKy0O8b8YL1AdiAYbn0PD+YxXF9IMINZ
ooXNVIpSxlJ8pvX4J/YXUhbnTdJhCvZBPPtRActeVYgOIHflD+N8pmlq0bgKHUxGfeH0VBQSzbGQ
2MlF8GJQHU7Zd6VcZO64eAOdRXczHD/WASizDuUZ0+eAknAKPan5Q9dla0eGVKIiLkGdBijfCwqd
loQ09lH7EoeihUfcOYWkqnHL2VLewfioHI5o3pn9K9vja6GErj5vj6DJuT3aDvVcpby91xKv31HB
FPjAMha+DQ5z8dmcDV7SOY+F3ByTHwbVNICGplshnTzJzIh2Zj1HVN4RlD24dZYJaC9Jm1G1BR4E
gyO+inKb6QDLarbAS7jedofBGTNNsVWPYX6oeNPdVjqlH736qJ+l2KwnTqgTf/ZAd3loWtz+MKmp
RpF1gZCo0C3Z+qwA6aSmnw+QHuNFQDDXRZTo3A6WjavodNkfPasY3QC8Bq9KTCHzaNtUk0uwjxDK
M8Hs/V+5pEA8vyRjGBERg/SKraylwW5bn6EftfwvxN3H8nFaTEa5NOQRBuBob2pKjhuOS6lWioNy
6VmmIrX+u9OjfXmBc+5wsRTfACDx88vW9tm6uhp1+m0jACMrKXuxfjYhMLwBw3EmoaW70uVsjyTy
f+ie/WQdl+8JHLHfu3VWYPAsWPLiPxyx0b2/V/iu39C4tqq+jQb03bB0QSB2Nr7jS/pdxxI1+G5z
RFN2RIMa+cghtv0a1JuXZ7dgg/LO9H7spwMMWdkIiRiJH57xkIUQDcC+Ci+mZ+gLixhBGW9q/C66
FqCAX0fnCg1pH/9EbbgXmkyKYGWAf6HrXd1z+eY3zlfUW5Np3HcrQDc+bxHMyRozWsBs8z6zNd6H
TzzgHicGggQndzzpLME+hh6ING3208IKiJKofcHbDz3+75tZj7IbSGOu1tYX8MwJleGcHF+JXRkP
byvGHqTqk9Kh9vpkfyFbVOqc73a3vQnTYh4lj2DQ+og5PcFRWjI6R20l/rR1L342AqNat39lavrh
knAvWbPcZwCvkCp9zSOnsXDOPCuBjjgBX6UVdokqymsReI+dLFH/OY2F3tjvtuMnptelgegwXA27
8k4T1o6qHIHULZfGQJ6Lh12zGTLCa41teXk+FSJCEbKsWCQ5gLlvmqHDB+7Fy5cQwV1+JxH46F6o
1nLGjEkN7qr+lIEluLUIzZUHfYajNvqjGQ6duni2mVwXTuLzVIFrKut0tGcryB6s5lSyJu59iFQF
FleGausV8VWsN4VMYi71sRCvObiscvCKn27Oq2T5RYW8B2NcPHq3McfVYfy+FRCpai11zwQUtvvx
J+kDazpLPx89dvXO5sSNH/0sXrCkA8gESfturcd3+MHNWbzxZchy1ege2jxO7T6HraXQgln0fP6E
DLE9msSu+s/C8UDsBGygOquAeXP8UwiIMPvZCOMmmkr803lUckDZwCyiB1sOXtNOVpMQYIlNTRhC
G9lz6P7K1EKHRaSGSI2E3dT1rLhZjJvPUO1eR8ROtZ4e84HATRCPreD06bBT/t8Nk+kGYsVANamM
kPOXACTpx2n8hADboB4OCmfoL+H3rlWmt3uNyg89A+ACvL9FiGQQMkBjJp02PvaSyYUun+zbWcPs
s4EesAEp5J0Lh9FQ1232/Thd5kusCbqEXi9jdmCjgANczlSF0xUTHeojh4AALs93Q7je0NatJtjb
zkV9sCflXfiw4fxmWGszScNzgYLPocE3rL6STbY0mscEuBc65L5zdzLBm42cYtP+PoB1bdKjs3X3
3ZeZkeobaE3X872cg1px1OIwFErOMx2gumelfHbm/njY7fX0xDkJ4rSoEgsZPz4Z2T42O3WpCZxB
uijUV/zoNqkwvNkdie9GVsyGPd7T4fcnbzJZe5xBkeA8YdYXR6U4ySi+MWK0eX6TZiOe7++tAXIZ
RpRj3FiZSqQz3ITOjUx/Z2bq7jAax9Mel0Fg3eJpP/S9bES1NWtZM6LhVEshLun5dIdE62HShp63
KIWgtuf240lePcA0xERwEMz6Gjc66k6aNLSUcjGcQR/+ipflCFUCJ3i6DzDTtuNT8yMScfvFSfQC
KiWQicl70FWddtOGWOrcmJYNVbfitPiOsT4p0h793L4BHosUwSjtIDL6OA7NcLGefREdOimbi6cr
V39YEQ/GrJEIBpgxuByqHsuKAkseK+hhxlEX8dd+m1AOrCkqShje/svx9/oPFD/oJUXvE+5MuFrI
Y7GBifuFNfruvMtEfv9jSiIPZF4qfm5FQFOA61De0XNGj8iICYMIZrftEsNmfhWLCQ1EH6N0jhSb
u6KQ1JYIlbKfMPbi+Q/hdXG56IeHmhwG3NRm7FBSfaRA+Cc8Gp28bfvrJplVLx2Q1e6Oy+MicXf2
0AcO4CFLWs0jYnDzSghnMG2gtvLFmJZXzRt6uSBkMT69cU2R5VOS3Ewtqe+5ni+JlD1va7g9zRgj
+BBMyWcXMTaUMh+49/jjnrurqAmENoDG4t4Q8W0RnlTzxpPD5N6YA8vY3aBlWw6R2BgvYVAgFyBu
Uu/HBrU6pDlxguzESH2ne4hszEOQNLjkChXqQKjDPkQMz/cJDOhcCazLfZ/FjY635zmSa0JvhBh9
DhOR60yEkAzTUZogznYTe1d3kENiZhdjZKCjZkTUQY0VxdGBJfesTYSoi0+w339LhiKdumacRO2k
nLDaksZIduUEihnhcqEZIdhGYeB5fhIpyEuV73oBvnV/gIr3btruX3f82BVPVw0eRBS8YpOuT8Hp
jP4x4oj7E/jd7zvtsBvVK/ACISDyZW6gWE9tSOnxehwIskHlsYU0jsECmmz642VCapBWB1rRPIpA
jryZ3/hsr0ECC9CvdV6ZDVEWPL3wef5r9QN+W7Q5M8lLuseSRVMSfJhg+fDdhKkQfNSgg7EBkOhj
Oc+czXMS9+Rt54Ts/lYPZUNFMXpCuqFq5XqWSXVw1zLp5eenQPHIZ4F4rsg+mdZhp7/Urvwp/XIG
zN7XtQphjwp3Cktq1vhMeN5sFCbkhmfwahOfUT9GF2jaFKNAG0Onklm7ulyOF+sPry95ktvG54w1
+0fU5tDvxXqyxMHbsY2oXBjsysk38oXH4W1SNjYShTr72/R1spoBKSrQyiC3U5h0sCSSXBX0LaP/
CJV9VFwGiJsCyVM/cXy/UwyqZU9H3GxIiPNRtQjB3EStrU0CaCJVXCu12jsWIro8pFLVrmNC5/vp
FpX7+KWohYxotC+4Sg1HOyfxUJI4hMbCw0ih2yrWB5HTEfDP04K6dceBmGXgt/9x2t+BpufY6xqJ
2T3/F2nSCtRXFG4rfb2oGq4T0/5rlEMaXzK9+HHN6k1/bFaFJIqPaSgemb/V0Ce0gkYieenMYwZi
z6pPzUpbXa4KM/5manx/oW50uqVnJU6RyNxVwzCoXxRfqWV/14EZu6bVXpLi/vwHKJcP6KsAUTLL
zuEZC/q4UTR5xMYWjFndq4A1sE+Qkw30W3KXsnb9NnIoC991G3jQ1Ji4eLTQdsD3ZGoAJPjfQZa1
AqTcfnq3Z4gCQcnLJ+SWb5byIE6rEFHEkQ46kyw7UpvfaGDZs897qmJ2+HpGMrajwNqgUct8AxjR
j/mpwx5NXl1GH4wHJWpKRsFjJzbjpAR8HzZn5eYb/W9hzVLw4iAL+pTSbmmMGNOcXANew7tDOawN
xOoWcExDkyS7kG7iBGwQrPde5lAgqXzLXF24AJ2ulV7vBbg5hvqN+HVawIVO5bv4c+lEAbF546Ul
NTk7TwYQ+XdAkgbCo81W1ZgOn68HX9+wjMfZnq/AXExelcFaDR4Q8Y7UiONTyARR+mqeaPEg4Q2t
ZncPnbwW/WxywpMHUSpoxLjcyMy9gjjS8qJcFHNX4NhE/W8GWYDGI6JoQFUcfeYbxRv20BFEuZkD
M8S5i7FanQj0RZTCi+g9tU894I3XKYO4FC3t9VRgbP9R3t3I+H4VOYVRSwqq4YZGW/mbyOSTp9LA
aGteSUyfT5lNjutGNQYairee2X2EGNuYDzqqVZSswlsdQrGrASGX142DPIHlUW8BX1jWKfZI3WDG
uCMg5nd85VkK5PCTV4opCRhiz66L5ERiNArVITBwGnp6SM5CCbPibE3a5cdHxzfAiEUmO3FzU+O8
pcxC9yKSBMqsb17mDi5xtVC0+32uqnouFjaJ87Yz8GpgDGv5LMh1SPgo7r14WFRNrUfWaHHpYmaz
Rz8G/dY5Of6Wpvc5BaxHSyvXGQd/oBuKf+V6aYqji4lCg9A5GknQ+hQJOGnCDiwWP63CbO7zW6+Q
C8PR49EEFXBy3Qe3KV81QMOC7o/r0vwa2SXy8SWTBP95liqxBWGbl1RN6hrtvPQSM5lpfHfFE5oK
iHwNXNzw+SEm+O7DEDtxVybdPjSvw0wEmT5e2dtiFacm+231nooRMzJsxjykqQtpjIfG28IiBaNF
cGYYfBKtDQLo9eXjMD0qRAQqV1JXJDy+z7oWa37o/OIytPcweH25HfBNqhf2QlgDmr3wkJzoGqvK
5sYv2Bt7hh/qvUSxa3eT2L4x3g9eISgKanjlGxq685G0O+bCYxIqLfSsfZUTVZ1ArafYiuCTGygx
RSsmtbpoDw+OGAVOho0B8q+OlJSEqfi/137yTWZXPnA4oXXNfQwnXC1OUKqJpAn3zQYMXJ8ZOgJ9
DDVKjgskW0oGaaj2KaoENppwJk2Z8dPDg4ifLNnbtK2qdW6Yp+2dCaOK2WU+wCSj8YDs57Miidaa
nzE7rCZcQV+OGNnmCyiggANkG6ybKJzO4mI/HPNhmY9Pa8zPMbH5FzA2VxN29836N3U8RqFADlx7
uj4rwzd4qARlV9z4CWg5la+G0+fvktSCSFMY9zgli2v1TXwN3yTl5ngQhOoIjSXQWfBxt+EI+MQ2
QpjABdkcuTRQ93O3/oAAEW1hncSSVUrVeo9uSa86q1yG2hKdXTWc4HjWDPlYvEuYM/Wi1feK0fpU
02BYfl2jgKs2Kf812ev9SpmoKr2UgXUhQQ4MTAr4by1i7r1CCuAHnJEnB25rZamT7yQvSjuxJnci
Wt9gHrVaeLx35eLIuhsfMwk6OEMLapmsmpuKEIdED9dETCFJC6KbhJRTR0AUX3XI9AJJpxwhFvvd
dTVtU6CJfDQHkxsZtVbfXtSlovgAdgbdIY1uVOjYhX2EN2N1gE/4Bp7XICF5X/4dZASJHb6zKlEH
eNe8z3YWMUgL3AZMhE3o0MPbk2wzIVrBreX7mZEp0jZaBh1YfxrISykEwUBlyH53ipFhLIt0J9j8
fiJz3ND41dmTh7ghJHgy127JeFldJO7qnswDjv/XAU+s1UCrrZSSQzOopHVM0OZCj/4fXVUWHg0a
DfA+W7i/AySKBfG8oH+o3J5h8InMLNImEkCthwWr1Ul6lbbUG3ztWDkKBvPmf+1A6vFCfRodeKe/
1xYUI8C4ZLCG8q2mUxNT/eDszrqTrwO9OVNUiJTOjvB/tUq9xamq2T+x32bKcBjedaymj/HeknA+
FXD3LxHOfKNJ+I+ej0OxvCcCKhP/mJTyaeFOt1BfSzDkRy9G+rcQ5aSa4jYJH99LSKphRNRok/mh
czJzBlqLCnwZrqWJFahSJAJFdVM71ltpXQcU+YU6j9k9Y8zy03zBacNfJhoD6e1j/XxyCFWhaWU6
zYQyjGNNuorYjwPMkqI0AUcHiDGMKb6xrcSfG9vuv9KJ2Rc+VNFOUlMF8TBwCEcNvB5TAggEYu3e
dWtkDHwTJHe997zXKVTsj4a7cB2DLpjR6OmXsP9p751gXt3bFSxwbgq6RzEh30cK6MXUFtxRAC78
cewi30EJ3VAQjLqImA62l7tw5lFjlb8+We8wh2kUeiV+i0/riqxYQWiFVwwAS2QRw7ljzTk9AHeb
A1mmGinAZ59KoeHsm1YebEL9FV5oAbLBdIr3CtQUAoMaqoKwT806JA8dxcdAKL3O3+X1c05qLtYu
Eo6fjez0IDWkYAGwtTLPu6kLYQi6FDLSf8c1SGc6Fej64vLCal3yuW1p/Y00zrxCcksD9IrD7juj
6qWsomR/DtBxJoZ6O5jcWcFNDBqKmdgaiOnqcAFtaha+rusS/Ue7suIHZ/LzjgJv/pwhOqnngEqG
C08+jxBkWiJU/CI/VGeSOySmU1VmthA/iWpDL/s5qLKbB/OyWmxwmC3g3FhI1XzlrhBmj9/bUxK1
twy3NUPVDZd78LWc1EEeNatoO+O9T5V44Nzs+5LoaHQsQrltMDn7xAz1I8NPxhMpIwipmvYfn/ji
5dQZdcVKpLUFzHeLL818gseeW4ZcZjAd1i25UXQbzTf7KqV/y8yuUb2cK2l+CfAf/CR+4ezGbmLZ
syeEQPJDJWCZ1EEbo+LVNwz12rriASg4gwH3CyRo7Tl1Oy1Mhg3+OqJZPjPTnXy0BEppNGbmMGLW
/cU91Ee8h1CdXjvL1R/snOVdiqmfeiSNJ63cTWdF+8nhX94veqp0/URscG4ofw9KHq+JVLVqRTP6
Wv+tovDN2VdMYFD/1Bou+qDkIyRCnTi7gpICC3/Xmzg4yj55IpJNr3zbhY32TzFUc/oclplMzEES
TXCS4vpjraMTooqfJk3pyPYeSGPa7rayl9gZeWEKii3S6jpiTP91FCprTRmf3oJ8lb0tg6p6s4rF
JditNx6K35UTQxek/CEQOJvpimibmIUUJXgWJI09A1SbP8tMOc6R5PzsLOu8mK48KmrK728YKa+n
DqpfxZbh45tqVXbIpaDhOILVAhWvvNi/yxzLgILDmImIgR3RvAbWxYCwHXqL2BQ7t3e7Zuj4aThs
VwNEs9T6tDgDRNzmMXBRiiiFuyffFeAR0ZNOy6E5Ole69l92EO6DG5LhfwxdgtM993ejPK6jRo4L
7igXKbTNZDTtqz8Ih1xsJm7tbbLeXYrG0kCLGq/3+9YGDMcwWXrBOPzHfadrPrU5D1Jw55UHXX9h
1paYQCkQRgAL4qETs/aTfEDjSCJaVk/QJarEO4ih60bo906dYbcUc6azocon/mEXQSIg5Ju+ow+N
yV1S7L7ep8TkdZSZGBML7a8JFNZpbSiQSx4JlKFruIkMpCfgJ/tNYrIgMUYIKstCzQu5/RXZ4EYL
nWBAa8yCQfXk2xKuEBP89iPkBSVOy73EFFYx+jm3EQRstEJJRG79dQrssqHhEiVNSSLbiMmr2YQO
NenpryvRor/NDiGFmPRQn36QPowd/5zT9pVF6EIMf4j8mD3Zl6IKHRZhapi4HS1EnVd+B2CC/yaO
OzJR1OAt0FruSGD0FbGluwKjajjJLdbAvNlFD7fBihLtzl1OCkV343veeV8k2WVofKOeHrsnuY71
tONVcTd/UZNKWwRh27BL9+Udk5bVxtUmgCXSxFLvwt1hBwvv+kVpfIBlS6cmpe2Gbpoms/FV2qyr
47JM5iSy397qKPmETOmbtKdWu7qmsjeoJ/yAKmt7e4CrkwAxTDVESk2yEq55MkN6mEKehj8pwOrr
fjAwTiza27hYNZW/fbkRTmt7oyOSz+WhZXGOvq1HyO3bDOvFhc7mKG2KF6lCN7M0ao1IwCOH9wVs
hguLx1GeMQgEH2X1w+jMCPmi9Ct7wbXK7Mz5FBbFjZMJI9EpEAAyQtC+LC3EEEub7AWPruEwq3+H
ErgCBjMBKrKprlXQn8Iay4YoAfErTChQO1elRDYaHqrt4l/HKAzP4GBpZxH1K8LKwonOyAaHA9oL
h0xtJvHXTDl7FGJp+Jj4YvngGfG1Iz6Hbuk6AfhbmC913dxXesNI7ckM8XgaWTu/iZ40qcDX2XPg
rhU32824+59gknc+vmuav83dye5urh5AeefyKA1tLWXBFeg70u/FdYRnYzmq2wQb/b9+O8Czn7Cd
Wp9qu2aixMUmfAn3bM+/mFmY946RdEjDcJdZXTuSk8iB8Eg+p7zxmaQjztzhROm1rzOw2tpamx/H
V6X8LB6Rm1wECLR+gvVuBmEqTyGz5ObHM1D09Fsq/fjI8KGTepa1VhFTIGLOdc5sRPoLJZfkW7J6
4vsV2XxTolUoxvJNxov3yjxzMhnSG5gwi82XCgrOufmmqmRvhaoishSO8R8qUNdfnggrUXSJ7BKX
hLKdW9S+ss0yMesX8/9fIpUH6pFfbWW/ApSGbevStj13AhP4jlJVVdDKzVj7tzo27m8asFK4x4Rs
Xfne5jzUnsRACX1aP+7XeqHhk1IOSRXFn2ynVf4/uBzk8wtPmLy0ZBvCSXvSAkxafqsRYySdshwX
Eo2wY/T9rMLvZHdxZ1vasIqtlgul41gE8u7+LRABg5z5dEdtFQ7ddOfUA6sDiF2eE8J/0RAbnV2C
c0AE+0JT7WkwxWqV8V+LSkkYKOW7gyGvcEpi4A/Ubbwbw0gz0qRtA/DLbsgRLiJDlbkLbUlI7kZT
C5Bs89W0LRWPH3+GgWinLl14jmgVAmilxk1C/+iXdrqQSKyhTshVLkaLXBbKKgRv6k4qcb19WHEo
v6P4dajA3No4VrPta3mOfFDQAzgh/WxhfQ12bAiXcuae2447PwGBScntHDyeQtjXHWIYfONE0X1d
DKfgn7hOak+oJjKOG3PqRwsZ1Y8ya6/HFkd98B/4qtMYi9T72AZ/24L1AlIkqPLxofJTvFytscHm
W0ofxiP/1AuYTOh/U8vOCrVaj5OpawhjbZu0W07gbCpp+GfeUUcReuFba3xBL0VSEWFqYAzWn4E/
qc17uv5WwexsmFtlFd+Z7xIu27iy/AtR9o4CGlK+g2Rby90vvVdfwSq8DFxpFVJPATkhfxq197fQ
24iu3ob2FnM2yzek3TENV4ECUYvxPWq5pKN/pgKRUBA3E7PuZVfjAIbF+YSZ0KxMrW8QDMaA0bvo
LRkLfD7AAN+cY6oje2frzNRg75C8FZBz+TvDiJchJg40kt59rCcXM25ZMNaSVRqVCCvI4HIEsfYJ
oAL4roKFVpuA0CDTLkgwDbzTLK4VtUfwRFh9vQ2HZghOMuBF//DwQtUYKsu79wUszIEL3HBWILog
j2kHqLfWw0Nub+yR7xM5ZTCIzcH1/om7+Da6Fxc9Xm5Sm+dhN2wH1bVNh/FnhEnojCzbZYOUzt7H
UX1l0Oa6SVtfOQmaIwUapXys77MP3pFfk78SLF/eqemM0hWUTNQlx9d0oHuOzDw/SjtAL+H/7I21
EvuV9zd5W5jwROs+hAWPA8APSL8fUGI/5w1e0nTkpc/VgWXxH89wFSMSVLRljYLSgn7IkUtHz7q1
4Gn/CtbIdlqvsmb/N7v9DlDNxyiPzS0sO/AHIJlvUJXa/ny5tTXTE/Szfs4XOKPNUvUqIKc6dfFK
UsoG0XJLKGb+tzehd0PWWoGuegqTh8sgSyQThOzJE8/UNdKuTHOro95w25CVdLmrQasM7iuNCpzL
fDpxz1UVFe1bvv4xrPJY/23uJPelz19i+FFqIQ3yJ8G+9+t0Yn2DCSJ2l2QLZtwCgGCFH3qiCMQz
X1oeJfVWS3UnfNzAZHaR6iM8uV/nJes0Z1EzaWNeDtYXKEowf0BZBuRPL2wuLEIzyb8kfgebO4yA
rTxXZtIMk3B2oQMMjOGv0pmbGjBZ6xw04V4Ee2eCnGwsv38KXlEuU7Su31/yxQ9bSvPp93R/HLpA
4l42kPaGMOaZgLizJOQwaNJXyFiV6DKDp0iT0CNJqyadgll1Sm9JOZQbNuFEzAwtjIq067MmPkYK
3zSyugVoKDI1xo7L0FbhdcaM2MSIxF5nRBJzxT/dyfQtkM5yEMgtmG98ZbQ0A6PjXEbdcMU0t1tI
G5y2+JtfElK1Jx5Tp0YHdc9ALg8iRFCEKOWCU/TMrGVmdzefEK66U3EemlGdkuH/QrITRYlO1182
opkNWTUKLNW8Iy6EReqMx5NFOg589B2ED4NxcstT78H29LfNr2MoTEL4SvD/UmOhsGQ+Uk+QDDGm
Xx/QT6TBS3Wxb3t5ljpEBh3cuH0XNBXjYup35KH3qaz0Vs4VJ22m8HO6PB5ReLJ+iuaYVqPfIXmi
vxx4Cf1l4bKXgYQ7pMP8phVX3x+qqauRhmwAFYsuSFmkp6vSLn+SaV/ZiFxCUKMv2BipylAw3Kag
2y5kTQkQ/pFnhH++D6r+ld1Pm1O4ZvwOxM0djN1iiQniImeuEliEZK1qfxpamXxRolcTha3+woQj
rOzA28myG+FCWRcTmq0us14R74q9CYV8B0hIgkN5lYObZr45LPexSBBjGVCyLcydYGV74xaq734n
Mk7NkwkhBjE8oyWDkwKSEa1h87WTED8ncDauCIcGQ0dR+DxoJjSqS6sxFbofFlWbiT3rJ566hRr5
yX+WaxLaZ1vmMTMTiWFE/mNg3J+U0bSdOGMqTPPizFSOUNSP5kVhZMUvas8rtUK6xrWQk4VxJSw8
oC4wqqQyB+i0wJJxA99/i+RwkWFiAAFcSb9qPuFTiA4o1mycQpl5PEMhZI/FxDwmspkGl4woptEK
U4k6XaKXuNRnIioHlLZLBsTLXD7NmBZk1/5WZPB4B4O25kyP/QzL46HmJktStURpr7sbyJxGcMNq
rTjg+1jlD/7HymZJltpWOmcFMXgk3osNqZbGNKOLgpDmSpy7qdnPsR+7BFzQCNHG7ZZAdBNhsM5z
2tv+Ict5GbeAKyHUcvHDFXPIx+WtDFY5KT+T78i4BVl67U1vaC/FmsYB7B9l53V43OPuq4Zv5A+X
mcjNPpykr9wVAJ0MgSHo/IUmQ3+P1kmuF8n+tp1+LPm/7pqoWLqKqwTYJZTEahjgnMO0a2794hXB
LfdSMCWe2gCsna4gvAZ/lcAnbJazbRHsS8/fTFh8v+lgHPjBTCFvsd2YEwkBBb0xZeHBRo2zKZHC
hUwAjvpmJpT3YhHKVRxuj3wa8OtSLySbeUkxR/1Y3MQji2xNFghhMR3Vbq61JbIaxD4bydrMWTnJ
JJz9nhFKx06P6Cmghj286NUEbTX2W95h1bTIDi6MszDN+/JjagRpXa77SrlQ4F6q8k+nsQbIQEvr
O/vmvB//qG5glrBWVHyH5qQOpOMqFkXmn2cyQQjSgyIlegszy0tiXXwgGJWjmrJLNEzkoWYStu2b
uvvX+mUHJM5JFsJIBjyZubPv8bti7ZAv+sXZfx52kWQ0TnU96GdITnckdVS89t+P5Gpkecam85gb
dEbDeHCC72SK2U/VoJA6Gzo2jAwc+0eu4/2HRpUeWHY9ZhjUB7CRGixetdBv8hBVH9DHW5+cRuc2
+lfpQOEKYG3QSEzFAwMmFYBdEOj06e0SUI6T00zdhXtXOsQc0B+l7jJcDXoCfILgIALOSB/wM/qV
CWZlccNqV8Yc8J54GI16Y/9RbpVj0Dj7QV4zLW3q58f6yoGQVY0sKQe/Ze5t1bj3vgRyg52n3SmK
HfZg2Sk1L9SkXY4Vm1KUqzzKRjpzzFpX5KIPy+Yb/mkeFygGesbUHJYt7PAIE2sbC+0u6YPNvBiX
SSQYWCg9nknjnPdodnrcWvmn1Ws5x30DEdJrbDxks2pEqTNv2q2Gd2MkdLkhQ4B3IU9HuBHEJwgL
AJ1a5V52+yvWNmFPghI9PXoqrCtEU3zPSNQqws4e+VMhG5f8a7VUFfC5N7+lwbLXTj1nf51eufI7
M8s83vR0JDkN7vYMGbn85/Woh80YoYsTfA1E9r85tO3HyzF9X09+QT1/NAg/cYHxxVAo55aMJobj
ProH2AnnnSzyS4TJ0P7mWgS9qgvFKU0WADjCYxNxbMa08NsHAW36160Rp+cuOmAXUItbYs4rFjGZ
wSLdksrFEsVQrDT5pdaJoxv5yrKac91FSOAwZH7uz25kPvAC+cQq+QbqqqWPKfk07xoq/08s9c2U
chlK4lRHTVCwICyu/X0Muc47hbKRoW1q6G4FyrkGT6XJy1izaMYXgz7AH9cqZlq3rzDeyk0YBb5S
xvtOoE+xTKn1RkQiIOIiCZ/E0cUrxzOac63Xk0xz6OUu4kbb5VRHD0au1fXS8OsMrvFFPx+A6eg/
AFJBGk/4hEy5jWDVOq9LaraoieAjsf1c9aQiLP67gHGVlt5VG3L0TrJ6sojzfruHY6is59gFTz0v
Kcy0NOlxuhiESBIFqxIDga7gv8ZHjPR+ZSNFCje+UGDvWxRYJBRdk3D6YitpQ9+O9xKPet5G9Uhj
j5f5RR8UfDgz5VdsABY4xgCqBzb5GkT9LFxTHhidoS8Txnh/al/BeWFw189oQ/ca83F/CBAe1z5l
FAd3ORo1YFUMTGdHxUM4yIJMea9TY8UZZexRJsmb+AVSUEhYEzSXIxsqW6SN0lecHhz72JoyDoV1
i5OBqowTZQY4bJUhmm95aj3HqveWPPddJ8cvjBV5/g5jR4t5I8CTWdfCe94t+cePxJHtdNv1HiMq
jYqNd8L6mCTI1ou9IY7TwIT4Q9RFnsdSjweMr9EuSAkpSpZek3ir0Ab4UqPT1VTpqkmceEVXrjN4
xjz7AomCcI5J7wTsZ23ii/Nzj6R17qBUr17QkHx+65J6FJdPZ0s0VT3NGzFY1eiqjVvRd2hXfs/Z
uC9sD9J61KzgDMS44FxTpi9mlSnv+11K6ddMD1Q2uEFlRlNlzS48Z+e174nTjiCyXBugEyvDzi71
NkQTP8LMwkdLJrsJctUcuE9lR1E6vNhWePwtTB6qtAGagbLnYy21fBUKtmL8Z4LzxAAXqt4mQyIz
ALbXxNRKXH6t/blLCfzclee2yjn2cYdEUkJUyW69JBgq6ZblNTYPlxv5KTGrAfNRsqZ5uoVbVlK2
ixwwXXuwywSKFNLcbqmbj2vIndqo+hB5TosPImDEaFbdLPTJI5M7pExL0x3RzNd0jKdBYXLWLS9d
DQTyBIMrl2Ex5ChfrRcIt1JrF0/UvsDUtmMTFGhF1Pqq2KGnQTgfbRtsrBgscQX+AgkinF1YSJfT
mwND7WvAOXdquchuDZYQKTUwiesWwNR1YbKtxpG1/rifBl0olikyhThFcIifpYFtxdhpqdHsurX2
NbMYtG2H6a5GRyPsJJ7zFH3EHeUfw5dMeCjbOSVnI2Nw7tt/ghmhXkGkDBMlYCMi7wbKELT2RC6q
mcLYt7aK/Fu5dM1fpnNELYZ/M/2Aw/BtRNxzpvJRTo7QkrSos9pZW8c2JljegyOGV5+rQ6Pv5gCj
HOeKA5DmlqQxKqHyrV6AoYWM7TRJoMtgLa8z6onfyu26/loxc4HQ6vq5+ge+R2Tz3TIqJVNKEfF+
It1U1tDbj57stJI8Lk3lLlANZhqOksSMmvNc97nU/9XDD1xwNw9Q0qkSOecEogZPCOtizVTGyJ6V
q7lRKM5dmkzSZqQuH2w3Az9CN6dXybRr3QGWwbBTQodNep7/4MqyV0jhOCd7G6LIclBa4MBxJE+s
+QrC0WqCGUG/lJjsVcKcIkk/eY/mOwP6+xb+xjEn3FRr6LSdPIM1lBmiugSguWqpb8emnqj5g6sg
xbUyuM3Tarzek8MxlUj1PT8u4jsxqqoqQJV4iQQr/uyMD61wWgy8bkJNPNNUy4I1O/xHVDjKLud7
RQ1rsHF2cy9AI8oudcDZhvVXQoIn49yl/Bzxini+C0cMJ3aOawgj68u66nK8jkemyftu7mjNqhvi
EUOUMYIwf2IJReBqQweGZlzOJVtckNmjQaTz+xtIqseAPrvo9QKoiw5a9/kPwtFUtJ+/AGEa1CfT
Wiyt4B3MdMR1lGRaJ83Y1noyH0/E7l/zZq84c/XpIb+Bulw1N0MZnNOkszw7ZKcr7VGoqmebISFG
RCT5lz0qCKIVZ62sxW/r3LT4qTwOUdpn2fCGtKBu26VTfxiRIyoAPTaxyd5iKnwLcpunhtjPpihc
5qFU4cZZlOeeEhK0AMkFItlnBtIIsR0Pznui/xceyMPETT6NYeBRgnYRFDML0uU09BIQX/HRDfkg
L4ySJJG3K6JA0k9hFQPAGIhjcrERI6hFrlUrYeiVZeshVpMBRPhQo+fO/LPz+eZIzSY3m5IqRrtZ
fI6l5lAnxLESoXC2Xoo62wV2ONn5s9B4Al1yBLDvbw5dgYCht5ScU8Cv6I0HbPduqnBWHlXkwh8i
cb6JZTDi92MWPjjVriGk9OFGcLoM8WH/XZfVZ/4vyq2Uz6QQHnVXUTLwFYvHxYitzVMD3PfsJv3E
QPge7VxRRxCPRhBTKa48xMi/llyYZdJDwB42GHJqby69/Ws87NgFa5ei3rbVczvhfftcOX6UUn+E
xUU8bL9BloZwr1sm905rHiX7/8qpaGm1GuXGVTQlfSTqB2oIR1gSm+XGRxOpx+iRAKWX+o7qgOTw
ZSgS1QihwBWy63ZRbmqHTyDtqAn8hxmPxXyjRdjyZ1rH7zosSGpml7oWCoQq+YNWtQoxAue2GKwc
bG7L60bbg9Jn0LtTHDL1fEvVlQBSDx0/g9Jovc9AR/FPvbJHJ3902i2h92JyGhU1zpjA5Acl9RO+
haJD+9qa8onLkCsjKZLvlooMPap4UgHnCVBVZNPrR3Wg4iQO+qremi3w1LImGp6ypMNyuafxRED6
ZhCxWubzoJoHlPa/XGxN9lh6Z0Z8dpuRybZZdLepAS4zzDkl3c2OYp5KhBorRROReLFT6iX7+fyz
WO2V4+rCHiqC0+LAs38Wrzy/jV2bT3dwMS5Oq9/ohDu473efJUIzRLkLL2xMD1cigHuj6JSfdO28
9bdoC6tcQNVAvr44JJ4bDV6oHl+OsctO09wIZclnElp0FLe9RuOqtGEgnx+Use2esNwiJkOf6Z5s
KlCs2ivFObTG0EsC8P3b6EWTqTtGG/N4Vc8S5wKlO8x6ioMsMo/TIhCC8ND1uG2U7NjDUdbeCFEm
TFkyQpY9FUy6107+TdsQtLpuYkdJF4PEWekgXSmG+2LGfufwp72Pwi9E7yfEr7qjCIZaeDoU9uYo
Td2BzyfR6EnrKBfKemJkqSVUSRPdu2UAO7S1oOt7npSVYc9+2itM8XhOFJOFHRnUoikAm6DHB3te
/jUXhmtsOnlCeBcPZoOJJHNZlmZKaUeKRN677UGrAKjlXYzB3my+bvybk7uPt44ty+zi5EAcSr2H
5zNj6ZT8SB3IHfZznUuYttEdVH91jCAGQnOcn+l/QJkU9YPrWyEfMV1Fpg+tQeXXgeE11Zs15KWw
8fpTve5qFXrqHec65u7O/8cwWkrja0KgEge+54EZiH90bkPaaMoMIoySIF0Iu/xRdI2cwHsIz9TN
ffyJQl7nFlPEaxYyUjQujMIWhpRp4tpCUoKKw3+ctWY+cQPEPs2+tJ2q/Q43WOYeXD6r3eiQGk/k
Q0yErqshMYEMI7GuyChO446W/90Xg8RIoOXaVuBtAwRo8KjHj4vq9I7SLC14Q6O0au482f4jQdSm
r0JAQ2dUka9pKQ4AzhbylETo1TI1XP8T5otDMPtszM79wuiFTsCCqov73jgUUT6yobz4aEJCRMN+
g2OxCVlEtgLI0xjO9d67aJK4+F9nSlH0+7g7OLILJ1X92AOQQ0DY56ADtXX7vg8Ick8oUDViqfsL
Z9oanFWo6323J+qeMc4cMymHOUk/C+Tcojhf48mtN/xrjR+kGPT4mPZu/osHCjA5auJvDrzoISTs
x6ztxP2ClbylurEhl+NLoOWP3JeKGqpUpt4EdiGfXIMkIWWnxfCDAwhbS9mYYVNkI2FUzYBuF2oG
DJQ34nvQ9JRUCD0jPMBoK9fdn0U3gz0ymDK6TsgF35+eFMh9tcmlOh8KSpPabl3g5xVK6DThHOS/
bS4izK8Cms34HPtXndE587X5aT9dnFwROoBNVNa/la1dMWrPJIwFy5+RtczuRtIVSLWkJaT3MLP1
lR+2f6tMVRmG5jsiS4W0gicN0lxlxbdxnJUROcyFbN8hAg5aLOpMg1zh2q5zBvQmTuf1QGBUjuAI
mmt2FKNKRQgqceno59NpEAUCd3AEYwUhy1dwaIDcc/97zRJNf1GpJNFnU5NumDOxsgZCf1YnYKOh
XkjxXp0J1XddDKDI3thTnoRMu78UmBi8Wyi2a7sLO+mDp7XzbrabnLlVuB7UcX7LBghfuvDbeItd
ONDf3yrgtjnkCYNuNqXi8xgmuJTwVnM28tp3leSz6yDuX9wbLFIwu/xTGSmxqPdJElxaHL1VHnEa
RTeyJnhdCN8W8nzbJLkh5m05SRIHfkwj7IyH4eBaF1Wm4rHsNlCM9jLibZsmb8lqCxWMVUiv8c/l
wGacAaJwOkkXGBCjl/ZvSDqlJPKF8Afn+35JaMfhQ1l1T8HEiEcxRSiox/YvOKGfGwXrA6u1Hi1y
czhzf4TclWdlrXso8MOSl0smd/5Vf8SBpSPzu5ww1VgNRz1r6JQyl+hUa4KaKou6nfA94LGu2jgF
wL0crxEtJu61vnAe2jMcGxqkVTD6rlHlBeBoqrmk6iOFZ58vMK2A7lRsEYFDvPvIbpe0U28NiyoP
IRIk+5eeunAwP/H2SY9QIDpfNDjYhRMtn/vRubP3FNHTr6ydLZ2EjZMYcZiVgOzCgZxGYkPNmTbQ
lmjsFL6CLA6oI0t7TzCmBpcPIR/bgf/YPxFlep/XioewKEc1QJhF85lS1yuujkz6pXF1OLmOdoNt
SHnPfuJi9N9OMJR4B66VLhFKEpAwP9em1nSjWngu2FhO/PnT+TlySMdJGjmg2OcBbw6clHJt7Mot
Mtq6KMmO/SyrhmwRK0y6MuFXfPl15y+eGFUhVs5ZZuUMt5fSRi1N7l7gHFslikup55GKTEGFz0u7
+Vk4YWup2YZPb9YV6z8W4uHpxmMEk5WbQWOwcyUSqVP/p8jWluKbOEegmW1cZKR1h9scS4A7E7uC
bmCTX8rnezKNzv1D+8ogUJnE9Clne0+P4CeKGv3HQSIUcmKMzyJztl7vFsHI6GEbFJCKpQUVHNJG
CjLptkZewLE2fk6cy3nYANniTQ+bN2zbworHhk5Cv+l+i+lOAXTNErTtJGl8xJxWRomTDl5oKUlS
mV4KFzWnUhSErgDwA9QCdzBYT48YrflHJsvuLMKvIfMeN+IRE9UYssq8kfhmfMuJ9taWCCO05dAN
pgufrv8AUCnYLM+oKgrJH3/NMuBA58EE1w+NSln2IeY5GPL1JmW6xd5WQT5fEhqRuFdpD0/I1POT
iUr+XDci3fHjQBcajmaZd8nM3YvctmV3q93tJNr/4bBHYINnYMEc29Qn2RkCfFg8m9HvNQvnBDE6
+4bF9Z/uXDpDPy5I9v/DqBGN/QdwJJ1eXYaLKzls1vYFjP4dh0bZ2ZaDkabFgwcqigKdIldx03Ep
srEznUtHFeu73aduKEsYqThjHmus5iTeG4RQr7gpfvWQ7AriP3mTFbVMP2W6iRsUKnyyTq14RWB9
ujRCSiA8+1yLsWZjPQliHVP6BEEKtHd+TB/JJsUd/F+VFi552UnogIV2A6/ZO/z8nWmTNF9uITdQ
37J7d3HCh6uSZzvDh9WptWdj09POTd/7PxVSVmt2fDxZOU0ce8OwUpGGroDPUifkXvbpk2izKGcK
YxywD5P7VLue0hAyzo8R0iGaf3U4AMSJp0HSY8j1ANVXcu3VwQl6SqCQgBiG5cIdF6hTAlcqua5g
YU166tDUl5fYeFXyJRhBb72STvLE8RoBM51riZwSJqVF74R6IZNejCRmfEO4hcQOLvrnJzlCQzJv
A7I1VwV3EqCpkYpO4uru7C5yJrJPxXLEQsEFwUxvsjSmg1OnAiPHMmE5tpg1gFMfO0wN5wUmRtsE
tOl3Pj19mEN1sB2EKNyC7JPej/YSHIHYspb94v5ku87nD2fVWecL2B5q1kJA32xyRmJoOhN+ILfT
uP28uOD8xvW1+m82Nw64ez8nF9CaDh4CWwQEExVjNRF4o/gQ8Bl0OWaaoXd6cEs/jWm6uZR5IgHG
HZDtK+Ht2CtJ5HkQPYru7446oYNyu1ngw+qQmC0PSLTpQSe5McEWHhYSqGtAJuXIpGH8qimg2kDK
V3H+QKF5dGNYQjrz1Kd8ewDYjkBS3fFhTkmMx8sOKceo1Z4S38Whio+wIs3UYyfUUaN+KLI3MjgW
S+LWgDBzyvTPteE9UXEh5rLRQRWuEqV3KInPvUPhR7fy4wardF9ogm1yzC0FQdrp87VJFwTwECIi
qk8wMs002AXu9sH5VDgbtJQwodBySyP3BSXLccFzQxagL1smmLf4NPP7WbVRZei76ORSY0CYdPeo
ZUdh4YEzDFL5phxOhUmad0cwMeZdReqMdl+EK5SJooSs2WfCKiC/4J1O02Rh6GfLKjhzUy9GJ4kx
JkFVX6CJppc1w91PTxrpFouy7wm95Ms4W7Gs+WZI+QRFDV01hO8tDioATKuuc+VXIR9jUCFhkLB1
rZ60LIyhzESrGCIYVpgaZMy8KwuB3eCggj3A5qB3tUOAV0VeAKnXOvn3b8QbkJydedQ35pH9mOed
rlyX9DA3FmbGKv9V3SHjOjvIOKvm20KyPr02sxW2DK89VnnyAHaeUO5NbmvQSHxsGli2Y3GBvZsW
X6gTjTEzlYWIhgcgxCF2IvWR2MaUsFeP0LZxC0s9AXQ/B/7TUXXVmj7zkoZB2raXNrF3QwmQI/RH
Nc5LSYLfxsvHh43glK+rHTOf5hpp0ZMY8djDA9nxZ10bckn6rq2X6sR7cy6Qwz4MmFWPiesTe4hm
81yFKdxLeLpzZ2yHdD3tuYwNAFmeMT0GEwDDVUAGMXjBBWhnLwo/SVxjcgtfcRifWMXlbHvMKK2X
ZW0Oig1WAinnfEV9XydgSxm5IYZ388KSMEwVohbx19t29tUJe3vEpmjX24UI73I5i8OnxM1Aqw4m
eMxr/uMngBo+UtBZEXQFM581MbAHE3A/gPlyl0VIADa43cD0gXRCcQKrxLjqglvtxhEyO20JvbgF
JPMocbkri32I7QY5WfFx3albK27OoqSiZkjsSywXdzpuxfJFNyEVihioAT8yURYnW1qPOdPJOGT6
0ADP8gXynRlyTU6vfEDuDv9YC4oQ0B42Hu/wC0bRmy+B2NG6lAlO24uT7M4cKuMCQVJOZIpIfuiv
+sN0ng7EQwk+mJy42jcIXJX4DmkIawbwdjxepAIPAjMyWqMygH7BnBJ+Fe9Z4/qHqoy/0EPQBU2X
1i8nFoTQi3ppv7PKsV5EQN4OR236fgCEX2KA1GfXWzquWMxFWq2xSO4sg+3rWqxjkkpzZRoyad2b
ID2Vyu8NC2i8MdPpfF7yUVeHEXDgSlpWfmv12WF9HOnOzdX5XD0LB2jm+UN7JwpydUFtOv2QA3em
8EHrityD0Tqro7ynHYENJdZNqMq9NVpuo2rJxNZFyE2TwkUexTui2TP7vWS2Ha36DDCVTpNwRFy/
uAD4v0p/Lr+KI5wDSrBFy9UNQIZE8guOWqlfnt2nNN8LAJF46QzNMfTOGv/D1ljIw6Q9sEVZ29Sc
krG1Ghd0r5aRX/TQDGgKO3tF5nF+1aA+ApbyaAqQJJ9sXElM5HdaqnFVS5GRCv8t+U6FYRBA0b9A
hEZDXL9zOFxcDOzAQAWYsFSY3x2kpXYSc9mYDYfERo7zZJkJOqX293ePzqWCXzaRflxQuf7A3eu/
ekcikweevVd6mBgnfggdwDpj5/K54VKReQFhyTXdKau+yKLPOkK3uX7/rObY5UzS6cKtWq8wY6sa
GsUiOc5rVvjNXJggzjPtGkYCz108XruHHQMArpG1RvO9QnHWRmK0aen+YxwHnZ6BkHJM2bDIzIRI
q+lBePXl7YIyD/Oay6cNPzii57FYa0l/KuqeFMNzhZGlcg1ZpqYx3FtpN71t/cQ50x6wr7l9jshs
C2/LProX2ttWde5DeDtrUeXCs3CmWIF0jBihOZKeWxqDkPLzsQXUx/H3d6PQ3Fx2lk6dGsxaWkb5
W/4KOuomE36Ja3RZbQKnXddkx+HZtVnSbqPoPQqUS7CaWA0uYuYTcOJFm5aM3N1d8gOSzJW9kPl/
6wbig4D8F4aREl74MX4JBlmg87Ub2kIXBslWFf5aWxCfBpewP0hRhxWUxONvzpDw4mTamaf33ZBL
37Wd2C+teVkIcAmiRjsV2DqmQUGfwDTnYz1bXW0V5SBBwpa1VT29mwJS/DCdrZpeOzGaEUxiwv2J
taD2CgpG92+wEMTgtOIDsEa3zxWqY63C5Zwh59nKTWxnj4eDrcrVrTi9WTmh1epwLDFhdWs74/V0
0rF2t+JZCheoqhzG3HZaTwKbTpIsAsNlszLxUw/878Z7CH//iFm3yaoSEDJC9sdKKtv04ghFuCnz
0mDW/+f5aBX/d9li7ukZ5ESSbHs3r1/Ji1uQnpfzOq0ZRzXZslDomV62UJwTcNMeeZlPPwdLrfmv
xHaVqtl2S1jABKxjJ5T1temN3l09PlYOVpS3PGP2NL9TuhHhhGQ8YUW8jgVKOCnYFRT+T07C9eFq
VDiDotRSCEcArMkrtJERbiz+7Ur9h7Nw5F+ozB5OYQGJ+mG+aCtZI+9AIc+9Es9SoIdPj871KWus
cgvKxQBXt4Bo4QjaHidjTKJB/8TLl/vGRQhwg/yeYyrhrcb7/jJHqMBkfnTkVwQcqU7SA1yQsSCS
rdQM/8gStFqbjDqjlMUWUH6Y6/QQC9IQK8TDBsN+alnVyALrlm15dCc8vJfl1IIBkgA0Y+a2DGZw
t0+O+933nKnjDjTO99kQwl9KcIlo7hhTR05XTHNn7lAuaKgHnuq/SO7r5R/OzEJayIxHGp4tU8lf
lhcWzRp0LHNIey1ZiRzGvPlPV8vnc0aTNmXrlBzh5dlUcANATCYTNIEzsLjQOYDNASkOcK/6G8RP
W68Gr3226o4/BjNhu5gQoWPKu0voekG+YMzyXO1aLgmbNH/L046MHKR2Og+1V5tL4QxOCnvtkhPD
y0rBX0LivcTVX3MyHh4aL3nLr9HlYWzOykNgk4EVO8f2OLrwnJuiPfkpHESEONBKUjeqyQNiXd7Z
Dmpagf6KHpTmZytglZShvpa4EERibUhUp8WzAeK6bp5yMkB4+T5ZPXrplBLxt8wYZaPXXz6Zp5jk
x+l77JSOqqwy7KD1LhjGaBqa1BuzYKVWmYPz57YT01u14H2A8yy3FJX3MYgM+7KMOiYBHpmzm2h0
9vj3x0rjLBkfZIZQwVEK+iwIcmX3DsbmSyxC1BjuVTu72fzuBZgM1fC2vNbtlCTl8gFUI/FyAx43
C7C4YidqCL14aIJsGUj/BqyYqbr+RQKrP5NidhaujV5/t1HaiJJna4BcbHO78rpVw4j0A45m1isH
7OUOmwahu+buOpbW03EmsjVwGE/L2NLHKFAPvVpXjcpgJ0FvG4ljh3rWVh5rf1z44fI8Mev7z5GV
8NXL9En9XptLftrWHtFY6Du2sHCSFcn44d7RFZK0fpLTPOrquCFVpY1z2Z5uAmlzdOFfDivd6hEE
uTa6MA6awhfdKZMhmqfHkNHQM/6KY8SWxbsAmE2I0WgiiO9ubZ4UXb2ZfjrKdkUNrKm4AeVUdPv1
jVt/2Qif9wi5xTWcbL2z3nYjW/6krPLrL/6MiWOdDMrTW92eTQv8xm5jjO7xlCGeYnXgnfn2DYYH
l3wuvRR+S1LESo+3h5TYiAYnt+/tfP4QAw0iChFLTKhMdbuE/skFoNkvOwQqAz98SCc3FQm4yyXZ
opjHNV9/OXNMXPpgfNFw+xfKPIhElSFzYcOTFzLzmjDslSQNibEYEnAwV78hGOzvxQGuWr3bm7E4
xRV1qInI1s8PIGd1RUI+vo28Q6TZpZ5WnzSPN7dSZsEh4O+yGDP1LY8lCptakKwqrz1D52ZwCz+7
qwmWq3x8E9moYX6PM/lyq+9oywtHQK6ujnOZydUS9O/eNsG/VtIbzSXFGJ8qMdta274n51b9RkSN
YT/NlxuoX1jnwnogWC4iqEP0AnKtkIzCoD2qowthaILkaQKtV7Ufz4+N9WesdQtS7Ah6jYstNOGr
Zo6ANrYrOEQV/7Jz/X8NRhaPQSGFZvjHywlyCKdRiv5KkkJlmGn+wUS1aEEkSCuZkNe1IrEeURjA
Of9sq/yYM/y9UlS5abDp9vF1LtaIcZMAbX4KtyOx1zFVozB3/pBrZOsDtmdMXRbRclLc+VRDh+6g
0GXwWRe7kpvI4wLcpfupzdm6NIK43gtkPtYOSP+j9xYtWluLNxi7+aZCzKblQBJTqkX2T5Is5MbG
7r8KVpZda1AuSmXENNkQDClv0IkSj7ev/Zz1RvjiYuzzFeCnpfcgRcqz6pW7hb889KsNw99Wk03l
dPWLLvNKvyZMT8CnRZzstwOwM+CnGH/ohDggxQPKnUBkBR65B5iBDARmQ3rQQkqYDfSTSWFQLWhd
Sv3apcqsM1mkldnlQrXeOs42pX017A4fdxndmNnEkofRiWqhL3q0sxn802FYnPuMYVh6pY12w+ZY
CBCp2JmjNVKs/cL+72nZdOvZQ3JgRtjoIDPLo5j766OZNe/x7q9CbyJPyDcMNM3n8WxREEw6YAC3
7v6+IqL28GTjjlWms5B+o9vifK9MRV3jWqmCkE0722yIsj/azi+JVkpdo/UETdoOQ9aJlVo2uia3
2JTzrJv/yjHBBfw9ysI1bp/wxrBDHXRUTnDN17SG4/ARlHqiXKRJtI9EtKM6TzBon9cOJ65QaVrk
TjuuX26JASk2tm1ybFQKIQZI3CegIbTcH4S/LqcOkIjZcwaF3R3CbM6gP2T5IkbmWuEhXvay8YJb
paa/LwJbAV0eGMT4K8ghPcV1t/IYB5Nlswo5ku0cgNkTky1KpJ4F44ShtF89yA7/YViSKUfdofV2
KWWw6WfYb1fG/HsiR31Jeubl/i3ABj0+jIFGQnywdaxU556Kggy2m927rk4xHyJfwY/Kzmhq+Cio
rZ20+LHQw0AAOE+oIUVmO59cKPSG+KLdq5itvAFHLVsDFz2DNdAvR3K/wPrLRzt+ZOugp4ATmj3C
ghDakY7m0NOcQCp1nbO9JTjPE3QX19Jaoo1BLkPmp9Vs+b1AQ37IZ3z/IpKz3V2p/WMPwFP2mYUr
THzcQsjN2bazRhTLGdTQ4Ku1jjtJUPVSKEyQQYA9koX+SNynA2/j8Ul1pY81B7wt44XsG18/JxSV
mNMP+84sP9XqYWlKsZMYm3v+liTX9PTPLNT+cwuRaiofIRURmVLCiKm5yh2ZxKee3JbO7kDCpqbu
mylD/o2/9Ma/r5ii/cev3iZHfLhTiP8iFXW57fZtWFa9SSvjPkQqVT5pFnBnCQi4n5KJDZ0a0vtP
anYyKPPtUCfMhtYktum1LCAZ+i9xho1803JRR/3kv+XtIvnfO/4/mXhK819vbdRr+cPyyvhamuXE
8CUIIVXIq29pb+LAY1VHCHAG1tLTfpy7iJhlzxjHEGzz7YkhGScNENd10abNKqgloZ/yfg9efc7s
OtbVdSzZhS5eGVIasNeSyLySo7RSx5RAb4BoYnFiBDL8xfjf/o692212hvIhvcxnb13jCFbc0tAX
7020EBFX7/NkvH2RTA9SUi+y8jBu32vHcNzyQ5yQNv6gY7bQnVd6c04/0xabPnragPxGCtl8BFFl
GW6uy8+M03EeEeTJTvVGPqm0VQNwGuRHag/twJQ+Y+Jx3/XdZE9i/RSV2RC84BjYoeOlADnRbRI4
ywAUczuZA8OpgNP9PfJtZbSRzh7yZuqDIX7OUFZ8GbDwFAJzDLJoPy8CmjIo7qH5fsmi4uPHDRD6
3rYdH+1YDnvSD0Claqcph0yWn8zBGe141nfNwMgX2ZGd2CeVSa/rf1+3H/d4UxM8zpZp6tbnQlX6
xn2iiHhWfySnUUIZcd2TAq3kD8k338zkZPxAzz4GDgqV0iSH55+zbX0AbG27MrG73hcDVV7oGCOt
Mo3n5HDKH68JgAS18pmyUzUKM76MkGy+cKNkGtnwmQgZX32iNLfQ8bCXWW0DBYTg4/1s8cMJNBm7
YBkNyAI8a+SX8yUaRRiXmZcd+gvxTrW4eARPY5IvftV5c6fVu0YIsGyzERhs8WhTxMQoebMIhdhA
cQ3k2WJuaVw1KKVzJ8IfmNe9c8PRFCs1Tz78fHDCmGzhf8Mobelh6YM8FjXa+E3H/dZtDG7E8Ju2
sUHXjTFvwguZojMM75zeSwB4fWsy1WkilqKxcxrp+SYF5cKK311p08vRYAX9nPpAVgFQx5EPf6Ow
PwtGAjzfJHMK1tmvRPWrPgaDsupnKqq/5SGLtrJc92iTiuG4ZR8bznQstyu/fp+2JkaoH57YRZWz
af41oWE9+/v3cm8nbeBF2Yrsp/UZUh8H+9/qJZ1OfV1007i8Y5p7AeWpmxdqLb9ITySrhRij8/YK
IIcshoqewC64t/n6FenTgD8y36pa41JHPBYn10RetoRLEmjHQjY/voOkA4MxwxjYPbLoldR1TueA
cITCznKJHSum9Cx8kvxD8W6FatlCny5WnqtgbgjytpkeiueGR35eGh8rn9FS1XGMMGp7nyPcaDqk
jWQ1nc2OM+3NtHG9xchSaxrQGeSWr1+gtQekUTuOA+609hegSItxLhuWjV5nztunLjUOkGuQi6cV
8Weh5Ob6j4jG0i7eCeQ32Azf2jAdtnKdliaUfmZiDQUMZddD1LIXs5OCZi4UgI++3K3HH35MNtK1
OxG0U04BRYZZXyqV2XNzqeSEN1H/Fn/z1mWxR1YqmzZzkTySIFL+mI393SAJNP3fq19U62ypUS5O
JnTl4JEy7gX7vJao3i1EnZ1qcYuYWnCZPAwEqCtw5+2QFM/d6ac3W5WwuCXqir0+iZKbg5xWPnKk
ibzz/gv7yYPR7AEp+b8CKxR7BnAbTQ7nhUmjuyfRsba/KJKmqAuqjyvOEGPpl5EazAugg0+d7DEw
X4Wb6hS0RPdC0YL5bkEanrvUp/BW2M68HaNPinG4mGRI/JJv2UqRR5SqF4SS+FmjXqoHsjOjSRJg
MEjYpA1pFwffxURTazdnY2Ns7Dzfzb9oZKUY5rsYZHOPaeHoJB1ZnobKxx6geXzD4aK6q+sKGVw1
UkC0fUqJ460J8CvzlElP5J8HzY4a+OKRsJazyMc5iSD4dL4Xw255h/sUJ+asO7PTYpB285jc9e+w
SVMV3UkZxCKMEPW1GN4EJAzYhtHiPfnqiHSet0EXNPOYKR4k/bOSJiwi9O3y2zl5xmplOJ3x0VZI
ZP9nFygN0F2U2Gp6BdsOT+1iVgXmq2cC5aTbvBrTAO6t1WmPDPOOzE/gX/XaQoloC2RYLx8mXpj3
PK4hHB0TZAqTqU3vpZ7Zixtdx7aFfyqFoCkZnuWr+c/8orvQPh9KGaMh3AS9GqzOMSUbrFr/OQAt
kNE9e3zrcvOUomUnSNswpiXFayUDBCwEpclR7mpi2UuX/pLWeBoPLFahedgaBasrsuaVDvP6ztN0
mv62A6BEfEfduBpzlB4cAOWxEaCAZIMYDjXQrjP3/eWGgeM/iFxfFTaZHyVxx/EJhvXweb3IyRda
H7BdxhNQzUS9BJyJeSUdeI8ep4RMAxp1YVp1+YmIGEkU/eWtkH9pTmdyiBbbDYCjI671+CIVUGX4
EuJzVrjSIGigAUiRUU9rvylAH5flPzx4Mgnw5Bkks6VOKWrrOmc/yDh2da9hFupl7T2cWX9kORrc
oU5blpJ2lqQAUnOID+TGNgveyCMJ81VewJUTvGtWaEUGU4QVWTVELFUOqcPmdxQEl3aMEJCm6ekK
aucv2ww9uhWoiQGsO2Y/l/OYFtSfbhK0KqbaHJw0DrYgWRSNsaI4/7Z3nqg2Gc+LT/AMLyJEp5nS
p7nLFAAwVuaG7Mis9WoP18WasmMGWmMkqoBTYzchGCu0payM/Lk43mMRV+8B0ItIR6AdCxSdJquX
bjHlf2Hb0+dncz3RqRCAct/7MFG53m8gfjrd0y9z7m13frIikUjeJuskw7sd7HOCyi+8sERQGGtJ
xMa2vPjpsaHRwDBKB6feP6T8cYPXitLKYL7Regdgyn5+ios36hW6WBhyF/tsqXkvWVxQyuk2dBja
7oUbZ0muqe36e9td82/dN80sK2Oj1LFXFnAXEATqMR4hWwwHM6zYID95OlmrcZdiKhCl7/xasDw6
PqU8DrsWIxNMlEAzlTV6YJMRZOs0gcKBmiJ5N6S9b0Zm3iLV6CP/TwapZ5BrQuI7JbWmaqneBnoK
eh1x/ioPA5e7x1Awk216siramCVSJ+zNVgTEvYrewBHUR+vJLF2sHoP9Ayv6/q/ItZN4xZrxp43i
1HX337waPgcKWmcSJ6nODi5aXp4q2vNF3UKNRQq11UWMAQoYxurkaScjTejSct0SJ2UyRZ1gEBwx
ufaxZ9AnYwEQg90Q8f3y+zgbXLSUAevEZQmZ12i4UvJ1OYY6RLLEBg+CXjgUfjjNXpoK4HKpvMnV
y8VYceJ70qm6/V+oM26e6lgJdKCWs7nleMKdBMC3YSe2pVp8/7ze0jmc39SlvVlQf36YBxKh62cY
9Pqlla3dZeIqwytsNOI439++cIvTpJ41lPkcYKrrtBu1dbJUd92d+HHVPHsvN59gpv2NnHOCMm8G
zlwEGzyXXTYbck6ea3eeSX5qSIHGUAhe3Jyd0KwdV+Zy7+6wVQCGgfaxfSaGY4ecFO09ufgW1F4a
X+OyN5nbiUSyQGAuMm1btQYAkNSQrGOKs2pJvXw9affAcOGEktXelEi0uEMIH2cpxFawSCDODYoV
lZ4wMmJWcz+AXtnetWC9I8kB+8W7gGB3K4TRTkzoK7Fg167fI4AP6QYDSyYXioJrT05y2iwfxQmK
tCgzP4La7+kfZjEz5KtOEfI/AjfZstpbShQ2KItWoV8d7awa/6kdy19dcbl+Ls+CmWTdq90ZQyUe
nvvxRv3xI6w6V+4QHMPW6A7YJL7wfCpNdip/5/Ath13IeHWNtkfJSDjqFISYHcs5yIuUS7R5ohpN
fYtEZb8OJyBFhKqEYYqyi4RlwuRujkbCiwymxnqTytvGs9P0x7V4aU/MLVOF7vm+jrF6/50fdw8Y
UII1j1kS/kpFT8joQLghrKyB+Z79lpWnfyTMChI2Oe7Q4jkeXq079eXF8wIsYpIb/BKqVjmFtxZN
u5fi5WsuSyhCHn/2boFjLa/zSD4SiSgMh2fFacw6BibPIldR9YFOj2GPku7QU32i7+5flhKdahJG
GvGcVJ2Y3BSZeEdPxjE9auhwis8Cr258ZA97ekXnuu4EVm9eyFwcxpH29PcGQ+hZzXD9xQDzYb6U
hjECqCO5YnvpNXpKuhsvgYSl/99DuEA+HaW2tOFevjLMNWnv1z1U5YZSnCXEfn5nLsNKS3aAGqH7
5WbG/IZ8C1eTAFVTyOCMsgseU7cKL1PMbwggWW0OWvbKWv4VseHewJ6yZ3LTna8LLvtz58raij/L
GdRXsnsrD9UaAvW4Ah6jhY2GjI8tk5StvqWivoFHfUvpNcqAKGzX44K0PMDRj2xniyzIGv6V5CTE
5i1qj/GZC78sjYcYA8GYys8ogq90TBMVbeg6WKgTmyFQTQ+5LzpTAuFRK6fTrF/1pN3nuBNDsGiA
TaoFofaS3RY3o9Iqsz3QX+qrXJyPM4xkLH8u4MGW01M6xLNqu6rqhghJ+2H1/yvmfxDp0puSSdyT
ytW4DhS1CUGKIeqDYpGInBesLl67qAHn6Xe4Cfi6yV0zwTJ+EeBj8xY7Z77gn+RJ+i6QVh/pLNxM
MBGTcBSR883Eora0es8FjfqvAq0ATQxf7FRDKjk9g/45Oe3yL03dzVJRQIzBh1gBI/W1pxo9XyYI
DSig79QEiJx/IrNa7OtclBn+hdvMgjR4gOnFdAmvBSknysUF0IUb7UYGS/th3Rb6qiSJQeVfo3lM
UzT45C7+88ZMbAdE+4oYDQTmjTqAAsI3ENuW24/sz88sfkalFrIaS/Q/ZPoW0SPdjvon15f/9DhU
NdJ7tgpddTJDU6in5dMZrmmgC9/0Yd2HEGPBYsKtC+DbAyN8CY9Wn9UX8j2naX8Hv1+GqmOBEYq9
tBc11KlsOxXGklhbd5niB2Jq4fQeKz7+8BTr+OsTqfR/Ngcz7g3bnN7S92qyFs5zOxMzyF2y53Jb
QZd1stD2PTGayI0ZB6gW5TE8OzfAupKPLkrgrmpm1CK+4cEjlok8R9Bi2KZ3z2c33xaVCr8Gzy/B
oNlaZHMqO+cQnLEXGHdcfLP4Hf9YS8PBUUOc/2VOCBP7qjcPK/3dRlClS52LoNorxQgY2WMmvrsy
2H8q/iO0a7tHCfDhZg5aibZXf2qU/2lG9T1SVrmV0aYZCIdn/fhGGlKStrXvWeomAANKSU7O6i8C
91WQxsKiAcpWkDBh8ZuV2Y6rKkvkZQhfsIpdeh0qxLIL7FqaRJvk8L8Kb/a64Ycki7FXateT6vNy
9J3rJGa5YMARTJsPIfojzV/tUjW/xFcN8DS6Sm3xMsyIu3L0VtpLC1NSLqxhZ1iv/eC0C8h3aKzn
8vZgTfD1vgmNwKzS+OpWQtITYO4zMsgv6x/TbuMj3mzoidkTeFFtmb85yGEiWIjdekJZsLEYW9S9
GclEKXHzybfg4ricBwb5AiPnjWy0gF5EPgXVDNodZsrj3Xn0awn5s7vIg7sjQypodBRsKwYogHS1
Ce2i/y+z23kJplPpQUUZ642qHJQRuU06Xf/FYHc11thmCnmTmRTEsb6q1ngXC89T+QCsk2g1siRI
m5RjGrM2zn6SzmWuxD8TqXktJNOTyNVeNIXONLzlNYmzM70g5BV5Ro94EgrwXPPE8bcO93JAcweB
9es69LKOUSyz8gHFkPfRrV6ORwfu4OUmoAna1MVCf5Xva0gUzVc0O5+IX9wKHil0juEqVkSiYtm2
YRBLdA/Yumh3/LB+oNjwgu4cxd/s6/Qnt3wcIuytUYuKmMmw02SY6cAbs6k/apGkNHbeJjQqoM3b
4lbcWCUV0YCb8UDpxhzrlsbtJM+ci26QunJLz0JomN/FYz9bcwopeD+TyClFjcojqjTv0Q2RSot8
kk3HNEv6H/OJiIkBj6DFdnlW8+1FMNZc1TArTKSsyOZFwawu+fzEJy+maOF1SPKa2Q3iOrWgtno4
5jX6002YVEvEZrQFnt0f3PHUQssT49x9E9PAZa9CRaHexAjs2p7WIyyzzbfBoHLseXAghe4eLnnz
nE0RfrJFR6E9z629dO16Ie/RDz9Hzg6KuVPy2Lc+5FeDI+LWnMiVb14IKIjFrcXsYP4aEhuVkR8F
y44ZZ/tnGHueE2MB/Y4IybU+aX0KgWqy5uAp5R84uw6iSbujHxAYUj6j+xtjGUivJDRhAEdmDsQf
LqH3nN+4HHAcqL9aFnKKdkvh1rZG4LBlzjANvPIRY0hmXhnx8GxV9yaUrRgAQj3aV+Y5O2AcE4zg
AFW9gB2HoNMQHZRtL1RaEDemnNpq73K5qPEQ8utXw5gqMm5wta7E/MmCi/O2yNtMO6SSyzNNivFt
giIV/YZkQNJn/cPLmIWEGGPR3w9R9GtoEkFmFD+ULar1ZnUvQyz9fCM4KmQvRxL2PUVR/EKqyQ1n
UDCNvRP+cp8hxY3j0qpFPtydYUOBfcWzAl5QirMkDZoRBiO1Y3SkubhAMsnBr1VX2cV4LfuBMzU3
/Mt9I3I8QR+9GivJmIE7wbMQdL+L2cKxp2gs2KNEvaSfiOITs9kohqwZNR6OGed38gFGFLZcPEoS
SBYXk5XU4CREapSKuMaXB/DEppRDkFn05IM+d2jNF5J4/dL2SnUQ4kZt9tMPSJoSxskzxMp7Qod2
DUd2n458q/ZTG7ozFSwVwn1ZEbG5Va/Ryv+jiypu6ewhj55GoWxY2ngbZnzTM7Lf3Nw0KoAzSscg
UfyEU2sgtFStUripcPJXZsZVMRk3VGJqZl9cFTYGNTuaSbUmGi6W0F8asUfeiUHcU4cZiTi+xeL+
leSVUSBn9B3EanMI8TFSSJK2DFKhBIBgd38E4Kbrbo8BKiiFd+MuKlGsyztPmy/yAftpcDhJAIAV
Q+7L7nPpxd+5kccgELMPJWftBLZcjBk4AUMNDIMX/fQlz4Vpp0uhXkXtRavSi+JnUP37xuyDxzTs
ApaCWs5TrSkHpcIBu2FSit/UD7kThM/fJzjIGtjGmRK5Q6dPW0WaumOmGP6cSF2Iv6r/QDKTNgns
xzS5qlHQHtF8TpnYUXtBNU7ercoeo1h5Ula0bc8fq2AiYxwN6rDA4tsHpHk6oavqQae9PrKacg+/
ZdOSvxmXi0ly3iqrplOAJJPQVguURgN8b5aCb+qYzcdC/74IwEGEbaHsHHkabSWK8PhEW/2jsteI
n1hKFIrhbeZ5gIykpPcT134UxY84dVVLPZyxZ9ziow+UsQZr/M3CQMq3QLuCZSWwjZqNV9dR5Sir
47WfzYZpqKJbVAla4kyyfPKsgmsl8S/icArUYplPj/r4Y9OOsWbnLWPmnGjWmyzXi2Gnb2d9b6y7
tfLtgYVSGNexKu51bVMvFnS3TjITckvBuQ3W/umbOpYfGjWJnifVrPTC886eepBve8tcQjIv6PFl
lTb82M8bdeNE1szbIGAuNWGMG6UH8JXWy+TSklia1UEjWnWPbqD8+Pr8FfPosvngtBP3QulnyQU0
SFUN1CAD8SzjBIwrvBjcoOsFQAg3XkOpvGeAj9B54EP/ibpmxKjUbB+LVjqg5i+q7iena5h9VOrF
K4XX7KCapoYpQfZSMOsLJBK/8xi4JcJDLB0X6/kFGLrMAbV/XU0skQZE2ToZsVUl0rd94Hk/QDEw
+iKS8AD+z45L8E8X/kTOvKA6trl/yyy81vgisA7oi6zN+7VE613MeddsAAl9soJQgWWUvUPB01mp
rEmaWtv8S700Lv+Q/wqkHeYm03qtlAjdp/U4zRBurDgYX3dVnPGRRZhh5tFsjjjkJ6rEkwKmqw2N
deMYLxjhnoHnuWslvrq9k5oOyNtFFZGij/k5/NJc7DimLTVqB+a4/jw/mtbp3BI7nduMaGCZgwKN
tMIzMU3etEyN0Yi1DzMG7v0pjqsDI5WtSkqwxQwulp+SuEhFpKyRE4Y302xc7qcH6oFSCpULJ1sl
I2KlmXZJkxyHHNNwKxgSbyO0zMAS4QyqC2G4ITpbZCwM0z3w+jsfL9FaRr+0nN49NusuLlvucI5G
Whw/nwj71RGlLw5CgPDfVdM0+nz/bFHfO9gCorYxHDy7z9alQ+NuoXqRWnOTJdDSxuGjRdInNnu6
DWDxtX7Lo1ilkCngxasUYDiE/KK+Ds/O0R0o26kMWi57+usVdcAaPZEhsZG36/proLQ3jNc1WF/B
JN9NuiITAK4bIlnOnCX9vYiee0EFk6CWrBB7mSgk9uygLNptu4zXkNCtX5hbdVwHPkmN184lolSR
VnoXhITPsXoCXGpYa/bQAA0l0WPJ2/9iN8pjgeOvNo/9ztNnb2/scB1etTk3hQmr6ktNj7Kp/r8G
zn2nxYbUpc0UYMDR/tODkZnxW0pOVZrlJ+XUOTVRSeWX/sjGEUq65g0pAKnG6tOz2lnDec7Gew9Y
IT+qUrrLBo4e2JUf2K7m5AixbDVCU1VijW9QbVg50Xm4gG6VsUygj0RYeJnUiZMJiQzKDjB53EGa
3rfDbzdNXEh5VTw3hmdYLTAk+uQpwx8SS3qou58HtZo4uuC4Zs+Z3SZThWkGwqOpT+ol2IWxVfjS
CmzVGbS34ojMl1bnP+S+O7iFZ9W2xlDhTVVdHkd50dJdfP//X7Il0AoAaDJbR7V16xYURw52Xjpq
HX1IqloaXhm3tp4Br6bOdxGblzdlkVTSJen/xEAr1wVoFm58CRFGRvOQsfe17yr1RoX5s939Usx0
NKvvVY+XqOCQMUiJU9GJND7JAiyh9svaFlUDco+G2gLHo4vu8bRIbI6N0HDXmqA94hfuFxNKpO3j
7u1BLaK51+yndl/Kjd9F5ZWbRQrmGg260RqYRZcueXZZbG+pCsfJlyURlmyIfkxV9Q5Absk34gBS
MGfhTVydWHGR7WYQRvG3q1UPQ9IIldmNsLnhZ96Y8WkDmTF6lI9oE1B6maUCJ8TS3DVXFY4bIUMb
lqksWlf+WQQoW7Uj9Z1kiAXc3OjhaVOMsAucNYvgDrC3iHJBPSnS4lU1gJPSaizT87zFweW1kKDG
Rko4MGJoVWR8oaIJ0Vx/GDW6egG4d6hJvacixdXhflMpkPJIDdkORwtqgI61Wi+UdFcBPZggSrvB
xjo5Dee3L+UKzsURCck4A254IPvVf7ltrlv7AkripwtX6g++z0iqMuIuGbmxpOS5NMJ0husgNwEZ
bK3l8EjrvMenvtNnYhxSoqqMIPJFk3z4jvbB8oqJZNlMx3yrYz8mAaJwNgEkzvmTS3kNJIhfXmgs
Xlsi4Ns0kw+NTZ3Y0CYOlwwt4M0ovK0UowpjSB7ise2rkk8DPid/iZxf0GGMRqHJHX/6LWH4iDb3
7gpDc6SRWp5jNmFlUl4vhRpz925j2ITfYQTOw+ysbg3KD13AkfLDs9aI11bmxVH+pLRKMoAo7io6
E3crX6X39CH402t2vue2ZDcglqynAdotMyCT+eZeQ52/bM64mbAxKXV3V1toR3Kfg5BbtJt1afe2
U4t0xeKaN9NA8+dSg0omZ5hhAlPOiMDZ5hhT9SIVZgr+1Vr4rrlJE/tCWETVSoUIXCzI2Mh29T/x
P2ozQni+hEtyDbii6vGcSY9Mvq9vns4jFfa08ykiJm7MSDiizLQU4y1uthLOdGajqZz6e2GeeU5u
jyqhOjGSW2wtuf+nlzyXqG2hr8cq3n+A7uwUCemmOAz0tRFMqTQtqYI514DxOKlEBUGvX+FxlBN0
8g2LJkfqdidCbQmBcYJitlskm27bdH7ScfgcI7eUgmgKlBtMusMr8WKQTMBS+OBO0xK+BSUPD+SL
EyfcEO0avOEN06nTGs0jpPjLzE50CSrLhqkJiT3l5ahvxBl3fpsarNqN1YQywFYSU+d5mBfb+1ly
6cu/xQ60LzxFu2gWy8mNDxnXh7kSD5fqvnAqRHhM058pIMOu5Thif2tJ1JNtMu5RTlsC/KgpQ20b
spxfqgJSMQU02cidgWrF+ucL1KPM1daPFMza27maDnby0MmfZAK63QYH6qCqk+KkX7FAXFbQocVa
yMMyw0wcr4BAyQXb2/m11rLbYbVKk3isvv6yfH09xST+dRxq/Y998+Gq7j+veq8pkCktHQNkT1VO
cQoLiuJSvbu3UPmpWGATBmf/65EEWkeBQuqLhZt8WwrbFO2IWhxpSMSW5u5MMlWFAun8z+hE70kT
fJ20mKTAektjepv83Jq9ZDdo5+DCkVhJaHxC6GQ1/LQGSA6nGkFuEf0JYDKOPN7FdmpgaDrpH1Ud
jCK5yOmcwwWZ6J6MF0rJHdVCQ/txAHtOGkrp+g4JmOP2VrYnLLN4hsoFLdk1z5nn03yT0/gFi3Ns
Ry0o8ynHbFmoaHTcrCKBKaDdOdvIvdsNln0M4nSnZ1qsBFFHAH2+5ZBcQTyAz5ed7tgaI3OlobEt
wEFfiFwdfNiJqP1vUseenV8/7sWL42XBz+5vBJElYdSGBmsnW/78fmDNBYXtTELsGKfhxupWfiUW
043r8B/L0FqeMvbhfxPlLETLW0agqoliypCtBWjD6umvF950cy3w8WMFeXsnVD8zSe9AQX1Cnr15
gOBtrjBS5uu7RrqsCTqtGbs4U7msCRxZ//VYEyXCpO0GDWwVub+FTRpGPluRi4uYSVEnXaHYaD0w
dYYFwUK8RiWl5T721wd/0fXaUeYUrcgvEda/cY2nCwPxY/2JNMcD4SOii+XohN3BEHoChYLXk80N
SD2VRym1V7Li5LyA5ElkBHRmyjM804UitiZUQOr26mZOWnF7NYrSR6v3APm/5zmQ7tu0JqZfTPyW
SStfBWPHUyNmo9LYf1JXNMAAu6Wxky4itHzBL5JCM7fsYavlbRv8zotSLmJ5cG5ygHjrva8R8ti3
NZ3hLeSyeihanx3x9R97ULDCmIAEokw4TgNRqeavoL9aHqSz1FWJvc6PPzWL2DbeHsWnEN/DUSKX
X2d51dAAuP0bAvsY2U1znsrMA68YZn7SJ3WIyiidwh7LfcrRh2F9Ym1wYuLQ+CUHcAlR44FBIxiK
BKQh3UUeI5e0vm5eR5qRxjT68gc7KGa7AuFlujFr/jsjo+OC+lJwo8egfpO+fXmOQvnudgcSKIGu
07Q1o79MoKk/wSh4vloxPTdgkjWkD63SbwsUHP145555b8ZS8GAKb/BG6jtwSU3gCzr3bfOFAVD7
vVvOoFKpBj22VUfUz2hC5oNVq3tT78t3nDKYr3aieQYFIynBGmZ9TtXWYHdpPnlLXCvxO3/4MHNQ
q3xiSncubdiKowwnF9hqUFSy2XQHN+tG1zsd9EfJgHQ6lLBMPHlX3ueges+OyB2ZgP32YP0/6/2b
7WkJno+EjJNawnqPVH262xN+VNYs6TC0z1IzD8hN5DSchtere9hAnPlqP1zcW6elKGUebWeTKdR6
tKT0fLSfun/YbPwzub3d3dK08eMSmjZTN/5UzuNuNz3dxKBHiJMAE5k+OcqsHqn6KeRnLEMJEaBF
jjBEUW2ZNMpj00SsW9CW+ajxzBAAjFI8MGMlaiyARBm28XacejTYonZdTgNgmrZc11FCF0uYndGx
06wdj36HOXqSP5PIKj+CrDiFZSLHdzpQDvNE6tvapBkzNVI2rIVPMTq7q1G4dXzZC86qW6Z2pTIk
o+Q5XwjQJKsT1LyFU45Qlut2bK2Uo7xuvZz/1QohNstZ1sJUhsuXybn1Vg7Uw1omAoXDWiegHIns
MGCKg+9xYiabAIKgh0anM3Ipkc+erXEivIUieit0rbWtxnt9XUbywxVxgTs18mPucyJ4PGTen0GL
kzSqpkS0MtobmTSBwU5FeaxGlITuCOlmYHS1dcqM4gErmyOIb/vq1sPezqnCgaYde4Eq5XSelLz4
lcAVA/PiBhtGW00XfgJCC43qwlLHPKg1d2AL0GPAP3ESrJSSHz49OO2HH0GON7irEJL5F/8ZDp92
M7IcPtVTW9UCnrw5Vt1U3zyU3LR6WKnCEbvf9nxktyXkbmF8zuH9lgpw8BVzQYvTH1FAdiSGL6Nm
Mg9yew1PWaj7YoYQjv/LBdRkOghbTT1RDrTxNE93WRZfkov3SzVusQh9uYFCQHOSYceApWXgDiJs
9mV3h17pZsxWSIOXboqtZ2tLm8WOGI9d15XAQEWunwEBSUCu+Ymci380Ha6L+x10XXzClfdegvTk
qrVhQpGs1lXFlpwcw4DpmEjrQ8dPRbnwzDFGyJqWoql0Yhx2ZLzNh5Uuhw/HytI0cW8ASozxpVVx
TaQ05zpM21dbO2AdGqCaTZMP1FcXrSSN8n5yMeS2olR8XFxzjGiuOcFFhmzpUwmyQQAtIahPUqyP
+MiGw7CPwyRDyuPj7xUhR7IfiCvnlIDDGKJbMByAYqFoZccjWMIQu1a7M5pjNGSfTSVNDjQ47mZx
iJeW70oHcfduexGVYSDOuYHBKifoXUbgVBF3VgqCgacUDJv8wj2ZtBw4CJX1QiKLBeAnWb7BfwXo
AIRE3GQGnKIM/E5WlNrSaI/c/7oUNwVURNxhjaXentIjcDKLYIiWCjFDJG4Dnbx5/fbdb+uQu/dK
vpV9kWH7O/dNkOt0HSi2NmlPe9BMReJCtOocepMdfLOvIr/DSTkylJIKUl1nbpYmyrNRW27DaUpl
sn8BCcTxQ1KyYw22ABsjEIIjXVY3Xwcb6C7gpRehp89NKhjHtkXBwJMRwxs1UCX9I5rQ8y7t4Zlj
ks1MjGOLmtaJsUA9H5L+HeCEMqZUWofT7+Z9RRkmydytjsHFxBizuNMKmKBsjImkE6eb0hUgexNx
Vs1B1i3JH0b82xGWxT0bw7Ag+WGcpUz2ekO/tK9b6Oj9p1lxjg0HNrUQm63139uwxD2/bPLNDH4e
aldMoa0CFsusjF4cqKiNJYiCUTRAqwK4BRttw0w7uR+aynf4guATnHrSfVLTdKQ8dbI7776WyF0p
9WfpVqbJAGPLNr5+uR8ziXY+HNY4TNqUs/eFzw15bOB8x7PFSbe6ezm2e0wz3pzma9aZP4P18hpm
WfNJbpbsAOD6lmYwzrq6rFV4g5ClBz7U0NcR2CrVKSC4FwUuUBbXLbSRTEVzfhAIms0n0BAdvEQF
GA3AvrTs9S7e9CQDLEMq+io7zuS5zF1YVo/0tCBOohduj25LQCoyfndpyPc83fgis7XrCw8HqNe3
xNtyJjoq9cXb6XdTDbkRFhT5u0KOK/eeDCVWbIyU2coanYBFy1TgdL2HwPXIDCUsJVdSvLZi8EKr
TPE4Wo3XFDrT0LqLEb7glV9Zl0mpF6kdlsPm6SFRxtfYB87Ir7U7/PoqXTGNBQC9NeL4Q/9/P9nO
1I2/eBGgW7ixeZ1Z09dEU2R7z5JPvWbNfNHZ3XeWFu94/M9ZSpTU9MCZHHg2F1HHUIfpYMq0gWPU
3Mz0MMHdZCIhCcmD5CcmSImk0NGdXj3ZO/63H3QtZpxANqyNbXM3kWu/uwpiTsz5bdgrrvMibIZ2
sbdyOpykNDQYiJYirm6V/WyPNShG/TxA3kgufWJ17uClBPB9Yby4D8Sd3AJw7rr8Hvy6ffH4cgyH
W0ZBvNqD+v31rvQeAzq6qSkk1pQCm+k8IUig/oHKBoShITdRx4wSYmwLXKpYmPUETe3IHL0hl92F
vmjT14HcEivhjO3ivrquN/o2CjFEhmjfb0MYp1DzzNWq+An2uEUwzD58LHTUmitz8a+Rw9BX3Nqf
LSJd+0QQt1i3W/TpvE4JxEPZK7qDcndfslyTjheDn9B6gdgkL1N3olD0SwAtsQpo0ozMXJ/MDN4H
HiNOIojVQCDgM55wj2HRPUExkqmOoNIIbfUQ5f+FBn68AWmQ93MtNGKyeRRGbGH17+QNZbhrQxqz
ygFAqPWiRLrj2Y0dRCA44B2UsycUYaOFzrfFwaUJz9NB3efWywR2ede7XEf/0GUxDvxZWmV34IHL
08mk9iGkjo8i6YEpOgCKekYSKfj+kyOvGfkpD5bTfW/bvHnCWOPwWsYYiqVUhNHVmxLNXRoARqZ5
2p4AiK/IyPiLpSqIvDeRuPfoQKF9iRNgYOU5YxTRTtP8F5aproZH9f2TYgt8hOnCE3OnF2qAporw
ZkYxKcYjWvAyB9qvKIk9k5a4652IURC6c5uSmTHwaC6XT/a5dI9dBRuhUH2i+DsFhq4HaQDdpRcY
qT1mw4P3yqKp+LJz9CxEsHFw4uufKocWrO09LQYTsnPPFIHi9ThfieBayflAi4GqfKYo84wwkyTH
FELRyeOjW2uEFkv+qMDYqWZD90XmCzrUeFgu7ssExYY1GPSolEC9kMOlWRTNQePvEvzsXkTIyiFX
yLDkgsqTK0vGl61RINgRQ/fRgcjT4yIqtivovYByuCnHjXDPh1t8EMgBVP+tK39YeX6WVu/I0AxN
V3i6qKcZ7kuRTuqSJd6iQp4dWeHU5RvRnuAfDRFUnpAAM1Ctavkkc4iU6ziwjagfpVj5tnQpRRYq
ei8J56GnrbmPQKrckVLXdcpBng2qfbJTFbfkc6km9Ujt9DT98kGqcV/O96vq+rOjNGxjZkmp8EjJ
WUPr2myFAyVrT8cFHD++t+GZQFff+jOlAknW+x1t2TUoSPKYycB+WKD/O8AKDjSMBL13F6vbVbgH
wBPNINmX5nxN7mxKIV36OeTjrm++WJpRREuxP6z+BJVOS+43tfcQGEAlKJFhC/DEhP+7sfm1qUSN
Eu7v9MATKw5S8cRqJ+P3Qlufi7OUIf7VCZMt1abpbf2C//BBEqXyR1qIYy9eoHFsIud2Q2nH0YRa
DOSvoVE/5WJlwgkhAeaVeisjMdZCzJS8TpxqX8Pw0ogsZkFzQq1jYqf8GbbizwSSu547GHLeatk+
Ku/6SBxwKNAEV7AH8C9wHLlY1NGG1SddQd+RIl4qAO0cYVOOXWDzPz809H8WnZXsy6rOh0oRqABY
yrixd3FAcRY1vOfscH++2hGz3VttecmVgUx3ngo3eP0U5yR9xYJMIsw7zu8pX71VLWSUJlbunZDs
Oc0A2/7yC8C31mNd/O3FIRZWIy5dsoPBQyRwQ3gA3CajxBEteGE4lgRHw9oMuDF058DoR1dXR0AE
ofIKIPdV43nVcLNwQgOZVZOGROb4wg6DkCj+2XtOMr0yqPzO07ZBEqse1ufsX1qmC3RXMTC2Ff3r
6AGgap1aHZRqEpT2A7V/KJKXw1t1LwTuRH/U9YAIDtlAVbE87SPCdcNKKsAEFR5Tlk5E3PabNUvC
bSi/GtPIXRXlnmUsH4ssYDxXQFtwNkOpwyCcwFv8uOfC8WnSlfcfT/Bj0cSJi4+dt7x0m7VMlqWX
1SYkkJzgrKhDwOF4hwDsvJPJbK3OEl+ZiQeJlI8cfnMyQjitDTWdWxLgkMaXQWCXzMozfEG9MYUr
nLOiBS/DWXQaV2up9eTCL1yjEkqbsDccQYU39K7KKxyWlTCw+Nikplp6w+A5JceGoPClxqeqyqTu
nle8p8sHO+UFOwxEePw+W2wXghEEhcvx325p7TwZsHjlkiKo9phzz6vlr+d4OwABcuSdSar3IzNY
Q773mm5OhpxwJhVWIdK5XR47vNLhZCPcfiL3VJ9sMQQ5H1FRW26oApiIVKn4xVuQgNOGHouDdEwm
VOiO1tj2p+u/3ejQa49JgrkXn6TwUbQDUumPlJarLcxnlfsZw0n+8mSRPcSS9sbErxntmtgSTUQy
rI2mBaCQABMCQz7v/vAynQR9kHr3bNYC8hv66k2a2kx8r1GPppi4I+Dl95GTaZll2w4vTo1PU/0e
IHZwaUpLt+7d2ZOBV9vBs5452yihtLCLmYKbAlMQ2Sim2pax2ZhCe3oFSYSwKUEc+5xfnSm+fiBt
rraSle4vsRtu4JoyUDo5nM4JswAg2uldGk6KA670TQKjYR7DMVJFuEYNzT1Q4PPEQdVDDcTlwWcd
mau+XUYOjEhoEE/IyNwXkKVPgIYbhBIZQd4biyqbsCUGyWPYrr5Dim5ZqWd4St40/Q+VgQdJBN1J
50Cacj4KiQpfoMSEbQMUTjWJ1xRgAqdm1BmL3TvtviFO85u38GOzYEbtUzsXqqmwD6dPx49CGccc
kb8aieQm0n82gC07pqCTBqAPZ0w0BNayp3p67c1S1/S+JqZowHadu9GOOTvHdvVme6iaVKOWtr2N
xMn/nWrW7Z8jtvIE6N9VZPlFRYdc3EB7CrXBEgGSf3BOnYxvMq0JlkShvkL9q3Z0xitNLnF7ZHLd
LIcI6L4os7ZAz2TIZNTFCq7VAvxV3JKxBRIhRcdT+O9RxqrLZI/n+81ZM6ArtOkOqEP9qLryNuuP
a5dXEmpRSlFwigi0OebetAgL7b0748jo3H+miEPq0XIaPohv2fYNGW2kdUgmBtOqES7F268HUSPs
q5kVvSMQvrWvNjmGnWA8XslJGVigbYarLxaOdTOcvNikBGe5GqGnvCdkpcbP2e9rs0DmTZNfNkAj
2kMoxpELdFu5qa0QMEiv99yVSbazd33XR0CPsuEyPAHVl2SDLACdI9TXetBDFOPuDMEZSfwRJf+g
KSnkTBt5bX7Er162XQkhLq1UzZfsNJN9KDab7aqcvhGQbDhDVFTylbnx+6RX6DRS/AzwgFCWUV1j
S58nK/RIanEO+fXxtwJNR5SCKH/qmg0eGQ2m7hgJKPGjorhiysgGltRy5wAQKkkmqHP0kSTRFoPU
vf5uFc7MjnPBYeMLSlNvk/KVuM0MJzkTrWqmcsBhV+spI54u0ft+cY//4FEemiUGIwW5v/VrKVq5
Xbbr/Hf79IVfpd8aWtHyrA0Y8NGZEGQKYpearLyYO4K44Pk6XCFaZ9TonF19W6/vVAv5Ik4wJHkF
VtI00HNJwXodmIv04Rj7FHbveDWmGNuHA9jO4hhToZ1rvM8jqCg5RajMlIVAAN/oNv+dnL8cz+7O
LVedgOELR43sSMLwp2qeaYbChGODD6JmpHkGrWireGJAxG2cAWtLgqKLJGQNOrWzZByAwZTXC0O0
CzDwv/c/XM/rYx7xvDauslFsMuARvtEQll4MByCuqIEHQOIUxRd51AC9dZKlq0AmIPiBZ7rqL/rg
4hUNBEyl67Hq4N4vVQzQV7uzjzlYlnzGpCLdk2gtDHEKjyjo6ReqcZaUXKlquRHRabCQu8RxzFu9
6r/EAzulWq5cbdmE8TdeitmWc8tFhG4n3ZTfu2zVCxZxIBgfog9gO1aZUzdGxXU9h0yClGcceM97
c6/dtf47GXkp+cMlfYLtedc5IgYgmIjN/GdVWROQoTpHpo2kQPxG20AiM6jSfd5hj4St2xzB+uWR
ATcm1g3lPwzrj6j5nHWZFS85TkiUoE3uLN/p3gxTkSveF47bJRD0ZeRttGikqfJPIcx0mlA4VtOX
D1MBMhGiSEowfjrMPLlTysf4yqYimV0jvInkV2yyzTZWI3nMpsyBQM6XQypQFWO+1Thkt4map8R1
BuomskoBd0M+1N49Fr1zBqTKO5PbXfZOLqX6PAoqX6YF5xji4AUzTKp1B+XYxDG8apAtCD1lr2xh
0L8gLI4WFtBD8J3PfQnaQoOsREcp5wDhsm25Vb0pyXXQcWZoUpOawn5gbLKLchds0VJlTr/dCnI5
47aVqdaVneJfrAnzJCz/jWiNmHqZcKXQu1wzh+6VqBOIZD13TmWR2AgrZOX3HV2BgYxEmPcL3+kL
cdbeVYjqB2sxBvU/ZunLKGblmC3d2bbOgZsoy9QW6hqDEPNbvC6o4SIOE2Chl4roXiuR1LXHUFw4
6JJS04tkgDGA67yYEWYhwVtVG0oWfI7gC4bvKoBfceYoU/Q97oQlfhR53BmLuyi9b/Zmh6rNDFtd
pL+EFSP00NH/ZNlZAlqwhXVRGA8ISN5zt+QPwmV6yA/QHHWmOMDwP0gHIH0FDaBlQMtT9QB6OVM0
lnNx1cGgtI05A/4CU3LMUVYzbj2gWrJyElFPvUFqFwLXBHza+reOtcFX7o8QxkAV9nRJLHQ+h+bE
KSbPfPeex2gNmNxjKX1q+8wMUmeSDCuGLynIeZJP6cetxNXYDHuhKf5PZU2Ave2+JV/Hrmc+/AVi
iPkIcylzyyoVHc4OiEHBzxQPCI0iLUS2DEhTrIjoMZqOwDLvuGhB1zFZiFrbQ+Lt5GLB1QsA6kgw
22rNpkwKAqeNk0Tq7oBT42yKcKSIthoHh2q9SVCzzYapr6Y+1ksaVozLo6iHdAGgUbhhbfOU4wGZ
mA61H5G5tHxOLrtbY+TaOoA5wShIhiDpCq3rDA7FpabSzXAxkNsIia7plNnMD+KSQKFmWylN8M0y
hxHfDY27rD4D8bd+9wJTVPymKUtfxL1IrxkVNnregb85sQoBX38ysjqjxTbbyMex9XOhKgPO9K5h
2A8gSjLe9yvqO1VVJ4jOP0Zq6RnF0oqh8eq4VV73b+4wmlIisqr8S2hB5kcpKkLbxiopcQjaYdqI
YngnvyCIUxNa/IInUnnf19WLdTxoZlZeOFGaBfSmyJvXnLGKSNY6e5JDMCVUeteXToxsYRoer3AF
wfcQh0WvNXAkbbt8gwN1h+4P8Oulmh0s8wdtJ4g/ctA9qOhiqzLqB0oc3JpLGLDl0QPZ3mBcffFh
eguvP4bLzts4h+F7m4Oq+v9oM9Mt/XaCzP1qo9Z4qRpl1n2YQE3CJ9TADkSZ4U7JLxYpJyJJ1WHo
J3nv0K5Vzo5cA6wXZm9qATY6DpwJbXyXchd5/nC8xBxS3Dm1/tUSh6K1zLLp7kExOJyA4uP1Ewcv
IvmAb0eFOusypZzDB5e2GsYrV8yaOZ64LaqVc6qOohwmv+rcp6F6Uy/j4TB5cmS7SGyS1m+xaJkR
3VFGiP0S87RYUNVAVWjZhbDZI/As14M7CcfpqqqcZ0BJwvtpwPJiOSr+ye5vkK54sVYVNIUB8zyH
DIJz+OACzFIv++d2v7AcCRCYzi1HwBhl8SAD+RJC59zsSj16cFXIDbQ+jOU00gYLN+AxNvg6qEXm
zDn0+V9t02e2P7LTbIPKw+h+6YZZuc0H9V714WxtAcd5RxJaPsqwj16A2iZ1VKwpeTc5YG4iymsJ
DQ8a7aZcHiK/D/bPzVyBUPdJrdG+r1GqtFGPGCu40BhkYDj7ztIjbkJn7RjfuEVdCqwzQp4cJiM3
u0inZ6a5+KdJlWMJ98ySLngGZLkGRBf3h6OAsU9arm1FomRkIfpayBnPy0dsJkujYFjYzrP4/o9e
xR3mErGRiwHgZ9Ok94vnZ+cq4x7gmX243aPFLw5Zj6e7LBavYnlwcRlyiZPu0Llwgznl03AjA1vq
C0Ex5d7jmJm+6BYIhY7reGhc+Gz4ITHna/Ce3r1ZTe0+GrsN8zvFVzWrpW+TRv2lZuXrGo+z8GRM
paVLZdcpk3sJ3AwA96wufdhP+MWScwUxPCye3Amvb9Ul7sS49nPqAe4H1g24vjai8ND2EZEmR5W+
ytFs0s1DnUYpqOM+19uQXEDfkK1Y2OtXu80voRvYeTPMi2yL+SKs1gjSOA6+3ppLA6tdX5/m6tah
M2TBzydGlvUF+9YM5joea9vjFTBSQVx4dUtvYcYN0uohzmky7B5HbaAySNZwPs/zefJN2kIR/1aj
vZydXX902M9IMWhEF3PvRAHtz4HlbX8FqoW+VVG+Q6adTEdi8x6dzSZBkElnSK82EDRI5UNPgvOi
jCxV43J/hoGYdc24t0EKaPVP6164LRIIK3JJAVblqAaeGw78fCq45mSxJWtuQEYwV2/W+OuuYE0i
ZE6NIYlPns1k+JK9T3kK+EN4q4Qpd1XYA5CLmv7mKhloyLqZry7JR7b+Sjw0T2PgxGVY9mHM+rfT
oFGfsFgHzgZzqZCoIs57eZrOCLtxgJCSJNWpmQRbMZnebHEvvrujyYwaXs0gkCRhhllDpgDSGpwx
yp+G0HtThOu7Vb4uk1s5Fa4y846dFaJSiz/21rTm4gjNiBAHeyfcgHzWlhUKt5pvMYfOqGMJdScX
Twek7SGU4PdU2Vzw/bOzCVUs9pe0jwZVfPbcjTKHgBLXu/DCWyKcKsAL1OeUwQVzl/yxI9EfKNni
OsIzru1X11NwXAdT9tRS+XuBAs9Yt2wr9zbOZoI2P6WXrAThx8D599zi9wPu1YNwjo1B0t7Qb7x6
CruQHZHURNI3xBaG6dTpYOez6H66zSCwfhg9h70b7t7YBeTPdS5egjECepH6DeoZJ8a8VIdAWLtV
1yrZ0c6I5rgomnbKiGuA3H5DKAELiDWzS94IJRF9X2Jek3acqBPUFVfnnMlgDyrsZtnWR7Odzmeq
uSQUYVGm11itBlenDS1afyh+g9sMvgUiSfUap0uPomDgwa5HZlLC7Tw1Mpqz85IWkofwl/NHfb+Z
zMTZuuj7uhO0/mZSnoLKY2f6c/g8UwM5qmB+TSH4xyVrET/+LBFm1lbe2EVoX5wfgL85ID5ddrkf
OBrGg2CulwYMHlwHYI2WD0Z2FDwKrmMTPAwV9Vz2vKmewIAfaDTPinUMbjDpR7/wDgoSusyfuRGl
UVl2L9pSriuU+t+mblN7KmVMcJhHD/jY7owPCaOV/r/0pa9LuHbnSEVxOhz2tSFfYP4mamOfVPG+
VX5N2nDf22he0QlNHz7P3sFETM9uvCUSYYaNkVzfuvogmBH+DvnptcWLvFywJh+RVSHLtl0etTkq
Ytx9/wUccUnwnrCTbDjd3R7NwXkcNMk5Bau2xdCYJ1/UUvUVpUuLooh+h7UddY6Tuk6izwtM3epN
+NEtm7DJk3ghc35qY8elX+Vqpsy4M3YAWo8egqVPqby9J9Qwv//s6Vae9PZ8IfwMOpHZIhNi49pu
7Rexu1o53ZzYk1HbhG9vJ/eSq0SMNoVnE2dSNKTf70j6AoO6T7dxyqf0M0Dn89ccMCefPk5ws0l4
L8+/xOgsKOvUD/xbRHXCV2drcMIh11AClLQjVD5ZpRlVBkExtirp9wEK4ru8rhVyXAaKujcl3KN1
n0b1l1IioeInEt+FdkrKx7kRH2/enjLDcvmOLsB8aUdi2ZOVe/fd3m1sGJcWOiOTRkqayPERlGeD
qHVXN4QWWxM/pVbXxt50kKLCoPHteA/sX3wQtIkyChXov/7428w6fNK4o+EfoSv1nQ8Oe3I8oVVz
Thvsvyxju4zUIV8rwFyDtWeq3871VHsCnVr2T/SKQouS4hnxjF9dTBtsMuoc47LkAJcN9t8/FGE2
CytzVk97NgTra5i154s9qkhtyb86M9kSyIKUCCygU5XDnku/L24T4Wc+RiApN6drE8yvezpP8vUI
6W1H3lppHdNAQSG4olXApBF3pPUw6scf5eNHA6+iQSU+IIlUGCc2mlOP12dDRSxLJqnc3CmXmVH5
l+fbVZQChckWAlYrvb077H2Hx0eSRlJh9cC4W+JaM7fYEHePP+088Yvn3k7lbZj/UHch1TVirFh+
zjAtr1lWufGYNVBlDvck+Zbk3E6qeYal08qkCEnIWS5/dhco1l8IO4TvhRPMxZEzNcpkhBqcnO4R
r8uD/n8nUkz+f1QyDtUkIXAisJc4YpcOvEspnq/NYY2mc24fUo28aWOuW0byG6QT/Tl/eDwXYmn6
5OZXwJ08Kg92vbXMI6NCr/hNiZu2zX3bdKE/qjnWJCMnhixafqR3Qe7JhxFHYedeqeZZ+a0i4Zxb
IJmWJ5A4AwawTVT0MU8zKuE3uGm5PgX0rsRTtmAnyO/KStA3bbdDXyH9BNYqWxsEcL8os5obYdde
wSrP9lRNUFkF+O5JthHna5uS6fNcofyjiphfFazu5j1nlP5V/ZYvYa481Weqr5+p0VvBr4YXiO24
ezieglrMKdYoKWp04T4koCfXrh9FXMAgL3vdKGZTgz7AalpjZtwQhXqg2JyiAO9DR4FZVpqDRprC
QvChcR0rZr5jn+Jd7b8reCtVAM6qRlR1/AY8CaFDNoE2LRcoJYI8yOTWyV5h66F5gQU8wca48mOF
4/qaEKNnuGpSW4giMJeBRNcOiigjydnCK+oyoQ4I+SdNfHjz0C7hoBq7Td4jf0MHFHkj5athxqvY
TpldHExaNfSJO0ubc05lMdsHsD4w0IiMwkA44XTlSF1tkvz63CO+fQJBLDi4BW+PRmG+FfDkZhif
3h6a3Jq8auZY1ec1OHhyLdNdOFqjn5FS6VVWZN2bbGcX6hNW+bjIobo3g9ZNYu0k6aNYqiRa5BCU
TffzzcqCh7efOD4kaJWGMGj8kCTCJJC4WbVyVAmVcFexO+dvXHDoyOFtXBi+87XnrjqHGVTUVYNK
yiKA+bFZM+Tf32sQIiK1KIGF+6kPWp0mVPrC4pdy7Ajr5YTLVCDMHMUx/czn+f3pJeIQQOtiD5vU
xJZwG8I6mJHznwkaTLsWg/mN98CgJ10Wt2/Gkp9U3O7WnMmGAy/0QoYeVf9mICx4xBqkVIs09tRK
tSy7SQol6m9Qrv+e1Uy4QARsAIgNjPDt+M60qVl2IKkRejKb5BE2rhLGwFos9h1nEhOVDmqxSaZQ
Q5IvXdqkoSmGdc6QWNHcJkbHTLBkvbUIZCWSktavKIYJOIvZREmWoNcteBb6l4PpWGbv0o6Sh6Qz
L9ioqbxULkI+fxwNmWVN9Ak+FfGEyNdenIh7zsU4rpEmsPxhoVGqL2LEoPeH4GYVIoTpkbpxXbfF
6rl0jJiXHakVlsj2hvTdnZrbCUPZVBGgTovCAZD3ftQofi+GVjVo4bvadwTe7uzx9JnHj6i/H33H
G0H4P6motjM03a+H3ZqGVSAi2uf6yCAK7e6PwO50Vc5dF1ECE1O18ixMOgpOf2VoqzanJnE0gFfP
fKdLvkykn4EBlHt5OAbvwaAD+IpKDZTnJjuZRW6C8eY9/+PpQLU7z2QN+6e2BdOjc1/4hzHqLcHx
GOkKZrdUeW3CYJeJsMOfjkOIqShVNsH2QuCmtASJ8e0KCk9RZMUbnPG5rnc6bWi300ml+ZnX0sUC
/xIcpBAeMj/wlmXP/lT3jgbx5IIagd3JCufFvhMjGRo52IiCQ2eknTEX8wO3PPO28TUQbrZQMBmT
/hi1x9XTdzdia3mrdvnLycxJTD2Kot5acV646Ou5tkl0gJS7oJqe+MrpW8pXvD8BjVFGT7BhXcgh
ueGlCt4e//KNNVy/rfmzNZ3/lTVAHP2KV0o322fl85Ts14rr9vgV+CG+iL58xFhZMnvWwUUCfd76
cz017SCjywNid5hCP7pfkPECzBcbiy55WbaGALyDUOobawg72Ugc5aRF83iHebhU+InjnkrKJABS
wdsJLSTrtB9AquJu1kopdY+JFBwej3J10aoAYwqg9uGBb3z2XoTnhFeOevwb2sCe169HaQbTs0ZR
VLt04/91TEGbO6TnqPTq8+HViSGhTUuACNPG/OUiaB8+eM3pC/4PdFX99Rj0g6O58jRfSv2wbm9u
/H7SzyIgRvoM4K6Q07mbLE9H9/xb+gpsBAx6DEI0Wv1EoLtCpd1d49mKvg2UVAQ41RciBeckzN90
4JyzqrE6vaKYkrBDDAlvo2fgDma2PXDyB5jHYPRx5PEYD8MaTQP9d0pKlRk0zQgvuXsQ+5BlSv+9
ktgwPLOjyDz+/C6d6wlJqWH2R3Aw4ixwzLHy7GYwmFiVIN92Va71/NmEmYu3r8v8FJeqg7E52AbB
8G2DOSUWJUaitx71H351u68OiiGkPIr34ItnHVAYdHqKk/x/7S+ZDrpvaSrPj0dAdjej5TnCjiXy
EBQZ+88QbVpSfV0rjmy8LzgQJnc9YZcWp7n+jMo5PvMUzJ0pT2WFzI9eHswBODExfX2qHfCCyUa2
XGZnLOJ7R7+wBGhYDQsrdwcQhcJUz4u95pdwHM5Sue40YQsXEuBPzkEKdln+vYjMPITihWVsBgzO
rc+2WpSCCI5nSLDKAew0clM5l1iq5xukV3eLNSeRFZreR3jQjbwkr+JWeVpD6csXuZfeuDGCST/2
2rYpNqUVeQ6KgNQhiKCFR0nhyHfypAZmchjgm//gQnLcwwLPZI+EfdWdoLb6yLMkARuWF2Q8zrHM
AUiAABXbjh36mES6lkMvFhigmI9UTv6qI2TRHzeRaso99iqmvVS2MTgCqBZP2mh/sr04S9RAPQ8K
h+BoMlaF//4Trn4jKEaIdVTI6gWjMS/61pzXSrYIlv2jPqcMWZrOhq8qeqj6E8uvPzaNkYneYRvg
MAAp3PSPX9MLlR9ttTHJmqbdRR6UycnvhyJkfcpt55axPW1hOgufH+J/c7jecvzdgzz04mD3IszV
1Kz2cFRuhqs00GIzEQWulOcWvEMa7v1MnZXkZPsEy/4okhK9q4TVJZaAJLuf5/g0clyNKAAobuRT
iauP4zegUn7BkxawKzEWF9sjgKa6+yulhrRZ4wUz7nze3Hxk0Fm0xXV9MwCGe3sHuvIM7Gig67wb
bvNY5WBocY6680Zt55T6GgR5h46M4NwLV1Jy/MvJ1Mdi79IcAGqfxvuaWQvpo13ka/A5IgN5ARPO
ESzWe8jW/7BkbHsWG325U9x+rn8q1OAH1yYMIe6OP/oaqHGLyBlE6n2gG0m8/u/hd0KnK8j/qEjf
gpawCUSeeRSFvW+tPr69dsox8S8CKKlSbWdQouJcISB6oXJfSDRH5cZFioqEAB8pzrV/tKBoYtqD
QfTE3YxCDydSenkqCxH4eL/6QHrIXNGn7rGY9aoFrqd+2Y3NH65MDqH1OTTsL6CmamvCH344V4Eu
FF0wkiCCurTLhw2/XMzxLyf126PvIwOzdWJU48JYXQOtKWAhEP685Zynh72FPOxpx/NNOlBqEKvl
e2Ebww3TmLjDi+IvTBCXuo1HUYgf4NT+JX0p6IwLbQBoue4JKeA4VP6DF9R/wzbuYUnAG3JGv3ZT
jI6zc483oOrPtKxObEYK9qC/13qyAYcd47oYy+MVmKkoJYTd/tgiuendvH6aBwugcGqpMW255hd0
8f0bpC9J3zUeDI8eT3zxr9WCvq6F0rrYTDLyLH6kgI+KdZ4a8xbIoa8vnRSraC+cu5VuRQG0EhM2
Zk0KYAu0bn5+0sq/W3zgMnJOcCDxed8BAqRMU2Rfznxwgknc+DM5Ywf2Dwt/oEc2EaYBKHG2EngZ
g6y/3AG8y3Djzelg5sCJ8H7Hp+3D/0PVAtB/gPj1lPXwf5KgX6WyE1FNcEJ+CqN1dc/Hd6Hk7sHM
iUDGJcGFa0+wDN5pn4c94ld1RUgajDtTlCE5kinzu9Wy4C5A3mJICXvNv2CI2DhLg1eEwu1aRVNA
sPS8VLOBCZ6I5u/T3uAySUJG/GBSYGGHVQZF1HUV0XBEV/AQYdcUIX83FJ1i+v95qR2xnCCJG0gU
OoEmq8hHotZCV+57XXCWYL0Oo/hpsdn+gwPyg7COjwAMMSNOY3f3Vt0DSjvh2QiTT8GqOdm+9BYF
7MLkUxwKDW7QEvrlfBt53KRpdjSk9sD6GVuFaQsLA5XCDANNjd56u/liFyGNLjppeDs2AgOx51yE
8CTCqvNJq6m2D12E70Tt0p4WDLNPFDEjLTJetJUkhqoQcmIGwQk1gJYY546RntCvYOP68zPdU+No
aPyMtJ4jpMHz54Wrbxz+eR4JcscVPabkOgtqeCMrz0m3TXmTsAH3yiTdlMtQv0my1O7iM9X8Two4
w2vtInGP808tlsMSt9ftTQlWO8CdOzWaCWpgB3cuGF4nX9KQa2fLlig30/zBVHuzDB/PPsHRjj+0
3vA/ocGsMZnomaNNdbnfa6/BiE8Ip4Il1o48GfYheFw539MUVedU5lqqOS84MbRjfc1SgvFeLG/H
4g9IN+XjLcat2b3Ia85lDDXI5WKzHJCAlPWihI/nRClWl4naJIuldSC6K+KPJwgJmJ2dwpyCo6OO
XR5sp9UtnKo3yOp2ugkPCYpdk1NNd+i1iZcIVcyOVGOiEGSnCnK987rZyYaSTTcpF2WGkkGkya9g
N0NNgMxOTf1fR0fvQ2rISHBK2AkFYcp98/MWNGEVWJJKu8O8C2fzbEJbT4OnQeXpfEmbCJ0m3C1V
AA4QwRlrx8XEBv/jCttwnlCyimLHgn+Ykg79VFLROg0GklZASXrOsZVWpzMgfvBAQGNxPpyIiDRb
xXv0qghyQYfT/pag6UQgapox+BQHVfz5X6x4V89FLfceVbwZmPZPTevJLfwMv0MZIUJh6PE3kCmE
06wWPkvsxRQIewU16a7UDFXufDtdaPjFmLaofajHzkg5Cjy4U8x6Xa+E2+em/D6exfxwQZDo6iPs
GL1J4i6RY7/2F6UW1MDDtkoCzNPX6KrZwjHl88JDsuewTKPTs/zrVM9jvJASObdrYkfSJGc+pncD
2tW/neNpvaix1BxyK9SCAGcSIH0w26LWfCycSLiQuPZdLuB0VIowCuO/YdyQ/wyJ5kI2BOJOBjlm
/VNPWjlFz8zNUBRtBltSdqeipnjcyy4N0YirVAar4MOtZsBD6flYbi48OyhUODwv6kd3nFXd3F3K
7KTE8A2bLkVeSNsg989AuSoLuXXaks0lLwsvA7rul5nt6SQ5NUgq+ikL4EgxZd3ShqvUXWikpmgH
c12DXhnDVB9adc92HE6g0PmiutYeyJiFla5d9uZzt8eSaXabFxY7GCZHIbAAg3OY1Zpj5zqV02xF
lpcwauoyfeiSoY/RLGFFLFWFcYRavhgPoVeGFjciIl4N6e5CYxFaOwCCTYrbsiTgMNx2rWFMx+ZE
OOYWVfQtEpzK7a/XSTtxrWNQdKtzjO5DtccWz/cBAsWuhNdEga4Q7lZeeC/wrh1yjJuGgCq5oxi/
B0Nce299/Y9uM1HM1qE2u0aN9H9rD1r99jxkJzcfMMdZ6moRi+XQDTczcefhUHQl760SD8efGz7P
ETPKuKSc4ljnBgygyuJ2Z/9+nR66hyFfKoeOqXwHWPFJs9NScV0JzJw5QF+UqaEsjVlxrbL3n4BB
zVPH7Rn/M5PMJOOmYwi9jrYad/w47r1/Q5iJFreIwjBp+ibSAxQQ183DzsHNvhGRMlu11UHVQOmn
iL+iEcaaR4kzm52h6RjZcAQHH39aT9zclyzor16z5Yu0TzEWQExM9Xr8OC34ztRlvq8XirCBDfRH
IEheMayxUWIIC2MbFKNmPlNB8RM3xcEMgdgdD5M3ASTEBH1zT7bYHUvv7XVfr9gE20NIYr2eRtho
UgBzdw5MdC4fYczwFXMpLhZVrZYlc3ja1/i9fFoA1MPlqtTCs4LRgrMcqkRDDG5eDhAMWPg4M8t1
klFLIp0qNrEnVg3rkIRoRx52JZOkpjuSpx65hlBqH/Qyr80vXvyp2QAbT71SV9NO9u2QCIo6CV3y
pqYEmP2V2IchwNwDHIuY6ZrPy9+EWbSATZv3g8lZb6ZJ3hyiF0OLCXQBoznWAApC0WG4Qob1ObHu
oNUoaBFVPrFB+bd74dsXP5GcPq9Ijf2IpSPS6Vslei4Gj+a8H6EoyZ0n41OQIM/Qa1T+cedQjYwO
3ufdnPDgn6yhqd7qxpOdjYLc88XFYVhDHJCHxH0ysRya3dpzXwp8hpUZ9jb6cLQyGNv6L1n+F+21
rIPeP8QFGRoYfFpfDJCI47jtQWc32Av37+MYcAYkS0GLhbxauMfB1c3nJWZEkZ2j85ZcJDGNY4f9
haVjHa54I+LSbqr4yTeCuINIk/LfJnLANPfmCw+/w5TarjaknLSTVeHK1nyBKmT15LaH/iOw2RT2
8i3dtjRK9JGMtGMAItkSPFLzrSgdxxuLUpIAOcVpio0BLwIRsH7Fsx6acppE/167jdIc5D/7DmKG
1pC050KbOL7oGV5OgsxY9Gxbb0X3QnvOoE8M+EMigDSq5ZP0xJ7oXesGyPAxb+9yFF7ruYjIe/k/
snr1Y7I+VlO0j7SUadRJeYsIbYqZs395cqAD/RIi3PkVahsLrOIufdyJvpA88Q/i1CfvpQCKRQeW
OVmRQz3mK/QFAZmawptgXE5QfghPbd4t6Pq0Y5MY3yvYT+41YetFXfssH9B+VcJXxg47FNg8K1UI
jbt4W94FIAQ39ARQ81QeavhJqSLKIgXW/rXJ9QHKGT4koYUTitteL8GqK8fVBjsASLRY5Lqbimu4
15YFW8NPzn2v+PB29vWTu4vURYUsMqLkUw3Cw4srRhTSap8LCgJnChE9ROctoWLHXMWBRZx5upBF
8cPFuNZ6m4g37AJ/OLe8DB+JRxt3HVfXNsn56PNFG5ZehBgJEHseiBJymLclhGOpJhLP3uU6Jzfi
9utj+/bEOxrq9qblx/bGs4Tb4ATifDbcatRJq11I9sDxT3+t1ubkR6SJ4pNotM6tREPTj/VuzhkU
2+vP3+ilW/JDThs9PoC4/fer4iwqSKBPYIGwT0EXU+tFcu+v1E0TxSuXkTxKU3HbEARJ8jb2IY1v
YVS1POulWHgfsyiCfffc8Mpj9UmAKB5y+9wCANWXYjaEe+pQVXOmjgIsd/flDELQualbg1Fi/xTm
gQ0qbH+CSfTlOeG5hdYLvKoICzvFgLqCiKIyJY7MFysWi43N52SbVc4Q+n+R2t8pPqSh1j1ETMSZ
u/zvm+7UbTMywFVBE32+QkJW3kzrpqTkoBEswX0JXDA0++sRWr+RPL+pg89jpN2d4d/WZgkfs1Ax
TD9U8zF9OGKGe71Z0dZH8Jt+X/sljMsXREpAHVLqbrZKicMN/4lZp+bPlN0GE4+gESHECEn6eb5s
7EnWJanA03v1fOioYyejpzPQejMv5N0hcCsGU2Q8N9wrUtwpsLx2G5ssbp1Pia85p5Zv3NyRC3OA
kKcqi83oQoT9+ue5DgMynuRoEVPqhgEsJqQALmwunzTf5wk2iBazd96HMHLEkHyiDdDDbIoFEHw7
5hFEDhIncuwwWhoJQCXl004asnyNPYegZ60tBes45M5PxRw1ieA3SMPMhQ6oslc0KQMnV5Is+o07
Hc2dVzyEmJjIKXvah5SzT2w987Pl0xStOAcR5dF3wLsHqMRXw7uBJnZmTdh9qz2aKMZe8YN8cwHs
klo1T8Jcau4q8TclGxyCpD/rdMaQRIhPPFXzz1krDhGaRvTsipC87EmG+B7DLvhl/PkayK2s+RMf
Rpcg2h3cSDJVeNpLCz8cwLJ45LAer+1WnQSEN9GoKjGP4BKE9HWNpqYE9zTG/cCd1vQ9Dy0ivXlu
S0W+RR/6kWucyA1+MdEqkfJ9FTPIvVIFdE5jlJa5QzqP0/pfHojk+SWv95+gmUIF9YZIH1UXf3KA
4Q4LlkCARRZof2a45VtuRUCHNsdw7DVrTJ90paGfxewlXrqD0JEJT+vMMAjXgZnsxDZyQpnbuX84
2mD1ReIbvS8pwsDFKdMhMBmAqBRK/XVxklznu4LEo9lAoX6yIY20/L9zWPb/7cPTF+gIGrR4VRYQ
bcoZXr7n1VVWNyQiSNk60yXvPCJGyKC4sxoUtBzzShMs0gnz85rIUcqslMYxvqWKDnZ3Vze5KTGT
HI2UkDexpKQV+NQzdSLg+QfuefUxj7pdvs8vk3/A80yuwb9T1fyitSqkzhWchlaUpVzR2E327YcK
fQCL7Q91GXGAi1hdO+nOHXABam1w872y31aEKW6WFS0P+V2cnFDuWeGEREsLpzTJFjSsj4zC/Xz2
shTmO3HVHzqvrlzJz+tu2dA6/g3KNKVEJiWt1MixXKRa0UsNSdnRvWFLqn7fhg6AmbS7HiC1bJGa
LTAoDJ53r4kjjtYokhyX1E4gl2wGzHtQBz3IZQ1fRPsgc1ihawtrbPzgf48C3hdtFerMYibpnRuz
xaaTOuXbtjoMtVG/bnkoEabQ+jhFE1VUB6ujZD+ii3rxAXfvnqGUkr99Ltbx2fW1mUIKdHrMs+Hh
xQv9GmYAkELfNAZQvrXYKFdrFVozPv8wXsH3R5ctRKIb6pHhS0lSxIabcgnPWDtTrUtQV+B4jh8g
JagdncyqY/qly7jBd673FIT3VrVsuwD1wUaiwYy7eKdAT2j9xGEJJhcrOVNZsSXQ1deJ8SHfz4Lg
sKpYC9Qar4UPJdGtlWiuV3YEZx/M1yBt6qBkpeXCDv4IaF63MK4py7F4+9bPI9xg1w/FPpl+tYat
rAxS6LaGu8g02dA8afMLntljUmkAbrGjw983RNMkf8y++sY1hIUps5tlIVaf2qQhFEX4y1TbNlM3
33MIpSvLC2sv1hWH/kH8wIxJoyjqVX89ZLrDPhS3VuPc+NHoKj4JbB/obqu/5qyqXUnPANKVc4hc
PFRUJZ1hh6eIBtfS8YO9GzcfmR59C857lc1pEMVm1HccYYTSBne4Zh07cnKieVgIBsIbP3GgLqpg
DGCGzdyUoLKM/md9J1Rrk/RsXzCNRmS0T4ikz8+nYQUlFN/NN2/95HOIy8KG/CdfVnMIVuAIqFPj
7pJVSXg4K/oiCMwY/m+4Hd55yuH4f2P8i1ulQ4Yh9gMzAMTabMKknZie7UN3GAEptHxxXf310WmI
z+llMVpzdcgorTm0zHi7bstL4Uhh5HLx3yfh2M3ABv2/9wGFXUtA9CBT8VM1SxDlGlhFATTM5pvj
v+ArIvtAaw2iIL62v1h9XZ1hDn05C6OXYORtLf/5BaUYNgpY3JRSUhQJ336cC0I3UG0fpXdPoFK/
1UwJa27ZfH4wRWL1EIT5xfvqrCw71tc3NNX/DUGGSwNM0BXX+zwgvWHhK26+3RSyRZdhtRWegczz
02wYffel2msiXqFgwdCzB5yZUVf+7I0ACQ9Gmf8avoIlarL8n9nNhC5SySNcy1G+8M887mdzMgt3
VLN1YN2CMxd7q5uWRqtTVV6bqUrBBYtRJjjUpmpuJPWiaNAUchh5ABaS3VHpYzhml+pmbFb6bZpY
lFg9/tIlEm0VrjgtQ1/WOOqbQ6+RcNGoJOq5W0j0VnDkv0nc7xVV2p5WM0avox2EIBOnP79eywKs
MKvOpfOCExUsccin9A3dVCQxNU7inSrtCvOWyX69wozMo27n3C3NLNjD+dJagU1UtR/jExCz76Y9
nBB+tqoALvF4rL0UYcfpcPiB6r9rPclseR+l/cuCBKyFiUInHaUaJNVsMYmxdthGr/5NgJu17qfM
0sIvASGAWl20+r0husebMM7lhkK5Ri/ENGdbKyQWVjxQWiVhC2lwYpXiAJcVNDAkbUaWAg1OeJuN
iwdkkvXYZR24rpTAnpFL8ibIlOlp7F97OecmIMtVFZtrMZkhcayXtakueE57U3wTWBj2zb1iU6nA
14kX3Z8BGjLwqm59vaIgejfIkEF1eAz1fNcN4IbA5IaV0RTG+4MsPhPSgSB/OsOJkmXzTI22AreX
VdVKhwleSkME7vHoiNZs9BqfIxioC6tuoqJBBhibZklFtnE9ugxkhd/kyTBbRs3G8eYKgOZ9sFSX
nhDGKJ0w0u3GC+q59vkws6hQuyjvFcFifn3CHfFcmJ6ljLJ99NRkDSexvYi1lvBsgjjrT4vbv1Sa
OA76XxpbAPmTOX0nlJq/PtaLxuPmvcMbgH/axrlBw0mIF7TEsS9/9KFIGDGYB5lYEmupo7z7Grqc
MnzWWW0GwwwaEONmdow7s4gDuIPavtzynW3Fu+AWVRGZ6JkXPwo9kOhrgHXVH6GCErg4GrNbRDZ+
LCHKZPOEP9DwV3RXj0CXvZ5nyX9PpTdUCXpv/ogv4ig3hGPISVWcmA/Iv9yCZWsyxvo+EUxR3vv9
7zFtFKNnGcaEJwXb7O5WrpPWI6zT78I7V2fx/rv6wYogr3ciWx4qgK/fgROXjgIc1tOAo5V1otKm
IoKF5x89gOn9r6MHfd1vZ6PEU3p6ZlVwrVm9z+EojHpvgFxu+2crh/uIamUwh3UCCJrNZJL0mdSP
wlEQsghNCAJJV2nFngj9Uz5Ybk32A3K8sve3dVwKrKQeDxbr/06QStd3uzNtXX2pY/c5UIoG2qt3
0JHRNk6T8VDCSvMmRk5pumWwlzxXpPrVlw+hDi9AXhoqSqN4QQtKnu1LX/tDTHvQN9ioTk5MAqWN
Njo1I1RyBU3mbgp7bgtuVXt0tqgFdniG+LBjSS2407HeywR/VbX+AkBzvxOwjvaSv1B/05EIa7KK
ccJ/dHbhAD31bDWBuiCCTSF0WPyHDFQTpqhHRJp2TSYUegfkuud4Mhq0n+VOBOOe62BCZT3M3qzp
jjvpbrUuqmiZx0vcNV17M+8P6926Kg1MgNVyGYzbdw2415YJSo2AbxQ4+Gx4lZ7l5Vvjwr6dThHS
kCK4HSQcVXuDxuizvdGScU0HUMMBiGxdXWvyo29kAVnbevtFAYpp7MeE/U0xiT6bxxl6p/WhxU9D
gDgvC+q7ZmEeoQgON7tn6soDQIOULbp/4auv2/7kPdkG+Yn5IIdik8P5NWUyrgsTvg+YMjbOsCTC
HKegNyZEhk96s10ypDHAJ/hPLB6M7NEfZ7l1a2rbzcVfx+E+SS6Ln3JlK4HesRhnqIDG6lrs794D
Afc3zHY93KQlf54dB8s5vH9N8jc1DS5A0Nq+ZQr8h3YsCCeDxFAHBE+l5IJ4MEPIDvoTBV7T0Xto
KbdWt7iIgLtfrtlTVBzsEKIzekSwJTMiLC68F/6rPeeHbAYf1Sb7lvOVyybtRlgPm6OQr8bB8yKA
4eLNi/Pmn2aLrWDrXL0fbNC5Ws0ApJJ7/LjOZ8rO0sxmNv3rhOSD//VQ1AchaA4Feyq1IQfSbDNF
wJh7btI8tJpuQWmU080ZyCC+YaZRs4z8LeyeNrRi2oujsMPpgB9bz+okfF2MQx4y/3magtEHWPV5
gWBcrytIsObP1dZq2BydquUaGH198CjIqvqHV07AZb7KPcrMrDox/f6lZsOve+DFZK+Wc0RVSVjm
Zdh86sPLS0MeORBaW25OFjxg4GSRk9yS9Ui5iSNnPrrx6hHnHHrGGi7I+m66u0Vn9Rj/pk0pxP2v
KdpFjjWnHPJtz+GyDF8lrbbAg9GdXEbmto0lyfnxJsCTqgtfxUqXc6QZQQu4gPykQxaYjRKQx7nP
jNY1nclaDRntUr1si/XqBVPG7KA2WJ1jgszt07cb5Mau6WtndZTDpOlltkN/QQBAIckaXQKeLuJr
vIAe9/1YdVxehLjYcNotAsNzVaom0jn5LwNZZbAnTnbTueuY1onNNCZJl9im0Z5zhbtNvh0c6kYK
W7/Etg4MBXmFDtFcm+DXiDQxJbc5KIbTOej+J0F6aAdgIS7cVGf2p8LpeGw4AsjlLGsruqDdfkjx
gteEmjplfL3XRtzoStLVyqrlv2OE+IsXTGHymp4/+xqMFoeBRgozFjyqlTOZPrDGIFZhjGy/18oE
mAGkyN+ovwwQzeem/gf6yKZWL8sfF8HHmKTJ3uSG+DFiisrGyz6BzK6qZ2WZ3DZ/150lFTF91GsK
77kHhRYUxeE+b6ARf6zYTrK12s+6d8BUxOD8SqH2r35Y1xRDPwU/z1mi+9iAJrlWVqYQQ40xVg2s
iZpoJDj6DDlgzPEQhoJr3puE4mXRSzJT/ZzdCfLb5jwfnA1kL7EB+qr9lozA3gJAyQo+Da3VX3VQ
MZTKEgjL22kcMT3+uSQ9F9qqCq8S5U6pOZNI7tDJbVjaYBpO7E+YdWzq9chOPPu2uz72YbeHyfiw
tmlDv+Yp6ZvenxiDncNIP1OW0eIf/bnqcipBx9WwSRkraLOKtBDI7rQvda0zx6Y7cX7ejGID7BOg
VM5Iqx9zleIUeXChxNnEgtqhhXvJvtvFd7q8uLAy8oTQfPYZk4o8CPn4NJMHyH9ipx50C9p7AUkz
y9yIw7McZM5zfG3BiktmfQ3/rKOPmc3i8KmQpm7AH6K3zZoQTAvPHYUbvpUp0uXuow7Qpq9wUO37
qG82cyiR6U7ouaKlZHrlLG22Y1On6OAHufpr46dBnWycS39Uqx4naaYdcwrSKpw2HK6CcaIAZIjR
8eLVRa+Rk2vrzbMwiTcF+tg+563ZY8hID/RDlwKA0dEyDIYtQYHZRGNgZrGxGcGUBEUEWltur5nL
LE23XXbPFAxZIBYVHCnfkCoLFWK8758UzNOTFXKRn8or/HjQzNMKaqCgXXCOkffu9hwkpqaFc7MG
3To7c/BgaXQ0OnU0aiPMtJX9zJxvHU/oe80pV+B1hzrIoLNHPZNfEd4/XhbbypmAtc0XsvQeBnsz
b4P8Zcg0ArQVodrw9yMbPH0uvM+pIua8rt9iF6eQJw5HC59CdvhnQ9SKyZ0SP3NS0T7ITXsCVz8D
/cHy4yWt4iaYRphv4Mxhqc0JfauvdEhOcxjibRDRoNoTh9dEP7YICefAU4B/MVi/Jesgpel9pWRw
RYe9CgvvKvUjKw/UzUK5C1OfTskB49v5fZnSZQZPVFuPiPCK6f40TNoxugO8slx95aj8eMjVexL1
NzbNTrLIC2RkGv/Bl5pCZUq/WBi6u1ZfNmIamtvMCWzNR1ICOHSNxxQhOZx567HDBiaMQemVoNHU
RXNihW0UrIbAZea4oUFbSbG5kKLKbyxasqukjoMQolCVjxB+Lx4Htz1XTH1yHmisWS1U1Y7QRqGJ
YjiXsupwzd3rZW1tB626uXKcrM1PIOZak//pTtzSBQEka7j1/mg7ZdPgq3zTu0/XneHaHILPHIKZ
boezbmA1Xtic87vEHhmpQy1v4NVKPhGoyRRT6y/guWeyTYsuPSZToYSAXpRfMNOX2Bnm6Ba971MN
lJF94GMbuh60VzVZXZcg8QizU4W7n5KtTmlA0zra0UX5GUPLXVXhYx5fW1gyp6wnJbou7R2y/0dg
gOIk83wKW5grBJadP8dbyugudIf9i+8AfsWM8brLWOpN4uE1wzBh0um3NWvuhZOQefondS3IQP1X
thmJ4RDNO4s4Iz1xcXBkhRsRXNQlvOse28QCvOXpr1DeEDjj/E2icryhRGSp+tZwdXg/ow0kxLxM
o93xvIROzQ6cH8s6RKWviILvKT1qDqZFQOE3fW3rspJgHojpizKW+ZOXEtTS+4zsKRitm36oDK78
w0NyTM38sylM6TkXCMEfJoqsaYaGaipUtQ1DMCVKJ1fgs7FuQ55wZSaBTFVAlkH5riKDh6xLIg3s
teT/aWlkXPaEviVXPc2tn/z6riQdZlfSE5FO0R8xq2AwNgQvTFBDimRp/4xWWYUOs15PVGLkDbB3
95gPZ1ykUm5Kxrzuz0C1sTG0gHyq9Hbicrxfsh7BYfTfl4k1MydCiC4Ef5mfA9Gow7iyB10LRU8Q
huqo5l42/W4ZJXt+24HbTAjC3FKVJS50SiJ/obw6LoV3v7jycRSH8wzq+igGPYAan4tvLSnQiLZH
f/ZYLI7lXyRrwWDRL8rFVCdy5lJzGbXmg4tcvTnbi+8PHAvxTuU2GCIuxokygLH4j8GX69miYZ60
Em+055g/fsLVtvPbpabh9qGGtWDbTCX3oqWHgL6VfQdU0FrH3Te2c6ah3UtN3Le3/0/3/Emx89cP
mD3hcWzrtdrEevT5BRZDIVGD+eHDcdFrtODndHmSIBK8NF7eQpdZ9EqagpaXo6G8C0zQ9rvl7ghH
D7gDoU48R7eLIUfhR/6J3GUoyREvgtDxIstW8OXIeJysMjsGDLuBoMpUjTS4s/8wjVpz11M2QYzk
FYnJMdXSVQbKn2vLJLgKudD4kroXz1ont/CJ4kKTzK5DkzaTZdO5bQSgrRM+rfyQF8HdRD0MfRUJ
RE+9qSVwBqH2Op9eowWmOq3VZuSFpzw0HY2XTHVGjlpEW4xI2hGKmyIw+stj1rXs/061VJrAvI1y
G5TW+au3HOiBXJhSXFCvnAoX+MKw15BiIhuZiqdiG/jy/Qe36UGmsJGAGFTLk2/yYNa/h8dbz8qQ
rYecEFDZfEGyMkDjHWfAeD2Cy7eahyE3Epy2/wZ7WKIEu5Fz3OGIt09II7mkMZVdMdZD/jS+xxjM
5+nGrk2p53CA2ULOMCGt/2Za3pM1wEBZBajrHzeVIJ0RICOn8p/iv/Id8KW/0aYBC1ZJg2HMDggH
6jn/g25Pz0ZFaSNTiYRs+hCqVBWvU0ydtpyE4mNKQjDGqyuwScRW4PpZt7k/6v3oF0DUUSckqIv6
931QmW7O/QyCdXxHmBuY1/02OtqtQ5RxASOooQZbH5sqfhhUQFiX5dA1ik6eYYXGZ9vmP+9LhMnL
nHg6KlDCvIixGLZKg5sNpdgimFM+BLWUK58QJvSXxEcR03tS8Shb64U0A3hYOOQMowzeqnG8sr4X
q1mUa9cne74FI1DCcrt8VFeDHDFakL9a8881nenfNtrgRby+DZ+fst7zqcr7v65Mvo4+EugqZtL9
YHAT4EbsOqAhlbS8y9npcxBWzwuC6VD5cyf3wLKq57eUla3EpW1IvgSPccFLZXBTyPzaxgySoPTm
UhUZ+Ml1k/ohpIWXpBeK3id945CTLnXhcF7QNbi4ju6X8lZE6tH+0P6kYpWoXKHJhZ3ot/hx4KT8
sHIU7VSQctYuh8NYtI7S6dQsUGCYsvmBEoLRAP7Okj/J1OmWygwAsPwxPUB79biu2ZAkkcO3qseY
wi7sJZn3+6Asx/HV3lWzCqFJ4RkQLb8KRYmmVN/EyMrwlSipg1ILgNUTWOcM3QNeUcRhtgDz1kbT
tGMSdM1w61SN+I3dTwAv/yWm1+Dr+S+nwtXHgl9TY6wfqyHZN8HIXQQSTP+WEAz7EuWUXpE7xuRZ
GcB7hv0lhS/lXXKmA4kSKrnKhJoiypFXrrKQ1j7xJTeC6xum2sIhOH26HHKOjC4EvC1R8Ba8ECPx
eYTE1+y9dmlGrm6165G+qu1QlRzjQsMpN6wvVphVRH7yh2oyIp/xNW19j5mpzdM/Su0MJc2ssF4x
ipHQQ46yZYdE0tpRJVt39qvkGCjLoGE8ihc3h8mYFHuHGwdWDktMQwn/vK2YMWEQFWQR+vLX3UaE
jbxzG6ULlehVrfHSGitrhnB10G2YAH60l0jC0Wuy8syNi/IKWy0SyroDG1M/LxQA65vxCn8/+U9a
GZh2+yqBS4X9VIL+A6RLoWNhU/s7ZlBRncD71NjR8J4RF/0spD1gVItifKrbrYW9Nv16vW69qfNB
rFucNyfRcH2jVxH9+D4e+x2O5Uuo46BGWoWMTGgrOHvgQgyZdv1RR8G1Ni8xm1Ldt91uNJZrc1aK
imsakeqBCkln95xM4whK2NbJKwUQPZFg+NQm1ugADa1NbF0xY5o/vz65rPjGDs2XSFyTpUxlxt/r
ktsYk3hhI1tBPdpcPwq8/7BBsK7WAhIHe+bC3pN/Xo57JYpAL3Ga3ZZgN4qew+D6LCEwjmLS1Sev
1rq0WAo6kAMSxG2OXKg5vHAaknERfzvlz/jYz+X/NfeLtEK+4b3j+Mve9zjMXGp779BX2L4+TiIu
7xv8SHC9XaH35/P/9ZBFoQiEjMUpV5oEuuBRLohqalfzW/hl3AtzcNA3WpiSlGpXZdu/84i1UiRo
JlrpFbN6MEECt9Djczu8qHXd1T720Br856Q5ovpzyHM6jlrx3sX0Qiu1W8REgnozxJsAAbla75yV
+u0u6awlM8lQuCQX5eZAxCOCcJKoD5GpkyTrfPpFvmrVznrhgMVh0hvKg1sLuQch/xInGjXpMBpA
GiohuXcGsvl59/yBwpysIN8jKvaree68FkhiBvZtvf9k2uur5UHOj/Bq7g7AjOravBfcnZgDTSCQ
SL/VjX/odA3ebGcwOqAlP6RrVovGNdHO0tWFuHTpCJe12MhdjOo9TG1C8U22xgKiLcqH9cK65/DA
rIn1kqQLipclzd+Lw7QSTRSQ3HqzUTV6XHTDqucOse2PfwCgwvevxq3pQrpdV28Q4vCnKO8jIKlI
oC6F89BxHzyCPFErnJd7V8E5rDnbv0zxGvpGI2j74hKq2i5siZG+l+lVjaE9IanJu5RhumZkzbTu
AioIfaGWPmLzOsvdG23nsfTf13rW5xutZjrDzO6QlzL2HTjQrkni3yHgEta9CCsNRb6DNnr9sxvO
yKtBMTN5U3ftiC0DozaXJ9ud+sz3zMAE0dd+uc1Y3tBgsdlkc0e1xoxEb/H8OKKOQpo2pZ1UW/hC
7CmtQv5nHrPF7piZi0NF+pslNRXLC/6CSWQjy+6hCXOK6UKfarTzVcWTT8Zdm96COmDMgLN2okXy
y0/APOFfqg1vZFgnybcxnJmjd24elMkSB/zqEFU5UMMdaBV0jtUyRh3rrLmlLP3HqW37iob2wW9t
7Ly0YEaS0Fhkjs6JgwckmP5seJFbe5cq/qKmQXHC8CUCEk+V7rHgylFBGu5Bqid4tmsSvjOir7mP
EDsrBlogJikrkS5a1xtTlofg7ZQbie47kw1qz0tXs4awR7hB/fuqC8vEJiz9XYAijDxUxhw1t1Af
fBJrAU4PQ7Hc7SUk3oImXdM8h46e3IgpzekwhT5FyDsa7o7ygxNtIo+gWZI1SH52uxsaKHldqic5
k+TTIPbGZVu+EZHoaJN7cSYM5o+MOBQEd8mwTuze8BXZl21rQkW6k2oQ+E78LfZpKbkDnuinXQwo
nw2dVaGeM4b11OTwj4Wbf3d6c5EzD3e07pSGbwLD3JrDzV9Q5cIglPO1FCT4XQT6qzL/5d2qxs2d
axduBG1KAf9taFkSatxjICHCmPGpm7Iu1k2Q0vR4AK7QVoimAOEAcB+EBBgxInijTIFyYF4/qUA7
HxaCePWUnT1voXNwEPYEkZ7vzR9f2P9WSHTkaiOGpo6ZnFNbC/tRjmbrWUDiUmny9Naadqjv87BT
QLiTeW2XIM/tLa4kgVDWesrC6NyogGIXMhpTA7cMNPQAMgirDWzAI8LIAFD7PpEQoeOZH71QiAxF
ch80TpUNjcw6xK0mP1TrC60QTLthghvoiFBziR0QgoBr0M2P7xxRVQFBImXpLSb1ScgI90Talb0t
tArF6HoB5T0z9Swc4hAKUIe5c1J7OyeEklqRwrb/8D/nLp0Hf4T+ZKp2mMAoUbJQG7cmaCSf+Me2
lsuTyIkpIrkwcrPYZ587XiAct8lM92qEu0sPjRc7CHqw74pPmMIAG73apx7YNsNBTYoLmbS6XtWJ
kTURtcYAtJeozudtkqa0+qmT9qZ5503W6m26j+v+gBnMzJmOtc/lLqpvtuIvBVbQHqjHyPtfj1uz
upPz17psjle+FAnswhCN3PLjj0yt9Zsdql/jTHxwMHUppMwb100HP4MYpoIjeGYB5x4/60/b8d8B
Qa/7ZJ6tbTes6U60e12Y0KA9hlXdeU4W5+Q85cIWCOEGp2JJjEfuyjAa0A6Yg0sNhg004HqmzEq4
HYa+InRh/GMqret9NqdOQ/9c3zq63p6/NPHt5Ppa9prEV1up4yEy3Y6W3t5T9Hyzmgutdxw0n7Hj
oRRymvpqz0JvgL81dbMHlF0T047+L9jJ5ExWtwQEjyY32JvOqpAT5t/UPe6b5qegfOeKXoi86n73
R1VKkdIi1v3lt9a3Dyg5WrMwwISKlHIkBSfINgaymgwNPWwKjz/uBUX1eYsQNgpC/8AY6ambZAOO
9T7Y6acsVCS66SQJA0RA6kcRqFfZDpYOfm7SazaWRJCXtlcB3YaWP6Z6PYSqHvmX3TQgmfdRNpRw
oE0XY3HsC+BPzSGpOnmgTq9ZABsAAphvUhMPWBOVGgm144Ocy/t52xbpK5XVvvGdDxd22ScpCOXp
YxvjdEHvfJ5pD40l2VDS9//woPZaetWjZGX6L08B5AyNatGenhrONjqyqxmosoTU//mCfmtb3TXy
OlLaREDv/pj7dg2X8F4Fk8av77GaG7IohfzITjiLRRFAjSrs8Oq/8896ubf9hgt7NNKuByrHWK0u
IiqOGSv+ZUFLYuR6NbvYhpyZxsKOjNGYoSCY1YsOTNk/HEdXaKZ86MlzOtB1fCGxjI7UCTq/ujAW
Vd4RDcC8fSX7dadJrNT2DQm/MnrckKHOKAWzciUTqXVwhkawbJeh7mSDNy9V+c6/hf9ZDQYSAOsK
ZR1dgdl6pRvYOpIwbZD9SC67plL1pjZTTdFFrbJdPLDqYIrUrwCDiFLH7XHVX21xbylPX3F56ltF
1VcM1RWa9Bls34NVIUlfqNCGvfAJ6jA8p6lTl0+F1h0HXW6ooAPpSO2/6TUffH53gbWJwZjI4zPW
mLnT6myzM+cF8MjH2TmX5+MVlSnFEQ/GROqPooqyn6HRlu+NMFb7or/uhH+Py3xNH8IAJzixBdCI
0apRd6xfoS4gJVmEcFY70vI43MrmIqqTDoQnovUmGRIRft+7Rlh3eg9HvB/dUGe/OD5qhmxt2W6i
fDSoHgf5GQm8rgYJDggprKukedzGpn+unQ+i9rb1tfz9xF9WQ3pQ+REEn7MVsVxE+wf14MWCWj77
LAJsQsG1LGzbmwlbbS2XdEKFAcVhQCFnut8jMX52ZRoVdvj+3zbEjjFWEKR4dCH98JiwySOwKq60
TlyyBY0UxQLy4P2uONkGhY1DWXyvB91nBIQ/GQjqIt/qxd6Mn7Dj2xdsASidfAaYDzEApvk44wpB
jesMsT3Bl2JlO1FZg8RpB0Ij3r5I7VnmbiBk91aXQTIO+mde4C7U5KNtILefYLi+1xFZSR/SIZF+
2v33FDYtrSPG2atA551CN+vQhyiDUOKUavt5a3PlN7yBHqA6XeJqDN4Wjy4G0wNsB9s5PZ8wzUKi
mTEE35TdMe6nBAjwiLZWk89o38U5tbTsDLL1ev4s8Hkn4CuRdM3WN91rgqH6ugnvXDnF82hk/kd5
EXAj9hyMFSWbDSPjF37WgmrKwsTbFtWAhL8K68JsPs/6qhD+kfVx2ovGKyM9Pf+hUlMqbDPBtgw/
71PkH1zpLDIz4ahRSTfhI/z1/eDYFjnXiEtc+V+pyUos3bwEXpdFgZt1Zld6DFh1ny55fxPAx9JL
++aNEkcgQASPAHpfXI0SlnL2f7VGD87Si7+gVmP8VoNArAbG8WbUKqjNfAD9fh5gkLckuUxT1nxA
qLv5kKFSduchDVfVyRHTx3ZKEK5pX6Jgl170ZdVV/BZB6HMhVnutr/JAAlYvyjSccnGJTS4piTdP
HBUTQPXxs22pCQ4/urOp42DiOJBVvPqD0yctEX5lglPDv/M0P/ofbDIq3iwuOVMrJakCcMDV4QL0
Y497DnG7l62hgEePWx16b6GHbVKoFvBY0M6lNd13vdC1ltm/IvQUSsoBGuG2SbyjhosqjaLVX//t
Trv3EbVEnaEJ2t7mIXUt6abNrPGgm1FAiDaWccoz9h158xwqRk/E7jcYYohuFJ/jN08/JpVrhJcN
HbD4nlhBScRj6ivOKxevkg7Vw0bMT9RHTFPpsPwn8kbLg+z4wl9gw38cMfGgML8RvJEnUXlbKzH7
xJL5nClRyp2Y2O6W5gJUwmc3pbkeiL04RWDOWZ3gGur7a3haJVT8SlgAPHmil0jgT8HcN+EQX/Jh
Z/ZWCaUYmo1Wp7MwSvzLGyY0wPmYBweQP+ZxRjxkh10dAq47yzFDJP6nYvfx0/uzdFck5xsI0JA1
z+y+WfpY1Z7H5goabhxq4vh6EINJXw12QVc5bismC3mazORpgBxGptKnXhu5WzBCqL6Sq4wIgsPt
zcdUut3K7M4jXUe+qCnTaG/ygbZp642ASGPElrphsEBECuTonK+sn0qlbD7ihoE1W+KFWcQ06pmW
yG0eq0KNBP3770cP0EYQaU6D1aPqyDs3HbR04SpfFJNJZNVE36xRDQHY00+Eq94USQg0VETh+f6n
dKD52USdmSSflvJfVynf+VxEGpy+TJ4lWU+1fGV2HQpFS/ppju6eP6XQfTjyyuSqPozW1c6FZGvK
c2RjmvU3b5GYcY0CuYc2i9iQLLwSBqI3hafm9UVUDCzRmEvYZkER+ujg2SHeSBDXWZ49Z4JtyLj3
f0IMNls3ib/tDZSY/eIXS/2iuJIYBY9sa/OObMqQHGhF1oP2MENqE+PYvnCHfBjm1+ewDeJA5SpU
h5Yef4lbdeDPbIDwFE4UAyj/qet6s3Rmapgu4KvR8+QpLvFF7oz8Fv+jMLaRrnNEJ/EMaepXjJLC
3j8QCpVy2slso9ukao5kDobVvLtNx5kb35E0lV1IXA+PpiSvepdrLJalqoUV5AaLPHgz2NebXAMb
tlcdF/wGu5pd4WNweLH/OYdf3L2JcSZT7B7qjUf7WomuW7cz83a2jOiJzp7bW/P3FOpxwaS+RWr+
xaXcB6qaduzcuAlQQAwLsFdpDubkLJ7sN6Gr67kb8tSHEZ5EbjLSkHjLzyq7WxWkGmJh7+QmeuIz
QWzz7T0lm8Oh9r/QO1N0bo4KkeucP1tVyvjCeTWOWY9IoJXXrry48iD7C/t2gHjy6Ks18ehowFAI
72QeHWqPG/qnrUK/ogEUxr4XF9F0KCMpWkKZfSZ97iedsvMOEfY61O63jqqwTODjMRfH7QYzBKZ+
8NMeLbOtDUERDBRPEo3+yhnULP1E9uGAv21IK4cXVVQYdYus3DMr3RV6gyAgxd6oHaCgwJ+SUek5
ztPqxg/FeOeIv5YBTkJsYXOmklffe11U6Tqm6d022P5VDoa9zFcjGFfOHY69FSTFHmFcOIp/WeC8
O9hEl8in5sC/jQx3LelxhAQrMrJQYmoY2PnhuQGCjVOY5GOyU1IfaF+nPy+2LLB4DDUxlExD/C+k
KD0wG8SgbvYD4nBulTjjf2rCZAyP1MUPpCdUxGc49kJB112M8o4DUaP6KVNy1S+jOPUSOZhpW3Pl
jbnV6iD2ONGDX2dTeWULVLSuhBloQnAf9uBb2Vjxr4Vmn75hnEhkXn14fxBcRdz8i4/4hYOhe+Up
dvp0M4jsRxgQwbCuMHn/plb+3qCeDjkOCIws+gO/5k860UJ3iVK/37BpQvYRYziFmZ2YKP46ypsw
o4iY2PhOYKOuHPV2luz01/6dogYtrkc6x41HbrDQm2/1t26G2XaMu6qurc2Sn+F8BpcYGi32rr4v
hgD0KJ+hcaY/Ui8b719lV3lS90TFxfUnjlSnsn25sq41QpzVT2t+iyDM3Ifx9OdoaN85eOjm4mvM
eKfkIh8A+KSBXZB+ojyemPxK0NkQrk6tcE+ZnkGypP2faK6vSfNzWHbuuhn/HUUTii82ti7kKmC6
vg+18NVLDcCI49xmq6885WZ466vwQgm8PIyv8SCsvkFZI/ZmI+k03gJWZTDqWp3MFnBQhYVDb/yY
wpNzLtDdOqYNSTR9OXv+VVYM0aU7y8x6OQMb3yngu4uO3nSx0kvs2mxiCLTg7pU6PQPy7oH4Lk+9
qAiNHE5qoGPfmsMtyZoN1Kzf/naneAc9PunDuiuTFjuik4g+GLo01UuaqZdCmcAviyru6NKr9Ly4
SVeSYxIeun07KQM9AqlJD+T/CeYARf7/UHG7Aze2p3bomyyMHIS+b2bJs6gYLPuoQXVzxOYkSYqN
xx/hdTPNbYwBvnfpdryMxWjfXpFvuS+BES7BelOA91TWhKvaQW8PWV5Xud66DazbiT86f5j8Zb42
LOYavtOlgH9EoI4sZIpSV2LEsi+e60fqnTZuaDUo1ji1I0giRDXO+lx5xWTVR5Nbd8yOYLKBqJLc
IVPm8P4GG5XC4o3cPFpLr+QmUFb52dBVQYT/GzW6d1uDwv7KrNMYIDWiVEQ/p70z7SUGunhScSdv
Qsegu9JLtu3DxbjBUTbVB6o8k5YORx41ll4pXZmEb/KF4FlWBDNJkWuf4s+vjDcuew5Xk1vgEFz+
+Lfghsz458edv5TuNJpsiJ0AXZ4KHlkn9hGyhoxNztK5q47u7ATSWHNsmegv+gn6TaXU/bQui2Qj
LWNmAnCrcH3Rtgz/6Aj3GQ8o5V3W/fD0T+nldzCfSgeJ9mpbLdlqw3dJ8vECCov9Wb9rkg8NQoYN
3xonx1d2JOX/fGVGCnxKTFwV7xtxFoyw7b1nzuekxm5KqQxDr0ou68c3dU/h2IDXQOvCnspc0/PI
ddsHWeH0N3RRxvGc/LbJdbJ7HFK//lnb32bnwEpFE4ceZ3JSBGRCz5G3eael4bOn3h3aELcSoeOz
147ZjYolzSrBTzGPAZ3AruI0Lp8RER3O72ryGouZh1PDahpO1Mv5/8wtsEEY4XbbsugkEvPhsyAL
5qgtTnmx+dcNkSQJ+8PESC50ZoFJ2lyXdGtUBXRE3ATGv6/8MzYB/61zrk4nE1hCOaRQCgNXPjdf
oFAPzi6cL+/RTSexXg3UiGZGUNzMPGUij6ml771XJomDoj3nwpJ9U1JHcznKCVF5LeM3nTPV0iPW
1R7q6RiV6tXen7OXNqzMGBJ0di5g5kzZfvcBLrx32J57LXE4AL7swAMQ/Jk2p/CAbGj2XXh00KxC
WnDCQbYMrIz20A4l2mg+fOqshvcbezvmXopwDFYwZcfRGZcDv8mPqx+ungFbN4fmDOCRKsag/oYI
6ANkQOXlzacNSUG2/tUbUJnXL/VSVgSIsxW3CN6VaXqbrkyiPBpas4PtZmC0b46efLVp3grfppuK
pL2FBRCW/bEDE2BXBmxnCwFssXonjx8CXasXCFtp7Id2PUnLTKMd70wZEUKv4bsPXXsebB4G160X
D/hQLsf5XeueTCXv5vuqG6CtcG69Cyy4KI17Qi6rqJnAVcDDKNrqiQEqhestfF5uT+q/PqBaSyBa
5+ADhH0r7uj8EjYOe6TyjVuFZhyF/C+ji306ej1cPw6aBk3BK9CaDHIhkk2kBlQU9hpzZLu4H9fD
h4h3FPZ4CISqJQ54zEGOkP4aqQBjn+QDAow1mhGobnUrf7HXozOexzqfLA4+q8EAxhSDQsmaHnGI
RARZwCazFmIdWBSaKOnddTjuEvMl13qb3g3DtcjDBrGx+7pEG+mqMwZBtKZfKG46LJ0IfFvXIOb5
9tu0sXznWl8zNDSG1jpNCAJXWYF9a3Tkj3tYKKAapmRE85mKjQkGBJwYPF5cXyp45iJpk3lIDeFJ
HzYHDlu92OD3f+58AlUN888SuoFKVYxzL9Qp9NWX2RQSBk+wAxTGvmY+MwEIz+JR8RCdqrXOgrFs
692K5205FicQHjZvsMyXKZtJdERnP4tj8WLwCttCxgj5wY84GobVUGdrDWn8EckUUTe/eeRCb2GN
84bYPK6Cwzs48SmXcuuiGiOfGOBD47yCQMsxd+cUpfd1gGcDCBvCKPEx8P2bCC/m2Ea+4TljsN9B
xXO1h46l1Za50XimI90fLxHyIAMSzoFJ8mb4tV2wUCxvkIou9E/iILfjDa5ynzHEXjgaejzojYeX
AtgAWXMPEXU59B6Ox2kLN1cfm26Kgg9MY8Z8rIGCKMnFqV9YqCF4GiilpItU099bxJjkscL3cRX3
wvULnsNGOrRwb5CYNuavTo68TxF/aEdiP4hYeo3zJZi1Rvd5hyO3zQA6IUZedFlDdqPOs0Q7mIB6
OY5xg2kXWtVQkNR2Kc4RLYfdqSLruH2I1nF3IHDOj3mQwF56awAc4+gKpNSjd17bS+a3zuo6waQO
p4yzMv/C5JxGpOjlpTXoMFz1dXfYYDZYz2KQjHZY6h4OGytuD0jG9J/zZqZsWTNX035p1H8ouOTY
PAe9qggBDABT5G2mBRGdk/jrR5T43K93aQpcJXhFAbbpUkp6fxLiS2wq+R3hiiuEJ1bT7XtBJfqJ
0naQjTrh4nLqeO/ZvDvmuuPtcbHy9yXAiVjnQ/N/WA9M1wCuLwogaZNx3r8hR6yaW+5AD7vrCVvR
1iOFAIM4GCZFiwGAZAOVMp3BI89O5l/Y5OIRQj6lB18Smxbbd8hd6stoP52qh0PowiMhBCH7UHON
I729l3Pz9DrJv0q8FwEhJGf1MFSNtPuW9oTYU4naEmJmrBZyQprYp2FqUeGYcSg7i58TSFUKBldm
xSrP0hluyLVUFRj2iIPZu+8fZRuy/1mGwlIAaJmKhd6HGGMCOwkAKGiuqmMSY9VFe+b7Z4pUXapj
5Mcdzl4BOcTHBtpVczzJ+2o1WeSVq+X9vMBENMKAf1JLs7votYICnjQucT2KyoAADVD1f471poyw
C7v9EpT0eiVFn17jPmIdmnX22kCvf5l2U5yu/6bi0YeF+NUvsyAid7TKMd2zJLd5IalyXG9jGnf3
YFXneKnTBK245hdj7gHPHsq5+tgbYfisI7cjDArru2fE94EcSQ4Gzy4y8hgxlmB/cT/hcANFUCsb
byJapCZAZyhNM1ppZECLXwAArJKCDG6+FGUYDKOMyfDmWk0va6s7zNw996Wf6C/aa5H7BXLEwky5
1NamQrLjg75A1MCZBJrm6HNVo5M8/97WxhpK+o5U0vNJYxTLFsLucNLss6Mzi4q3Qxhh0TwpF05x
lbSbdH/JyPfnNa6FzyDl5AV4zlMf29mm9SophLFxkG5TT+yGoxz4iXLY6PwXOST+F7t1xaCC3hJS
4MOwZ0lUihqVuEWfIzi+pU8Lr+qA0xIt0WmQ7IzLSxV0V8AXqqjXUj+z+dAmC0Jo5LNcU6uhubxj
HadR00hOOMTxrRrJFgXNFoxerYFeEz3lcbXTN4sdkzKnlPHtI/fQdd8HabLQB9E2Pz2LwC1AoNzY
PXc5ndRf0yGNCNM0m9zEoRmliNlY0s6GIThpUzZuXwpRpV0FLcXjscfk1H5LKE1j0WjFm8+6TVqH
xrq/rOOsvlQ5WxXFlFc5zO7BA7YI7eB93jzX7VTIOvjZ5f0kkD6Dqty8tNARK4AkhF+x2JLWHYCl
CQkanyX4QFrxkhWScWUuCWCpcpYAznMl4h27jClrQtNWtOMDeYmFeHUDbZ9SzKehTSjcf3lPvibQ
pxMkVbaXhR/AuwoSOTMSVRKCdq4ueozoSMAQoF87T2LdWbwiP0awBPge8BQ05fF0UGi7homxdvNS
tbT48kXUl/DbuzfFTQBLB7mMhD06kjjbdW5D/x6hSPV3Rb4Ngt9Q8C+czA+wRGLn5sj8zz/ubawz
TABWE0k+33lTfIgxUqveZ4yS54VevF4d1ZI4VK9dSaMBjSim/D3gtD4x2FiT0rauZqa1J+NgwVcC
mqMY4UrTUjJfwF8wJU306J/dIpEa6AY/abwHT/z7X5porSlDbf2Yhc4zYFEr0m8LcCQT8gDZNYLq
+Tdmkc20jNjBIrf1FW5csvPW0FhkAc+w5qCFywAX2p7Jz803pQGrLOpUHS0zJpi+u4XRW1c457V8
pt18gcD4zIxhFwL6MvXvUguUCzNeafNMc8JGgUTtGG3QDT53s+wGGtU8qgAHXSSkZIOPLvyg1HXo
XHEi3SSW4eFCb6XuvbP3dfz9/rjqnaN3IUYHKZmyyVLp8/agPUaQhOk3CLZcKv81EacIacYXvosa
9UXnnPCA3iX77fOiruR84m05FGl5QXZ3/aLVSJhwq3lZLzLj6x3eEgVE9WlBlOOe5kOXBAIWhCyH
dlie94jxPaNY7W0VrQ6enCUaAqjS+SZx6hQz10MARppLEDF89Dn8Xk9EIiNJqNw6zn4HzN5nJRzy
b29fVOgfCw3CWeDlKU6HVFpwJlkg6xh7qWg1OBiTbEdNXIKHb6qtIiq9WVpWMtQB3S+mVQ4N6290
LKa7PIa6EQ29Bowx5/GyabSihIX6ktU83MVCGLX6ofHdlpDa0/s83nl77VS4bS/IJChC0MG7xAtF
QdwCL0ZkPn7BEphRGduptZqN0Y1oyFNmAawrJWWfUqYvaxc54J5EX7cSpAR2H4GYJLvZgxUJ66wc
l44Sww5mN3EFn8RH1d0C0Opd1qTGHmQRMInUEHKjNmFc01L9zt7DaD1eOnS7VR9oSdNqqT012nrH
+QRD0SEVXTZXz6gfNWyxIUhUufDlOka1Tbv/3gA1EhZKBUrul2YzH2c3WbTIKOhdLezzLD7PuOOC
34K7ASKMtopjXzBM7PDmjB6Nw+zZ/y1xjKe8OYtzWFIch9eSxdE7WeEZjuZMjSdarJKfcstVElFn
NvLuJF241qUFu9krJ1Rfgf/fi24OLQ3jx5qd4tBHFOflnOo4NoJMUvATuf9twa5ZBbhFnk56sAJ2
4n18Q4zXm7ZskPGhDSF9RcawB3fNO83Ip9lhOklRwYJd4Afvd5p+P3mWF+tYRA/4PxldlNl6HJTp
umJy/znldOaYenKrhMetvTA2CqDWglXIBcWD2awABCGqJ1ZWCV9OkHONQ30rb8W+5NpYMPcO8OIO
vluR+/juu7K0BmXezQbFvZjK4m+2VV6i3E4ZP7R1RpEcZ/Q2nt+ieWo6JzWB6RkYXzpCxhamnHLD
eu1PhO+UxcpOv4/ADB6JGIS1iAU/BArCyD7PiUW4vRpW5eD5RsApVxQu0bJXHnaL8tHtwcJjlt/Z
j7mwhlThbS1KP9E/sHFbLrgUjCfkaN/b2Q6JcyplL+5cabwqWEEgzKb3xdyndbvnssLSwKapz+/5
aGXGV/EJzmQbWDZAvRk8RAuNRlzPdL+qdJI3HHVq8wdG6JeTa2rz5rmCIYpmR6RDAbxtoHBQYrDV
kBwyPtuvM3227Vg2e8FxLzO/hv68oCATrPGJ6MJnsrlXu6j5wsjruoT84+3pjIa7RNs5Hw89lEBR
HuEsJRcjkXX6JKZS2y+B08lTBlc2dxFjWx0rWOLY+Cvy3dMwrd3lYBP6DeagIjyvIsVPwlXp5sTO
0S97S/tz1m4PDtrLPjHVaPBzfaVfs+hRQ9ZSdDGI8hWYWKnl+4Qms1RHkFRcEAsKrW9mXDZiz8c2
hjxMS0VQW95ccOrNcsLR02oVI57czgpkMFKgDrRiLtoqx0w5W6b+UiZUzfM9+LmU4aH/83xWTkwW
ZKh6qVqQVDO6lju+XJZl9C1cMphNLInu1FpNTnyGlrSqvcv+9WcL6uRikVRYhvzju8ZTJ5kJsp0v
soWU1ww3VwBrrQvFETyFbZHx9j8XuMDCKayyf+F9oBRLZs7UL1leL6++z9zuYXj0L07uv5ArhwJS
xna2Tc7Yv0rXZRqGNvdYvXqwx0aQ0kMrivyUUuRjwHJGHueVT7cWjStYuUiNv/hMpEXDA0qpCxCx
FZkuW5MKbxEwSsyEGMKYTVtC3yfnyHkjIt0v2I7E6z3CMvQcSs0lUY8GruwSHWZypKuIu/gsQzAa
uhPzgBzB6T3tHoXQ1o+23aB7Q3JyU0wN4psjSuK5MTjge1n/pw5Dj/a9JEJsZLzTKm5y2CVs2DW+
U1Syo3vkeSy+4ON4BkxGmrbO3QRPL/gl8aKFFruyTCONkMDEmOYZQwEgOaPuiAsPppk1Q1GmbWUl
MACMR5Ar4s/rNK14dBj75QclLTL5Qxq5JyaDaTTPraghrzBO0ULyg3Nr8luLtPtGLO7xBea4bCrn
2UEG8mSKlQ2z0WSXn+CEyBftGCppht5uzHZ9EqkJyGwf0Aiu4osb+6CUVT0UghkW404kawBtiAe6
nZKaHoT1E0ZXYnNK9bmV7eoxxb3jshOp95JMT3UhBSZQz4PEAZGdpO7F/tfL/iRw8fsMb4DJEnHx
gHmzJTZ3EwJN6gekwSSYKA+zO6je3c3gp3M3P1ajbTK9rU51pGTE4VW0Bz5EDvVcQmDXDAYJ6ge6
rtVRlzsEozwhjaQ78ZIq2Rp2XEx9UOHFuOgKDJO/KDjXqY23bGF6Ee3fwYcVQM+LY7nSB0cA58ki
1rahuxAPH8lJ7KnhRfmxJGY7e4hD/KRMOnyxjzOZK7qAH1OO77bmZ3U4TAqCLbuzG3Myqg93f/gO
Zj+RyaAvyz3zDEdo8zBLkR6K5ztxLd+xQgg0WDQpXExeg+Z826zfgiMGid1eK8f5BM9aesDyjpTa
uTBX03qFQ54i4tv1luaJRN9WmMGLcadHtv9gRM9kjn0FIlZFUyPluS/Me2uCsmdu4Yj10QxoJReY
6a6WI8u4tCqFjrHVaOmh1HFcPYLE197bBVGFMIE8fsGR9ahOR1zEm/kTnkxB7xYeLxm2nxTWz3hX
yUdDWPzyLQDC9ERL2Mk1MR2uQU281e4i8XfXmEbgv6yZaeWfyPN0Iz5OZEg5WD9mHipRCQwBww/A
Uv1xpvi9jodBxgpQppAy9F7DOsYKJgA5nvL4w/bP48wZGDLCSpwjzxjEC3EcLFmX595r38Cm3IgQ
OacCOMVhQCLpSDSC1eXnzTv+8SAOArEd2avPXToeM9DgTB+Tw3wyTDfNPyW3aVMZtxnhmdFr3XRn
OjZtQc52Q6ZulPEv1FRsDvEV6hUNr9iSXayLpae4FMPW6j3feYajqfttHruPFrcyvx2m662LNI5J
nrWVBpsrhtRd2oaPFzdbZm/WzFrfFhYAtDMqKKJIkSHvBq/9Fa8A6rwJ/zB8mMB7TrQAewifBSZg
zs8qGJomXtq3CW29bpV3bpVJww5tyKKmfAz896EjH/62ams0QWrgqPpKJZ+KCw003ZkPefNy8E2B
duokv6nEUWZRLjqvdo3JAsrEtQ4bkHTIArGKnfA9e6p+S+z4we/S0VbJJmqONIPi5QhkCnmW8tTg
LeWSF7aYwebBjHaKENsizKyBD8/RSmjalUql2hWozQ9pusyVO/nCWqCRz9yElC3Xs5CkxAY2lxg1
bODvzozpgfOfWE6on/Zm3PIsPvOZiUgVOeeuARK4nkpJYwp5ameMe0+/rCmo0GUaYn+Gw6VBWU36
gKaxI0XHKBpqHm01BoOj9oYhLi9Ojjim3lMW++HrPDHWLd48B7my7O0c34Ozty8jVbIggT5B5v0+
Ogg5XSL6FpUD2iN1aun0HAKbl1uN+lO6ZkaVcRtgms3EYaX9vSd1ZvzmcSAlPW7Q2fYBqgcYeDTb
QK2AVuDU7hLiLGCCAAJ4sI7TwRfcMDpuCz6bq2oq3vfh7FzBhcXzbYAG0FhnX8mItvQhwK4nrmWn
j8sw327buPuXc/7hvPWriq+usLG6jlxUlAkpDB66OAYwIvJH/pA5mDZk6g9DktkSTFraGfDujtto
hTNU+XIzJCLxXUSAXMNAw/zVJa17exNGVUt6YqgYmdmBdt+ZwHCu6Lp8d/G2qHudCi2VVyVvub1M
3vy/e1phA2UCvLf/yD/OwlDsOj7uNP0ImER7rX4OIfVU84ZGi7m32PJTRl+b8CQHTtwrFB6wC3pf
EyMP0qm7Bpr+wGPdirnSXnPfGLtt5hjAuJIxx8TrgAwgYa6ZrKwHplAswjCvkS+Oao25E0+kps7z
1Gg7Zisl07ozFQmA5AEDIRbYVcZlMK8rlcr1rgAp4PtZC+iWTj3f0YSzs2Sz5miJE2EVIdkOcni1
yB0ttqHm7ActJc/FmQxeCZD6AReHvV5hrjo2qN2bVsjOYTF/f22O5JExBRM4yHl+EkkcyW83SFBO
ZkfS5IwRMgO46w3nLzwpxYo/HgEhOj1Q2pCf9gwBJP8XPrMj4H7Au/9lGAGbirphsDFLPXT/geyA
0BROqdm7mY+Pt9/8NOUP0eLO4upIVxN9FE5BTApAe8Js7yyPX7u3AUnjlG/xfniRxTYevPwhn4if
RPgGbYidwQnV3aCEU1R6iEqMT+fYxgmdJVy9XF5SmuClBH81/1MY/AxCcOoSy9IwinLiSDU885GK
ngIL3Ir52FMNAygeOo7uU0hGti9bRqNAWSLNRZCldEnOnpGjPtyMDX5IZQMAcvSrP9MHiHRw07nC
KZj9AjDlU8/EJ5wjgwvCtI+qb6ARJK9CuNnQoq39deS5c1ArKWXL7SwFeBb5Q/LnFTJ8JC0B/u9J
VlSesHlHBcWXRMHlZuZgR3pfWvNCFEYZV0wTtRAkpxl7kISLdtoyH19SCWdiG/mNTeeZNU242J2c
gCWe1liapP3SmtTLgA75dJpgAdQwNqXw3pyDUrsWlIWRYu6Nt7PEKPz6mHjJsf/KQz2KVNEzgiTT
l+Kqkr2aFfxmy20DmJ6qLM+lS5NQy5dU4WPqLoI3sExzg923+1RE1qMn0giKWNRlLVOND9mGts2+
6DbihbDi5RVLkR9wZGseVtVVN8HOE/r45+4fCpzmBKZq6OrptkRJ3TCwi1bmgezizhOUjS5iRXJV
YxOpP93gj1tp+YOcZfN+gJe3e7Js+hM+YUOHFhnzlKIFfh7MrIu3+vOV4CHH1aoFbIihri27T5gT
tUTeGgh5Um9LYfvK52nlEa34ttpwgtr5C4E9cjvqrmlBGS+UE+xf8c3KhUmRLilROR/p1EmoEVO1
9R5FcNrvZbGfqVS47wXrx+ogZFHJ04mz9TH0z2pZUyEdsRHhLnDPwHLDOlUugSiMR+uFD4TZorBZ
rTKVZ95XaeoiHXqp4WVCuRQq0Lyv+DH1aWWDJ1/RGmwUrzReQv9XbqjRnhNhbYAn/mQFOwWBUeor
G+mFUbJF+oMdatNUegWPfE+t3Lcm7aq0ni3k3Yr2M/i0+IpvrNdublpfNf+1wkj4mNQqlhMiIDUg
XG/E6V2g/0tw4yb3TRF9U9UkGRbN88Gvd631oSkRPOqHRsdopuuwj6AOWohba2CNnTgiQvVCe2NC
sqp1XCWF61sbTtF4rPjj/a3a4s8zkBYxEWSfFH7qjjdlZGneSAi5eVsC/TZQhjD/HpS4WrZf5vZA
WTtlry+yKU6llL3QLFWDw/SlDvTibCfGoYSLcy8RzxcF5r8MsJw7zaB4lEDDNekQnIgflC5P75Lh
BkV4CYo1XwR9lLxg9nIozmVnTT60IMNIHsW6kyCDy69YNrqOzaSXMWcHe/slCal0nPoViffQaZcZ
DPLYaZWjcq3vUj4QEIv8foASJXIbUfBWuJ7lFLDK+dGYpi9eX89sk7ydATwHMwzhla0GBt8rRAYx
oTU2pEyfhL0xrRE4qGTpqBfEpHGHm943xypTzk6xdxLVXmrheQFcvgTRb1CTLsRUal7TkrXgyYjK
kVwEi6G8Pa3Fb1uWVS7BtWVQZpYEmOASBwleicIGBCloevVRPDuNK0d3CiUUg8y/+wICoLO8nMhV
BFxoFVfofQiLGEGkJ8oCJPG+KCOrOzYsDk37ziAoU3LQBub90D3GKSuxEqpWfzYxPR7gIqnkV4pL
/eZOVZvP6rMY7KnoGR4fdQwgvOeLJv61kpRHlN1FwwFfNMYgLjIdblXL/78gOCGHhcahri65e8tn
OvcZA+d/lfA9gI4ADp4R2hSWVC5MxOHL9oVTC2Gs4j5vLuYbWE+kKWyzoWc38y0lY/HvOzk2/udN
trZa7Zz3nt74xBFOVpushW00lJ/2Qr/ZGQnrqCNmloFMS6BN2FFZPaIT+VFgBhgXPgUDj6VneQEg
+TtmNFX8pSm8KX0fl6jhU7NbWFECozSSJZ3wiAP58HCMmYiGEQpCpOZ+UbVesoGzTJqWV7uatsuJ
oK1c6KWCHWascGjvEGrfqlLi/xyRMW1PYZXi30usLobIf5J3gACowEtddTlOVvdTygO3kce5z+pk
/NvkQiAdZzcelai41ymEiGsDlQCwGuqfRK78Jhi1qzuJzdSGb8UYmE1DftCpC0J4ldq907Wpo5Tr
bsjbeqGQBGKn1c2GCDDs889jRp/invSiTV4V1Vq+3lEItyOJh32E8XG3arO2+SS9Fn417wafgj1+
T8SWaqgwFpmFF4cFQoEw++AryzF17ziBEAkq+WJ888St67EVEQg4AOvS51c/Aw6HqMx8U8+34FYu
UZTu15dUHHdWI3t/knQEFkLbBmj2xTquXRcvtQobqnQoenreeqKqcZ8XpXRaeFO6lAGHbb8qNeja
QkrFLm2pW+xm2XBxaNzuX1hlfoYuj7kSHWu5vdETaFUXV6K+yAdprgJhP4Bucp2exnHZI+JdhpgN
Nrin+eHxExQIcT9jOI6VytmuFUc74epI8B7a/vRC8I9IwKKkLw+m3HK34uIrdGuDrpua/kbC2Mw1
1K97xYFEmYwsoeTGWwdcK++1GIWbLoRo0hcJDwTroD3S6jQbFcGM6oKN7g6dvwnKMswPMCcCe0pd
/Wa3avAde7oPfWqqUCW4GkvL3Y0tLgwQFpTCf01NFrTv/kiUaaq7d5XanN3PisfYHgnhIpJJ6OD1
nXSa3PqkQ40t/BOa3dbkaZfuuZpDqc5/ATHm5odzys3JWzmZ8MyX/m165MSBZ/SX+CQG1LFKtJO2
MwZvr6GeXeImFDndZFveRJK6H/MoCg/vYIGVR6rO8QM4sZIigJyeMm4sBDX8QWJngvxgN+aIJvtX
XfaAtBVO5GM6frc0fnlQ/3+AbrxOBF1f/jN8FPWzqe+z+5ORBJnE28ZPCfkgn0oYHSleSz6KlGZq
6C6sU9psyLmtebMVu/iBK1MpN9ICwDHgxq6mPjetp3ZPykMdUPmwu40cqUCGBOi5UxnxiA7e0GmO
pbX+1Swtkb3TzqmA/vrMJRqK7+VLZ6xKRCaXRxFVAueK389K6sr/UJdkVT6taSBGO7gIu36incHs
D1rmVeswfTmA2PvF6e9/Zwdk4vUGwQgNxW97NplhbqsbJBIF3/DxFg846krGfYo6iLLh2/McZsbt
jWrxCgRo0wRfnEwBl1/VTVBz+wyeMlMzTcARhCcFHEnJAi7r8fcaaU1NVtZEtuBdUHSzsaGB38Z5
NXhsVuCfYUqoOkseXztSfbJ38BnyKmQs52ED2RJpdvJeEKxaWpJ3RI3aN0UR3Y1bT/g9wAzEkdvh
5chR3HAqk8pxY+Ot5v7i7pcebmjc3EL4hLBuEloxYam76EF23HOdS2iOcsgv1ce0X3UeEeY/8OoK
z1s210XYFr5n6om45lz52XQBksBzdCqVjWH3vzBNXqOaEOWH0ajXX2aXW+TejdnIRGU5VGwEP/Ot
ZrW2vb7An9hcxFbLSuNUKegRYCyEvSL7Y4T+P5izD6GqM84LGM04cnGdtyI0ksxKsP8fRQe4ByO7
zcX7vPH41PcY0csuFVg/D1bKGWTjUbIH4Wz7ARnKgxOj4wtmiarJ2UvMDKig/6ntk8cjoUJnM/oP
jHOwIQeBMshEfnUvSzXSLZPrdyQC03yT5qc2QGRXD62hqYdrNZc1EdbvNvi7jlbhMJWOoPs9jhPh
MQ7dm1kPupeYtpIPw76j/xapdVKn4sY+ZhfCFRAVTsMwlFVZpwMSMqVu/6qeyA/wfbFRi1c3OoRW
iJyLgXlp5FLr0GP3JeDOkCjncUdpFy3Oj6zTtuzJ9IvcWXSjqnFRpkrxqEBiYCcFW1Rz+QGEAe65
f15hmUZ2mTsT5jkS7NO2NY7DZJ/W82i8AYpI7s152IRZH+3S74Nf+Hia/l47Ay31z/4+eKwarRKg
D55gomZmwI8oMQzVNIDlZGI3HUC+yw/fnL2YDEaroswQHjh5gmmIBjwJI+dFe43WMiFjnrxdUCYx
xQA2qzLQMvqDnHoPKZGvA/n4bnKmnxAlk5PpvxxqpIEOdvt79tYxBh+Q8XNxk5Pi3E4MrhFNBzKX
lI1wsqTyBX6RahZOlqqWoSqJR2aydTNZRSLDHypysQCXi6OF24gEIbnagQAfr8jNu3FSK4MctUa2
sVAkU3V/90G816WHgBEPyDTBxeKdWwOD+qrOc/hH1YlSh9kII62QIpoUvpKMMob9as1FAhv0Qes3
4XTXg4csAdxLxNzh0wN54dLhOklFyuL9GH381FODjBF8g9sIvSLTvu332Ezj4YesEBFTQ37vcuCb
O7iwNVSesgYR5H9VGRQcNpXy/IuwSoM9ZQatFGELdnX2axv6ZSNnZ5e1PyBHuY5rEZKale9k1F0H
qUfghf1aPyxKGfSsXioknMjSfDv6mBHcQdB0H78f2kI2Oz4SPJkXiExBghET6ZWLNXMo038d4s0F
BoRZSFeFNeNzdqZFJbETAaUL/OJZpHpg7XeLV2bYXiH0jinTJsoe/FMqCRCzPMVGWyritIeZYKK0
zg/6PGREcYw0upP3jZhB15i1L9uevNzTCkPbKk7B7Wsj3sLYxmGk93JI9MwDuekGJw5vZKL1KPkf
eo7Hh4BGe4lqS7TRgTV+1sBeDoO0W8UFdhEpCoiRInNnNC1miRl7SMKswausBSXYqGUq3r0HeIOK
aFQPRkpLn/LH0/W9l3p1bhgrXRcmH12vy5+QoSF9cK6CiWWtUKDoqh5w39lhzy4BufXxGnTfWnyN
UrUVk2JAK87OoGUAyXVex7te7WMmVFzYJMMVBrYmu6Y/zfhWS9zvBfDLbUPZZJwVH0fhGWoFEQfL
+lVTVGbEKkjUJIttqk7ElMNC+aVlTDGoEPKXrPNioi7WYlTfvlINan6w9UYGBP4K1agJT+jVJMRN
Gq3xpbUh3nzPN3x0lyqmZcP/L2QPNpBv8CboWydwOwxvB5IPT1ptOQPyc24TlQO+1Pj1ZvLNsDeP
mGS+DLyB7H2zl28YQPWIN0zsgAWWATa0kOE4nsmPhYfbmvXnYYDUn2zK4YN2m2vJQwtHSbQBmft/
mnEVcBVEhAhUGT8xZM63wjW1o0wnRG5LIowBC6dtLcoj2p4uIjQmnF0nxIxNxMjun2+bxQktbf2U
Xfs7eHXxjj0CNmYBi+ejl7URrZH0mNLHQPBdDM1sBa8iq9djGJB/nxT4ODqEXI9OKgJOtAN+vnml
4//3W8pb11zAaGTUHU/pgjJ+YAR33iulrSy0DCqfseBqjE2DmBBIYPRxt/y5TH71YvNgzwbrGy99
1ArV7o74eGQBr7wOe9eYoOpj5i/d2pQ+Jq1SAqv6P963SZ/7Iy3EKyIDB+vozT0VyRiw4kO1bgp9
/xySDShmgXpcFOUUbm0qLJ/IyKVIwt4eEHPQQXHD5RikNW3S2BSSENeehHApcrlSodWbF8Zpoy/U
W59aBGoEzEfanaOaIb0QWr8RW1ULnzGVfxnrIRVnuH7RbosCYOoLManCJgTUB6KDuChbOMqkftWc
KhMxdbMdM2IBJE2zbIGqOIyHYDwwO3X1sOxoTWOo+K2Yzd5OgC/1SZEpP7YWMNCfiubd2cClKMrP
QMlgUkFHC2BYOXCZ7dcWDAe3Yj6JkpiYyLfjk5oLM8q/g0s1q46IOz1kBaiaR63Q11aUjIFJSe0I
9twLfYW2lu+1wfnBCz/z23OxHrIoAC1u6YwUjkCIkex+Ic0uFFUUwh+31o8wtpVNBZSakmnL+esB
rF1KvVZfFkgE9MrRxlgKYhGLFrSTJMEBknYKLR7qVLTvVJzB3Zk0GeLPExUXr9vAU6NooneiAT6j
jw1swhl6gMUeQjtBo6CjlZ541UXW/JaHzDYpMczwJK2zUNqXcNLVLE2zpWxq3v5j7gB5UCwWdtKB
ljI/guPkMX1mByYHb6qtPQ11ropiGS8OtZQ3/oE3jk+wA2ytxwW5SabDX0eHcuoX58ynOncrF8aW
v+iiMUi5J167Ri1yPfk8c7rNIdp64bkolnyCOy6AYzPV1jx0IFQlYhjTDd7iaGA0995bzQUDY8mI
kXVtktUfUednuaejEomCIylypMPkWBjgUX8twyLIJc3m3nFqgh7+kHbVBrdt+l3VJORwymOnRcJP
nREw/6HDPJwp2HJ4aGMHWvgZlbOfNsCjziodLOhB8jVk2P+CQcPazzIiT3ZINN7S6NPNAcaj6NcO
pRiqoAbS2ZgLmNnw29J8Ezz4CQQD/wXV4wLAC9a0DeoQhg1PT6t+ogcQm8oIMPQJRLLUV/QIwNF+
lMTLoL9i2pMeKIVf2ia5dsECSFy3QPl35eBwJ32vPCh+nFFKZEKmx1xanCTxKM6hWQNWPzipMRoQ
Ucl3URRay7qocSCWWl5HLXfEYzNaEmDytsFYot0ZKbpkk6wgrmjYiVXU5BHoMyJOnoWDAogj1aC/
2i0CS8PpkkP7ZVGDXuOn7MTyzZxwm3Lv6PQvv0ta5Z9Sq4O50KHgH7NGU1Y2SyYE1J0uy5txrQbI
0OATn8NQpxG2ePggTjDgEmLoquuceFgS4hzoHYPWKKQeQWGw3XcoEn+orUM8rYeUCkopgk+uFEC2
/EdOfCAghUvqDR46P9EB9FKElMg7lJwaJJwtjqtJO60wLXEHlDIlmiZV1132DJYUO0N4YQjD4N8H
r9Ej5lVsY4bqb2P79iPjLusnIzvBcjwdzg9i+SVOigcJexWmG9nRT3+bNA1/4mU8Pc8PdvpMrvWr
FA9+iZukdT5EqWmIP7JcVWb7TgpLUVOB10nOZetUQuPaRwEICE0Fjc2OQtX8wf/zrmaBDrIB243f
Skcyyjrf47W32nq/MacGW8wN+1a78IXO76WOAFDKqbEN7F/VZVjOuzxEouB0ACr9vnZk/F+jNx+C
gHps1EZmWYrSiubB6w30kxeoh25zWnLcJjidmA9bQRfaA49CrLFjisVSr199PlZqisF/Vse7aeB5
fNy0PiSyW4XVognBw/FRj53jz/NDbgD1gkhtS/fhLhqYn/zNHUc5RaDpybODlfR24DcYTycc5n+Y
rGOevPQHI2cITVY1LPz7qYsM4RWRYoCFMmE8AEgaNmzn0Vj0J7/Ns94ck2Va/fijtoOh4p84F7KO
oQK7868hw0LG1MhgBCaZd6OqO+1Sn+bcRKfhHU3eFVo25SFfes72yrZL9QGBTIIK9JC/YnPZ03QJ
WvzRBHXE+3ioanEE+xSUkCvhuTuAre2lllcEAXXUZ8xtiZ7Y6vTt7Mj1dnUq3rov58f/8jqSRjCC
ZWYigrsB9XPiDuEf5ibyLcwmuYnCSRjeUOg5wv1RT8ijuzkP6Cubbj9apa3eSY57tkJBGY9H3X3h
FjjSazPLj/Xotgky3n8ynlXdnIbrzC2ycautA069iD1oK6B9NlzCizSTwnsg6g9WHpxd8mumcBYB
cu5nKujg+x8CWHLse783EcjGEDzvXFjkQ22Ujq5CNUOtWAKyJd5BsdcalUH4vqC9/HAzajqJGSu9
9T/DHi/m1KCtSWlTslpVN/3HcTFPsffZ39Ysay3/1vHwPyYUtCKUwOmK1s3NDhVwME6DDhVNp5jR
LT5ixmssaW+Uq6JDyJRnIAExjAHWCF0Q5KXYzMYrKQiu4inSi+ooYBFHoHvZ0tYiaT1FefL6u3PW
ZDI3SbPJj1WJEl/Oe3KoEgg5vSl0l1Z4DVwo1BR820DFavgvSe+om1PjAvSSYjCDHIZhHhnM6qth
6oFGVdhItuD9VAinIqVKa4ccrhGtQWFEmnSFPREscnyhHWbtGm81y4d8SUWlj/FU5E7HQRGT6JkT
U9IGZxwuyafT6mcUeupcHzoa81nmQ4J2sjKkZiLMhKKuWOQ1nQQmSvcjukWuuRKNjn+Evf+vY0zV
aoleBGvdaiUrFGdS/mNm+JJEdhkR3JJeHmeQYxvUzmZdBsUsmXGyRm1Azr5/mSRL8HAccwlOfqwJ
Xo+OCbfoV6x94+3/c3xRha4VMFksauTth9IQ7AZ5abdExh4iZCsRF51I1zgg8llnBJonAgWHdi5u
LO+1R1n6uj4NGoQdlymq0pmDF8nwNToYL8s/TAvoXJFu2wvX+n7pnKIGq+4B/o49eG7jxbGSFs0M
CSHtIttUn35wgT2dBa79bfVKgNjory1+aTTZKTTBYtFA0MH9M9rS3lOUvsgWSGHKQBIMohxLHxNC
CUC10STSnSPMLlc4J5rDGoruqy8kRAFV/NGg9WFLJoLuNbz1CpG7ID0wL1uTiVw7ee4An0jRbQry
EglyZY0/egRXYFt3gz+oIGP7W9ZUG8KLdc3NvT6GJunzQ0kkPkNjx1nQHhjA4A3gJK3jwgwOEScc
GmNFAQjeEuTn3y7YbnwbLmO0699/CvXH1MWfAfYGdOc2V4HwdU+JYNGQem/qIp9jOn0CpBq/ePdb
cJHUpF9C4QenmJLdwIR7eK5qbx3CLwxJLIzveOB8BO8x0O5Mtu+PS/Hb8JQlgoSMwuk6TdQBMHkz
nFjA1Q1HvJhAd+2//k1v4j46H8O8by+fr0//2vAbLPFGwFLx77UajrYMfvBzpVhXMasKD9R1uk6y
j0QJScHsVJyZ9nwp7QnZ5pBvizudPPmk3f08W/uGoXkM1JeM4IjvNZfadBjQom6ggjLmK/N3s8D3
RmmSl4n9Qb4zC4noam+K6np83HryFVY1nwk1yAglp1G52xt2b+csAVNp4bdfcy3ezbp7BNFHvCwm
8f6m2WyDTz7kv9jgw1kWpZHhhch0O5Yb8cDzNlBNQs+habGFqVPafRccXmPRfufUxDv2zTG72oqJ
ydMbhS09eDzXk7DsCP5MwEQiM8QUvE3AvcgMczkO+LFU2cptrdUjgVLTksSQHQHDhvohrFsKgGOk
U9pHxU92H5DiI4bcE8ym3ygGqTWLKUcEsDB9mBb28mtng/kc13o8DnQg99XY6rNIFXYkgSeYewfI
xDBo0de31gxBpd6MoeuuMdwlKYLtyhSCNMrLlqhYgIGa43+ADTIUbJeiRepT5jICiTXhJAHWHL56
iEO3dNzQjfpgL4TBRtJx10DqvKz0mpTleubsGjODxW8ewQSNonK74tdXEngUYw8yvdiTejohOTy0
t/pZcraUGQdUB1tpMTp6oz9Xp3+tNmOlx4riJEadL4/HgdRYVSYHo6UIwoTJ5+Q9MJWVR8TAZDt9
0oDQ11839LuIz6ds7sJxASt966Vz5oBITR1QXd2lqW9C9CxfOY0av8Bn318HKktbpCUoXeLZ3sJm
k/9tCcGMg7tGlpZzYPo0ANQkoMNvg3/8hjvBXuELeYoAfOhAARKx6VBdkae8FpfP40neZdeWvCnm
csbITTl5FxTsJXISrsfi1JFAE9+b3APhNmByZXdE1VgmbO6h6L3CpMwfCjG/xJeoOyvtDKyGccFc
rHoxK33myebM8cJ8ohD4gl4PxnPb6C1jY1Fj1YnKX65ApvXuKeykBk9hs/oLi+7Vz/W3iHVpQIXv
jsI82FivBd+b2Ag4QlTRbxYW831KzPYABPKVNvhCj2g1GIZtQSQGHx4iZarqbBIEl3kPxCo3HUGy
3YgboFTjfYecvVkPJP3Vwuq1J69g0u2OtsrBdkec31mo9DqGgXhxRC3GCeUkMOQjhgOy9ZJwABBK
FirqI/LepKta73szO9wkwO69f0Y2LrzbFIx9RRkGvAcTPmhZg8jwh5MNaUkG2Zvm5Rav2SxIxkU9
JGfhBzi4AbNktROdziFpzA8a36OI+LE9JWERRbpol02ZyZI6NjG4Nn0reVuNDDih5JzzUiNYHOah
THqPpOQzXboegvkZ7rkzcCvOHYqvAZosn+0CGpMXGvHlC1WbfsNWT+AYjX8OzYKvaBqgH6IFJewB
mKWP7wKdJcAt7isR/9DQxMlmEcsfd5+PSxWovkUG7GbrIO96KfmtytCkSNAlA7GciILg3uq8scXy
fNIQ2Ulty/d64o2bOEDBAZtFRi7tb4D7+/BfOOrSzUkxM1UQtL2Sa/Q/Mdn+11aVWvXZH1N/7RKJ
EX+6sgeI26n4i+F6zZOE6wgD/KvyHyCK4Db6PYc4+zCklGzUDhsKIb0H504Y3E5/pYCIBVpPk1S1
/r4T1g0mWEywKAfJNu00uegdnyvOUgnd+XCAVxGaQ56L/EDYnMeAM5/lOhcj7/RYZp79612Bgx2H
JPJyjbD++SNHoKu437MkdaQHxMSVrHAc8g8spx+NswuVH+MTEOMqmOb/yrG1cagjAnqWqjcjT+9V
jKLaZNaQ7znBhpebbeoVmI8Y70V/Myt1kYOU6a37eRPSfNGQK8aE+8bfoZUpeRu2wl9ANq4hsruj
xBJwRYMeVOu8ZkUlNGsdghZimHJE7UY/srdXU6arkHtscZfcwxcOaKKO8hxDyfMZMUZKnxF41UH+
zxWLDjUgwA665XPoPhwv6IBJqi4gX09IoLvyaj96TAg/VYKCAdUyuNN4aexKdIgPKIltxz7Se7qm
XLpVpN8vgmL6n3uWBr0EQEwEbi0OHxSP2xdAuOosAA/ofGDhc0LcVusLxdZGojQUUJG2oK/J1BMT
lprcSk5LKvnJ1gTYEpE2guGZ9r6xhgrVlWN++Yyt4jciQqW3IXCIU6kVD86jnm5HLFoZVgBcEZFp
u+/OIjv2EurYXATl7Yn1ovhGPbmdsrcqooN1yWgFhlENJ/Y3K3DtDBs9xo58uljdEQN8SqYIMKhF
RRJlK4TRIzTFlMv6k4VeJ81y8r+ck//+Ucqocej0k7fmKpLiy8Xp6AzgJYgrBJ8d7HOBf8iyoMvr
04UkL6VgBVPhnA2ZXmuDFAgSxD8bLZVIJIRrZ7pNKf4ZBZAI4WCs0WAL1AUqXdgqtxPO9XgtkXSL
p3pc2offP45+ascuYw62WUN8qb1nb6/SNbxM0vrq3/TR14tOcfLP6sthfVs6Nr3UBZSA3stsZZaf
mH1KxWWryIq+ZLsIsBdH4F/vOJPQe8XTD7cj24vPAjSlSuULfcA9ttnFYRAwMr77frGWDvnYNX0u
6rB8VFjY5bYOO9RTKTazzVi1wjB1zXUnwadbdYTAoTXlKdRNctvmiR8EipoPDPaxAgkABz5lqnAK
YshItbuq8Li9BExL3WcO+vn2ZocJRThUFYxpdRj8eML9YvFuqCLhm5DiKPE5LINK3h6v5UANmNQu
4EYG/5k4ttLqqPjcKUnwh+FlCbx2l9dQ9LYlzMzrXqDgzFexEh0n9Z4x+RfVNNSvlw5ian1cIbxv
vOzgDvNc7MzXe0Hp3sKV5KUxsfaHcUk+1KuDRfYbn1e44shA/xOeZdvUFQ00J64yyhkETf5a3kTJ
/qnXCeaL4zOKp4wxyaGq5MY5SrRJ7J89+tWThPh8CwfAlSPj9d6mzTYcMz/hQ81GDlLVLDgTj3nM
+xzPjfWCFvNcfVi9DPCLGMeDoEZaWv0MjKtZ2yh8ZUkYQ588wRJed7AigdwEhm5T1Gw4ZEOWCs/T
D91o4ShcpaFgrTxPM5az/eDRar+1a92bVBvAiVJrHBngYIaZxk3aMaMKrDE8TiAQlE3dFvFJoqD0
TO7TjhrjBCCZwcWnu9ozInQsra9Y7XZThuxsQPAUwDnv1moK5MUFS2QOUkIkn9R24y7qjUT6Uh9L
+xY9n3Hk05jvWZOV1HD2JFy3SRtgu9ej5KlO/WFpc/3tnbl93fRD42iyUDsqq1azsodbEhXpwib8
LKxTphpYiRqanog3axAyUB+kHwAL/h95XYKgrknkrGKHWhNUVxjl0QY32p19ETGd3zwoIz2vHARt
J5n2VCtWPpe5CwthNwrQyXicmrFd1EVd7WlGXMXL+6sFYtoMgCfcoG+Ax9W2JFqdQnhNOzwjO9k9
Q/N/7+yECFBF5yx0qiNyC5b1cR24HT7tDc4007gao82MViwdku08T5YzhzFsfgTatpGAhcjoJpe5
x9FSbXhjYlRtT7Rk2JrLpVdBkuWWwRnYyGU1PzeCRCafi1HMm6UyYBVP/Bfao1hzAXWRDIia+Koo
j5evRgtu0TZHKBe4okR09RA5nOL5+jdKJTRW15mPujG1SLK8nULAFxs2y0Z3jO1nCvnJrtxROPeT
i1iHRI5/WsO8Xz0uSLA2yTRgC5gBqqlkiiVDvbG1ByfjEVZlsHT7QCSe9i4pf6r4z/IBDHEU5YVA
GIIZHY4ZEk6EgrnDdiNmtTYUM25NZf2B6C+hhQ2gjNaD8Tj9vE+N7gbMsIjtWnyRhUqNlTyXZTGQ
jMKN5nfwVw/AVwhZ1SLLGyIjjeRIDbvB0X77QYyUIE0c6o2GG+P8RiiAwxUZq6Sert3RMcz1MyHK
Te2fyiqscFurKG8iP1flJU3H21IR4PW92AeNn4zrmtXQrNLxgl5ucQIthik6uhLT8qI03WklYw1k
l3huNobCFGDKLcO/fg0y2H3Iz+3Rea1T0e5vFfn/2gLPG82gmzn0tp1sNPHAc9CkQGpyqxD57+fS
oAlPHcgBYg+ndiUWMcNRHrLb6qH23VTR1z3XNv8lDKRc2vSUID65Al7wR9mzwMkxsxNaFM/h2tfO
pCajp/A/DH8fQcmYOiLeMbBmB4aSMLwp/WjskH4Npd0/Sy870q4z1Ow/l4GXD+nDPGO+SirPQESs
2crjlp0ePU/xNjEFzFGGs9V4bj1gshJQguF+VZr9OaypyPYVzHaumIm88K97WjT0dCSn2wpk6BRq
rMCEHG2MDfgVYaJfSOKuhAEMyHNvhYwVIH2J1s/PfVRCmdTHDTp9K9ChPtfrQCBhPjVYaglzJYRM
VRdMpcIP/7oNnBIihCR+9x2dQIi0p8WWIV2O9vU32QHj670bcYWlBp/tyJrvmGeg9GJBg3rP7Oh3
6vKPJWx74tBnYXgd4l6ndD8FaVKNgZ1fR0EtZeQw5OfduIPfDri1LuXZz6qEkzo6fpTqmJ+RVB2B
o/9Y+TvonwzMYkb2fsvxORNKmKRCdZnc2NGvN2+S+TATq67d8ABcttOVaL6MqqONBkxZJ6KN5vxe
6MdftH07tEGPurzX6MXNfqPLGtLWpoQZgoPLkjIU7UzAd8K3I1t4ahO3+3aLrnkkLJMqYpDp2EPg
ET18gmXpCUH5Rg80FchyBSl/VoKOeDt8fWxJssAOXFHHOTXz1rZ3g3f4C6YlCp/y9xYP+ETSZpIi
ANn78S8MxYxnGoPcg9JENU757gxTtt84l41sZrDQ9rryVYNyuExMy4oRTqBhfLsEVgD+ABcbEjGU
tYddBJ1/XxftTMvxQfhun7RImxnTzbpF3nleRwkv0t7t3G+rFaN8QHjC8OXDnuDmiJwzM6yv0Egu
mtH7ydnWUHAZKr5m4vKT0uII4tjvDFEzMXtr/2576kwjMhEiJPpHhkPqhHeLarAQWqzABMVuALu6
sKE6oLhvxG5gWYoM0IY5hrAVddv4ksrqTcNT7ODZI68hwzX58GGzmI7P9ivk3pPQPqt7uZhnxRUw
VV2ep8x61MVRfBD10zLP3Yb/K904z2Hxump8H6++hXNH0x5duNgzzFn4TzFPrHQnO4ySP90CiICA
Wa/0XIh3oGNyXYTb+q0q7SgIfHLh1VyJ2LVl0Yk1PLShqoTbtAEh13yH79LQY5VoR6Ily/raZmgw
S7A89YbuYizX/uE+vGcqLDce9wXAkptr/UuouVepx4d9Rum8xjzNvKU/IzQptHPtXtK89cK/OBsa
wNMJvMdcJOQTh2565RZrCCUchwZb1ib6eCKuJ/+u6yCSFeGJL2wn/4PeQs7ApkN5fp7mW/aNfQw2
g8lce6mjtEMCPihpbYiTV8ai9ADPruAHK2VYj/uuLKu0FvFTXU3RsWjQTbTGmzIB26D2UMzRSoGr
i7Hf/mT9BLYRG73sf6oNwK3EB9+PHsT+DblF4+teuG7aBXh3Rv6C35P99krlUzqI0RDDDmfudgYI
Gu2A23hNL6uN8T1Ty7thoEC91DqcRGJeMBrnnkPYA2vnAMt1kUWW53g9BZC4hh/AbCSNVp3MtMan
gXfgSjb9e5/PoS2z7CvDYdDOC853xIuVOqYiVUKgbAKADPLswI+ODvE7VGBoRaPfJ+xlxkVqPv8q
ZdoAag0RyYGZxRG1981iyxUKvOVv0DovvlPAIOxVsNEiLkCCoh38834X6AaNT1bW8tv/K76/Tgo6
fxa9/0EKoLDyASAIcNs65ewJEDpKuHcsa5N8YdS7+k2dLTrJ4+XKPha8vLQM/5AWtUxgMWdOj3L9
nhd72AVhBKjd0dQ8EougINYWgiyU22OLR5PNDw3PILRB7UrtrKEMfJcbLJa+OgfMcvCwz2432j4d
ZoT/eut1gWb3hFERS2xdYGP5tCd0B1+tslzBsbdfaCxNS7xIcJA6KK2rUptw0L7kvLMctqXiVbPh
Ot3ti5bspYAyK5XqjJv3ollvwbqXTaSCNb0rJ2lash6q5KM2vA4At2MAow5PSCep+JcIsggM9ewl
usfCVIuAB2juHIfuwjt2BCS1YxC1u47w+OOfH6sifYGtoDyuXrsXpKskyi1/xUFSfgdHiU715+3i
s2zn91S6X+/fYOyqyb8tNYFFaTnBiIiwvQrocbJ/924VcvuA3XCav58gVyTDUDaYD3im9fK4ziM6
x4OrDvS2aJRDAM6N0nX0R9iCELrYp7NkRugLRuDl4ngQIgpDWSkpU/2CtZ6IMwwJ0PSJKVu88svs
CjIf16Ir9TVnb4pUI2FW6EeAifgsuXthZHfh76uPi7OHPXuUVyElilz0rhbFkHSfJsDrFr/ToeqS
qG3waGiXjIuSYQ4Ax0rNOeUiXw1T4URzuCUN4RdYWQnoszFofm300g8gW55JY6TihsN1WAOg5XP0
13YMDsI5I/i3aoZLCYNsxfFTNk7xSjDBrvxOQf4hO6/JElBfdBm/ZM4XR+9oATNr3EZ7iSMlfZf4
AmQFaMNRm4/uZoKWrX+ewrMkf+f2ofWNAxz7h2iJx0JdTnVyeGl6Kl5HDRTOeQ6RJm/ESTv07xBP
3OiwIea614V+llpF+Xh/GOwRygTYc6Q4msIKjyUxmv8OeA4PUWrk/7pkBmOstT02+tMfEJbi4Sf/
TC4rWcG1MHqfzAjvlazcV+NV1wUp8HdqykV53asSTcvpnPYIuO0CddMeZnRUomaIJBS35xXB1TdQ
n+0aAfZ5EqUrLKacWHKqmav2bVmE3iZUqly+CyOixritYF/f8OiWWub1YTS9efdZHsOBJQS6s3Ks
vTnQoFAv9FetK16U6DwIEbK0hglV0+WvERUf0HZU9sIFYIuVR4d2Furiri6VpttboMZDd0kUJ4hg
/LRy/41oorG4krX3GQvIB0GpZ+gWrKOhyfA3PtU9oUaNNYaNZbbZFrrRjLPCdNv7vF71cSPwSS8P
PdxldwHaxk8ZM7nnezGKwX5h+ZHmeBFBPqPzX0dh33is0kFYPtMEl4hRcJ5B4enI2iv6PyUdO3li
dmX1XTzCD0LQzWNlE7J43vbMZGNGaejQqbyUnMYv2M1+Ynhd/1e4YNKw+CWk3oUnSJ+/p5JL3L0w
CpZtIJUWyLg3h0hw1rhyoBKYb/ZgOckd0/RB1kvT8hmCJm2U5UlAKXbQpQPQ1tBIzXENnrfuaR1c
Nk/zN/a3WwCTmJYc/XxCC6VkGIFYyaiMvygpHerCKyLwgUbgmCbeQJicf6kJApcckIGvogB1vov1
VS3fdG8UNny/YK22HNIeHHv16Xzr96E324Rsj3ZJnMQ9fp8zHndYsEcbI5tkK3iPL3/J2mTwihfx
673xEmpWhvT5UqYRWn+OorUHB7+YSYtbamloccprgcLyVfmGSfuqDHQvd8sN+8tVYrB6YhLunzM3
Iwz5I2LbvR8N2RQMyeZhe7K7U2cctxNJ8luzsSpc0VIJBWX/rEdjsn4ZKDt8+L1WpLj3s2VOA8wF
b56N1b+/on3tOu9u8TTGU+TRMvHaU0//bOY3WAzMR5dFRIzfMj/nPZy5op9065GzLwhYaKiWSpyc
65W++sQjQTtn7bsYeTuqt3rykVnDVuWdX6C9DHxw+1oPQjC08YKt3rfQUkupr2qQfFWEnJbHRN8O
gjfNTwwK5Q0R7VY6NvhRKzJCi25GBNf8YfoD5OuxOkmFkv+NV+ZX7ZCF1m7yxrjSKKEVz8i4n7Dh
eFGrxiTBoXqjb5f1X7c2JRFXRz1c4k5lfISm4OwFrMQVQPw/yihhQpeIZig56ZwBRDR+9L8EJguD
bWQcQM/f6/Tcc5CTeA0OfJH9fRTlk9eGThZDZXYNE8e/Y6lqA1624UM8IOhvu83dXOIlQedvT2rX
XU0+DBMxU3nIT1oW76KPl1m/DFktiMAGOklk8//Gy/fsKfzzeNgQ+qtGr/qpEc0TOCM/97wDMxnK
4/f48yXJQNH/DiTicRvJWleETf1Aew0CFp/fQsDmWfLVxAjNbAqrPFz/I7sfs5H7UCiMNkyiNePU
8XLfqiTzStItszAxv4dggT+A7LlSFSXEI63HqYUnjx7gbHHL6uiU8OQdovJcTTheDq6V0xYhLEg3
t1vi8l4DE01EfkqDRg6kY6WRSfpFh9Fp+2yT6QhTMlQosGaPkyW4JYMhNLR7x+x1wgvnl3wI81Xd
VSqF5ADj05hdw4j67Nidnt9kjk5W8sAzQvyqf2Hi0A5LEge8CrvrwhnRnKKu0z1GOZPmOE1kpgxn
XuNwzyguuU3lyRDx5INS3FcQ6IXwZGKB8ez6SqWqUtEAIOYBywDil2gHjJfoyX9WyPmBMO2Q/WT1
q189Gfk7rV2gN0Zv6U9imvd0kCY4mVGOHk5m6zJaTpau6ixrVirDr79PQO7lwK/MaejjooBXODeQ
EWq6RFoM4VGDZwsdd9svJFyfVcTsPZ+4nSGrnhx66IONxqAmHI/G52/TMFiVXdMTRAIRFdaO2Vut
l0soc6nNpofSZtI/gHl8xBVORWj23Dd1nY34bDs6kl8cNQkxCePlDCQejwWOLbt8kbz3fZakfGhC
ZfzMj/m8diVzaneKacaN9Mljy+aRZiZU2AUJEqgLlknS0zuiN+fOjw2hBhEI6MQ4JexzPSwcmr+X
+0swuf4ifEToDov3/mdVzlmyE9HHJyMRLmrHDgAlMpYCbZLz01H2ACOTpabdsUrRQnyQL7mhUpVy
6kRa/kSPoRgMAnu0+LZ++CZTH+HXnHpfzvo64TIfstZhoqw4rYzNn30YBzB0mMuCeaOM4aYBv2u8
N93Mik4FQV+Gns9xb6DXcYkuVRlJnW7tEXW+Cc5gjZoO3Wp/UHyANWqIthDQE2h+tv1SbhccRKqR
MzPDpJQUD2/Vd1WF1VU6pKNja1iXiOEelcqJpVbeQ8Ss5LZ1b8ME6JqxTce+/hlgE6O7+J3OdaFm
4wGwRSfF0Qte/z+j2wNNt9SDDfXGW1ahWs+pOX6ETHEWfrRk6X6Ij/DVGdJQIfa3MCgpBSfGQK8Z
h6umJvEJQtmlI8EcLWriUlo/8jWZhL6XiQuEz2Y+dFAodsNMpmhuFo5hIB+XE+W1iLw45NtKcwk8
c20b45d3F1aA9ExQSPWrFHMJ9ylCXtYSHZHl6gzpR77TBmxXZjrPnKNIQC/bg9dhJFb6NA8XXruO
lclmu4ZF2cv+l1bgj3bAnHQ1REBKyXt8GJb11xWs2ph/3hWNuF17ofaeMzTPeC3AUmIaQ2AOvolG
3PS/kS+v9TAyPjG8POpuC29eprZWlzfL5bj3JrY5fo8/2i2enJWRYZlPoRqmAQfikTgdIXaQdbBF
FzjieEiq88c0NGgtqs/s3R3l10RQjBeFVMNCdsRWBzdazDYe6eO3qCqXKOnrm8P2HPHrRg5iul2O
N3vs1FYjd4B99+uLtu0tg3esUJdQwEdU+5TwqKLjk9a2dAEoPmCNrwyjpaSh4d10DjHqkryfgjRu
B+UZo+XiEbSa7DgSMeYSd8C7g3PNyPKJVP+NLxEIt0y+MaB4PTvXebiUm7W1GUrQbsCCVtX6+s1k
Hjg8RTntC38eFGjmuj8a5qHnsJXvpMtHRg8/1JmnsvuMISOhEWXu3WvebfgknDOcty0vMvpsJopu
9crJtEj8XZ4z6chlGifPpwg/vbA2VeH3AH5O3D1637G0JbIbW2ubzcPexneMHg0VsFWh2e6y5Gqn
44kRuMkEx/Sww0Wn8bdF+oz0UqGw76MPr7jPK5iqAnitzqEF25+xQRLz5Se+LQ9wX84rix++nU64
/x3SFzDQH/l7ionwrjpWEUSTYmi/4RLYH53msrWPqOAlEk5qBJ6ovnYw+wFhGyK/A619+DMpgerK
5MYifx5vkR3xxVlpu9/95mMP/IBv6+/av5hnoREvfj9EQhmfxEZHE1YSJWjl8rrmVYf0uLRBX2g1
0DAi8JG4KyEsVTrGfFL3qoN8aoLddJh3zFYh7VDvBxVxeh4l/zFxIaHqHCFgJ8a+25oPQRWnOtP5
c24oOUvhxw3pEqRzILQu6iglGTpVwjYD/gd5qSxPnYQBcaXdyGNMw7fTUcE9aRzH9AvEVZTcakH3
hNIUxI2IB5cJcSujfmVaN+dAaMFv+JJFB+a1f9c8iWPqSinOH2ckfXGUqnmhtI2RhpymrJLSqfmv
Q0JASAGmX8f9mTUPkTyJWZf62JGDaUvig3S7hfxJGim6JCc+F3e9SrL4Jw5vnDPHWLH+EABZCKMa
QfIZtxGpJqfEHfd4fcLhmgtEUZhhJYWGkq+eNplGnV74TTrg9u1jwb3ZFGHQW6+d26xugOaCkelc
8vQR4lsYHQ3+SWmCaLIW1qCk8D5nBEHZQBjCfAEBMvj7pq43omLUWNU/VkHUhfd5+3UkcNv9gtWT
jNpiaLqX0kmKONWrvQHX3zV2EXU3IkX4a/EbAZklU/ovxkpO7En7Z5lcDcCt6zOp9/0xkZ03Jg1/
nH/vQ8IoZLUANUiH+VPLt6CKvUp/cFc/OcIfdP0SfZUUyraTyf/VOFDpOdBVufe9QL8UQtb8PNug
SBcU0HWxedSgMHnhblntK21zUQ8egT7acDh7dojE+dO664cMNGoZcnn9GvRFeh+8m3Ceg0UPkei8
LB73AByaRBto5pABniNLCI8V8fxx5LQ5VPY9s/7koqC3pROMJWWO/g+iIiu493pqSrEx5vid4hRP
/NjruIACpftWfuoHKuPSOxT0vntz+ha+y8TZoLzfS6DjvT2zs5GE3VgxQKv9eJQGlM92E5EjjHKj
rR1cJp4MeaVITMlX+X2C3V2Bq3Klm6VjTZxnirIQDUp4nSh2LMz7PW29+6UoxYvfevMLJ3BCld/8
ovJa59c7E+MU9Z9GgOFvDhTR2JatD26Fe+QE5NN5WJ8AGL6SpPkvh8jKs1QNXNmjwv53WSXcKtAA
fuYUJoGP4GjYsW9PJGCPbs+xpW8gsW48gkJi1Tra+Atw2Egs0EWSeKpwb8q+XS9kBjKrbWCZ7iQF
5Fm/Nza7eSZiMujSLZhFO0d51jgcgBJCe+0J0uwA14pkauU7YeXkAgbmds9snvsW5NGjRwWsXrjB
QTsm0B7syDTS8R7frhsE2+aIKqWocHm/vjI5MaRcN7Nj/KRy8Fn5EOjB8CSo6EZ8ZnaWJ25Ug2Dc
lxbJOp5iaI33mKMX/3UjwunqTESaSrC45F43Q0nTYRFW0NLs5dWkpuLZcIRUvoYI8Oi3t8JRbuyu
ws1kJdGuDN6oEjsnUi8SQxQlB7Z1YRK9hgdWTRP3SHDsyoemUu/4DgqlyGBAQ7YOLF444fClPcyQ
FSls+87GFHlTfpVFbV7t7Wu8XqfIuPNggOGG7CX9KfRsQOPt3HL88iyQoxjbJ5F42sa171a5YWbe
69qZoysX+VXY8oXbuOEqPNJIcOd8pS/TzE9tM463kMc9pDzwhsgs16N/cjQ7trUu9VvI754PgkAw
NkbrlRAYhoFexXjopmp9NUJeKqN+TJ3mn5+ejIB66u1LDajCfkRM1HSYNVuAqQ4tQv7A2zOz/Dcf
RF+kdvuKq2HwTe/7A56Uqd7Ivm1FkeNNqYBC7m6E1tDivzZyDrtPhKgoKCWugJhlb0jdJpo7q7g4
HMhzgA9m1Umk02MLecQO/DhDLWCKZvRyyRadvbrmhlG/FkIiZLS8DOoHve0Z+zQIYFQ13fYt1Fb5
p22pb5K72H1Twvu6A0WPH2+Ng/PHPzNXc57pone+zsk/EUyra1pzg5JAAzte6v7DexyR5o8+Ayrt
VokQrhA9MHRUTZLBzyMNmw8wkBzrL9vPCdTPJ84oHmOB7RLVFLv3ZxMuaWlnUxKwny7UsePH5HMk
TeHhcSxf7+ALJq6gwTC1MYzzcKKIiXXX5SHZsfK+OP/LUoW9QPtsgSiqTJ9pUAtWUs6tmqto8hj4
2YYU5BdHjFPjF/EWCX8g75Es2L37nboFRlmtv1ajoFjsz7ga9iOWMe/JIPa1UCHA60shFEqkTp0w
EItGtbS3wT6DM21vkD7st7pVwPUVcrTx5SkcKSwoFWQIxE3iUtkNJowt7IRDQvvudS1ZIRZwX92H
rQ4JzvvGUp/uQESe3QNFcY7HteYI/hguDdP8mwYGb9jqLtIDu6D6xoMH8BfFvzzZkVAZsMgEAy/j
iPTtxsi+LfsVApBOisfXWJW+KYUffL5Ua5v3admDGkq63a9SEa9S/U6IFmDeV8m95EpPnBiaiNYs
Tsa5UXTaNbInzkE/jzpAKyDay042o0ltUtra0wd+SuHMKU+cozQ/CEKyZSyEuw6lVn06uasBmY+H
Rs2d0jUIFyit2yfocUHUq5st8aBhTmF0j3hmh02k3VxMsNem0wo5LkQcx2blOskIe4J9lwderakI
la/jB6a/F6pvPkvQ2N58GYvpYxwbRl+F/69nG0sLKHJH1bJKK4YfQ/MnbW5RId0Kp1vBjrq5g7Ac
nbV0Vqcbhc2V6GohXgXdUCH+TWlNXvU8ypdYbhdb6oklY/GbZz247FFGOxg8c+KAz2ZzFoenfE+x
9/Mj39kg9rEaO0MtejY8HZtk+g9cX28J8aAi4zaGD7nLqWRHAJnFyMsvU0cZdiKLih66AopfwsOZ
RRDYbyVu2+NZKXEbKiknJNuhc3rNitd8oaYXv9JiBAGQr4uzarJXw1+FUu6/hRHCgjONj3ib4Vw8
jKezfT0TroRw36fRmW2tKy9G9jpcIZfNP7+H31qbx191gXsjQWkhvgxdRX+DRotP/NFoE5CoUm+z
g3/sFzArB0MdYcPf0INw7G55eRGK5rOr160FxOFSh1xgknDXOymriULwxAV8DzANIlEB+5cv30Ln
7AZk4+JuqY3QO5IcZx9agy1vgMslqYh0AlUkd84Mbf8e1JI4tRpIOCcbviBw12tYZSmHYPSFxyv+
CwbAXarSw/BOIz5tsqlcHkS94BzLzQDCBFHq5LcSftJnbjkR6fNSPY4sqdGmNUqehTaXCjQeD1UV
g6SIRcZzgJgutgpTJulLT6DzIey5lLv3xOs5+NEoTWg4xRFtINwGPGDeONEn4OFjzuzt5EuuwyM6
m9ePqjzj4D0MphkGO4YbGLfoSrxMR0rj3zwELZjoaAOEcCbdVzSx50u8/lkVHXsIe3PEd/iLs3KZ
kQva670BRyLt5+JxC3YhI24HcezgzjWdx5QQeir9upYKeTAt8n9vQtfYDppJ9bek8XAkmQ/CoI4+
jbuQkAfF6vVwpX5wathv6K8+CscGtOlIcULQvCLGrZ7dH8+welItiO/HX8GgDhV52nZAhhcogryC
2/2A6IgZFdwlrQLjTpBXYnu6kJRUcY2Ws3oTryFSs1LSSfUhq7JlMcY/Q8Q6KKOCFc2WDok6aUCg
k1mJi8sFM/dI+sqdBi0zVio23ZAuekXIxS7fjVlJkBDlJTohDOdHgkBnA6wVIaN6Xa73K44SJWW6
GlhBLMq6TjG9qtoaPgO3IKoVduzPQ5tX+72mnEUieciCBbARRr8dbde4xRK1xDJzBaiQvk6RZ5RL
3kDn/O0WBI+uxMCjTo+w9LeftymQq3B10j8m5I+/4TBfKkJcmuvndrlC92iEXEcB/XguZJugfKxz
eNlp7rNhHnLl4Inw8h6RrXnBzGgP/ZEkz9HaacgY20iAIGGjxia91Iu55CJiFRWzRlcsgAZmOluH
xWDPLUYaH4dAlasPLMVKGIyLIfmqMw92VynZaXpq4B5QEIkPL0QeoAHAPK4lcwuMnIkhvICMIWgX
5nJ3zTMGdCM3tLwN1zCTZROO/40DlSkTOKnxPm19iOp7It3WbxpznMnmOBPr9XGRox9AMymOJQMy
NzxWXPHoV+aF8s4MWFABOtATnlZkVskw0dBqf0sj+XCPg7R+B/FEleqjaY19iJSKxhA8l5UABVEb
E0IW2QGI1T23SpUsrpRwwbCZfg3ya6Ai1VdxCiJpN1KEt4o1aivEpa5rQIDA+FVoRCY1KboDIp2q
1JJ3EemeM4MGTp4k4Dz1Gm2lSNboi2my18x4yJ6k3Onaf6zpIFE85zPuvXevU+yif/ZA/eseeIcO
BcCQ6D0Q7fpeBmEo2lneEqKDMOPwoutZlV0pF3eRH0DJjTecawew67FUtmMybXrEXMqMGFdR4APW
a4G6UZeKo1fVXpgT8GKKVl0NgNMxouiI7SdeZx8u05j42IljEgTAnYHe1w/Dsvfq0E3+G2c//3Eh
5oA0AH1JfdLqVLGxEhJq/Nlasvmtxn1Rq8Eb1MVQFDJkBVHSZ9/fFsgh4kMnz89ZvCfr0VROJcFJ
FSRG7TBqpGHR3hXf7qcCCiErImfM4BtD4z/9nte8iihK371EbBlSA51dxiL0lmJjlCq/pjcEIn+H
tesuasTc7gc1Z1JYyQc9jkNRnvhKx/dYWLJkXGqYj634GGWwzKT9sTi7ASMZNqkodjaaTQ62FnKq
Uv9ciVT3ovAWwNMOms2DFv1DOyKWWo/Gxi6Rbn+Wv3Udr4nwz6q9EvoouDZlgTC1dd/8KeIF1D0+
NI5OENNn8dfPsJB+vv6H6MREWn3JXtuxyvcWTNUYayKFZNoG8r4FfGSZy9RusJ9VAEA5VV4gAkZr
kq5uMh1zJeJItKRH3sUOeDJPHFH3LWHBAN6k6XDtjvhSUPR6EEretfbuczBekPuPNVuA2i35VRP4
dutE+LGXyFiv9286jyrEjRhmFw5s4/9G1fMIQF7XiZIrkVxrLEG5xdxrruODUJe3s2QpLrf1WOFP
c9mZg+tzXsQJmCzM8DXQR+0dmT26YTz4lMoVu7EQPKm2c97pAa7I1vPuW2+mVyzTMgj2yeK38v27
9ujEdsXIihGLA1YKFLJo5quGRdA5zN1463nGG8CXnx17+eNZDrZz4Nik44j4uE1NV33UKdn7050j
bLvD4g9F/db4uyTtLprsVfRovz5M+IBjXhgaRPkHfcckXcgRREFfdQTgbyBMaeKymh0HSVNIJ1U5
HlWHvM5gU7sZUkV1Zv99rOZHjs+Zmy8mrkcdBQw1brBoY3rkLIck69flaCtPfjVLi/8aPCMTZBxy
mB0eCxxlBdBPC0Pxk9HQsUVBVs699NTGriBuhywDjwrN7b4y6ycpArN98HT5d468hEWB05/JeLzA
ZzrECONP+t60+Z7aXs8TcwZoZNDUiWlgS+ic7+BpQnpLz/mIk0hCU2HnfP6riHw7KNY3Ver+wEQn
s1JmEF3/cOvMTlFYOyIC84UglUOUetXviYWR4U/6IAmgagYwmRFJx7BErG1cWz5Mrx2XdN5sSxRf
OOLB4kBTFDNpKcntJ+58kMJjch8sjIz9h+I42NvvxZDU4kvaBL/rO5Xi/v1kztZ/zlOCq7zm8Stx
jbK3aVz0DbCjFaeB9LG8recfE5ksTxg3unnr1TXvRP56b0Fq641/EKgVYkiom8qv275NdbMfpz0a
ZHHlFxJYx7iAeuR3wE7WxOV61brYrzE74dMNEB0+j9TB/tthvztNY5MWLnkpmtpb/LeOsCuIFSVH
Dwku4MjS7Au5btf58P+QIcYXrEVrGM6lFt/L738oF7tI7wgKf6M2wc68itPhZG2byVwa8lBlxqTo
xVbiKQLgbcUFk0ASk2rDQW8wWsBYv0LXEjZW7E1MtRn4zoVpWRMD4U5irAzpJP1eqy+0kzSO+b/I
VFtC2szaxUculmvsj35N5QruiG0egMyesMs+Dv5VnFeBP2wv5y+FcKzR2ILlblT1moudpl6H/GXH
E+0YTf2lwF+7aGiu4oRz5vaXNkwkW8D2OnKkTAkb7myQ3Tkjmjz6OYtjejTxY7lnJ9B10cHJ0nOv
ZhIKqNx1lNT8MXR9FSGTc59neyJ/mVaA3RlCY1gUnyH0Q3KRNBnoEDPXhFN4qincMrfSPyk539/i
xwErRj5IWPNtScmbPkXyl+XMGsFmsm4zeTWhhR5fAJpQMdKei1f/1VTzsmxrYgGmETpH5sGKG+7B
1Dm7UwgKiseNo4urovcqg7T+tt07P2Avyuy9MVwl2H3w7AyWq/AW0SVKTQtjeORfDn9NLYU/2uCw
3OCW11W40L3mG4IGUpkAKpi3C6BeEQEyxD6pIu+vqYeIR0HUXRxPo/p4UThet8S382BC1FgV002j
Pe4KFNXR+odNbiZdScOSnFsxErvZKQgQ4xRhdkruVohjN+Yccu3LXuPwK0Rs4GfrIe5BzMv4PHjd
cE+tHdUPuGIAfCpTJxYUsOVRI4OdXdjN2YY6S5qD281OXeGpSVEwvH0JULKFHjr+QHOJiUbS27Q9
4ZvHdSY5KiQNzzS0YNS8altxdOwJzujSdspmW+gnu3CuhXnwu11/uWpsh8TcJDYwGm8xzyxqYbjX
aT7IStmtwOmauR2WBO/IulfxmK7PPAcNl5I+/2ltOywmHZx3YtWSM1GmSuK/f3IymD6uwGd2kfgn
A2fpcfB9Goc2gu2D8ZPLBKi3+cdHDtBLwjx9FqAOGH299NgNPDzwYjMnX4pCmoq8Z049yzQd5Ofa
eNbtWQjLxvn4MZL1VEu44N2CUjpMVWMjLt0g1OifzzqVbD0ehpTMSF4/5o/Vdi0KDKe3a8sSYVPG
outOrGHp4XK58zUbs3U3V8LlH+7noisz5DrOPR0FXd3+wl1kcF01rhAamgN9Jwnfl844FfqYoh6U
HR6KNeoMusep8yapZkxRZcN2jes3fTBtFaf/ovLua2p/T6FY3/mvbQ0ZNW1d5p0+yNo4Qh/Z6yI+
eeuNOfEDLog3bhKRS5Xi/YO1eGtoxK9HkwvHdkTmCOIzdIvwaJiFEcaGgn0PGiKTM6toEpL4GpEE
9YHDLc1z/ZXGQ5UFoE9sL2e/C8nxYWO7CpNRf+rQUNB5JKLF3ml4T8tRqKOmVuGysJtFCNnLVrd6
8CmcUoWLeUQ7DYMZrBKVUmYzUYRqmWW86DQ2urfcFjYNqnJL27da03U7tyI+m0nnpWOyOjtO5vPx
taw0RhbX0fPLLzqeZSo7rLQLWmxLED0PsvHGWGFaoRlWYJyd3HhnP42/ngblaeanD2qZPwRjYv17
btl4/JasVIY/XHz/ppVj5HnHyXVnrdYSwm9oIvf6/O+upTY01ag8XmSO+qE1hAr9iLQxFtlCct/E
BBxCqRO42GTAgBd2oNokMuC5E6RdTCEmFf7xbSkPsuRy56Ex3YUY3ELWZMcn49x6FysIRYCEkx1p
pbM7tNXH+sZ/CKEBlAhLF72o98wUkJQwMDEHNXOep0RYA4IJcP45m3RJqwuZsnnBqi/5wheKYwzD
zt0TRIKN5510o1y0JpDWGTcjYb/PH/oBeyE/8yLxzgJ+qL+oSDd9US35Ip1Crlx35Ey+S3Gxal9p
w1+Z9VH4z4wuCcEHAKlTCQiriIZiQOeRFxZT6uScBFyeOrTohAp8CJezTvZLVJMmzTlhmLQQBZD+
CsqTCp2soOcWKJau0DcSn3pbjD719YZj4LH2z+9PnRrryq5soVb/OXsySiIoKI5XxVEnjfjQdypV
88xAtfeGte+xkb+0aZsWJ63fwuwRiFvxUGI8BwtNaJ6ekifMf04gsX84ypQ8FGa3/cvdpEC3D06M
dumP6lSC0jPOUGvxxp23usS45/aM4xSvH/OZCsoyMBU5xivjWc17CsDmOUEF/rRSMJ9guyYq6Q9J
Tnd3xn19G80t9gAoiLIgP7/PDCY8UKs2OimdoIY7koce0pKoGPMIR4SnW90M7u8iBh+cguWshGHd
YLvx+OWalxapjuwyn1ul03sFKCh6jr8tOX+ir36QX3N59qb1O89rVy/ekWADYQykEZskISk2F0Cj
GF6ARyBeRpDUF+I7b+L47xOVKXMOHxK4y0khEJaY11cCW9omrNH5R4lm9/vvDNeLUFB86fXK3ACO
+vQ4xskCig0PJrms88mHd7/S3kNgPdn4m6e2da54wxtNzHLUeSjQwMf6zVs5n5Kea4X/RteTWuB0
K50aBzph0e04xqoKyf635FSrCy0xZSpnmDHMv/feLLfwAYmY9y02xFD9NdbePZoerrZmfb7nzLFq
Rgj4vbYvoEanKvYgtJEVbN96ks+e1oo9OYnX33I0CVKKm1cyvStw8zqsUu19A+sQYwZKtkHZluW2
bLRRJSZ6Z2w/hmXrKKTYcG5FX+lcpwrifEiUxvDD5hMRJ0ArOyAppElgALU19hf14o8PhUhRcXU6
cxkVHx4oy5mQBS+z6e18qZdY1kOafYRTnfU3o2wBLG5kPYOuAHBGJkEQ1Kc9LCuEwsdDCFe+8ywe
Q+kSiiRIJ4sDLu+5LkFGk2VfE+CpQt4+s4bv4OelVBUSI81J8TIdP5B4CfukDF4W3tQFZ/TIfuVq
2HGMqCG0OpzDbUniAgnGPx3pU9Vg5FfwvZ2EBVn3H4PL27cI1tnBTF9I8cTJaNpnj3NZZo5G8y2P
rtsSlHEwWy/mXSzjZ03ycrsVPwTfhGEl8L3N5UBJ9KHyHdPObQuVTwBlDvcsEI5G7LVeQocU8hzE
nfLRyYOAQLe4FnW0yn2sxaOIjOQe+9nqD0vh50WFV8wrP1MyizDJbXu3ojprhURg0pqZhkw6kOOh
RVVJuU+Dfd3xymfnECTFfGhohiiHLnCCRm6Lsw82pRKnIVPIBFlrcWd+/un6UN/dJOs34fJFsW5d
HGcCXFe9jWYsEBmbhSAf8uj6HvA7hagyeWMV4MI8blXXlYNrhTI6FPIQPksFjwiPnZBl1CCx0ouo
ZCm/70rzVkS1/8bFNGFhvrn25vJ5GtnCL3U/aJvLwQCBtczOi1sqXNmW3RooGIYIa2U/hqxXcwOW
NDFHu493q1tnZtBEIYrpTVgmrUqpmcPWm+NU/mFgxoZc+UQPJuNvyke/noDthMClyHVifW6FPTWR
kAsbTGqJWpVFmqV6Aq8xg2heuljPcuPVJoYjf8UVZZuBpSwpEzp11IdcufDPpKULyaynKr/Dl21e
YfSYnvR1mzG/Q7AakktA7D4i0GhPWCkybdZrLzEcyQzcle02WhcOhn3oEg6N6iaT9Rb01CshA4DE
qxJgZvTjnMzGiT16P3JyIlSbHmScr93hK5OHbGQDF9XJ1xcsvLjrsFpYOo+xY7vMbMLOA81jAoVE
ouNwCM3A915P27tUW5S/iW9FuUa1A+aVfjSK8JOCWKfcmc1rJDPa6iG/oQ79HelBT3aAiWSa+Nx3
l3rDZpWiqaA3pQ5JlOaXGixwn1/yjNv5+YDuMTbYJwhA6DSJsNbHKvvak7oZd5sO9xhd1RIvpFeh
q9s9t2cg8sO4TqM83rHF3jS7Lp1gZB1KPzk8LkMBVR8IQNpDd8MdSReQ9HEN7FIkUwLz0jq248O0
kUFuFGbltSmiWHXA9smrmdGB10pZw8eGlRrhzsT8Th0389v8M1qcTFlzaPKJzJnBOLZDgh4qmbRY
sfBNifqy8KiODrlUCCIkxzWm8IGDju+rKYH055oCtEx+tg8Fm+4zG2BXQrAQJBvbqKQ3PKN2Hgkl
s0EaV6yybCgTjVQUCWOJ58gEVmbsvngkO/lgedQ5Hidbug1/AT2ukA6Pf+R26nB15MmgXIvg4oJK
pVnEWLDr+FPtBChbC1g/50GPjG8oCVh7csmk631beerBb5FS2yPRT/ZKqMGeErXtdBnCpsmYQ6eX
9qZyBddAcrhJJ892r6aFq7P+sGzGvBbS4C3uo1IMIEhiHC1U6vRdyr8mVEaA6u2Fy8oUK7pG5Ddf
fspia0iavctnrO4pBu+CwzqiyoAhK6bpabDG7n8e5/R5hNRwlODpPr+Zrb3sJCNmz/3ZSgwx7CB3
dOj3zemwMO6VCOghwUc9BRto2g4hkR7xGvwNs+KuAeTyFl23+UcNMNialuaHyXvc7CiJk2yTrTcY
XBADXkHNHQZ7poZR+013s5YzjfmTW+iSoXvGBsddaoC12AN+Nc2zdXsKsoVN9pbFQf3TH37pAj6R
zy5R+gmqP56o1/Kmhe8d2hYCblTBpT/6VSZBcxtcEp6N5h4ycGufAl6V06AxEVA5051zry3bsPbX
DlUWurKkfjz/PBowevC6YWpYMfjhrlmE8VKo6MCGz5+L+VRDimnnDcI9WhNp9zKQTtVEfbq5Yv29
av8IJkkU7ze9PIX9gBmJvwneXHm+uWuftVmPJoeMcE6FqFGzBUF5c64hTdMgIwwqgtRczRN8sp/P
KLPBcsxDxE8/wefSTMfwWN58ksoy7lV3lMSaxk7tZDCDowMJKGqDjGuv4HmvB7KxKQYQw+KTWMo7
WjhEI52eoQl3wjxHRsM67Wxmj70MY/WRNWgXc/JF5GqEkAHgJxR9TK/J3EzrQaFPChgs8w6qi+QF
d9EKCh+J9cSd+PLrG6kkbPq7PoL2c4IiyumV/pV5aV1mENnKkfWvpXyoXqEk+V+vGeiA0zcKFHNJ
s3zGneONged5kbw1rCWfL944RBglUSSLb68gDTOrx+xkwsni6F7sJlRPHZkqbhp5H75JDHfy3d4F
q93i+SpIN9C3Nvt8TejEZ33N9omlHIZ/VfZSsHSx8i+i/DW4CIy25a5CkzHSvxUv69l3gift12DR
t3T19mx36+6/9Gnhozc9EmmErMvTMnGugLKJ+y03TQnb1vXBjf48mMHHrB6ihitxlY1fAiHICpkG
9IIuLUq+e+mklRfbb2oBwHFvrfqp9MAz5c065oJDKD9SEXvm/4cnB6QvGYrTIp2mJpmCVFl2LlnA
sdfw/2/XYY7O0zY3qjmsTXSzKyBOGUgwaxclx8bJCyuGDPMPmN3MwCLybkk17Ny2YehI2V5whRSJ
dN0x3YtPEVQiiksRueF4FPzXxVuSqYihqeR/qstLaV6LhnvnXP7hb7bsg2tIM1LQrEcFGv/Crr8X
xAFHgxVN/XXRnfVV4HWifYNld0Ao4k0ZPP3ILrjPq6D59OM8IJpX+MV07oFvtEsEry1GQ5uEQOC0
cabbBfClBKb5Bvaqf4TajxkdgQSOJsdTs/Z8EDRzr5YAEDfefK4WnEDwiRbKSRW3wk8FcOUOmiWU
uVy1AKwGyFYPpZ38nTDdofUrbyf4SWAvjdrQgPSyLpMSjLkkOyv2FyeNwEFitmVp5nb6MOhiQKj1
SiHyNo5UJq4/3yBZayBvi1xHr9zCo0eEDWG/qUybaWXyq/u2/8J3nNZWfum2aSp6FHqAGtx2Bodv
fXyr3u5HcZxkt2I6Ij9Tr6z/JKTez++KJXIT4aNG7569BWLwjLawn8eLbUVoLc/Plf2Rp6PYTHha
Iau5Z8vSQRPoOtv/geeh4DwkhFbJeKa5sa8oppWmvHI4EHbO8VWsQFhLei7mLJPhfowYo9C+3Az0
fNuSJ/jMwRnVJCeS6ttzg8jPpNtF17oqRMcL6M5AMwki23lfyIjbT9grChqavOMqSMNKurIS1sN3
nEOE9IUTK5C1tUtsCLrShXEuH1P0cb9TmkedN/qR4vAX1z6N3XHUE/Xq3wl+CbPRqGk/YERRpSX/
ovfsuKLrYYxvhRvZkJ4utG633n5WPtBRcwA8eA4sA7e1fCGjBAr9POWv2HKuhmK5d2C705Xz6pOO
PI8UrrgD+iwk7EFKOUMfAJNtUy1DefM9YH7Vo91JetLl+ylk5Do6bXiAVUQh+aBaQSVqUHwUFNNk
3+eE+sblVF4ZU0snRuuczTeKYzgWX7uaED269Iye8YnDGxyg2vbGhnDK1KdaUTMBDNnfQbixtMjQ
CEYOjMqqMv+T1vPSMIdR+RY5foW9qNIz0/dsiXYzTmlIwqdCd+NsSvARLMPdK7V8++Jj0OpD1R4v
6ub/PnTSITvBE4Sf8S0hoGlbBPEJ3zIO1n4meJvw2zVxLN7wv8z6GJ5KMf75Glpq5iNmA7bEdwd/
W6R/TDzeZcPS/HOPRb2KxSdv5dRRULh8nYc8Hynn/5bpxfxUJ4T2s7NLGIkkjUWZ2jNn1uhqv12R
lhSOSvFp2+i/H02xafrrhrXqszhG1/UhQFCBmNPkC+Q0t/g20E/CFtMIDxpHvwrkqdybC1GP01/k
0gd1z+YqFtxbmZbBlRgiLXMQsxc8angIbJeNH/AGuuErs8oACJD/2l2OT6EwhA4+VYgXqhuxwteX
h6Qu9ZM28INxCgq3et27drU5tFSUjY6Iptx+xaQ2v6pALY3sbPEiiYuDGMmVQEWiVaC+QTOxaWNZ
BP4ccmHKnC8MF/0LouU9Ftg4ZtdEly2zlg/AoScWfHXGB2y2Gh1rt5GOwkfgL9ZWd968ovJpJKqA
6ypqD2rEamAePkuQopuzjndgHK4PLkh6WmI03NJYhxiOt9WpqEI6i45NvI78gd5KiWXTL0Ng0ftW
kJ+WIBCYBDbVhrWMMcFPQhnF7uUOY1bDKgR707MkxJ27YEe0VWRuAm9hDm/D6v0DNjPXDhU5pxcp
C8Elkrsrxp9a3bNI+TWYanAdxDUABYneIFQOoyDSRjDUvnLNV8TyniFLO4fObeD4lQuJS5FIhdUe
F4Lzd0Oy0bnezH/2T9NxjZW8dUIKV6enqNgxdUA44Ax/4rDA3vxXaV0/AtB7qG0ORCmtjEkq5slr
GapgK1U/O+/g4qzOfHcqmcsQkanhFfVDgwqOW03YKbp6zzAC/kOjdc7kV24ULq2CEzgmUrZDbd/p
pDHtEIVfcJMRMFY2UborwTaVM5UGb/UD68B+4C1pk5jj/5U44ZF3DStqSd2dUmkTMyLnJps1T6eB
m8e2mp4oMH/LqwVXDfNNX36SSWbvytN7QvBvHKGaMvhYxu+360eOOmCwJeRa2Hd+ycQgyVvpO4vi
oq/7P4GYVw1bF9QsbhLfDzdqQSDlcST6YYav4Fqb+qzMxeqAmG4cXNgF5xOyVN7Q2W+Mf70f29fg
N2KFMnIDjqW3Ownwl8e/pXZMak4NA/z/JdiPK+uo44rEb/FpZ3Q1DZ1e5uX7/cmJRh3sHbhd5yhj
WzjU5VDCWFXTh+G8/5WrBtWbKVfvtT/hoMgGIUq3+53zllyMAZxxYkJqG7ltFlyBg6jP5N6ioOcw
v+SnRlXpMOp0YYiu3nxWhpJQyPTtiS7On5xKPfN/tYKcUmAGja4qAOVzmgKyReKpv8tIVWvPizk1
mjpPbTyNJML/V2yizPDbaPWHSUvXSU9LxNktxUPidTBfkt/YO2FeJZ+WAFE8OL9nvVI5uepUj+CT
SYB+cnRVjL6Es9FDIeDLKhxplgELT4qHHXUDrOSS5FR4z2jvtsD4cRK0TureD0aQ8avz4uJCcffW
NIW1vxVP2q+hkQ/OAwbMXFLS1MdfuqdnS6fZh0glFjvxjQHaUsv3603XTE6YIJHjAErRRAujIbtb
dCsx5U0nI8TT8Pt30igiDSEUQDPHOjcbB1aFfB1Cd8tA+D7ukvMMk58mRNwwJuKsHV/6yTYINnAo
yzbPmWUVteAcdpOsJrgVDjFkPKgxcFIHT3yDNxX8CiAXhlrF9b8DozljHTXrWvNIj2WMkwtQZ5bK
6Y9DztSeiXjHqC97NpMydTofnJ9IqFlLuWd8A1CS+ctqQFR7vOYcW7y8Ib6NpzbTP2gxuFYx5KBz
ocWvehs/2pzEZc/VQrR5jeJ5S+iYlR9pWFq26tGq6GkqQBKnomBBrPPnWTvQoY4eiv84Zho2fEks
R1jc9nP6YQYkJCwA6IzJUjtnVZphTnCh2lCi8a8o5Gdorw2gnSQZes24BZg7UopLQiM5n01XsdYM
1mYQT3kmoeqeowqeT28dK1tvSm/5H3DoARK2ejKrjWBHLoBNQPXe6LUrdjZAmzsNCIPX0Yd+kDzw
ZgJc4r5idzkGLINpRVQ1aMukOG/zHmr+z4hcaUiuz7qZrYaIfogZVZPzzeUNRxvxIRSVHnAj0Qmq
0zaHYxsdIGLpd597pX8D+/PavxQUVMqeDFbvhtvHunaQo5frzQGgIOCyYmL+1AW48tKI3EgmF8Df
Ckc5IKZ2VQJqBoNqOjHKtPS62wfoXwcFQa9xLPfD6qPWIbi199ev1T64iwOaJyneBlD+znLvnN6U
J1QDekLXmkWBrs4l21nhORNDsP84pWuPN+Zh6Oki0lhfVEgv0TZGt8I3HdgCY3eZ1p02EJZVV+EE
iIU45XErZb8iZtQfhgBRG2CkQvUIhLfDdOLwMigijiQbMZlv5Xgosong4Q8mNGwD3mqGpNqHpiWU
CVXtZQfY3IRT2MQkzL033RQ6JZWJLJzFWtQkkD7AwcAcbJejAd+g0Xphqr0v6e3AEShIBIrHuZmC
SXf8CSqi3zYNHsX5aZ1r5YUsg7hbcY6I8T5xmnhI8R/acRns5enSTQCLRxRHvlELIcqmX6o+zZ3n
EH2NY98uuupF2T/B4vQWK6QDJIE6UZF8u76jDWM7o7hSYskTBn3MHoUanx6pN/8JP3F04Md4ONT3
lNsp35frhf0wz/GoetDQNscJiI18hhvGRGXqTadAFLzT7nrMudzrVa8wPx+43P91Nw1yLfnNetpb
u9Uyzn8I9etRHm7j/vR3E1OYSIW31y22Oi+hN+yc7WK9akTeR2xyYEmh2//sUjYKFppGNW96z2C8
0HMVqEshIT3kp+zwnafthyUiDWyH6JkIVOiBgIXge3m3wrGeeyTTffkMURWJIdLGIDRHmJ8L5NbW
sVreF15M5zaeG9CmlyKsQsesVflst4Oku4EMF0xoA7zX/XQpJwEz3TkwRHRiNHFDs7/j6qsSoYlV
oJO+dr7wJZbfkfQ/y91JStRReDG0S5zwfJZ4pPNJjYKh/9s2og/L75CcISV3rLY6QXBNvkK411Ob
x4seBW5H4tUceILM1icaRFyVcowxqrxFz9EQ6XhYoDWp4he46UOuyxhpvz3XYWQ9MphnW5VvKFUf
HgHvcUrUm9iOuCtqyOIad+sc8tQwGVWRM9OZM+9i3nXLt/bq3y9KNKfCh1PaMzfPn7pk+JvGCRYo
dbcIzpv2D0bhtDcG9XQFrn+sCRb/WImoR0wBkLAHUSLzVytERmFhdYqiCe5I3VQorsqAhKGa7HFV
k7+Gw2gDJYPnL5NShJlBpordBiEEWuckLslgsTrtkwRIyQ3ahFuP88s3g6y08TXwEGaeaIYm9AtZ
g/cBCxW3pz2RtQqfR5wthSDLtgQZjtvlwfkLrswxX2wiGSvdUERSIThcDVGMGXPtkGxzjt6u1psA
KH8tv2x5ocFNG7+Jhd/L5CJEFnIKv6iylxAeJNr6NXj3nrGRhd6+VRQ35+fUD7N2mHhZelUUJjCZ
VqnViSMFFTxd0fNtxs6RXZO6DnZnJ4tVVecps04Tc+w5IqckCbRe7gtg2CNVPOUBhTrRaXNQvTwS
zlbJ7mU18uNeo15zlIsaP1PU1aR+s3RpUOfKg/9FpTNqgcDmNgcUWIS9YmOWiZNOWvDVbLsJ9Apm
cj5UExwD4EAlP/WNJgNbImx+NwKKatQ5X9o3njwHV09LAGQ77aFBwn2qpLpp+GBGv1ilwXObL67S
IvKNJOewK2hNLOJytkoKD98VZ9LQ0YwyyearNfFh79L5s0++ORlfAm85eEPmBBxhJ55dm3FzdguM
FAfYQQpe8FrvjUE8nxCC+kRSi9RzmA7G0SZ9YAB5yUkSVYLQH5uhaZ0Mwst+D5f0KP8DUCK7VWSm
tGPWYMrDcbV8Bib/uhyZbGhk0nihyo4tWoot5dB/YKh+EyopxxuJuSpt8ydB74IHMF6K80R7YiP2
44KAypaVzaokqpcjd4JFRwtWN0tvst/NM0eQOp5ahzVOEMJWkQJdGL/6CdmsC2CBmEzJ/1glW6DD
/IPAS2ZAc4ARpfd6tjcrtc/LeEPjLnzZpd5vxIAWO8m1B38qrL28AWNn+52fsRECYLgWmumd9wYi
2m9sFMB23sKMJBhNeroAIvahSJxtHCsm4JMmhoeaHQWDi5u1He7G7lc6iVUECw7FO4n9+2Az1pXn
0NbiTKKjtylm4HwxN8W3IDdJV2LRKrlVCGc74QbNWO2clyUqzzB0Bj5fkUW2QGrz23uas5Yd+A4X
IyhX33KL3WAdliaaDzfQQq+xHxXG/9JN11JqRLMkZFmZpt80BQVphCFdVjXDjH+IktddqH4oJItC
fEbFJPtUQGcFzoVLP6NEjgb/oGDIoSCFJm1M4T8Mxi2BGBS0K1LMwmv4ONadepFGeZ2hENd36qyo
aHZgow01xTrunt66rRkIExO93i30AeRneg34GIHR0z2dpWoa8mLuZYIzDOMEAqIfPvU7YVTo4VQ8
GRjP5cbssewLMoptk7GSQ1F/Gx6E2S08LNQ/TUsfDSGD3/GddmBzXqXlNdUKOFyIvzrYmGVx8i5k
HRt+0gOrmreonqAmjH1QbTOB2nccwP51mDvITj7unLC0JwQ04UnVsXRVfC5Ct3clrcqOgdDEchLX
XH9c4ChEQNu13NFzYzrqU8OPBqMKxqhHxw82+MwaO1JX1PfW+56PKrBuwiz0UaenwqNvjloML9Kg
dTBHV+LbNIoNEBHJVbgIO0z2OVZAe+UvCH08pq5W/s2M9F92Th8V4IXPp6EnsDg5gFkc0XVmnwK9
1nYMac5PUO+8Ca2voDx/vJIsMRDrvXf/qGAxrrQWNjGUjiz7CVYNQtawHZP+AyVzwNAo+rR7wQ8Q
fmemEe/oRm0jqy9lGe0furMDQEPhwuwFtZmdZMko80KPhB06VNFSd8LbgCjJXQbKftG6Uabmt3nL
BO3uPRcLXqnEqnj+1z5MJAKxdegsnhVP+aGH7zl+ODyD2YEez8ImenbLOZrIlVpSW7vo1tzc0XOP
LAV3gXUWl8lLGAZS1t8DM+DsWS8v5dElUXfOWyxqI46aPCPpJFwMCZBp3AvIfentfA9pVEL7gGka
tJ1Bf46cCj9k4geltIJYVCGd2uZIq2+CktIZzpj3IfVsyABlmmAWuJxQZC/o5V/sWkK1nOCA2XhZ
j0+nuI+9urIedh8q5MkyjV9KQ4QiH1FMTS6wsOaSqMYkMHLDmY1oboD/9H9h3PnowerrGdFBv2Xb
Z6kvM1Stwe4+EA0/ugW7ZEtOWz6MZnEy5zKO5/ctNY1meVX/O/AAjZtsPtsGwD3/5W3GiBOOtlY7
J3zvOWEsZ+7FSv4OCt3N8FjdZL6SoqezVDgyn6FQGDoCcp/N49/ZFOjw5aP0n+VDikSiqmyc9bQO
kSYA1El3JAjvhWiK4+oJh3LBmpi8N5MNcQedCNV07MWIK3WjMelvQC8PpSw/VlNa+fCt1oF+u+Xf
v6H3RZQ+fWbazysmG4MGjzK18JkFNbJGFZQXcoFePy5AkJp8dpRPLBUJFSgkNzYVdrJJfiLzuD/S
HZJUgruyZ0LDzzlmq1XHQl7lisa4CePXGTuFVbtgfNMvmNwINV5FA22SoIUmm9aVmuCQHFLEdTvq
bvAO0fXX86CbiY6ceYP1abeSOI001e4HXX2zX7Yb1bXSIemkRaASSzqo4NvafGuaFmMyFueKiAzD
jEqcz1ZHMK2dBuh8QuvgRPGbC/0Ap6quvy7kbhrc8xTQ2DjISRrQVfWtjZkQPGBZI0kwEBK9ySpx
h6Ol0uv16dWUYv5gGdEtNW/8youBnT834DY8bIluY2rSQoH/3xzIgocuJmb6t9rVy3EG2qKjkOFv
i5xwv8i/F8xKcob57kVTYl4Vbwzq3LVhirLfTaAMnSf2jtosP0CpaIoVut9O1xImOHEtm7mQWm6A
+zNSfALWp5HdKU2ZCVWcInUUxb/AtC+eYJvl7Nf+w2YNe69WIgcv+BTxNKmv1ZLRz3s4R+AOVaLb
V7Xm5Xc1IUEYGXnpUgLKtsM117841S/h8rjsXSh+1QXd6VQbYH8pjIVpPD3a4Bq5cPnsGMghx+AO
3AZbOpGUWAwno1v9n7LBp0I/S5ilr3KraTGsy50tsfAS8Q1SRKb61kZMJsbWWkeB1tBZudO0xPUl
vEOOplmchAg35ZvYvDrqqndoKjqf4C8nH169NYZY+hX/D18FPJQXe4qYC2suJXIUpPBm7Im3QdOL
ys02BJT3JHEvJ7R6Yc+BYi/yVezFJE3absNhaZwMF761PSWnLzlt2lffbv2WpRBJkMHlLV47FEL1
TPoHElNgZzcAxsQdPhyXT1Jv57Gpkw3ZrKjvtEkxwvxlNt+sMOu9Gs8t+6CEnhoBx4KTAUbN5eiG
pxQgVWyZmvQoMuvM+b1E8OcBNYEdhEWdtZbLSc7RTxe3Up1egfMUs9HBIL0TRDH/8pTE9LZfIayq
boPUA055MXPgEbmEtoDQXs8asEgMt7pptxYZF4tjUJYtED+azA3zheiExAYOl0INrDUkxDcPh9z3
cudvI/nWmnhSc+j14NBrxxamT2l4TvZXDcgaZdpV25i3EX4xNsBBcE1z/1VzXVE9BbKVZmE+ARFG
IS24LsVbE6AtIhNG/P0ZfRSIrXEetq3nicyD3slVV0oSzD6kJ4y4HsESren+vqcEY0Y1aNLs+gvh
3M01kL7SXtsN3BkPeArKOtyXm3KqTGsy0cqyfdGw3EFMmXw3CQ1C5TDTkmUY51521787k/p0avmj
YBMDEU/jNBkC0jZui1Of7YMUkHCyTLUGxDOf3+QWVM7i97ehy+/UwrtqCtIiOWcotigAOQ+ByPXw
JccP5e3hFylSP4iK5HgiyfuPJzI3jkYVTejPcQ0/8lGoYSzJKY/zfsvK2SfchmstEmzAUE/Sg5rY
/tj5EED2pITe66HUXe1b5YsY8iK8fPSF9s3zmxf58GR613c6nlShSUB9LoiSkKBu3KEMW0X7lKSW
RZEE5o8OpoZQDCQcaIdYAxdJRHZVG2dQg63EbrKJRfXgP0IXWD7LtCEkaj+KG95MkicQa+R/35zt
P2gB9Bt8r2oouU7kxoI5j8lV/crCAhTfqfJa6HyF5xVx9CS9nPFDuH9I2pLy95ylRoC7EVc4luCq
M3iumdyU9WKbxlo/OAFbKIXiB4k7dmDxaw7Nf8/ymGmUKwBffdlY8OfIcoi0125/qcxEekI2w3B0
L3TzlexPZcnbLg0DUVlisnvp3wYz+py1/OWcVrvLEDZvWsKhT5dbJo46HD8zjAPCV927I1txqf41
ZbG41Vs6vPyp4UXEDZ9uCwtFqCDJpEzcFzBCgx82M/OxrpLG6pT2HiLX7Z8tjuLF76CcuAMouTMe
PqYbjOq54EtdCThoHgYH3u0SO+cYSDNp/evlox/PAGhVEMyntEPsqzgViRekPgeZ8hJbAjTExFlg
mZ46OopB3pWAGiJY7y7DOuaLH4IzZfIiWJm5EbZlQD6w8LDNZFGLadbgNpn19tBmYAeQS1f/5qin
zO0DulZXffeM1nURfXASV/b5B9oLQ/OHUXOwruChRTvchserp85R9pm9bo/ufL2Uyi2V02TqnSXF
BAFVuBE0FOIAe9OAzmvS4/jxw71UFY9T3ft+OKwnAvbQRzrZ1gyu7nHUly2H6Dg5cY67rM4FooPo
8DE6I/DEX4xBVsgVY4k7PZDktim2qqnvJuHhN1eO+aDsfBZDyf8ElWhEY2dalHBbLAGaxXtBv2FL
Yh0hq6mmiXt5AFJgxEgnbsgOmSgm+vSGqDxT7Ck6brJVNAhRnA9nw34hBQXxGaAlfG9lTG3XCNqR
F/V0dwX+ffFaWS/rZSrlwu5F4RaKesDBCNS+/jyegngwnLsc5n2YczHx5xNxT0UmBuBShoKRqHIM
ndt4J7JdNDdGP5+3HSX3spPVNNPBMMgGCEk7xaRNyFp/lvo5aHIXL596WhfvHFLgcEpZi8qwliZg
htOBXsoDJFTrn0Qbi1ZRkOZwCoiuwINVVdWAv4R3ZA1ycWk+sSDpn6yUnrLdfmlNzPYBODY1/HLe
v+xjPZuIBdZI7zet/B8Fy2GggDmMY+8ZPTbwnsVk7zPGxKeRS+IHfBiLHdKvkjK083v9Cv/sElsG
VWfHlthBMU+j1kYn96GMlRQvC5rqiOU4YqcMqQX3UV9Cp1A8bZoCdJB7ygSeEXBH0XB/QaYvGaYw
JEL5Q6MNcDvzJgFhOsI8N8Vpvp8C5oyEiw06iLSOIxvMrgwn9hoA3Z+AQuynzNhexW5nv+ls/50E
Jnrs0Hs6KYFGtzKk4KQ/8dub7pKq7aZGRAGLHYFnoouI6i64GToTt8j/sX5k/0Eb4paTmcTo9k41
6sEwCkvB4p3H3FlnqHkF1K6A17YAlJIxwiEvl5/NAoFhjCsHAKxSd708G7huijOLFkWjfMUNtm7j
XRYg7xLvRKY+Rv2RggC2tU+t16D0i3Tgsr/LJ9r1ah4YnErze2IYjBgvkePZrXf0eE/BIRqdIYCw
UVTAIuOSGJmi5UWiglXRsjn4j1X+xhlgWnoBzgeKC6IM40Gvnbhnd5z6sMJluaLlIyLvDfvPSMFZ
Qm1XTOPURblGqTFSw+Ik9xx7uYmBvA57gBmzXbd2D+sPLYcyTHioVcGSzZpPZ6UnfUW3PRDndAKe
+JQT6w7B6M840BBStrakXb5Taq6LLeiQypqT0jlug0o7AgNMElu61JMuPvLQ0DXBCMSXf1GjpWJ9
emjf3QEui+9YKI3q2IQrrapVMcRLCxNdN7qs3FSNUMo7tAGBeKNeYQcN1W+zEVhJlBPohpJqrIVz
UrDRuhV2oftFIgH9yYOKeXQ7aYKZ3eT9LvpkACyZzJr1e58WgGlmSu1xtE/cj3HltBEPUBBqsNtd
PCzpHnGvP6HUsZB5JNk5MfpXkKgkoOugwSYnLjZtmibq2bJvK0SzvVBEOI7A0mXyJPsAQa4kzAf0
H4egsgTN6VXqLblxh8KOUaAhPZKPnGtoAvQ075Ad/oRhfHbHyre4p5SKjbBXq+4JR4sjWMJTJNmO
ohZp/apKlbkUtciJDJn/1eOKXgfkYvCllKq0XUJYIgv0ijcF6Wf/QZ4wu0EiIZZECp9IyImbhKR1
3oHK7/oPHpVqZ+MtUfmY0CP1aSUD8Qej2tj9nePyJpEFMKvdK7a0hqOycrID9p9+/9hC2bMBVyog
yiTmYDyElTkB+CPc9NhAR6uns5MQgMuduhbilbWcv88kd7bfZt8nN9tUD1qPwSIYQbtULipETFu9
2feU08ddazV54Hmx91tW8rTrtgMh2jhWuwKzkCCeDN0BUo5/XJJebAdc7qNoN+fd/iNhow8ktA9I
wknAV5gb/6Ha7ZxMAhf/Qt6vK82WL/NxQLQrtTvF3mYAISRbszKNzeD2RbOnu014IlWvGw0lSzIr
wnCFKGqDhCq1pOPvrWl9Wg/OlglxXyZSlN9UG/U3yn9WM7+bfjJchLlrOowBABaZswtbF4swC0OM
FEc2YXeX4OXd+c1mYlsZXXdpTflWj5p4M0WVZ6owlpFPsdrFoYGUgNOBySO4Wti3pD17w9UhOeyP
0+AvRfNTKIJSKDcZkgzt+KfIM1KE8hQiMRnaLHjPgq5JVyDH8jiq+O8mG/SVT2kPWUc3vf1tj7Eo
N9OarfSDLd/QVPOd7N0c/swdMMYDo7yg+lsYn2xsMKkKlf+bdWCG4TonIQBG5gjqU0gMJzM9P7g/
d2p1SCokP2ZXEXXH2em2TbmQtwkJMg56XqRQUWxhsRoV7W3F5Gzj/YooCE1E0LcTgfhyHYvaTDCz
Dibr0EmPYGOWw4yJHDnA9iJUHcbZwmZ7Ym8+ZCTpZb4ZRmX8Q3RFeaic4yrg8NndkSuEfK/HRQl/
eDJ/yMD67M2Veo5htpTf28pMJ6N77e5q9OzkNa2wmGFKTDLYYiZFjb8zuEkRH6OwP3KLVTBNbOo/
le+ZXAyEp9TS1SCbFd7TUfuZaUK3AMLCaJ3PuYU71HhqgsEDh/kYm4gRQMtjvsolEUGHEqbXyp5f
1PGejHF0ERIcYDr3PF2OufiBd2/1I3mc0mLCVtlu84TjhPdn5MU8ymbzMEj6VnWHAJwt+GLwM9lX
N9AqFqlifyF1tjrPDuxFRHHwN6pH2MiEphP+OyAOIbej4ttrM2rzO3Td2iXveqY2sq0up512J9JQ
QjsQ99JHoEJy3pj6YJ6Feo1ssuC1wYYPB3TpWX6ysuiLfvJpyIjxfoZvubNAAUx2qiAC/K0if8CY
xm2o1WQXY5UOlZyL3v7+IBrgs120+TkGSWRn/s+94Pkc5x8Jv4hYb+6GL9JttVbP/o3/AtaTZDtC
J1Ft/mWU9KwyZ/NV4vnU9EzQH0BkLnGtFoCcFIWZwOgs/aD21RUgtv6Q46u+V3Ws672dzTuwGuE3
s8TSojawMyhzCMyeek1zYWcyUdjuBbwewVsF5EGTBEnCceSg53gEyh3CcNLz5RKtEM/VO7fg/+9j
nBOE/vRbzPJCryVDt0xdMdVseuTneLlZlFMm3a0GcfVwrLIjmu+EGAB3JsYhgTEBn/wwsfsmf4FO
mQkFaZ5hPp3QdIBi5euBnFl4Ob1LREv9D2367yNWtLMPVDU+sz4hC9rRwKUp54GzZO7r+Kgc0HBD
vgS/P8THXsH+Guz4/HIGAjjP6+vGrQYz/iLHvdHZy88nnvBIp4DpvDmxVAOoqOrqIoU0gT2kcWmU
a2XMTnSGVQmybm51RAxnRkX9GsfALki8JkDpRLkoSUSbovAkj/Lcjt35Rry0m7TSLL9rWylwJaHp
+9zLleSo/ljj3iGJuw+D4TZJQW4wnJlfm6BrrEZUapQJjpnPM7rJgfj4R0/5PVSIlrVwVXvOuxZX
u+4jVVH+2jqGpn8ejA/TGj9ri4ncV1P5rQghIEfLk1Tl+6laO3NnZd5tVFAcTmcv4NSG5dfdUUHM
cJ2/aVONx8VQ2T3v1UWxTNliDt+pUHZgmr/3hhyxKmyv39xkUjRoO0XK7lbiGhGzeoyAqfTa4irA
uYM+L6B2tVwvRnG6N0jM0EK5G9s2h58jZY5nXexFAl5h3HcnEqCfBpeKo0B48YyiW+wxnQaSmckC
RvWKMpdD+LhLJli7M1xvKf6fQB90ELA3fpW0p1fZpGF4voxdQHmQr3XrI9aPM5YOZAvyKgyi31bi
Eay4G6DMRKfX3CLVgKQngCXaG/i/HB4rJSmpshn55HKH9nShFmWnDaIE1tvPMJJiKiuIbf+Gv1qE
NJsTaCpuEl8pcfmb0LE3zdcMuj6jSf4OSnBTZAb82kzhn8lO08YpV0ZWRjozdU/VhhG7rq6Qwsi7
CPqsOTcOAhCOYgQUmC1oXKeJYwAOCnkBt/REQ+KS9xLvQqSeNIO3j8q6W9H8fA0pWstUci5FjBiN
73nRoLz+fO3M4GGgpLBn3SZSBziSdJTsZov/rbTX9VQbPLgCMTilxdI0gc+n7UDAEG2WJXtbO1UJ
/0ba3WQEONSYXfOlfTBt08jPCEU9lo46YzpO4ZdBO6iFBYMi+pILF4DKS/dA+wS8gi3fQudYqxZh
EuLMNlTiVmjk1EpI7T2zu8PJhyowUyiiomNQaWp3sONO388Fr0APyU8gYFUQMK99ts9FVg1bOkRG
DSNgz8DJTN8blBpIjwD2ATO7BEvmQzU6V6Xm+ESyl9A+SwP2tCQ/rit/l6Qm0TrivSQohIY04N9F
Rz2M6xXgbsEoXcbulOFX6LYf98R07PWkwbcbGJCiFL0P/gOvcRkhPZ3njngY09PbFZqAGC/94UJS
dDsLsd+iKydntHhcmumG+8bzAqHv9xBj3DrCqIi6khK0CIF0px2Ao193ORtkZECvUS2QLV83UFYq
UPurpOuUuwaKYK5nW/3+BkdAzU3nQZ3tZdKL2oN9dO6QoUC8ulnoT0MJfaUIX1tYfLIH2vcMnKe0
zukGwRAi+rEWSyJQJQdga+BeARLdOmfj/qp6mjR+Zh5Btm3++bSRSsE4TESGrKVvAAr5RiF3Kpz+
e90Pkd2z9eE725Z8Sd9yv82cTud56foY6etTz3bIYlY6gSth4WdWsQagN2sSYmBdPXTC4b+Vf/Gs
WxlfdqWVFPwTl8UHxdy3G1Q3ktu5eybsyN2IoXdE8N7gNBHAINv1spmM0mrbQCkeCyMH1ZwJKmCS
t2iD7Wg41/gis4sy5f3aM78Y9OY+aLmmz/gsQGMaVE8I6Fz1r6Em/9pKCaRuovlmKXKhl7dPdXKG
pntghDVAaBT2L/mMRTCvC+Z6y3dcATxr/q1MStqZGL/afyf4HRMAbDM76z1NW2ucuEjxSueMQ90l
dCBv0uz9gXKoVmvd+YaPocOUtCmbN3sreqjjVn4V8VWkUV8ymVILYNnNJWfi7RQcUidQStP+6d7l
m+18nH1h6W0UeHi0vHRtniHaDKpk3MgRodYOpEGTwnA16aQf8U5YBDXWL6av4HVBFx5tvks61i31
fifrMKwJFCgyfXtcwW4k1MHZkCbF2LbhMXonchiaBGTIBuKswnhzFTagy9APWgj7cRtwpLp4JDlZ
C1NVbYFtnkDvGJXc1eHcTuvmiAYUDHWJAFUiHbEfxkRqhsjnN6gDtEJeNUCQxlMRof8SFDbR95SC
y1QSH1dSaTBBFN4zgBMMauIYsBr/liQVBEIevj3dv7/Hs7uIFv4gHqa2BgsvqKbYDYq27EGIdZLj
zBUv8Y7k35cdif+xrRcCHlLAXG00SH4l1G5HF3ZgH5VSX61+zGbKF6kqgATpDvh1fyJvxI9OT0iZ
LLBWY4mKpZQd5PVh2R9HA+mFusYBd6WAqIX8EUF49vLgtHzHrSMwBdQlL3j6RBu2PUHMv7G6maxn
lBBI8YjJvm9yAk4tx7U8NVuUzIx0HFZe8EeIRdSFShz7Vei0rR0am6dEGCRYUhnSfZrJ7+9OQbkC
5H3HlIT4PURzueS/X0D29cbEpvS6CIpHQD7Ar2lBs6rlRfZwpDxGOu6RizYt+WNVRHxtscTxO8f/
W3P9DLJ8GYz2RvF+F+V/vNgXmIeMupCnFAdowNbEkT0XuA/lafAurK6zfvDwIxCUrnGI8YKUW6wy
LCEEKJrhJ7yVkOUAOEPPQScbo2TS9qpQx0NDzU5LYgo9xWJ8UYdI0dWdXzLVDUUMfu5aS2eVEZBO
U893oldtOH4XY+HqR2NnhfktL87SQgJcQlh08Ev2fcLlCZvG9D4KvPUJOlLBBd+lcjfVDfNEXTvX
d+tzvJOjbDE8v35hN9zpqR01cS8VxsA+WAj5J+r7xfiBhQnLMX1Xvo781ORlBg22b14Omuq83odT
kcjrHLELORkrefH201zX9Qg1gYuCd5xqMQaRLy35Hps7P5TpIaTFf4kA8ide8cFuF7Ra8Vz0b8yg
B1e6YqwMjUSxNFmVd7klWkGuqswUAz3yUkQOttN/e4fs1CG3r5CIP21TxzN10uAX1Ui9rscoZvpD
TdYqXhZnDy2K+h7Cm6aMcSqzUVBtBnig+JF0chf9sKegYAaDQpsA0fLpf79nppf2uOgnMfDiVOiS
agIugrXAu1c7Z70l+XwTdDhXUgAproEPUlW6l3PPZe0E7Nz/lpM/MdaCEkeKpEviyRwrnXnmdXoE
xDL2+gF3iYmnBAyUFUVas3x7oj2Rt4UWD5v0aSwDrregmJwnIxdUwQ/FJKRehygolLCxYiXAbmrP
rsSVXr8VpiY1UEeeufttRXFBVzlmtA8WGDyCqPOxO2PPlsUvvy1ENzEWbcJ1FH5LBVdm+Gn4BpQi
ndfPr88Il6FchTiNF+UNUrDG3EVZ/+sEKWznbpP6miMSmBe5dXD9KNBuZnWRnrqDqGriNan3AaXj
NX9W6ykMOLnmmEnEXOGo73OzXmFD/zspRu9wwNArsnfxk773g5AedqgQ00FOR5H5qgetFBq/VPk8
fy/K+R8SIlu0YOQpa9mFhlzPHGWcUu9joSZCE/Vgdtbt4d2agsqFSJhOcqYuEas2Cvk1CrRhI0tn
vxLqinyaC4nydNQHjKWgdo3yNFOy3juO9szF4EfDUDHDqd4UDJRWQdhjXOENOF2hzBkniH7yJJJK
D0erYNc5diY8fEfDVZFsYQjSjXYgXb0HeXPLM1uFP9rEe3MnDGnTkjW+buCdvWPaJGsvfcGOIzHn
zK/3aS57wWUfG3/eAdOGeJkWXN6Qbh2Q6nxgNXrw6NjiX4Fkv2H8C+aaFaGw1KCbiftP9q0wack+
fORn7NwYyQUfMsO/b5z886zr+loPd7XDLVNT+U5PUQytVa1tiVwjVIlBBeQHPAxpXElslEUybkPZ
hxiZBQ7lmqOxY/bv5hWvVGSqvE1nvMhMNklTRYAxXOc3LBEz7mff9/TY1W2+bPzYV/wyKo2lpE/1
PRHKf2Uf6bpKdaWSJwYNW4z8g11CuUYyoAwfr3fZsTm7DDXxB3tpf7dIZEyJ8nSYWXPz+OrKSF+N
4I+ZZnc4KhpUjeEEIjVAE7F1aKEGBdb2m7ZCGJa00ZRu2NZ9zbQ/XFGeeYNcJrI5+rVEbXvIB7J3
/Y5XcTRK894U3hSANb1SbED+JAPmnZLjO2QfL9Iy5MOIbM9Zo2mEAkdK81HQkJPNwsv0+8f/NbMp
+2Y6iuCR2ddLcQXdRrmTEEQp23Br8aX5ZSiPRZU3DSmnrdVyfbhxVcTfqhWVw2MZWqfLfbtliC3I
pJEj7LNVfGszVjibiSXUoqcKLirzoIxBbFIYbucAZKZO05Dc5kajTXvyykjDqYPwDOLNqT5LAJey
xI3Q1PmG45nwql6ev1P1kya6r0s0XWwCxVUw0OGC5G8Mtc2+rmK7rPHK+1IrLDhb4RpBviqaGDuG
IbkseBXB9Ebp+O/P+JaMaJQiTMgyuw6H8LHFpuHq3G97wTjquXzV/tvzTcnEGz99exZpAwOpG0Af
lPd9f82VYAkYGqMYFU0Gt+duFbhRfN1yhjoe4gy52mtV2dC8HtmPFd4mNUV6LT/3s0FMwYqiYmU9
82J4SBNVrilp/T9ikEr2I8gtLeaknhDMuv0/QCbfPiaG2g0I5DpF0RpAFFWFO0QjJBIXEUraWxE1
JtakMqHtl7WUwBNEqqyNrbFGIMbx9o2z/3W9uNvOTbvZBfHtpHBb0szq8X/VvVOLEXzOH5oPDlR7
2Uub4uoj+TgS/IBAAiPo5P8BYfrMUkTcp0pceVIMNDqqOeRmbqOFS4ExZAHgkhxJBJbuUVfaP192
4yNFNqmLpg8XElfif0AgbYKDbIMpmVeZu2kg9neTauySoxRTUiFs6HzT3m1rev9fqvlVSZ6sx49l
CsrnQbWC9HiQ1pXzX1E7Pxo7YA6rlzd3+nTSApCnojgslDIdO8nxANFIiTPtaAT9XrEb1pOxsBtT
lWPRW/a81z30u7wqvDmMYXWamVzgsjGhehF4QAmRMYTm5hfGab31D3Q49CmtWLr0ocDSETe0wAfB
/VUYBwt4CPbFgGyIfWX9bbwY3vCMN0BXHDdGSU0p2RR+Buj6bPf4IIBnajCnZvOPGGNCYB9m1Yv5
7zUQnqDHSWXgt0G5ejPTnAmPIN1ikiNQvbOJoTdL7urNm4xl0TUtK3PSQIdu+5w9MJpAFaR6A+MG
E+8Mk7HsvJIMw+4Z8THWB2Me+k3i1YgYKYViyT8OHxUGULOhIRG89sr3GAoUaanM6oPIhCjAWouL
9VjchgRlDaHQIPL6R7mqCOM6QFdKvg/5EPCFMtMvCA1zJ7yZL4Grx35tcMnfnl1UPvaTYkoJkBoe
YRzSBE0vlqVob8YAnFNfc3Ha/FCT5KW4VshMZ5itR/hkvLVv67ovGOIGX7UpefpqC2fooVVrFVS1
Nu7Ee2iunuyuuYj5X8jvm+ywck9Yqi+AVG/ehm2Dn9vR9/w56kYa116nEKGSpFzZsft4q5Goh4Yp
HVu37g4Evph7R4zeeeXSVCazo1J8mdlSjApt4o8dBN/5qGQFt9VBFwf639n6aOlcRnNvlhCTKA77
89JNIKf7H0hV2hrJe69+TVj5FMJ+Zt/R1afQPnsrnvngGNxXWwduXTfNpqTFiD3Jfb+N9xGG/w7i
LUJnQutFbymXZwR3k1xoOF0kRsNQF6miV4IcV+hJx6DWUDvAC0K9gj0B3qag2dYFca7Womu8rMlf
3qziaCK7qFPCWOQZpNcTQr+c3PxAkcs22y5nMZ6/ivRCpCkuU1mv+VJNhS8ZhfojJcQISJpJbETJ
dXECQRGrIfVXHY3+Tb10uRDbg5bGPy2CRXGPO1NQ9HhIKRmNynPf+/erqJYrcvHJWo6QZPLdqBiX
qGnAT1MHTO+B+/qG4rGEdNv5lb47uLxchqL8Sx5todO5senIPUJSNT44ikq77gpzWDPVGfLhjZxB
KRhXV52dHvvpQBwCsTrbhITK+RrmXQJSKvHMbsVeniCQJi1/7Ao6nTeBeDSJg/SE2RUb/to5iwxT
CBukHErFh3J3Mp/SC5IRUWvbBv3+ytYtaJZ5wUYpNptBSoSTn8Grcr4khLq1b3zDYIkNA/hrBld0
EdqVvHshqNktIiF4UrSZT2S+e6jRCPISz6Blc7IrzDDhPyScJ/lQI3x73ZmbceE0zK+Tcj0hpazm
yOvUJ4P0mx+antlac5cOM6nsmUHEXgmQ0+/ZxDoUJtcZ1UCeDK/Tym5RpGeYz6T/EPiGvZRqnNzo
Onb72B3ARdYDZZI4tpE18rWAPfstxGwyMs4SKbfEr1eM8HHo6w1BfF4TUTPqPDDGjd2uKTAyAT02
mHoXc9A83waYrkJtMRdpvMnZktsN/2imJ2I5TfiJPaQ9Cjw5+3oE8XyyWSr6cB0KMPmq6u/ruLRN
IXtxAXV4xzIu4F/loUvd8MXBWXoUF6CaXBqpxN+PI4Z+cBt2SkSYMdkg6DrlF2Z7JCkPGzqpDKTA
vbyE40lURnhyth86f419NHaGXDKj3xxOzUSI+rlT/WndlrlZjgZ33nlE/1a0wB1Cf/4zGMrTZKeI
HUGFGPP2ChMRUBRJhRGc9V2WtHWnOeALhIXkh7xvIRXCATkCFMA7Cj6Fpw1o0a6K54wvHvTMbPgR
ByfhV6oguTbCGWusSnJtwqz7ATsmvWtSPKZNvbM7HnNYxHDuHJextP6BMZKefiepJdajB3GI4Hit
92BDk0GZeIkrlwb3FoVGD89YIZ/HCTT8LyoTxKLkGpI4RvcgwQxdsWXib+UZqQJ3AvyMy+sMp/06
hJyelDFf0LaY1qJBluUo+T1HJxWa0cHRtWhwmP6PaTkIIX/GyGb+LBitZYVyFA3iYtPMfUaDtzPT
+hH3cG1oyk8gHYWTrS/EYA5l3gvcaiIYZW2wc6doE2256jgjFvLVNEfb1mJKg5hbMpgExCn8bQaN
fYCaKosZLqLsUHkzJ71JnFWux5zlftg3In2B8FQkbInam8rBrTZnACNU5cYQ6vPfGoxvpfESI/MD
5EdlZGoAaTl0Myvu1P6jO3tmw4eqLSaj642yC47NwHm9+6ix3AxHK5Hr4aiklyisqY23z6YkkX1t
LCopwhgryAkmb+KsjNOhFnz8B/5t+69c+t7dIRVkY5NOajma7wVPkk2gufuYH1yx+nt/Ka1mv0jE
3CfafyEuF0WlezXDCDopHOhsxWddZiHMRfGUGPOMDItDBGTPIQz7ZSZeMO/csFcCoIFzAEVmE4hs
dz4/VG+o1E/Ms96RaOgxnS7IpdieS0FOC1Npe2NUrBB229D2pzWkFen2+OkQAOKziklb4g88p8QM
nIAmERBc+2Ntdxllq50kWRhc14mcYSXF4hukAcvEGfIQhUwypy91XHXHRYvvkKRc22/Tdi1Xlzu6
knWFAlfBFWBfNQ26dZQ8+/5qUWLyEgA8Lbb6S5FvOK0yakHhQW4WNYS+SRzRO+X64SMCtw1BlqAg
5MZi22W57d6b6bnom7ZJ8PckqL98uBROjHuA61AjNq+2eX3ftSOfX6rUKunHAjNFhh7+L6A/clYo
EppBKfKo0fYwODR2XlC9izLeXjnjkvcNKGH1LWbydq/BnRx+7gaT1a7DljaMATUS3I7QzggIeAeO
2AtlBgnSxsMkqX7E/Y2bA3gEyeLWdVvBDUifxqqixkpNlMefBssAmUmRZ0OsWb5UOFDiIyREdA+B
VdT9kQxuWqfrCODG5SbwD2Z3nbnDRpOWi/h2oR5pttcvOgrdHmmvjPlfPxHFlgeB2IYihwWO6XZs
CHwj3JLIcIKjHKGC/rAWLQRQmFzQedD1kTl7bZn6hDWXe5H7yGXFoXnrDjmdHYDzu5B44agvxcJW
YwnQ28GCCtICXVXFoxMF90lem9eYLMckiSOrqe0qsBDDDZ1FMcaZy6oqMcrg8JQ7ca8ujl4n60sE
lhCOwko2xP9uKZ1lfBWJj1zoMhLdY10wlRs5NbqLKbGjN5Vu6JMFyVQ8bakuRs1cedSwThHo9Eq2
uf5qH27KwxqENyzwG9VNl0LbdigVJxKEfjdj0jh+VzuY2FM6ImtF2QRn5dRUofNg4gQyWBk1cbeM
F7EAaLctxqPGVu/jzft75V7/lvKHBaYC6KZjS+vAUZWL+TXXikuIlGdgQSqHphyDB82hUJkKqGmS
hnEIQGPMw9MYZy0M+Mnjzz1oJwniWiGcPFPnWnCSTopGygmyZV265zHISYVtL5kVHR67KBTuz/v5
27bgk+SzMgs3mnLKw8+g0PHGPJgV6xyBXLfC5rzLokIC0LOlYXYjovyRM64KoBUC7O8TEdjUU1Ay
0GsPjKmP7QCvZgukccVxnrSsoq36Hj3RXty3M5gwbLGCG4PJv3lK60GhVUyFqs704iNZ0nLhI25A
cDSHddal10n+tlRCmwil0jpRKW9SFOUAef2e76wwugt2gm3I8uGJ/ijfyhJ6kqpPjHWvgizImeSn
oOAMrcuPUa4wkfrJQxbMxOCoZorsgwa1WMIhdLB6h8wpFbM2MxZG4FD5ZKYKm9guvyGtn6bSbK1y
keLsxJ2Hu5LlebKuvJFfymglzeL5CtdcFTJfV1O67decaOfzOjCXyXY9ZvzQ7kV+JzryuFAbBCnA
3aCBMyh6ai4q7UHbHVlHhW7oSapfrBUUgC4i67WGnOe+fKQrgpoa3t/Fs3ybZ7klhDMyw2dUqt0+
hYLj1gVD0CdvI0hHQs3pgwhFY8ilqeaA8ZalnMi/cnzQ3JDTa0HRIxyC9/p4MR8/UB23jAWNxakY
CDDBIjZywIYbelDtsFlQNOI5vb3ZREHfHZAS9tba7bs9ym7QGplUEKWvfq9MCbxCxho7j6VrjYDA
tKxbJ//hXvqUvfz0DFqGAVtcrZo3AJzD0ZZ4UzNXVRpkBpasuu4epxypshG/nTERmIgGcp0wwmll
aPY1xcf/3USGRb+SIoAk4pvyIBf9VAsHtw7VVgxMgnzJt0GMu8t1NVZG8yvYEk6Rz/zisMcaZlWM
CduToChF8h+SEpf5RoQ/yUDrQh82Xq/iYk6z9rjW49fDaQdgzxX91wSDLWYlNInNf6+N1MAfwMNo
iAGApAVZ5YJfrUWKqmLZpMufk1qbBQgnV/BA0f29UjnacOJIm5/ofgsuq2x/4RCCJjlNEwIAkSK+
NmgEM4HaUUDKuYT3QxyhB6qtJVP32pyKIh3TQUPOtfKcf5fDLnOS7ir/Y3UN25+9IDmyqFiAMgtf
zSN255faKPI/5VD4DTFiiY8KpAOn6b/uejVtWo4v/PrELun3d+HdhioSUFOiKYeg5Hn9uWIpiHTP
nwAtS30AqPN7fCQfLrIj4RG0f7wMuPozywf6bPMtayuXTlhwyiJFViJUvKaJMM7aBPDxhmqb5k8b
R2TpyOQreE4J0nn9/AqUwrcgMcuxqEBLggpjAqk6PJb3YgEtMTzSCeDNluOBFgT5QOHs8TWcTLl/
GRZH8oMTxjhznBQkCfYiGJoZbEiTZLCGn4KMTON/6z8KAKoAfwsQCE5N3EK7SDB9jQvUUA6gUQFe
THpT77veVVPjmlyntb7q4QtNR1hO1wnjTQUvhT68tnXoAcS0I0amVJOODPfi7KgReHrhz4pbAJb7
VxwSvZflo5nahi+FAv6f4qTg7TqeG/obzuztyb8iCHmOYG7lrZdMHLz2P8kxdWSEPgwyZPrd422i
CvdNFfFykvZsxSmZSdV/TbmbJpBRJcymcqO/fUpXvNq7WUFWygab9z7mjHPPGQKW094ekF46hahv
auwy4aW75I6WMQL0fiiQS0AKcyulpU1HGz4EQuT4v+R4GbtvZP3S0Wxq3fmCzTskPREO6KLVQaVr
bmk5ULxsJJP5Gzg2f8R4683qw5/qUwCq6u7N3GrevWgcCxeyY4ugDEjIxwh281wnuByyWoCsDHtx
xttYh4tcMXFDBFfmk8PWm98uGgFMU8ptOS8Qh0SEZ6FVlYC26ZSuF1ZAsKbxiG6VJIOrUDkweW74
AqgzN8lSPQ8PQaLUyQwa6l6t7u88UPAwwJOol3A5Ff1fkR4fZ5ueQkYTEGWviCInpR+XJywVFMD1
kd7VRkq/VMqM1ykuUoxZqKs7jGKN2YjbmamBnVOfptxqEj8LCWeyf0HMzB4Ot37LazdNbFGLyxey
kIK0rSGlkq1i8GBvVWZL9HaNDq78zDyzVRZB4KXCY8G1uPxpQvO6bNXhbyqxW5mcoGpHP0Kmzj5z
eQRzPoNDLsIE2rPZQhm9Yv2rK1wKDEppRoIxrkUPQ09G9Akv0m5Mn903lghA3v2IL8rqpkNFWbcG
RVQes+uJuZXZc1V/y5U8TX1jfviWiYsKPn4nswk75dSsnlcig+D0WuGdg866F99S553CiQWOwwqW
0kyUzPDXzCn7QsASbLuBDUGx4bZcocMbknM04p/oJ/vf7Dl658uCBuhp067/o/shDGXwuQGsQQCL
gDoWeaVw7Lq6X1CN2a/bY1i9u0iY2QHo3ASBPY+BslGlPofvST4MAjX9h0DrkqyXXuoE6jORx40Q
d6zIVe0Or5y86t4sCB7ZS/WociM9I6sd0ShNeLClgeAvon4Y5+aw6LrSNGCLLwiRL+orNKOPaVAR
efXKKkDCTNhQRCBgWYq8N3TbuizSeOwhQ+fWxnbFUw+rIEjUR1dh3ndaKbrMcca2sKv0ysjKoDyJ
icr9o5yf2Sb+mDqWbV9UrN6u3Sw4jbxbrcs3CagTBg2riRAFkJm7yt841UDaGoXEN9i9V57qv8QI
J9JvJdohMBV4FYKWoCiTUe5dS8V+hg4KtZEidBLzENHCL7TzoYGKtEns4as1vlmtjOAEOHlAr2vC
IRmGwDFOMVdKC6K3wNtshO87NWR4Y6NZulkZOgKOnk8pHwj/iRNoEbjVb+B59LZ3g81gKAgE7VHM
Yq5rN1Q8zTTS4TtySbX59OAqn/oVjRJ1dOW9FX3bJtQ/Hlmi7Ep7kEdYsMbB3ji54CuFXn9Ffg/D
m11sGFXwrDFKX7Kj72Vkdi/A7K5evrVq/ma6rRPStUwUzyBLeQEjOpg+7b8VqV5Kp/aVw2HkdQCN
HQwWAFOqfFTBUVtXbXZBM4GIC3MXmJkjzQYowMK6+asv6C5729fNkZy1WCYIDnbjPFGcUrmkN5GC
lXxnY0tbM1mgst1VYTtsAiLI54GJFxF76SfcCFoJR/SSm89aO4TPPxyfDD6WGh/kQOPKCcZwrqkv
D71ADgjPHKalmKzYYRi44vQxZtHS1UKIVRuTYZsNEXQQEKFPPO0LCBChckeUC9JYSCPjMsnQa0n3
bkfA4KmN6++AuK/egCELq3akO2d38XmE1P5i0/doX8kf9hwD5WeZbdVU1/YUVlcMpBqC7VNrMP+C
Zz8aycC74kA3lGFbdhXHPt3mlPRDORfpNMJMI9bYGs6lOsUOCwvJ0UMYsz0WWlLZE1lFFaoP25GU
7goGervt/JRt5vE6/X1eMMdPxanW3Z/pNr/DIYm+rXygwdl/D4LP5JA+EXqlOZEc6hkYgsaUMQbI
+Lr0cdR2eDrzbr4jMSwiyt0xfU9eKK47J1xLXzPa2x9DGJKmgA1aRQw+R3VUYR6QsotWDoDhZ5mN
6UOTTvLLZ/rAC8FWPryJE2bdQm1lfs/UTO7pLICpFEC9wxIoLO9H1arz3JHzvV8S/D/hnmKuumSG
XVi0UQuJ9CShgpF27UMveATgfAtnpwtzoXhV0tga82Jyp0Tg+LDqxRhy06h7nADaVvQ/z0/qmkjZ
4zNKvfDIGBrVaB/2uMZL8KoiH0EN29BgL7GYlauqJpe1oFJkApGC6AET7vZ198ihsM4bE4SdMXeM
519xqZXL6r7P3usmunRgs6ByJHV9H7DeQ4ya2UOwqc69qxgAlgYWh4CglZe/furvcH8NxtMwUZ1l
vGOkOHhOUirJiwnrDCvei9wB9s2ylofA+CQ3faQRhBSSJYuJE42F8ZNUCRAaoYluKlcJGjwJ5fXm
2BNnwvvxaMm5jwGdGxJBACgg0wqUeW2/5QQLNh7wwBcMBvSzA2QWB9jPaIm7kFTtt3h6iF+cgmlW
/rtqYXU9Kwq2eNfcvgh5pKKkquSu1hVOauZyDM5zaJklK4ophhCGFs0zLH65qBhJI8rsxIpbckUj
/eZn+2O5FEB2hHPu8XM67hHR1/VKBy5QvCKPZkqMEQB4zk5hccvqMWBCr2JeHmSud+fSy7KmOK4I
39CbTFQwz1KoR6CaRM/VST+MkCqREj96/Ma9b+M0l+GPU4EbT7ptze55gI8EQGgUMQm9LHkW80nF
Tu9k9XWBiEPv22lFZOWG6T8zlpn0JU7D8n9OI55ZD7HewlNv1MZVg50ZEEfrIACA98dWIV1wB8+/
0UBwMKjJNHi9eSVkKO0E9T5aIzBh5+KuEXD15eTBadwv06Xo9NlkNzjbc8bR2Oef5Ljf1yFflniP
ofMJ0oMkTlrD7LzTGzSlBdCrTFDrnnADViNYXV6N9J6UFxh62nQ2Qj8NL77UDzUSbLo9RyDnFGD9
EIpr8iXtVo48T3OmFcPbSleLC4sKaOORGz3vUo9ZT0NmO9NLYCIlyAFb525IvfMyJ6IGJ5Zjp1DU
KAiTn8ihy6whp/f2vRZ+L91Qupzdh/HR4U4awgTqJhVqFCwUn/aVak7JDZy4mqIYBHflpM3Ex3hd
xYMI3+P1eM/AIrCo6WvvVrjCZjUypDbhQf2SDISdHZkEiI/uZfhmldlMI4cs7vt/C/vn7smdC57u
ufdXz/gxrQIZKwm7DH+1E9UOg0QAMMmDdxwUvz5F0DLyJUxcX0L1oBnxRUjC+dEJ2R0fGexyMdqY
rLnyxtDnhjrr7tmtfeoZjzYv26SkSmWpJvxKmh7zglSbKUHC0Z+SNDrwN0P1zCvHa5aZ9zYhWHoi
44JXR0Gwfv80JTRVpB5gjGXUzojRxlxj2JSFIxSJH3rgTa6GAsdUkJSyS3K3kzSdATooa9S7njc1
oq3iLE2IORlPSxmL3sdRuCG69t173uzLCQ5PscEFuTEQ9sB74W5lKWxIrWXv/XQiOeGznSpJZQxk
hBNDlaAUSQH2Bim6xHoH/1hQV3KtnZWfV5L0Dgkrs1CRL9qOCkTnVYmFOKhEbY6RvVopswh9db3v
zSgCFqecSo4mCFMSjfJOwGZYTo/W5dsvcYvaZdJExlcokYI6x4FtrZ7RI/SF9S2a0Jtl1INFqQWw
xEidJ8URBv3+YzhE8nSORMfmt9OefW9YBV0zCBKLJFbeFWtlj7I5MemuC1nbJqS4BeqSXIp4aQlI
h/e3Cr+LKOShP91sGBeDiGM2qWXo5aGnG3J3rSGNbJJVuIZ9VtyLx7FuoG7KYNSbd8/B5KDWPyrK
MHAp7k06ti3LAsz6vXa2JfndJQrHHBC/9AjcqM45evS9RfmWTMNmK0rb3Ze0xRQrNvqWFXEM6H70
ciFIplYvwKvm26io1doP3KO1vG0v6wXq/cI71mDkmJbQuQgPG+A9ZZeU2QjPR9H+0O6kNdhaovD+
vTK/7zfgOyJxmWsuyyEuH2gJ4PRhAtwGbx0AcNzOEmJlRqTVDhMA0ilYwIf2tXbZlFEFMYtRiYaA
41RmRNIlBfDQwxelEWg4Fs/Y2yjtLs4iYI77cQNIpWfPX9UckQbW/ikGfkzZ+Vnu2dWAGfYm+tTW
/klJQ4v4v6Ujohade0YQ16t+PpG24nlCx/dPbp8GpRhtupoF15c2L+oOUh1g0mRqMHDMvxth1KFt
LDsqWtxF+hUaGVvm3cW+dwkOXlpmmH7D0Fih8tCI+VoD5A+D742qFqwHWr9PLF0d0ZOakj8883Mb
qlAp2W1JVdZrKSLip4k4a/5C+yyJtuhmldNeChET9/nTyADsQNADkGGMWIQd+kYFagHAS8yNQ6hd
PjIroxAc2NZpvzCblv1mYRDD61Ics0jXMPu+u33Kp5e4ihCsJP2LYdhiqPPls/kfGwybPF1DmpUv
AsfLER64kfstFZU4yqDf08KnlrjPwcCZ48smQm1upUM0ZGN7VCRiYMhgL/3wdpAanv5hE2Ofr6dH
ge/wAK7EoD5X26D36hlWHgx5vvgtPTIRnznN5AosdAjpCQqUyKcG/vnOjhTFqpKvGJbtyZa3Wzpr
MbuSLKskIVmF3/pla2flXvL1GY/1WAB7HwrQKxPyC8A6BhmpBdE0L4sy+q/UG8douwoQJq0W4nHl
/y16iBvot9hwBOxmLrAAJ+Th41YDC6I/KDlWnQs6YOMRrfvF7slUKPyTwVARVWRpEHDKd1bo4/go
ztmACXLYmuoIij4yVsWbZFocwoXWNa2MrieRfgKS0CKeZC16HrwpweEvgnZ4dyjpsCNHmR6JOCXX
/XamO7VVSMCmEUW+eV3KcfXIdOqptVwN6jSqutd9SgOZ6909SKy7JP0z1jwl92yfnjIdzqcH0tcC
7xhDiRmX+fg2eSW/IvCyzN/TzEmfjTKGF+3gFS7vZfOKFft48r0xoTUc8pHZ+1T/e3NapFzqawQA
o4zn/bH9aMoaXZ0tmtp3ZuKZ6e1jOe6Br9UxyVZDY7c9nRTc8FumuXRQ4g942gOWh2j1zK3pAtTB
r9hzEnOs0VSgV+FlD2Op4DvbXgn+if+6cnisuOxlLW7OTTeHFshgmlO+Jhe9m1LdRWwa3KaDvRAT
z2zupkIpuuE1/vTyxN8g1FgHfvRRNR7f8jkIimjTU0YScsyosQW9FGvgvxP/zpCDw+9ALVGyvvvx
FHDD8VsTNB3DG5hG4E3OSI9AuO8mPeBgcWEWMy7za8a2j0iiBqpqwmgleOvvarvAiRST/O651Zhp
uphq63QC5nOclGrKvAe2sCQQouJ83zUSZCneZLxywqJPFar2Lx55HLrDPDOL4G3B4gHktD+jwCqg
vnwF952kbWpvNztQgnqOaBk4Tk7Nj3bW9B9+Ie1Ji+mYO2Sbl058/qKNDHr009XHDb+qO4yJKUnN
MU5zHjhA4myJH1Fou3MoWd10F3wsKRoDd6D6+Om6KceY8s/Bc05H5GI39C0xbXZ6lSi6eDQrB66/
Hxs4s+Peugw/1URRA834sSmQIytRg/2fjaTBddbNxDoxVWrc9zQsRQjHhLnaYPK/lM0KTyG9DmA7
QwOnBAR+CvYTD4DIDrZowMrfGmLikiQ6fRo5QwpK4ixlodZ2k06yvGno98qeFUAKyk56k/WManzY
GCmCuQpahupsMvHuRyByS0i7ud4skHE0b8gYOMVgdwpAQ5toXVvvi4G2uRiTbBBEmxLSu5Yy4f5t
SyeTagh6usyTMnb9lbivsbqDfHHPCZrQKLMAvf4w6jjNndi1MG3S9zBWVndyEPRRsBCuNt3MBQii
6uOGG1Eoh1qdVtd4/cUh9i5njNOsrmoA/7sia0uUIRjeDq58SRUh5mQhFU6hPXyLyzFwnDtzwMK1
6K/xLMrAUKBAX0aWEl/uIlGGJ0Qp2nLj9BJuILfujGryQCnLr1an5w7RlvWfruQbInygKKAK8Y4n
ruxFQ82h7waZgTznqA8mk/1PnSx3hg49zp0IMtyGRpH448Egx0S1VOxBrv9vjmJ4q12pWwHSeChh
APKymYbo58+eG3lTTSLiCky8qPIoJdU5cQtpmcYHJdPm8/jivxBSufMBsVAE0vqWtIeQtFRjUwq4
BaTocF8MEp0hWnNOXqDpfo75o6wu2L9Coe2gmTnOSv3t7sQvd6dMJlqiL7y1KVQ6FOJFhKMuJ5gt
GXlTyLn3hPD+EfYE5vN+ir1Wq2W2sFpxKkvCVVfQF5BlWhoKCTXGlihbvLOQ+Obx4mu5Cdl/5Wq4
u5PJito/WyZcCKqYhlxEK+WBAfxA7KYLdYdCh/T6JpQOdQ3hkWP0FAx9HtlnDqPx52J7Con3VKbn
Z/MixQ4qDm+mHrRpRipaZUTVKyA/ykE4HDT8eMThhwQolEPq7jzNbESHqNHIdSnCF7WHQDrtmJvZ
OnfgCXMXdPGCB2Pgt9+075kbOu0EJJU4bhEEj/zwTv/rus3HKtmd5GDRam+yKT0wHX//sj2fvUAK
a8aPsNU6jGADiIXfjgNrDUEVzfbQhkCUUGK9AXqh5J718ZRgTeZnThof4ON+yR01FIP8JMp5wkVH
HhGhrOHZF9WgZfQKMi1hsq02a3PJe343oAfd2uc/LqxlHgUebser2yPzNzG+/ZjaIVzdfCvMFVms
r+4DtnGmmO1zDZDlO4cDn61dVC0abyxm+CABcMQqq56OsvjXFg8sucfGrqPSXCRKH4MUqu8FKJrQ
lMDkWFB632P4rkb8Xrq+0RhFBbpazV+9M5lryguYIrIi/MT3D2fQqDCGAP6AX1ufD2P1xfcFV4GQ
/Zi2YpSEmceP9GNpPKdu9sWCaVp9kDJ1laF6TSx61QILog7mBD88LeAmqgiHe0cUBWd990Wmi+yj
SKhNbZ9e2HYqoPgv6Btp9XDIdt0KRMmE7vHOSlj8EDyvtd06jqq5dxhR5qSoED3VsfHQq1Icu1Ff
ZvKM3cyzM94hX5jKhGyGk8k1oiyhOpiM4yyeIFhZG1m3UGdAe4HZdJNtw7vESz2oGQZkUhiiEFOm
OdFpoM9aJHd/dNg1l7TmpQJa67nuaeUTfKPz8uOtUWiLX/oXXlElMkXGxKDvZt2a0sYLtBzzrI2T
mxf8yKv6gKBs9+mmkIDz0jieXVtNGR/RdIwYuGwHlQu/Wllxm3IaPGadc1090o0TXxOkiJVxL32G
kCqaWqTsEr0fsQmytmTAxQc+iT+VFtmlSl3VjQcd0CgDwoAkoC0MX/f8XJdLG3yt9B4Jhcx1931X
f1LLA7s+6Rn9Z+tMwk1AOMslXHgtD/YSFluKWvRfvJh6tSsSs+rXG3C6dXtZcB4/NBTpyb0TiEN4
qoUROEwwJUvb5vYApvmZH4XEApUA5EyYUq6QVb/uE//gHUjZ5UwgKKh97mFHbyDkQ3sPn/fO3Dz4
rsI5mf1rDF2J4VasYwcDUdeKwljQHLMCPvmoYmDiZhEjghqnDTcp/cVrxsfj25YXAKtfiGKEdngH
hPGUZY1IY9aLmDCJO1QUBPXJmB4J4cf2OZ5nMIgYqoXTRAca8gape3i7iQAtoMM/esj/0lEo7Fdg
XwfaraafCeQyqNatETZ4m3kAvvI1XrdzOTbAnMkc56UsgHWaGvzORGjpYMSEtSaHy00sizvXcGgR
P0y/8qX8VuZgbV1sWnGIUw51JKknhk0FvTX+QD2VL1Hi53/kMcJFvNNGOJlivtSplFPaP/Y0dvLu
QQgaAPwAwxKJArXvxO8VjLCAn6OqEhkY/lAu7X6tN0KQ2KEf+WIb6gySmQ1UpYCCNd+7A28S/j81
T8XgUOFGCpu9RLC7EhstqBvqvn4d+1qXyvuNWqjzDkTy4ZsGBtmMLbhhqephxBM5ZzJ4jy08Rt/J
xdN3ksmvIM+xhA5o2Oss/TI2rBhYvQYuTRjnVa6Jk4DZ4J/4bHtaxltQdUEZXLNjez2/K1Nj62N9
/Vfq+dloc862x+Q3eRYqhFes38yzLUZsZRMHjjkAn8uf63QtGT5QnqudK1TQkOecLNDDtNe501gw
X+ZZSa7ZoJnP0goNkhVU09aGU7BeZbVOXuGXdysGLzfJxvOsSKDWftwKdy4u8eKmdbPyMQg5M98g
2issb3U4uQWhuAJb6AE2aFKJJlgHsrJhgEXo3FMjGiP2afY5tGPpZwVtMhot1DXfa0LdsuVhV/5n
Zvsp47n7F9L8JlJKpxurD0JjgdRdEAIXxD8ZWnwTr/Iw/u0WQZd+iAGUh0m9tNipuDj598BTkf+s
XmKr4pmxgQ8ZqQ+aQWA/68MWZfK2gLIvADWns4FmaL5z6Xtn4gnX5+6CgFb1VSb7Pq5GxVcwtgXJ
hwzXtBGZhFxS3GOx02hqV1DM6pWYgXrEaVvwEIdsr0ntXE0tI1kx4xUchKqOT68DlTolAe9E5Ifa
ZQ1tuiybHSzw6Fznhjb4jIb13N6h/7JUi4QqF3s5bsY3QE6hShyO3AzL/0M4vofCJu+ll9eo0PI8
531hhSrSc/KFAbf7dLc+volSLemJbTHzNt2wjpY6Iw1CqHWPFpH4Z6Ks5eAqtqTXk6quN5QvSFG3
oDiYnMZGCZHXhylK6hcJsgis3vMVahgr7s8Tq5xUICRrHCFhcyMQMphrUaqjaBJrZWMp3Dnpq7l6
4H0TEEmjtal2vPmyXDuBkWLBzl/AYbjvkALegkNY/w8XWmfMtCv7T6j1T1SYpFfXFfK8+RqNKZ8x
o9naRCJ97Q/E3ud9N+gJc1zEI8zrljTaw9w2CJMT2zkcIs5piD/a9TLqwd73vb79QQpch9UViWVC
ECxjy8Lu5a1jXHj6Dl4UhUb8qjWrx9aPUu38M3RX+x1djmWHeKw0/44XwvjZpLl0aX3wqG6Dx6f6
nM9HZ86ztxPECFYcPd5Za2aIKjsh2wz3MTjjaJHCs8M2wA8UKpSEqUMjO8uKgZXORrCBEsJeTck9
0R+bozXv/Ehug3whz4kl00KbIU8Ak5qRuF6Tg66l1/pgARg6zyhGH9YGwajpgixeH9a3u7OCwTEh
oN31P71bf9FHoIwvKYq/9YKMYzD7gunJyIgcfCazgW3ZbH74Q8sjhl2lqmQkBtY26wlwZfViCvtQ
KHqsbnyXUy6ACI6D9PY7/6pWTQ4VXj8ZrCo0NWJQUKNPcOTF0UXeVbSEUwzLoHXKl+dkAbNTdP80
ZqZGmPt2TXZzMIhKSfBj0CrJD26T5BWW9PANzIc8GhOqn53oH4rSS1nULP4kLchOuAJKa/66gU3g
6yWixVCXqHhUgpC+F1EbPnjPtseUo++UkYiQqzuXoVnzY4+KPDjG2boqzeNeZN4zPqKu1zIUgXkN
BUFAIbrSb264aL608oJcZ3if9mtHmo311BDOXKwPbSp0h1iAfspE70xfDaDncZ9VplVTYn04zfZx
EcTM0Erj6G0E7uQXmXCBxkj4njR8ByZmoj2opWodLwfZKqEgAyH65P7GzhOufPCCNalBgsHFcHpx
FaNsUouGztGu3OWHixcEyRDTqHK/1BcFgZrx+9s3dU4gptVtEh8Lf1yHh3y3RkZ2Nw/hn3qkObH/
KnfGdvPUABsUnNdb29chYC3mXoXt1OACWU/atD4qGBQe5fEojW+nA02OawG058HCq6RvUVlrAfjm
gaUp6wDde7C0iRF/S767YSSEXU6mTNTcUHXSPz9esoNrbzxc73oKqcAOBl/BLNgJ5Pzau3Tk4mZr
bWUTULMnT8B2iSSM/JI42HesUhpd37U2h/MoRKoD/Y7ybtwknibJmb5ygokw/KL5Hn4cTrXQjXWi
UiNNa0sVfB7BC9VNbAjkZEDU4s6CCP08Wu8Qdxoi2uPb3PntimyTwfxzd60Bmr52h+Gqp2WcFWG7
4mL/R12qGi3+WT7LuBnqSX0454zsWELBHV4WCy/Ca6lLS2NUiSRh6v480wqEArXYQltDedhaDyjR
Db6xArgtmuxzCENByIPD3Pn1cAZkh+WlVOAQZ0Et71VE7d1eTAa7wZBfkl/qNjbRjQcc2FJxkkZR
teB5OuAVb8VvNeZs/iMP0vuicpJ6mG9MhrjWYPRC5mzDYmjrePuUNxHxFTCYRa+IVXL5/R+jFLFW
XcIldFxv2a7+Hm4rvBuJB3pbwR0dKCJ1Z4y/2S9bL5GxXsPjx4YETkIx6gcbRKqe6o9F8vbLDRqg
Ls+og6QB5jeizYg/rbm6uKWy4gkvMiTeAVdUo0G3ceg9ekTLYRh2ORQkReHvr8bY28ocemFyx79D
mhnHAzqgPoIG2xZTH3NzTaolTf0IHPE9/3z7RkyfNh+Y4Vci2YpqgJKMBiGoe7sWRH+gOK7K2Yqq
VmiGLYFn4hdjH41tbFO0fZpcOsuZptmbFOst5jxMg51vINGfRm/lALLinjcjgdnQVjLTlFVsP4zb
4ClHkpU2WEBsLMB/WGiMEHfbK5gd5SA1Oemyhr0K9sBVYelAfugXJ7k61F+ImC9mRNM40HbNIf/A
4S6xUs71/56dMBiMuHP/p4yOzv58aCHMZscKP8HQNQbffM1yaWSGgVd4qB19QMKDCZ9wzBrwuDQ8
xtBjSSAFw0jPAlzfI+SppPqOmV47jJVxL5LZhH2+OKMpTwMEEMPg1DSbjoyNUsbaCOXnSLhSesyF
E+gbK0BZ32MLF+HhZ8ij6cCcbcOitqbA0Ayag9H7Z190Vm1wq2f/qVSpaJLfPIsRyrgBvr+KhH8O
XATTz7vJVkm/6psNost5exxkt/rba3k6Hyy4AXwreaveAILNvIQszfvrm4Z5f5eR2iubtusWav+4
WlnfxrIJ1Diam/pIURtasi/AQHXIZickZo1EjvPXss3Z+4NU/pu5atYQ+zBDNfaSvhfNrcfIak9P
cpCK/H7JUYqb/6fjV2Jg8M/7jm6kz5ioeGQRC/C89hP3qJrRrqafypoCOG+15swEku0866rroWt7
cHKKrdRK2BvcQGUPK8YSBHF2PwYqz3SCIScJvVYzFjM4jWSOOow9QrmYDDdn6yNfp6c2blmj+MdI
WTDwQIp+tQq0pSw7sZrEGtC3ATWmXXrcBo5RZX9e6qT0b6xjOdeqX/TIAFkZ10NYeX1Ffh3YPm4c
4zt8Vciu8hSTMNvi0TelhEiKD8Xl2LD6ri6l4Ql+X9O2PIpaIH00VGnUNX/KPCfPlaa9p/nx3zAr
RNBAy0t3fIPmRUKWD1j7C1BSEiq6PvnAr8dWgVUB+DshsyGSHrUGfYJl7+VAcbofubDB1M2Ma2Gn
S7/ADZ6kzjtyOOwINWQeWQWLxw2597nfvoak2jrVkvlpN3ph/xyfaAoTLOkvyIgOj4TJcmh4a0fU
NZSWHn5pIrfRqQUQK2eERZFls7dMG1DwH7XYIvtn3Yc13/cRbiC3C9mATYvteJQjvMLuWbKuiB1t
7rqkXyMPcf+Ew5wsAYDzJocIfBvE5fT5Vl9MIGFLUMQeve+0D2hJugtJdkLg5QxwRySxXk2/iuUF
47fBjDOGgcJQfw0Izy+yJVBrMQo+gf1Owchbw8Eo95tgbOo5uHRkpuo4HugWs+vDky2X7xW3t/Xq
nXr/cOHiWXV/cH7G5xnx7ZqUnXWqNT04b4HPRd4hzZKaq7OJvKHLYY/o1pM0hhgPRoKPKl3z/NSC
aSw0kxD7WCElv57AuDe0aOPwJWuZKRD40cmoz72Q+4N87wAhXejgNiHUlJFPwC4zRjUIiZkV1dzv
qmA2WWf7kr+FrPr8W5GcAl3sYie2O7l+i5f9/ABkJMiMy0LqwFipHX8e94Q7by0x7f2gUvGi914P
0Fpj05t8EZf0RJkYxODYoPXg9/dXR21BBDTlkF+pdOOSzmIz6tjY3u08fxrP+Y3kzEh+ORWYp6Qj
oAfDnJ6Kr2KvN16vElVBPKIU2vSWww2FBXw7pPY1XWnqbwEj2M5aBy8l9H86sFs2U7PDoRp1WqUF
+VXlJjEFh6m35g3xTnP5lHkcl+MI1zh8iW8IDKHoqK5Ry7UKnvzeH7RsRl6JEDpuwlAEanJDooe6
p8uPO5bFUzHVMYz13N8q5g8XoO6aO/A2PJHQ933zyvrIPgdGR81XDwQWX0cPitqlupJXvUtdgYSQ
e38mMjCUGxY/IYGeEkEQmFhdwvHaXG888wOGNObtbbp5S5i4hTExqKfJX83bOUhbUZ/KsZ+EVk5j
Da1+kDm0VXAP0SlxlLmIlYKl2+oNguazAgggZc38GHdNV96KIrQOh7o73W0N1/dYaYBGBAPFZugM
GT3TqTw28U0u8ehJds2wxh74oihb/c9PE5pOQ1yVXwC8LZ7vqrTZU+c8bhRKHJgrE9YT1EDdk908
sdhSA2jxHa+AKbXclth7UrEkNAKPv45kK31WyrlezyP9usR+A6i0OJGSh6tGCmDkXAiXcV29QVcV
rs4NgNqPFPoSpS4cnRgUSnnyAQjo0wd74i0OYok91yfAja9gueLJkaBFxEeLX+WKwGM2w2Au5B0Z
Xu5eMRXq6TlnvXMj8mcbKcxvuM4c0htdDv7vfPgPU8463+2S6DROtNiQavTNpCmVGg968zIZXKo7
M5QFa85XptpqqaCrKCTtvPhx8DWsvD9WvnxTxQIlR/1wFZXktpZvoc+uM4XgCazCC+hVdEYwHMjC
TvsPQx9740859vpVCQ4jbLC8G0LjWZYX/hhcpU+EmJg9jgLSdjFEH4hIFM7Fcb3BEcOr3dDINc4e
NDVVmX13o9VGkI6XXKTuENynAlv0rQki/0Mytz4gOTNjpA3837ZBLjOT48uwD+GmrNyV+E/2mIuY
mbtp49U57NNCceHLJV88vStzceMgIEeNFF4IYwY/9fZbyvJtQ6bjcqI0sSTDGk9+o9/5imOdmZfA
mvnI5CrtrmfLCOThC3D62fMqvkq9OQrC7zyuCRUmU07REsEc3oLxo6A7/wHH3S/yP4ArD+Nrzm6A
txgJGgGWZ2Hczi7YKWOFGCQ7Mj2KjeRLZwC2CLKgrtXwb+2CkNPb8w8rrQKh/UcZPV/QW4D53Q8G
YYDaqR31i43K/AHI4KyI7tPxs2Fu1VwjC1JtEOy6LBCjFNH/Frfnx8PrC7csLWIx2xEp3V4v4AW8
FQzSYCfZPOIPx9+dCzaUIWRLgA/I9lYFXyJL5bFcA2/0PTAr/VcZT/9m61sVbFmm0K834Z/C0d6d
8A9zXj1XZfWe9oAORYvf8/zz0S9mWbTY08DOJglVsFgjtGtbv9n4A2JaNfql1ISqKLCpvpQ0JUJq
FI1wzpoE0SWsgcsfOf5efb/jJbGrMtbHMcPT/hHIvpfoXQ5D5HS3jGjxjOlTsRVSLfMrVLYAFyH2
4hwCaUuee1x4EuVIvfQs46UdhoBVM/aHFnOnN/u+SZAIQuKtzMcUfS0h0Eox/wXZhSXfuxQ+ZuQ0
cfae5lslSRA7+h/8eMKxmbd/KCag+HPjKcNpWwv76w3DgQggwbkVzhPj2DtSRvRWlsuX5h82TS1u
j4iBuWt9LHhcNyoYJ2zP24KSqvyTugI+hYY/icQEFE7LXC1jtit40jBoNiupFRcHfYZucUTscxwA
JNwt/9MuP30SYZHnDD+mKlVVtX0YhpdNu8d+BX5AhEGPhzbK+0vJCd0w2OWDdkiNfD2PIYU/YNA9
pDVSlEAZ4rDgKJ0+OASjbHAXsC33d9NQFV7rpdbHbhsfFcyJlxvyHxy6a7DeZUQk9Sn5h73YdE3e
LO8OB/fepHqM9WmBIT7h/gDmRjaNnWJgzgZcnzMp8+v/CRBSesoX43mgmQnHFrdf7cqkFapiHhWN
VpT19iuRNXCNflUSLOkTC7hNQ3cpqMIXc0144ECMiMqgbLZP1Si7lCXUxb1ms9Z7xCRPT42HxeTA
G74dGcNcdwlGH6NVuNNuZ5g7RjkcFfUfuv26Ze3veDWGJDkutoq+pF0HmcbWPe3dInF9QF6tLBOz
q9qOZr6gPIsJL9P9+pRVH/d1h6Exz3siU3cMB0sPOC/9ilN3aytJGcnGw7Mgx2Hz1qHXsbndv1m5
XhXxNapHlUj8gh7qkPsltmRn6mp0ZmdSALSleNTzlWpoMEZBSvYv019NnLfRefEuE3kKXp3/ztmc
o3AX5bEcdMFoC8//Ue8M/1CN8QO8F1kl960WJsmzP1Fxl3UJM7N9XBF2VSD83E7EkcYuvN9ugTpg
LkLXsNsgHN3/mjOi7mlYYpqo0mN0AgLu8O2+MDFarjiAGvmzfNRLjhIb0K2ZZAZSUhFn4gjhaHkS
Y99GBN5C5N03KPDKmt/++3s9jhB2ZTFd+OtH0USFIapM4Lu6OHkh0YmToxEEUaXC2GQu0pixCeqa
8gnlknOpDBg4TqEzWyZn1Dm7Z1RGkNBvkoqABz+TIPrzaAYuIJ/qvfVXN0XTovfBo7FCHC8lhAuM
8QD1k6qf/vl26I1nqK5d989bwki5tREx7GzqmmuMqSAMTd3oL53cpz06FqnOO7yxJIAwdPTOdMiC
yDLDlhEoUApgPOajEmI6Z0UCUFHyNpXSdVK9d+qZaushiK8gnQo5DwaO7UaeStgpcS9W155YTwZH
uePeiiv+mdGWy6BObLhm9jH1IjLNokaOhNYzS8hcLKLerHdcyssXuH8JweTsZkJtJ2seFMDMG4BQ
4k1vDZw62AtwnZkb84FxT1+abaFMFvADHkQuvLXnJ9EFT36wgIhnPHc3PoYlPomxaDH3BnJa03Xk
LdtB1ve0QVBbrYWu1SdYpGnd1Sg8HLWHbevoSAEKCFnBiW0CQnIOoVUdR5EQbWRo7ym+AAnA48vK
cB72oLZjqVaWHP3zxuXYAfHanIC/7u/12gq4wkjR80JQaRStCMXy3KmsGH0lLe9fq3PBqA7U+q25
YG7Nhd6mo8dcu26InM9m0IdZUIfyZHghYQy1rU64m5N2JRGMcwQ6+XBp2sVuu9jNfvsWsCHvq4VD
FP2G78RbwXAsG57HWzH9kYYhRsr59TezNgI/tGJ3r9R1O9++SGNsJa2ZqEA09Uyd29qD2u40T1Ib
fuIbkVSgEpoLEZRSBWUFVC31hmNvnmeL9aNo0Qz4264XzYxVDlNf4F2ndxL+32+bCOSXjXjB4cAy
lF2iWO3D2jpv/o3Mbm7QFOqwhnGQx0SbHNSxPcR7Xsa6KpUvwVdcOD6ImtFqc3KqWbk42AiZAw0g
1FbbiTxWO3FMt4emVORyMNHOAETeTdPx1jxbdj+GsP7CQuISSaM9s/7of1Q/yo/otGbxsWOUOfKX
HFdGPQnrY3Ly+wUBGKQ3/m3Bt0TXATVBovWLr4/OeYmeGLO30fosAIV4I4qHcj5JXgNmFK97T1El
TjdTQHviIap3MdfzOGLaBeJ9YkI4F0O/KRLxPf1vYiqQ842/9M4+kKoBz3w6PnQTcMIZqyijCJ+b
bBoxEgDlNzBlaEPNUto2D0jNh/7o87R08IBXJCjEjc7/qYL1aT9Co/Eo3Cq9GuuxzO2ZcvwFxK3I
AFroD/aIHkUqiXt2nTjQnCKqw3HtOtr+ohteAAZQOdt6jPjqdZFS0UoxkpibedP3I8LM+IjOwnJs
ejk/qYnePd9JfQ5RXMGnRh4J9fQyfjsdIg1ZkWxsayYvfndVHueSejuN26RGJ8FZ6dD+YZjpjfvu
iVW1MNEW7I27h5848sYeBn/gPwPY7XQ19IywPRZAak6+BXmenx6+tQmwmR93SOmR7vd3YtYTK19N
jZvzB6Joyp/HgORu+/1TQeDZD4mDjbzLxb7dBaXCowKORyVyL8tUYJxAB/3HNA+jGBxTA5mcrzQd
dnc8RGnGz9NoE/3OgdRt31M7Ym4fxUIF2fFvZBFZv2k4Q6ucT6apAxnxl7MuAuiHZeUviJJgqht8
rYsBK4gHl6pBPkRGeCYmUPUEKWi/gmrQQD/QW7PTAUGPn2trWrVTai5CtC4asRjQo4F5kpuiLeTX
6IkkLL8Jav3+Mo85Ye74VWB9xo3sk7FU6ELrkjFpyNpIwgapw0mBFnanMBm2jeqGoz5FCl0Ue6he
PzuBDwxReD0WeAxpgvIrti3tylGppmJpKVQfmi00rHX6SUUfGc80p1w79eMerXCfwFfCj8gXid1P
8BiYqJfFe6BAfD2vmr+7LXsBtO3Vk5DxjP/jxvvVfZZ9CadSjaKjOaAr6n9q0I1t3N0D7zUVSHoE
I/XQjTYCIY3ckHP/K+8dfqt5+a2ELya3pBwHuHKmKcHLCDqBZFbfaPZJhHbcDpcWy4CJbZPSBW9X
hMDKSlks7lZOKq00iKMxFhPU1qUrlyhO5HjxqzW5FtDmn/06B2sXIul70w7vUAgN67U2pTrhsegR
MioxAp+PnSTRQb+ADpeKArDKlYsvquD3AwsWDpX4wv8hqbkUdLFefgE6/inWb1DQMsX5lkNVYi9+
2jnOzzu/LkpWacVNeKRbWFTrSRvY46X4gxA3ojB7ZBVRe/F7t/heL31uaJecBxpn/1KoHDl9nhYM
wBDnGKTCflfLzX6hYk7uSfLfOl8it1QsBq4+hnu9/FBdU7PSEHriIjEJMc2TYudJcsNy/IsSKgeh
CslgeLWg/Tivqg19BtNNdQuSEXu70A+4mTbgDbhYfzgSetiHKFdkUvQ2BmQ+gZ091k8ccbbjGSHq
/Bt8baxTVeBxa0YFqA7SFKb+oAnMzrIheT7wpm91neh+YkyvWisvij7emQO5sfDfFrQGyLGUw5Vk
ax2w4Iq0OJOsO96wkZShS3lXC8e0ZIss0QKp0RG+mB5AAwZz3UDvKdRL8dYzUNbQLteMpPVhdGFc
HO7hdkHoDZonU3JUw+y7TVSjHbbhI8DRuzKCdz5/BvPbmIQEu9I57ES+UG1pMr19ocDCicEI5P+8
diRMPwtYf6CS9mC2g4SJm6FV3vA7kxJ2efAMrtLLRgrkIbI2Z+5/pqyFfgAELpO4UEnqzDYTTpR/
6nskSlSn+2UfOq5DTkuxffl5Ak9bE0JqbU0yTg9xZmyvPhQ/zAV6RfdOxrLI7n0XebO/tTGF0T+6
QY1qBsp4gYpJzysb5zn3phU/hgUx3SnWys6G7+D+QjBU/hVhy5AIoXa8YufyKmNNAiS87wpbEovA
+OucU2ljrD3qEB4rdEB/oZ2CEcxU8UyZIA5F3gAm3M1vqRshs2mWIyDKetbxtUu7sv1vZBAGPffi
BE/XfFmmtchhaX3o54amZGGTTOiEHYyrlXBoSLs7+jNzGqodp+JIAcYxm9wwe9qUHKTRG2EQIllZ
6Cjn1SiAaNNptap0nSLxWYeWk/73e58wptjBvlnM5CLcIugSQX6P0XyOvXn/sjYMDOy3Mfj3A6CY
9HRvHZipqaIEmYio9GgEfdS4LEL4qaKKxyUBOYPUkX6dJcHaLjwZ+dt7B/rqRzQ5ySVVj88xsKH5
nxFktTEJReOk+jKue5RkjjoR0e14AxvabmjgO3F3fEUHLQAZoo0Wjf0z+1xKo31s5/IvHRuPuOUh
9YkYgBBtEsyzL3xiFbBc17Rw/URtFrFQqmzMZAfILpe2d3sdGag5TK+/6GAFB4l2CPtG3TnAeXn0
pIeRf8mQa0xzo85Q/LlqLWm4kFeJpJ8/Ft9qcqJlBeJ0sdJt00zedGPmQuFWv1kY9QpIt60qYsLF
nvoY/i2r5gOWU4Zo1micuTyajX3s6imhCRDPB/8ZZFQlkgBWSiyaDGnS9Gu6JsXT+xRYKNZvgH5L
7vWzWRkc0gt5DVzIRn6R4FYtyzFdZvnxF9dB7gytzk3K6XFm0Qmp+y7gTtoNnJequ/6Av5oc6A8n
12W1QYU8BZhYuRdj2zTxi+lHXOvm72KfhTIw7XDhpNKP94PD7JDlRuYXOjTwcmR6KMgQYKubWWO/
DHFPTGtiz0sHX2uON8SWSawuljpipYe4KBg6YQMJCzWM/D4dw84oXlR02Et9VikZw7AWCYyLL0qL
jYb/lhnzHiiBjG78/78OIgFCeGlFts12E3a0CUzVIXZ2pL/0X+debqTWbav1FBJGdq0Dy46ePxTn
3qRxbgNSkmDhSK5Mehaf8CFk0qIiaCLF0fFZ0dREWqws0PMfYyuQeBt+SmaXU7RjfpPRwja5HM/S
ZKmtgbFPNntKQGgwK0MtDGlwVnNGywJgAOrsTyzx+8JspJXFD/IM/OWarH29VZWKSfo0d4P3v4D2
bZmHe72jdSgMP0V2qYlns4Umd6eGHM4rJkFGmYInC2V1mtyu5H/7kZbLYa/C8Nz/QcfjDF29LbPO
XcUJyNpHvtxfx/yX02H55qUObjBziZ8vJSGjlmzbbMZDGI5oUzU66EojSSAU3TItHPLTCKsHQW1Q
icHv8IRYd/w65ELW72rpQVLFT1tQoFGm00F+c4aLD2T2gNP0E9NH5a7JG4pr1USs34bNmOu3hZ5l
QWEG0cZG8YEVEFovDfi62+a/tNUO7gwzpMH7yBg1gcSTdnZuHND25kTMl+lLX4lYpX0isZtR69eB
N2tNKEgnZsNPpY/vO4jAC0osTDbL6cItSgHQ1aEQNmXJ1Jbi8r5ykwTwZi+/HXdIbpN9LZ7Jp8zt
eEKYg1UEJWjLwWQ53a6Kry0Zqt0M4GNz3fpOw/22XrD2kHpNc+d225rW5koedUmEbBnCrP0GOoLi
/rAmskOe8QM6VraAwp9d1LA9mHd7M5deRLl7lwYZ+bEx5HdTKkEvkGW6mQLoUUg1pSxrjIzsCDlF
CVxmHv18gGCWo4kHfhDZlPuJpzS7sH2Mwyy9DM/zW21yvrm1P22qYBAFJGZEJZxaNMM1BT3Z5CSZ
39RaMJiUUDbrkt8jJziTtV+C8tyV7T+o3rGjDxVb7Be0B6iV38R7vTOMtEJutDiiWEOosy0myl+7
ShOpj+5fDtwXQh99ixWjdfaedFmHqCPe+Ng5kX0OI8O0VABCZvdknqFmNjJ7cwyR5v/hfHS3501m
xkOpLm7iSHBXPE7gAn7JQKFT2TqzNxyt17cpu2exJzuryGUFM5p8X79R1HFAWuBvS6EJHNsaDh1X
we3M/faTWmFnuA/7lTrTANaNUCtYSZ6HoYOpd5rhdh2E50OKo3oMtG1g9qMmlloOmaAtLryr/icr
N0pNW0NHIoCWebKViLXSnG3dPjDcklRPfU8dkH0q0q0p/FSI8SKfAmNhixbSsdVmUZPln97dOFSO
FEx7QWjOJIcel9Zi4wbVr58aF5/mZLONXIYWh+Jl8v61LAxi5Ur0EHq8Y4fDebHy+BhCZgqqV3HQ
l//irHfdUgz3T4IWjTjMLde1UbJ3hGl9drD95dO1M8lNbv2l4cDFsYIu23C10DethQeg9lYuQHRT
ySDQN62lm6P2+5ZdsdIOnzrAl+Z7cfKRgnUHPbqeLmT+2POgbUL0NLStaku1uMNIHKJsmCd6eFYR
vL45wu8pUClkOUS+og7UNVZ/E1xjXGMsG34Te10BGMS+UPSM3JX4ACk/vjxllDq7WeNLiAeGdbYF
0Y28zdHs6NqYDRdFE5obO1bZ6ovrrVP88P8Sa3G2WnGmuBfzPwOzp4n9t7G+CE0XxefpGABqt87A
HTbnvwjqF8lkWvtHFRgBqrQzST0Lp4Y4Btw9ZaolBZqlrOkLgE/kvlvPJLeF4GXWWKlw3hT6KMqs
fAXkgZKlF3TR/33vZ5xI3+H/asONnEfY7iOoFhWXQ1ndUnjCUiO4S988HzqiwT9sNjKcuHuiPpvi
a1sV6UrVfKUnmxlTXjaIlzkzSuZDLZubnASdxE6o5+QaOGe5cx0bsa7Ef8dHmSk5XCZiNpSqHpro
QclA78WWcUgaO6bs9govbtCSU/k8kmMjnOCuF0+V7RXlj7COqebMjCOvu9XFGdsPQoCgdBe3J30e
XeNjDQMTxpWKeU9HdfOZ/fevN2WZc3BVUez2raWXL1iJAIoMWDEmpPDpRlrHcTY8SazeW6jksYNQ
nFv2zcuZARU67193sPM97P6gzdK2Plkc27qrWww78A0kzq46lH68cM7RS3/ro1ixeH0+OOGgonqu
+SlLmbW1RF+fFyIRdmMFBWLsd2nOoe6J1HbYYnqHAmt20rG83TMUKI2SenenvQKTPNgr36mdZGN6
NylNzxIfabMM/LpfcDqvj/96PYIYnvzXi8AuHQeDtCHbcc/ziEI11TOcU6L65yoBfFgE2RBzzVcf
DDvWGzZZ/kPfJsgm8xNB6NCyyjzer5m2qZb+F/qn5Bxpg3A2PhYbMGg6rwOz/hMtufkX+pvqVDB+
8GvDsl95v9revp42L6V/MDQe0JXq+oL5X/z021QY+TqWw1olMTfsJeC4X7YqCgH1XHEIbqxKQqdZ
g+fRWhvbjp4O+xyB2a+V0uxhNPNjU8p+Jjx2d6n5GsZDAWEUbdtreGQHwdteRhmYp2Dbis50TfLz
eaz/t5fR6sp8glYeYtWTCi8hrZUtyyXGcimZbRg2+pp4/DrJ68byHLIiwF4VQZzI/yNJHuZM9JnM
qfHmtPJ8DvjlbTvUeok8HPKypGw4lK29pTeAikt57YXojfj2idtZYGg5DIN8COEgbV3gWvOmeXaV
lhVIC3WiTInvi/99s9y9bxma+lm85eiFc+tv0M2kuHE80y37FXYNirdNSIIvkn6WO+tB48B76ex4
0tR+Zxje6O2OvgeWRC9kht+P5CIL2kCfsDSkZ8Kv5Nhun5Sn5GjuRmvdb2Ff2cEiMf/xOQarseA2
6VmhsQ+ov+64Ti8+8DJ62/g+PkFWRNudD9QMjKKx8vGxNQKbc0hlvxA8vVd7QCeQr3IkXMsOaE+f
tkMdih/4IVwkBZHpTcuiwf6gG3cziyJlR6l8GxoZ3jjbe1sUdt1JPoboxLWdLHVTjOd1pl3J1ZMQ
zOMScLm7XGmXh1uz6cMmvcsxK3pD2EWAx0DlmNjk52LBPhixMC4NOq399+dEtEJARW+tbdod975T
i2I/1aUjwm+4wlrNu/oFIZ9YwFuBdwRJD3s0GNcQddfCRb0Zzb7W0EeeT1vw1hqloO1FfKUXDFTq
QLEwASv3Do27XXQRn476/2EQUalvsmthKjrtI3NixBDA+Dw5T89AdmeVlkBmwl0r58XeWxp+PTVm
J0GCHtrubtbn5FROxZVjNABAgfw+RZKavmOTnlkwnmOpwNLBUwqkRXSv6qSc4a2Zxs1ZVWPAdffo
WOG4UIIJSI9SotlEe1WF8CZFLs7G4pC5doy2snVfZfyfxV0bs0Mc+lIru6tk6dN0gSNtCVKIInw2
3voJDga7CeIT9/2Q0SQ0KirxUPmVGKuMZ/5suRULi999aFrpbGBf9jVTINmpjmEGryCg0uEsHwxw
yARkj9yXY4gBUdBBXh4mj/XeaPAqUVcGOeYXE9Wa3sG1y6VRl2fN/YVGa6vjoj38Kjj+8GuW4Qs5
pAuqxMA0UR8EgwbwuzMf2s09KZTAA8ehb4mvO45vc9++VW5xPzolIvoMtJq0VnjuzAqILcdhsQjv
qbfFdEwNhihk8rYjkNzPRhNwNPNU3uevWN+DmwZDXq1hdWRtYETft4XH+DdH3g6AgGwqIGKd867t
4I9oeJp4QKb73rsH/1gOi3OmkeTbedpUAWgp6LtEmFrgK+TAE7U79ewgy2NNBMc5dCOgxmJdzV2b
RxSlUsjW23XApcfTjRWUhUhG0tc1iqq3mYGASahUkMWpmH3MUG071GEhRGNAXXXCw7CNkpUexKMh
pjQhDe+3Z/l4iRAUok72aG+IuS6b3gNelTNGDqJC2+Inp4HbTXvtZ4jmd6/w9V3pmvysLwA52MvP
X9YJVr834ygO5ZAaEqz2DaaI6kJOIrQJ++1ICmiuW40pk7tQav6Gl3Al1egCDw2U4FSoUGKosAIw
L0pDE7je4nqaMn4TzqwfIgG8FIHeZTVJbL+BLAfNLekkSOPy/qwdtB+gNCu4y1aQvXRS/OoeKp43
+K4ufR35+llFMI8PETlplVuVhyPCNhWxZ9OxmWvib1sPeTbkkzA7r0lA8CQ0rf0oSYT/HZmpjK6F
UWpV6b+xxF10FDv0WNIyu3z5kZrfHQdVxNG4/9JXwvu0okioYExO30KtjfkjBiP45MAhG+Nm6tZQ
djuKX/bkL7HFgBLgaXFgnSloshHoDvYVO4A736RyqjEr6TLsZ3tVPLbh2XIfeoVszlIiDaLDORRv
xMrgr6MPJwtCVaUj66aP7FfhswLbXj7fmyPQ45EJ7dEWGnLYNPctJdXienQs1gAZM9YpwHcTlHZp
gITIgUIF6IAPO8O8kLqwGq3MUdrQZbHDy77oQwVraAh2KtwyXBCjMDr6rxC7481nEVHQzdK9xgV4
a7xbStmNnfns+nAskCBZqe2wskFGCRAv1Q+sWUS/E2iea8oHUlg8llBD0p9WoapyK7c8wvov6a6Z
HctwugglCBHnp7xfzK4c7R0GOqKyHbAI47w7Mr8EV4PhRaneIZQ4Xfx0AyRGJZE0kLSdwoCpRXB6
DLXUNzAzt0dhn6ucbr6HopvIjePmnGZKNyjRv8X4mFiHWbo0y0MHrl8to4szMGtlcm0Vl6KopC/X
aiXsud+f+E9g3AhImf3sYjFyBXIeqMJOQEQz83wbKttmj/7I9vraRMG+p4nlFqp8v+MgcQ+J2QUy
snJeOgLr8VZcqNJrlfD6OHbOCI0X1tq2bqltmre9q43GEoTJBbuc5J7hdvBwFrw+S8OqVbO8dMUl
azhBAVLmQG7LXaxA+CeEBN9jiEQ2IHxoxeNE+CzN0/qcTh0+M3UlluYruUGfLyJjyoI56ovkXxQX
IPm4kWCrpCgMQ4jg2t5G3Hnfx2WIuZdowAo0XgnX13vHFIjtsnt8xeA5u+rxgyqJ2W7PBYGelE7O
XvF4LFfMQ41usKp91FzDhhFLmUdBfdti5tE84RO/ex0QTsAg7G89ZVf69ShG1A+iVWxZ89vrsOl4
kN8amR1+MRR7s2Ldqt2j4K+jnlcp+1L/9tKZDo+D/eqltCBl4dndh2l/WjsbOVs3avlUUpgZLqYf
M1hKVgFVV53P5t+6PSJ6Q37zNRk1yj9GIdMXu+vvKsJ0t1IM4wu6JmSoMgdIoUubAhICHDxgWlMz
q0PaY8PcEaWmFyZVjEEpn3LUTSqg8c/6WB44Og7NgM6qZLcecuE3xvcj+acC8LhK14vk0pmNni6e
/XIYsUq+T47I/WrRONJ1Lp1Thfro6Bf8GKnQTtonZAy+eurzq+UIvOWkdxeBvjKm4YAXlg6FZyx1
kWrXmHgjX+PATfJ+dPF0YVj3ptAg4/8AdjFVVkbCaveNUibKpnbax9HxuUyCAcArg1egK/J7+EkV
5A1QGI+z4q5cme3JG7wR4+5PiK5xrunEs3+HojXi+bN69qn14mXGMnzgUIi+b3Npay7BGWUF9s8u
QN2M+ibElmCvak2Nu8inqkpWUTX9cy33+P97O+ih+odraufaL6yKES5Lpswy8ivAdB5GFJxkJTPO
pSrIudTHQpKAI88EY2MFeka8W+v4RMOqnaDhsZxm4tXSHfhD/rymJ0PwNtGo8E6Vih1d0TWozhre
+GDshOD3LJ1Kiuj67ixTUBq/fRnaT3vOnZOMUlFv6Nl8Lpab/3LCwhpPejlSE/c8DDPYs6+H7X49
wxE7WdK8HiX8ydV+3W04bAKoHDbHRf/TSYYVPtWfp4M0UxphUVt7JcVIUx8WfiIIr16C3zsI6d7x
TBp/x+lPr0npCcCE+D5JKjz5D5YyLd2ZnOeZN1PeCw4pXwIuGL4L2srT+ST0SLJMfHM3DVsxpB7G
D1v44CupgkmoJp2RSe0P/75bOrbWyzUeMeGDmKuN8gWRFXfOHrR72LiMvTA7VzSPLanYYZoB7PCn
5tVyl6Dk+uHQlCr/yhwNpdi9bGJC5FtzejzrTkfFHMr9nibLwkWUMV0jQBJOoQ8lKbz3N0298PFu
XsTmsx3Qpx6DXSNBVah4JnDmgBGoBKao0RRPiL6WqvbYOl0HTEPV4GQGV5q9IQn/26VqyK25vBwg
u1VpaI0HiJFpUh16wKl+c2r4t6KKXbY8AryVRMmvv//U9i3iMzegPFdtq8MUx1MzYwYo4ONwgzuK
7FbX94N/yU9iV3i3GCT0vnpQFVoVkpFAk7J3JdF1pjmUiDHIrMc+SLnpW30AOGVK543FM+ACy8+W
ZzAcmm2OYwtOT6VUe0Pdeq5PkaVGkosDZxfsdJXZXbx+uPP1Q14BWZ90sjWbcmDhhAu2h9PV7uSK
MC+VfILWLzeD4D83NXWInneA4QBmCmPDbA6dP5dLIkhg5vyap8rlIOUn6eiko31zmhfiEgUnd0b9
Mw2+mqOwZOgMZS+EQyswXnGOT7Ka7q8i3aiRDr+b4tZnjYXE/WLkl1bKisvUygGmq0u5AKCr/tsL
DjcneUgkCri7hLheDwy05de+RBCvjZXavU11eXMAr2ATqUvnYIwaWJ48sYrAs2+33trvYjedxw/S
SP8EbkI3B3o96kUI35x7juiH8guqd+OWl/IZxtPmy8iGZOnca9XOD6+W5Hz1D4FGrX32JRARf3hO
+gNRc88XG+aL71D9RhEL8931tRONdmYUR3mtvHrffwvDFUc4Ul6AcbkI2MdrTUr8uxKdX4wP7a8I
O7lzkiqUNvrdH/k1w+mlrbmW1KSpKMgig5OrDzdznQJocNUy+rI5KWbrOmmqiLFB76o9rIFTP5X3
6KAmpp4u3tUO5RYAF45wJG0SVRTtVt5PLof2VFfmOOxx+hSg1KauI0PLuxo3yZx3vO+c2zN5Z/Ku
Eh7RG/hSWfXXHZ4YFiOQXrVk9oRrdFMkEO+SvIzRyeUHzb54N3nIVMHZgXl8EWpBVb3evNy3Im3A
uotEatErNGio3Z32x8kFnM3gWl/tLVqabClkQyCArFKtmX1Nw5vz9JA62RDIXJpFYqHzjuAfRRcv
9fO2iwNpNzWCXhc9lTnX1JdHqRiq4sLVjWIo+eYqpcS1S4b+HUFvpaZxMpvfmM7hDoZyZ4Jg7Qhp
kOQipoMyVODJcBcm2HsfSTs3mW4xazI4WiZyEOUYrIKaat/uP8tJ4GY/uvVir2uQH/UAGmaN8bl7
7V9jH63dHeiuMcKEJQA4rLWP+RJnBDumJ/g01dGIygzzy7rRWUlAYOlju9LHOF5pnDpwC3wmZxOn
X65rM7VKDClSOpCtjHkn0MiaBZmN3MpPFG1nLuMJsUGNQDvzfdqqktiq/sjOD4+Xoz+Cwv66g7V7
8ma1cfl0ALcIfAZp1AJdwjfCdrnFMAhRTrEwNDjaVnn/VNIM0yVwJZPcVT8DqRufGl8DN43E9QuY
7DEU28OLdD3hwtISgaXQIh3zlK18CbI10Xw3JZ7xHMNJm2nsY0RkZ8MqKOu+IRGpBCwJ5x3kKcZy
n2qoeCxX0DDSViOkmBX/v887vJU79RlQRa41afW8NlTMnCNpXjiXdm0uSlzRTHGtQzY+9g4ZOHvU
+jlvry6MJVT57+6f25GcoVaIjrwKs9uotl2MgmFVcuBCgpQ4zowIvlSrtA8QoxqEplySjZuJ3V3O
Yo7S8Hf7URCD6sIvIA+kjV6aLXKrw4yWuYfBZvgFJhuFzJWb+3XIqikGm9G+ZdiAFDVRB1LbbiQY
N1WjQNipMLgtcNvRcMykRTUxzYyi19NJHAtADlExGmQmrB7oCJXl5og3ajBBaReWVjwJv2smTRo9
GGAmUWLktdMG8LxwAC7zbDrJGLUtOfZ/JXpjorHaIMX5Px+NOvlkukXv1fQGU3cd7hg7d4R3flFj
a7mxeVtMzYhxkmnIhXQG8zerEYXSrdSylqx049oFUYZzlR0+Dldgszw8pi4nWyo9BR39rNRQorPB
ImmMERfbA2XMUuOhmbKZ3wxL1PfBJKzc0jikSSjrLApQ6cuxamGcrSpOCKygtG6TCsbI/Vpdej08
/biG34HTfRzhlm7jMCS8JHU+qJ/cW4yodKXs5Oay9CbDrbugZ7xN1H0T5hLfYAOPSJL36/XYg8Ba
VzW+kl416O6+ZkJiiAMp8NcScxC9PNpD05abRZYNYKSQJYaZoGV1fky/7pkvznkMhfANHeYUhT6h
LrJnkTniM8ZMLawSG8wGn3fwAWiQPTbr2mGVA4P3+XRq7ymKrd2SB1rCur7IFl7nmRKocWSUzJEh
ssxp/6JjYLzctK0SZcRiZ1UrUFYV0xJ+ePj8QsO0r4BQb2FqW5U+YxzOW29Wlg91Ph/8uasSnzKz
uhU2jjMjWWuNM05a7Hhjmf/rkxa5y3vDW0MIxssE/dgKAq/PursYeMYu6mxx9z7AspXzIHDq5Ctv
Ws6PKuyEm32/u2ELvLThcjGpSfau7eQaVXjq0N8z3GK7UrrsOoHP+j7yZXHft50FXYcOdP8otSLk
s1bGx2MZhP0iwCtVDjeFFmIaTlHFtnJ1oLGOrY3SV3rvkGK4n/PTTJvUxVjfImED/zHYa9LEiVwi
WCco2ovLdWvBj64uZ7IjzRg1FZ7ah+1YV6yVexy9rACoiUNkFinBD32i2vdrAdo9mvfTShMz2rSf
6+BGSU7AfHeQhdks25m9V9QU8Oh8CBWJqqoCKW6beCx2yhpzXxtRORgz/wrATRmVt4VuzrURwpeA
3kTWDqPqDcFQhjDB6BvnFOyKyxV+UD8r4lJWei4/32pT+5gc/Vvif6KWCsUUN9Wj1Dk4+wQsIf+R
4vNvsGALKLrYdhmJhyoRQcn1+f/H2rNnm0hX9YTm1DLUg+Y/f6Hacuv42G5ceuZm0ktRuamgcJSP
MqqgYEdr23fDoVmoCV5tC3+y6lNZiPfNGzh88v0JDc/aOL4QGu79ujSz+RoSqF+ZDJ2uE0sf9q12
vRXxFPslbJjTaixQcREEuWAG9Z+W4Wc0AuE9OoKOGEUXYzO11TEXggJkGFTR9oXfu5EBT+VUx+XY
6tDkBX29JLZ3u8a480JkL4En3j/olhkoEh1ex2Revt4mswlwvPuov0f+4xEdt0VvwNGdNzGT4aPo
XaFNV9Dmng1xPjjb3Yj8snuYfsa7tiGS2nf9DaWB9zLNGYAUhM84P/D8Q86ppUgszGoIdkLMZPrP
AZT8qZF9liK4sIVUcgYvxabUWM52kFfYaanK6mnz4tfdm3665XUB5VpYegBG2rL0iYKelUcwChWI
dQmWqF9xezNQt+dbujdGGpTo0Pbb9WgP7huBAYgazkVtlNrUBMkJyhFCIe/v/3ck3kSGHejBSgNc
hoHAqKvNSvBB+dTEDYSzF+iYpOJHNxVhY7AaMhW57Ljac4qqh4BDAsRWoR72Ur+4Ms4LEslM/Lip
LHIOcuM0USbWeGBTfWUtupaXFlxh55j60e5BP42zMeQw4O6C6fIBjQcTWN6K9EcdNbnaLQTiNMY5
DM8Dt4p0Ode108dOtQhwW9HG5AnQrn9DkJyMHib85lRMNLt+YVg4p2iKV2vUxCaODvFLlRjRLoy+
mpNnuDq5QG5P6Srv2gT0ROlna/ZDpY7ZSBOJF6dgo8+IRxK+g2MdeRvopvKFUIXPQCtl1Y2C+lYw
ijKdhYyf5O5PQEcD9QK6N80Aow08U/HKDpx/Jj33FtQB3X9qH4n8whUX4nualAAgi7WgZYA4gxaC
xN3uUfi9dccyJ13yLwmqiZkY+X8jpJ2JG24AO/gDq952Grwf6Qxk9Njl9FA4lKjXKztxaxL03daq
lNyIDtUqZdaJkCcGxi5GbsnngNHiMDxwnmxCn3tIdnJ/GqwQmIMJs/yMPH9CZwT1QF3FjHIXFrYD
DDwRBPQWj+OLqeSo2bilF9mxOxQg/ssNmbg9VsYjhueEdU7n2WDDHNJLYmyBKRQveKPT7rEXx/Oo
qfYnUS+uJFDU1eY7j9rWFtFU7NCg5/zYqG3XHBXuAu8iFZysxj8teA6ks4JTcqREC+FzqVdOwpsj
DSxXDPvX8naMOhrd+xU151JwxY+jSAkD6tUxikUdo+/RdPiItzGNi1N2WhKm+l0UPALjuQGHWYd1
XO6VwvTQDsYLAPKvzAOXdasrp09MutXxktodjDJOKo64neCzkEXGNLS8QUW9m08vF8wEcw8P+Gmc
dwwdDKgqKLpk7G2pmRWRmpFLy582O2qGtDQ6B/pEbhL1PPs9keH/bxKXQ3ZFqyfFcIDUWuvEwcaM
EJt5Qy/LzfNqYaODoqVliP/U1v1zEm9n5rJtqdvfMd6xgMb+QPfAvlxHunyPArkehnIl9Ra15C6H
ppoew7nzU8VC8vqyx1adD24Kzo88mcPwDkEnzYUXFfogL5eH1mtzHla0xicKmdwMlGAfJiWXq5Rg
SAnWmpYn/mJAPsGuyTdFBdRC+NeztbZ76lRDSxcnR9/qA6a286kP+CmenpoPoQAuhbWb4kVnwEeB
e2lKOL74TdhDKRhVuyYzf++N/0+pidpYS1DqPAHloHFkZuordTgfoJzPU2n4SltV2q0yjcp14sK8
wOFDoW+U01cmfnrbTPyJjB2wwW79gvAQHB09mofgI7WuIgTzKt8ZZE7u/Qb0T2iREio2m8kSgqx0
s3UMd3+35qVJZa2QVm3HmYNHs3vzrz/zSqx0mIZBr/Gd0sBSu3oUjQfE0iFHew+87NAzqiWC0z3n
o2pgmHgf1YyEnbcnMxmDxe53lesS/I5Dxm13kc+YomjQveCevtCKh9FBnmRL2Hlh457vHGP/CaVR
OyNjZydmHQW6iz1UTIeDwDv8Qz3y89oHSOqVWaShBd1gIXP8YI1mIpVIDoMkiPn13xkDKez6RKoh
aj99ACiRZrCJxfhIG5oKYknH+33y1tWwxLZKHwcOSGqLLuh/bllh4Gb+KRRbnIdfM6REcoAYvuTi
HWFAtyDRifYuB8x0sfcWF+cFBtiyrxKQ8+GIqEfNYTFQLeY+FXMzjveOGzIZEwKqpE70yZS7OFAe
ZAu+yCtS2A/IvOAHxEeElUF6QK9P2G9TQpg4xyzml+IlZkbFuvV3JrXVFvi9GYA1BW9C+gkytk0N
ZBbrmanYfAMUXPosm+T9RwD5YfogcQI68uainS+Shd6kxu/4+fU/uTtDKJcv1+HuLpJU2YvyUvbG
A/r1G1yUjdfe7ZH68ej8IZzbzZLXARcSYo0CSLndKMzpWNkxiOyzNKk0LZHHE3tKbUksl3PQPJ04
khKbQspfJoolW9EDCkDqsgFxWF0OUVq01aldni+v5GwNL7VLAE7AT8NUkjEKWiyLMANTcqfQmN+v
2CjFR1Iy+nImyA8jlT4Aibo9641Anliz5x9KQqY/aUavLGzFH2Do5aplz4QfsYns6gGR2gtVltCf
nw3m8OJrmz/YXeTcXYYrxnXmPPaEidcPyHDVx4HSQrlu40vAf2Uo2vXVyAnNSGVXVsFkQgGBGYgP
L75w+TGuIzrtdB2zlpe/KovSYBO9ejRXd1wyRq8XdXWF7l3MvgURYYXJfDb4x6Z63nIe7aMt+TqL
Yka/+/O463ALyw+6Cb4n5qr1z/VfSGv1IWtPZJgQyiHTW4RbN3ZoBBQSaW4LJW3Z4Ub6lhNZMpCJ
8dQ/GCuogPyhcBnMW7rjH1YCmZ1DPhD9ad3XopBRyNDjGo5lLiIOIVvzeFbTbps8A5qjwl9plLYr
4NfIX/QA9La5uRQlgtd3G7tenAiC7W7pYZOFNrL3TFTe11i3JaMMStvYMSiQJjmZfECJwKAojHFK
shManCQOoCMRCFQUeqBbFfK0i48aaB/g/Wksyq3T1xUJ730oP87SLYghmwI6gSR3nTfkGoDQSEFK
+Gi2JDqMBg1N3nZzREppL9qJlIlqLHoaWwKmBx00A6uZ840x2xe2Vcz9ARn/BtTI5QuK7ZhQdiYJ
e9FiSoQ3kNWNj1QGJrz0jQNCPmoea8hn22wr8en8TMjGefOfTSQShQXESfYKzOIxWldwkjYhN16A
zOAjpxlGb2JqHeXg1FceQwNQ+x4zmUzDUMYArBy4a6E907fT/yBSE6gjDhrCwcxIsC1FtHA+6eKr
sihliiyuzXQCzpWW0CTGwDdd17BUc/Z0kJ1Vdnz1dSSuQShZ0SCnYmVwxmlbu4eiSEtBibXxjGd8
BZZVnKmqQjg9wKV+yUcPuAOzvJxMY12DTy2RfwFRISW3Q3wERibaNeMm0/7TGF52qjaOF4fKnam4
kzG+J7N/VT3G0vDmihUWkIslPBGFVE3J5WQ7FEYe9d9PmZDe0FTcqkPlA2XCuhjJZfDMa7GDLwqp
JUMO/mEArr3hIIALecYN+DxiGaLEurmbEGctnvcBSSYvNd+Iq2OQX0XOUQ8jV6aaqu7YsmrRaSZU
EhwqYmxhO5fl+VYuE3cJuKU/3KgGwkewqWzboOtBZaYjH3z7RS3Mq0/l4fhmrCCwlcQnVOHaYVMD
glBzeUDVARSUwT8YJj1JX2AZMfCkh0yRWvOnU5MaRiTYYggIunXUAobXkJIu5zdhLo8SIYgFRN30
VGC12DQ9x3KNAD6/mw9npSSHbNA89oDZI+sXtnnon3sKfaJfik2pwepzYGYygVVvwSPOmBzNHQRG
mg7sijCT7B6lNIF9JCfGz4zVDNgink4Yp+o2R3H+r1QI6NabXWHY954oYjcjQsuZhklTlT1GNNFr
9w8DQ572Xs478vQTu9dGyYtrot3DQdrAa2D9AvyTahW/+NdZrfqzg1lHWv7mtVqQWECvJG65Xk74
u9ZTkiaJOs+Q+xWDn6cllntw9qnrtxlAKfV6Ao6cHAE/tNPgSJGGx+2UQLvXYXfGwfvo+2Ww/PEl
1t6Q9qdng4SwM65WUD234b1LrbgrTk+ay7j0OdWBuwLsz/JS+BRhTm7RcOal2jZvgNCO6NWm4mWd
A+FEuNlbZC+T8X/Rlcqc+iSjTTwfgFXkgoiuPJrxFwACmBcE3/zCrObNgoU0KFp9o8KhugAWPdFi
sTCSm9iVINauGHdj3lVbWGaPGxYgBgPwKL8evz53tQBoGOleW1QqaYvPqov1bsD3PfCCxRjKl+K6
OFSuYenIHVo1vBBysFBWs+Dy8/s2LvimCKxvyVupPy1AGBr1dgkowZ6FFDVP1+Vf3F2SAEqkSejO
4hhNvkvDg4MYu8w0izJUPWJ8GV4Msm1QaND/Wnz3gz9T6FvL+kDGbNemvuRpmkyEP3RgV7Bt5HAg
jUcr3Zj/9WPAXmpDpybqmcKJSK2p/xFVHJWYpbAZ6a/1zSBS/93PGoMz/1eJV6hmpHhMpP2NOMhK
CoJJqzteWMnrdM9FyLo2GvtZwyR7N8+VUDjdzPYkP3svDAEPsmhdLHetgpSv0Ymz3mhG+7nzTF4n
Nduba1c2b1nWNP3mTW6KUF4ZzjrApxI7H/qfcdzXpOhOSzFA9DhlswdCREMim23pwtViIRjjJI2Y
QPWlgAk0nZMsoYfRwa3rWbWchk/9wF2tFhFJaNc6YqZkqnrTJ3pUsE6LJUj8hqEoFEsqKBaoLxrg
BkPmxoClyLBbDNKdbb5mMd5QqGnywKzXR7ADDc8ZVEomQjUzb021YXCDc3dBoR0CxYUkSQ/Dl7/B
Z5nukTX1/lpQDyBu7Y86ZmXcuHF6aYHgbPrBdNRmUySIqLZV7cbdDfxaSBjCze9xvtseMbB6cjO2
lY6cAMTVUewWdaqyLICp8DkJ/WmqS6U59Zj+Bbt1FY9CEocwhI+lPD91XjjYu5Wnvh6jup59xu0F
k/rlsPdbdNp/8ZOjA9j5jwVM+36v+Nx/B8UNAKjsoAOm+Dml/wANyQI6wi7vzVQgwg/00ILNK9m8
LZKYHW2Emc3d4iFO9WgyB+VrBgvn+CELkmvtvW21X2DT+mZUaVz4CtAWBjBOkezRz/HVCVLvdMR/
9Vj8uw4lHjIqUj9YumZKRtTE0xSJCJFcIitobqffsdd23KMz3KWb2ZzYStPSzOc6pWS15NgRG0Iw
zARiJ7yL2iZL4iS98TXsL8tlCE0rc+VLeEN/v1ZB4tmblf86YwZedVNxd5ZH3VdZlfok+cdU4wE+
qqKpVqd01QTRahYKKJ1ZYs6tXXUzgQehl27kywvK8v8MSVhcLVjX2gW9fQPtjxgsxD2/oAOVpNpX
ZlsYHzNfETzk4ok3p+hxqicHajp7uY4HIbbXgJ0coxU225+84rAh9hzt61TYLNT1RfpyPP8OUf60
0GCo+mdXS+75t9s3DMemA0a6JbpIBZ8EJJ6nQx4GiN286Fspa3Z1lXcsNiiCGwrVS5OKFlEcZCdv
9F9JFxcgp+ASLFIfIxacTM2HLnryXO0dZVqhW2f3XMXmVzHFVWlXc9k8rJlaWKUrBe+4NcuWbpIS
VclyNiD0oWafTwe4vxwAvk5oOr02RnD3hxHRzToPLmdjdkRmsZCQFZHbd2eZf6sP2eLiCBecTkqV
nBaGzt7gMf5jhWwWPy1B1ZMayRW/VsaMEDO/Ktwboha7g8unWQAH8OwdXQZhTYW2cKIkUO5OY/dr
opd72HXgSdAj3emsAsY+qwu4dz6sTjBGlAoicb3ZxTUNg5Ihr14ak6xTOo40LbGelSn+FxNjTKEe
YP4oIfsWD9hDP79bsMTfMH3XdZxfxoa5mggZ4YPg1fGsMu2zpYXY61amXItHDA+32zFSFLcmj2du
ByqoavA9+6iD0Z6nJxLelTtTqnm3bOSUmCPFLY/xzC1JCcllu4qihgE/pdOIFjQ3w1nBYJwz+1ra
sQ6b0O6I4ulFLbam0eThhPbNJ5kni/HAnKoVOBngH2Nv6G8C2uy2nIfVmF2YC9WBBnsCRdBTezyo
4Ze0sqefFMgqhFczLnrRgwEXD4aAs28Oqh9ICHhUMkp+kL1RqYWPqKIClWdnhZBqikE42lMvUlWb
ImBYnEhwGTGfxQ/ddEnmzxyrx0wfwu0UxIKA8GX22o+UAkp3oO/tJkNyfmUNrZoQl2dfkkhmqiYA
s4nE/zIoTF2t8oxo3Q5AQ1Ibi0Rr2oXhVjZbeDzEJMswOihYbxU9iyLbRjMX0ktqOnfchbqXLV90
DrzlfCf1yWLrswps0qc1hLKsy1ErvXX2Itc4s0HeIzNUSwgmLWEJINydzyUctFTZlItj+woEmvze
DVQuEUkRYdmZSx9QYhA4FaDsVGFhOUknYxUEPCS3dYJCHfk7iET2PlfnU8xA25zHP6esdpjbH91x
y0d5pudj527RFtACh5kN9zL0lEs2KASx0Lu36TgEOf2h5THMdcPoXW94l67opd7zofWuJEOaeWMH
rZyaa3sjzFFgOY2snj4SBZpXoHc/RrwkiR5xXOXaqregn3is1OBABCvLvT4VW3QJRZZ5a7nvXLzF
8Xu5VlYdhW+i23Gyx4IF60z9EgAslY0mBTG81BoDkpnoeP1d3ctS9sjRr3oW5vulKtzHhBsLnhpM
XEGLXXCFzBHtFHVOZODbQU0G7lEz0nCeTxlwzKyov2YFmMQWJo9y6nrW32ohbE66Kz+dwwnU0jX7
3A+BqwtsjebNRZ3vmdpEJwGS4MbPUk/DPpL03WK9CqGRMPmztFp4QOfV8ebkZM3pNcs4t3OKAMxI
JinjCB1s1ABBOQ1T28C+xLwctyMhEjIwCXMx0y9cMZGi6/w2MEqP6XsLgbkGWRfTZDOVMbPljhFI
RbB7IljSn1k13b2LeIPJSQHXuifzF6HXhAN/V0g02xd1C5pHUxxMFlyPnvT7rDRfrTjU4xOdRtWS
GSS4p8gztkhh1MHMtJOJnQONGs8lllRz/3rxtxfPQXQTUDA0nmZLEjCSYR74Eh9jXDfZJWOYoQA8
UGuEBqP+flJx3B+VsPaBzfuZ2Wh366v/2FqAe4xUxhIus3al/SwITo3noG2GUzUS9Lm9koASxc4m
BVvGYsBdRsKpt0PsL3PS3RVOz7JfXVqJAI9ppAyZJHsQUWrcgwBTdOhq0vEQAB1snZOKpgk/RrV3
x0fNqyfsUsSuLlofHxtCxlX2dUB0qXNQ3Rq4oooNLRre32AX16QGnVdyXBSnEJUXsZvkJeguaWg0
AIaRjyjAM3BzJ2xYE7/BR5Ka9zqrLERR2POllZWnlMZalXhoDUJdZCvqWB+ReJDJp9BBN05Ju5qS
4WXNCD5+Gktc1Bwx7Mxjhdl4mdWVHIy0hBMfZawXBjB+r2jwVOfbkvUFCiJwYJmFzIZFz4fh8cRE
XOTKWi3e0qEcl7jvOK7mn/TEf6fC+I05svGYdrKuzOgzRwouBrxnas9tDrRBCGvrypVMrfB5A9VR
BCbbeegPSnfOC0iB1LIEcaIRCBTRFQSxJ3bixGUMwG1clT9phb+L6vLTwkLPu5n5hFLg7AgZW26l
JmP6N+ZFZA6ivd2ykPPPed7oJ867ka6I0//gSXTecZcVClkrBAMhyRif5MvBD87uw7F5+1AwiR7b
ILYc5Qox1Jf5MRVbgbvST8yQEB1vauwFeenAV83wRwv7uoHd6cyRi1A2sysZwI4N732GresG1Mpn
JlJJdFto89FQ6cKwg6yoFMua/zY+VdbK2cYOVZPo4wJuKZCwLph5meNSvB7QQJvgedEnXR5mHVU4
Pp0YjgYz2N6yg9vEytJFZupy913Woi3iu9S25o3d4f0VTjaxQhiHoO/HRgWOYn0Q1UGyfNmn7qqT
6PyHBzRdbgGj0NKTCdYtvYHNyPG2eCvBO3jRY/SOOLNmJyU2iu8+aoCP31uNEJuO61EVfEwSYlx+
jxk6ejHBHwnladw2qg9rhE+Ip4/ISM9qIdWnblDPQA1ZMf1nsmcaMySpQUc96YM9ZCsRt9JVwKnc
k4WMG/zQIBNo+L8yLXwSee2cltpOEvzKhC4NYtZ9WNEhfpqlYlBKUbQLF5LGD7baMjOXc0/0m9yr
n2jO+yC3kc0F3Mf/HkIKz+n4/u6d6e0nXchJ97Pv61mKlbtkcC0OnOe2pYDwx44h9I7xOWLTvgoF
IuMmwyjOU8cx45/h1tIbUKBi0Q5/DZW3ltQjW8KEjQkzr5sPN9aIWs/R2b9kNJSKcdD8XvpkvvF/
MRtHbccuHhAvKAWjHDxiOzzVdwZ0vEMSVD+TnbG7olkeiB+GvePSnnas9+b0XMWzIrhxtamGHChI
pOmrNtAVEb3WWu6kcsvDO3UFfF7uWSvtXURPj2Hc/7My+WTIs/anZC+axm4UN1TeuvC2qJkxlJyX
d2dU+VFNAJ697RraNS5KoZcG6FcbQxgbKwbSjA2gH495mPo9/HbSsfTNPy/fuUv4c7YF2G4vvo7D
bRPkWtwQILhj8verYzLpadbSrbcuyMjKQianbnIuaX4RzN+cxq6S0fO+U7RBQ48dkfvGYXYq5kB1
gPMnx9PzRBRtERUmmkmD6JBoqchjbowrrOsnyr8JBIvIVC6v8k7yBgaynwKvHOmXYBY+N8Fo+Xs0
4hkN8zve9kbACdLREHnw0MKP9mEPagfdQJFcpKYa4ljJH34vVYsXlHUS30Rd5ui5gKmfFX/RWC+h
RFRIwpEceNuXfNssjmLI0bVov+TrUfQ5O3n+MtW5aJ82L19vDO7XUdlH/oYMKlvX0RDh2gYKKE/F
G/JnXczMxAFoj6CXI7HvDsKgNn66f5T0cGpBaE7k1ajgTulQLGb3DUNUHvoL4sYDqm2WhceCc0lQ
O1Z+m+bQDaFcHTHbslzeQ1GKpzZ/qiewKO2wrFCcjsYZl+acqMwpw58vKpZ3RylIQljcofrVtZdS
ACme0nzFOCrI62+xEJUl5Bm8UAiRRPI8M8HzHWQxaa9SjruA0Ykul88GpSt2NUgBxD7M3cv81fB6
BQQ48wIyOnLfP7tGLwyiZN51eDeUOVI1dT/VI488QAP3niBLZOJTRq4j5/znEmeGkT1BXfL57DNA
KBJHeBLrR/UxJGZCMxmKAJ15P9IDG3Zb2aI5XB2O4ZTaJVbfnSmQGDJoHFKT/Zo8rPybXDy95pPp
SQomDoWzKOyEQaGSRj1wDQhxlHh+Y29L5igeZGGqCZn1ZcQ7SbkdaBkS0KUjAfqu7mgkApEqTQjs
kH0SsSZhsnH2OBGwPNfoVtJFhVfnzxG5FiAqmm5gkn8qAImJ7dB3eaKxdela9UDmaowtidgZefwo
FF4Iu41UyjGxshBADIkG8veV3fbMQkAujlWHwTHuF6jy3FfEdZJ/AZJd9gnnHY938ySNHW1uXtjn
VqTtfSFwFv7cyjt7Trr/FgHkQoELpL2hI8/nBVFMZh1ewsaiEg4ZWQMDXSztXenngZKIHXnKfeyx
57JtmrePTz3/a55tpQPiBtIzelnZPgzEzVyH8yjAJ2N7aatgp/QQVf2uWSUcgVuLrdMnxt1yGLkz
sNJR/6agcgnbJaNFZ8h708hQcL2DywOOJkrV6L35EtyxXfxoi7JrnwIzfzDsqawKbelIqAKjOLHw
8AFzW+hI1hE2xWJg8N/iLtawrWF3/wfbGTPaCB2DbeutH241qEi5auNByD8e1nlbrEDWUf6P+NrU
lyEt5FZqmndO9eNbVUPugITMTRV6Gsd/wiqXUZ3E5G/fmH9KOIy2zbSNUxLkyqOYH4yxMowY42Wa
oxIa7aY0xPvJasm2EUeVm/H5ofUqr0cxHJdEVSLSLLrWlu3a9AATY5ByZAzg60D0Iy8P/eOUiNHN
KmlcS6YH96DZUV0uI9D81XSs7kb/RawJl4HzTQ4nx5i76f7kkcQmA9YBOli/Hou/lb9Z5BNnR/Pv
HZC0TiV2I/OOHPJ4aqt5hRU4ZRfsuO/4ir8RLN8wpQt1iyPuZamkoghmwMvNOweKpOZ7FK203jd6
hDEArbDVCvs4Z8fTI5Hu2trGUSvIzGD9sATGu1t1yfyYX+vzR+SP5j/J39uV71tKaAeOLUYX7M0N
aakNYzPvyVUe2KKYOWcjqRXr77uLuWAVdsQmn02fcdt1Ii0Jpe6oLfqcy0d4PMTt7grW8rsGC9bS
PWorNl14h5mdr2kHGbJa8Az34rxk1DRuPiNy4TeKv5da8kfzo0BuQZ6FlEdZuSHQ7FctiEWyuMmw
XIkzaJfbJqZuNNM3GQUY9yCqY0F4S/DEbwno3uioBHo0sFbVmAaQ40j2RFLi40y9NpYbS8P9RIjS
Lu2KwsIIUZUSndCHdOlH9aDlPGmKR3XPSgKDiCijJTrg0bQ7RQL9YcS03a5n2qGacXi3URZa/r7M
OEpzwzWpaA2p8utIp/b4y2MC9Vh8obmYkJ5ySb3eLE+Rd2Q82abkq6b/R6BHq0c4dglMn2dIdlpL
H/85QyS7iPyNscOkRxRs/3TIqveAk6dYH8h2aBekd6oiO4Pik2PpLz4EL1MVgnejTMXi7GvWxIfp
A334SN5Nua4CoYrZ4NKrWGhAa7yXsAXSd+/FZpqAfI+UCwQyoFWZluD/wfenZHAp2LJU7L2gGMox
VWU/jhTJ+/VQJvZQHwwwk+lPQjnZV0ILDXBSiBAgYefJ3caAf/xDQ9aRHw8S7TjphvL7E+ig2fo7
l/qX2WLObG4AQTuhyqxGsm/s8SYh1HIIvCA/j78DvktXcA/NyCIdTbjOxi7b5MuHZgbQxxnoPZk8
B/qyKoBKJ0ay4pdyxXenlaaeNZ5lpgubdUy+4qOAD7vFNoMFdL4iqK12Cf6SGG0DBadYQP85wfqD
tHnKBSit+8QFJ4Eks0yqbZpp3NmW/jYqr/R7AdWD+TIIQKvmLeNlocszwCszai+M78YCks9QAR6l
y+S3Rhp+m8b9iFJlLRa5LlVcz7cQFwFeUl5V1dx8Xp2iSW1ROIuJRbPwvRinEQFUoU6kZrFOO6yY
HBI9MKp5jQaRHcYlb5QNB3w/LsPbUyrFWvP4uGTdqhnfcYDfFJgY8szSTP6ovDM5OybEO95nuAat
UGTgOlbFY2xdSh7eMKlHuCFoizv0M4x8m3MUNgixzu6dmOZqMmWEjUY807Ro7aCWYXskG0Mo9t1S
kpshVl1lZkWxhOBUGvWA/1PLTQETpQdugjpAyRT7I8KfvQXsPpFao9p9/+4/JZUHlEyTCKqAEvOF
hViaeLJvukueqXA0vi81Dr5wrCyV/dhRoLgYYUsa9sRvI/6pd9b4CN575hDx7pvfXo6cTbzB5Lbb
fNneqrBGep27meV/cCjXG7tLjVV3Xl3PudDujcjI1utGY8A1klrLFrQskhNAIxC0I/ELqX3JXOsu
juaoXJohkLYMNDvJapyODtusGGl5Xv2Txp5O+C9qsihND11SqOYg2AUJpeqCk3WuhKN6KVAyVzXi
/tW72+31p/cJHCNOfO8NOxLxmqD8peTiYeeBdroTMLd626dBftp52+WrWKw+KGJTb1IT2ENlco4+
QqD1FS7QJnhRJFkQOx1iK1nHeidpJ62LNBlBRr7uVrwDdRXlZWcUi6SOcQV2kixIsJKsrfb6A0bi
sgAGWF2nklF7rA0wccvHfCU5GWyNKBV/K9OuA/1a5pd4FveW9x9gyYHo3MNiHl8jPAT583rrIMIG
/AB7Ku11gL4Ta2r3ksBcpFfHnUiMfODi7Bk+2u6NpcEb+AAbL/+F5vxCt3QWXiUNJm3r08NvO3Y8
XsxqCzj/UqQKfBCxO0HtkssHkF2NcjXRDSxH6AFCvc17GVsvPMrGFdxl98pSFS1XO7pfG+gAYqX8
7KVmOo2gX/yZOMde/lhhwK6GU35xLIk6ecq5+CXrl/DwBZrb7vlyb8MBV1E8dbf+Xsillr40qcRf
VPjFGY61nJWp6Bn5PEhkSMbdCi9r2IJ1r9LmaYYWTsvrbgwHIdjMHMCZa5CkFwbIC2HFgk8GT0Eb
d2BD9D/cFAlZ4azWoSKy4kwWOV0cYChUmRwjTRGSV4fbYL1fIlUSa3NAvlUY320+8S0Vp/yY1dia
7vP3GW0fjkL70nJF2foaolnpCt9htgNJD0dGcritQnVlVD622DPZf5XFjsAhkWu8NVsAzWfkR5UT
qOQFLXmNrNc6xp/khdnSE1DqvAnltrvgRmvifHemHK9Ez1+NNz2I1IJuxojDCudPtp7yP9g22Dll
WzFSSxYbvy413YN6e7jXVeyGYOdcIzTO/ywSI1eVWk5KuKHQTGuvuiKoF1Ae8URLUp70E+wK9xN9
J3ePa5yHkrF1mrUY912hp8vEFmgsQPPWXito4W4fg4p06B5EFSnPH1iW9VYLYQ8tBdNBBbIGkc9X
JD77x8r0Imh2z74fcodvM/RmkH7f9vMZS9pj62HNq1VfB7yRywDFrM8nh+CyFS25hFbBthu8oeum
rMlO2gTjzs6KCk44bQYOmrJ8WygeeOHIZWiu/wfOcAjr9Va6ZB6UCTKuTLQGyfZ7rxxM0+gK2Vr/
tPVTTxaPEYVHAq0y/ZqLEMR6mjc8104T4NMue20BQMCIlR7ShLLz/uqIrjdAhfYK2+ND/tnAu1U/
44aZXyg8arteHjHUQHQREUE2D2Yb59wykiyRUJNbHl8rR+YCwqSDMVBKx90Rjhy6Z42t2gDoTJ2W
koEfAPTP8bLGPgjJty6dnivUW2DNZv2Cg+cFci0+Nf0t9LgngiffH5fKDp3/8JH64TFmZDsqyBT8
8r5qRUVJywgN9tOox9jiWhz6XFVV1YTsP7Lb20iSvQ+2xIlQ2EhpCwMGTGyApGnMzqIfvVtUvI+/
4CecW7sR2cPl/9aTZpUIOMy4jj+KMrzWzTx9go3iV9reiKU3SF4nxPJct6aQeZ4ReKs0ieWO9tj1
nPm3ondgjS2mOESJadPxfTCBgjLqykDHqIUB0TLn5GiXs5JrTJ07J6PcIjHlfk22Rah7PicBUhTc
SNoAaU0NeEhAEa4dUWZuL3gFcBgKq3rVrvU9f27wNapp4tlrgpmnh9oMG9PSsmSjSQh+gji6mpsm
BAwmFaHVT64fqJpNoZylZL9AvX25EcXxUZxLHaCSMP99Q6/nNuVVWnoKmSmxyzEylR/KcXTYMzVC
0gMxM1H8qz5pr5Bms2l28Ew5ILi19E3HiCeNO9HAej1JHMp+vh3JpTauyGQbYzpaUiLA7wd2/XXE
tOYtkOIcmzhqWvZTiGA3OvGms6fXMPTpOZsnMJXzpH9nZ23xAxwLGTHGQC6HTX1qDIRULuL4qPh1
0Ued6Al+DdJ5sZqqCEqHSRjh1th4VceMVjHNruPa68/KmCyiZjo6B9B2jgWJxkmO3PbpK6ylkRO0
5nQz6B1aWWqD29UcxBzUHRAGxG/qozVWUVW3W5QOC5NKhb/fWZ4wGWdZzIm2p0J/QOV6OG8lk6xE
VXqa/tQ/fweckre2Yuf9yI0Xpa96VpdOhTlmu8lEhac4ZxOHBijR2MQSlOJD4bRGFdmlvPUs/e5T
7501FDJCsXuSZOpAS8BdkS/lTM08jmH/lhn3m1ZcGy0vwV+3D0RiIbgzf6H+lNYNDuYD7WbwirZs
Zwpsgx2r79u9sEvT+AG3axC+rXApGs8PQ2QNlmHEX4euNqQPMpMTukp7EX79SiJZXgNOG1jKa7LA
9OwzEgaDI9LSvEeP3SGJmogxDGmhxQzIKdsnX7j0y2YcVSk3V6DdkMXfG2V2nK5kfKC55pP81xnu
NqSi9F8PUYw5ZdS3x9IrLyf2bV7GvADISd6tjaGAzUguwosVv5/CYlB67A08BF1PG57jFbVDV1H9
Z8awGeP2nEIPWS3A6mVfSZNXFjoKeWbSCkXiH8EIH9guxHf9NAvzAL/t0EDPooHom64yaK0O4Hfz
NzyeY0r8Bo9IGTHMCCaIwdT0EM5beRnSZlrIdI3yzjMxdQ7YV6lXlWb98Wh8YkfROPWOAoQZXBEn
ZVF5y1vFkTGlWZkt6JEt+WGQ76IFdofRMic7nqIHni/7RpLFwYenod1Zs9gMiN2H9rtmbIRndSzr
R8eSdvyexjsapaOW2GrwioGn4CmKnw5Bn84k/+9o25cJDC9DyriS/RpGkq1SttovrKv1v+x18GKQ
g6infQYjI/0nqrbX6cI8tlIT55t7vZbE2C2X2fMjQofOoFZl7b6NvjDTtloAxYDj7cc+26JwPXSw
Gzh2Xk4BeAyspuI19EgNYo6u4F6i9CbjWYfCDTiD918mo3TT+oew+W9bScEYCuBBO7UpZlN4I0Bc
5ui/BVUgcoE5SJA2g6TjSZ9RqQowqc6GqbbR0O7E0ghoUz2DsUAF99EX8GhoPwDtf+4lfPu4+DH8
6bJPK4DHbXVdbZQFMXYj+KknzeCRQ6cEtP1uXb7E8QGVC8w5caTbAOFHC+EC0b+KWn5VbmL/iRnW
d7x+fBCZiVmNs7XnslT2ABIHbjqbwTgCK1iaPoVNjj3rH2hUgghWSVO0xSrxlFcbjdgedxRoXEd3
Wdwukm10fBqhNI182/hSZRDA9AwOnhIe0jUcuMFjT5g8u4T6Wu/BRXwO3uLN6LyhkzkxTbbQoaK3
15w7MT1REtQkjyG/D8c1fAMLC+Xs5N6wnNmeQE4Wt/AYffKuNNNbV7CU19odfMl1rIENzxnfGFuJ
tdF0Jj9SxmOios/MFXPKdCMqQOm8Qs6kLcB7E0e53zh3H96VO6WiT+PvJe37g12jagnkgEn/TRty
l2ThLgI3EqoVSpqrdzEtmHDfI17eZcXawqN18zeFfCrPJd8/4ahBanIdJzGQQTbRtmgm5YizIuXd
YnKWiR7PgwyZ2Lnqy6VdimBdUYez2e/2XiXWNSi6FLUeTkSgEByoCkyqXpayh2rJnCmSXdhBXEFl
1UP0zfxiqyaDqr2+UcQlZXCAGKb9QH6uVtFPiHotBs03TnfG2yO94MmmQX7H6yms8Oz5akV0IOpr
x5Qses3O60uOE8cEGYro13vC0UXNx02EZkDaafyzp0F7wOalaA8S5niARpk+MtJJD4uJK30L+cSE
NAsJTriDKqkB6t+JxaeE+V6//7i8vVLWCuiQHlnhk3/++Fph+LUNhhSR1/LiI4OjRJvgjUwZWpNJ
lo7+TimI0mJfxAz/ga38Oc+jHI4X0uEuYADvrWgxXuYCTVl20qpF9+2mHNyEIBFwbepSFsf20BN7
+f02Ynw1RD5e2hKidGyMBwQFanMaHkYNKZhJtu2fmLJRnvKP7+AW4ktEpA26oATYSGhJtdfBa4nn
Fmk6zH6gstQdz2GYJQi28XsdYWyJW4PKBilvPb9bNLTNa91h8s+cGUqHH/fqNtpV+3lQ6uQF59xi
dorha8JZ3sFsn7dSt60kN75eERyZNjRAOYx6vujBrE5Sxrn7zdOWwKF+VPoqYtYpHpYxYNbVFnnH
mHiSiHPoMpnLaDrV/nza5GGfdwSaE3c3z2dpYk/XfZX+gYgahnmxqVUgnDGXOAQz4jmEbfUnnhHo
cNRrm6ngb3Mqw7ySigN5P5UEQ0zPQhgb0FaClvrG9WevHbPBMBjC0P1MMxs7XQhSyC1kTPbUmeOL
RvXQFxDuVJHAouAEvg2DzhC2DKhwka2KKluQ81/T8kg/dqv2LVoO7P7HoXZEZxjlxqUYI1V2KCKE
OH3aTBLzjfaTzTj1SXlivRVNIUmtFh6cR/FjThjUdMlDnvTlNCcbzfHKvEiAtzO0TwfbQm1jNMqL
hYTQad6JRaXVWolfOpUAcnhq6Er+dsGBWYP+DEZafcMbA75XyjRp8n7CAC3i5MZM3kq0FhFttCQs
xrALuoyo84E9+6JADT/pP1sGblWICqxwnNw/BOhuQfU/UlSmH6fAuOiwqHj6QPM4aO7qK2mjEdUK
ygd/EURf2IQgNVISUbPAsqt6DSxrNcKqYtw48A0sfIXyC3HaeJ4bDCCo5ah5nZR72S+ZNaNFlZ77
AGIcjGe+gQFSNUgpulETDkGwtIQVSCNUBGm/dCaS3D30YRoi/ruv2lzpOzeTEEsAYGJaLSeVBNM8
vGbAQjHTYfyET+fSInYwdJdrJKa0g2uHf7mHrDrphlOvK3QBqSbYLb5sPs5hqOfy+v22eXTVxtmD
DljDDE9VLwQjAlGQD+LI8J+mdQ4RX+HuVaWrHARVTYsm4+NIku+JThZB8B5fUAK2klYosvBUub7X
53drGHQ8Ye1vKSgvBNGPiwsbqIeDDpwINfycrrec64cdhdfZu/5SFDAf4jNJeRg2vmg4sz9kndcz
oDoesGGzQAjhzpZtANOpmO1o28q7Qw9cgPY65xLLrs4GSHPfmj//endi8e3LF95O5r5AScncQGRT
zKFeLkPxu02WVvxmIpo9ilXQFxxfmZ6cvEhyzEea+8GH1xJ2Q10CF1SwFki9UrwugbknkXc5YB/D
AQJ7D9Xmajm3zH/AUtw5mi9piCCINBhp6g2xafMtYtnj619M5WLwgaiMUHk50PK4MsOTLWp7nJdY
G25EvTiaQzFNxfVv3uzG0EyRg+YjprRF1g/C8IM8N0QFpqTPrsHFM0n4tYpogFNuEb42CQwxO3ji
e3SdmPWQ0rVS8rJr/z6OXb24HrYs0iu2+mg6vR/1Z6r6Yr9vUkMo+X9AFUj3nU9Hk9VeUvSDaZpW
AIG9r2U+xAZzYNxA/p9R1t0bp7uG7wdYaecCEJcMWipijKOt0VNYZrXEVDmSN5GdOI2vrRs2QbxU
rGwCaBTlT6ykrtTByG5Y6xGAvwaN7LWbbxqdhfXSaftJf4eNNA3mENf09r42S4d0Kg9lMnXrxLsQ
I85qqZ+z31HGBI1hX4y9XNWyeI0ik5ebNwU4/A5VKICOEw1DNeuHUACHV1IwFo/xeDvqYY1oFalK
UsLtlyQgR5O+aGVXHfFRoMPMRTOq95Mwc5WT2aOgKhXTg1xF4cg6e0W1cLsv2imWNQChfOKtNy+0
UcaZifDB/cN5UAcWx4fpShgT5Mabbl/wRmaVOP4fk19Bs9Lo3UO9qzveuVkWxGmdUM8HI8kxCYTn
wTe2LCpDkTxkE4I2WQpdjFEELKqKtKTg4TKDXEF3ugSb3pfHShx2J7N4oGxa3LvwLoScNRqxkHxL
a4gYmG38IKEV29+N0ZwzJgZZABnClz2pSEoecPIgwIgXahNaABktkx6w2JhKU+7GUo/IxSirwKk2
3PMfAFGyAEFVB30DP/9tGVxEdvIV0VgsL9f7frvTaGZLXuDMPjeG67KtDnjZAIwSinw/mZqorSWZ
jaW1XFjboJ7nrIWj3gTm47cL6yCeTWyLlmgRwsAqThh8R/LTbawt8E9cdtVYnADAwVBgw3QVsdAG
aUV3MixUgQzFdqzoviPLDOo2jjCAxaxkZtB/rg+i4MXa33YaA4ROXXL5jWYl+bPDBM0VMxDtQFZf
NB9qEjqz5y2CY1VOTOmvd0oFwMru1+le0AnkacXy3g5Rm5V9lZEGVpk/aSooXJhQ7hmJbCXrSVWH
tPzVj8P7tlRawr0H+AFHNZkQJaIKgAOvBiwfDOQLVhCu00CwihiO9/qM4o1/ubBtXFgWSv8QY1Iv
B/ZybrteR4k3E8GA1G2R3qliJF/yoK1/OyFqGqTI37SBVyM/m3n01wZYkSmu60oUzkQUzeRmhyrB
xKdHkFbvI5ee1TyDMVOX/hcwJqHN5stvQ8fV5TdCHzS4hEuWolPbOaCgGRxNMuJB3Y5LDGpdKG0C
UP6wGVkNaevYKcmmJSCggyc7nzqbRhHRBM4LaIVbTN04EarCx0odwjiH/M50CeVJ/vAdRQ5EHNtL
fGEzJnqEaC7K/77pdwlW4d8jQcFq9hSHt/Oy4YZhxGQBu/jC+7Jlez+F3W9WmFQm8V8HUPAfcryN
89I3lUMB3tZ8rWo07pJ/LdwRvza5541glE70+N8IPVoJCrQCa0endCKLTU2m4bghdRWT571ZAjHH
hA0jeBzPA1bhlQNuAVvVeZdyHFoxSHjADthQqhINJUqy8cyL4CyePpOq+Dy4j3xK1I2NrYi5OzC+
tA0M5FRady/vKvQLP3PZeFTF/tKYL73hN2q9rqrxhqHXXqZKVmgnMQT1pHrOZnKkSTMTc1j9Da1v
JSRq8drYHoUVGzN6Aul2IZ0UCWvUUiDqJe4YvwaRTwzfNlv1gypdHrBgfSW22LKcS8TG96xy9KVJ
9sqQ/5XfAi8HLshhNsCj2Bh8CsfD7HQlzF7UV7rKkxVywMBHxKHeIovdXYDQ3xKC1pCMKYV3zhOP
mTB0LszBz+qtfC/RB2GsZONBEzxQeJT8/n85J5fapsA2R1WgLoPQaC7GC3nzWQSuA8CWD2SYB5Lj
6HcNOY94qM1P93cSVVvnm+xL1AvBZcqcYCjxoWgG/viiGA3MRpdfioaQsr3JtxaIllYiwFHwqVyO
tQhYugKaStoJ/PDBIBPEXNGGbNod8nE9EbXOuF5ZoJNwrM0iJVQubk4uGoqTu8PkFMSF9ovUK6cq
PWVswDzXl9A91Os/HgqXvl+/aj5VJw5VhosmuAQFBPZ7EsyOAPQzLyuCOeOXaAJZppbVA7wMTA9U
SNBHwmA+seadIjPCO4YjdGnuMlUGL5RQ1PLYAEPlrlnK/4kvARePotY3HyvM3fGaqsH4sxko40XR
jLh6cfxo1PFMAmfssXViMy6eMqi6i9vQzal1rtZir3Q5v4CJtplsqHo5Ewu14UcpbLkLaO9g/UHs
QZZ7iy5Bt2U9rDzfs5fqWicDZxknD2qIA3gHYbCXMcL/SXEyFsPcewPaKJyRgKH7kRSMi+G748gK
3q2DuIrLdzF7uJLyo9VceyXKHAHg6lT2FVNOu4S0R60dZdSb63eHy8zAyqI+4uvVPS2yFOhn6Yb8
kpGKycUCFOPNJc/yNVr8lMfVt3fteYRj+Wy6rlrToPfyiKWovY39kTj8pJARVaQOtEIeQ7JJWqPJ
21+SYZ36gnVtd+oIpoO7Ubwa7PGbfY2ZXX8kNjEzmUXpZDH2zyI4uwZVdOCjudyCeyTq6kY6vvJZ
32oVwWMLav88wlbDvxjVNCE2WAezkeYIhKklQwvPQLCJeKQJZfBpWdvo+dMeI+OSFSpjIpR9wNu0
3Q2esooD2+5xnfpXJx20qKkNNXgDCLypNs67BYnm2a0B4LUXzh87OoXFMshezV6qCw3LH3n05MAO
FCTB0uxz3ibFQiBnDwb7AGpceC4bD+9f3eZR5k++Nl8ZkC2lR0Gln85p5U65iCsqwgj5HgSA9VTT
tLbHeB8dm+Efk6cyn/j6rnjEMTtqo4Xm+012SPo9OXiBGvUCpzL4kvTgtzflfzQWe3EFGSKfgj1C
8UlC6PggwmfJGxDFbaBNNHZPvZb3goW0+ooTaYNtGREZmMJejmakFcwPKkywFfbmVytn4mjRJH+l
7jhX54SF27VVWo3SJKBdT9sRHH0KPuqQkYSDTJiLRTFKVLS5jyLbtwFfSBSRNA/CC6LsW/786OlC
mqgKIGNEeQ91qzVm/kMuZ7XIpAftOay2q1oLLLliMgIiVVtqwJI+hG6v9ddg065VFny4kUSBsocC
g5LDeGu8FPbLRc0cOs5AL6BNm+lv/jbXIlNE5F93CwwbSVG6E4mIad0rjG1pXgTw2N1sJvT19+6U
nsZYfP1v4yR8R9UnrZOVUkkUmX5uKcXQM4DHGAVGZU1Xf5ds5dtItQQHvPpu3QOFYc0UTkl0q08a
oSbyflvkYeK8Z2h3vkXQeyM7YbBcrMuxZacST8W0Avfx/DDuUH1EJtXVZBN60FQBg+Euql+jKyFC
YwPh8xU8qa0YjR987ptaKaRUvFShY1h0FcWePRRG8eRHW8FWK87x7OYeWHQoC7stH0EgnXDCxJcd
y61DFY+WzpmhAeIUOU1i+w/bUZo9v7yBhby4K/GYtgssJqT/wmWnUFuvBFG8QQjK3WO1orghyLDR
6rBbXxfvRKhhIiuL29iSM/FjRrptm6XOVEK9Kuir+0ZkEM4TmUr4Mrf0LdXwMHoexoXLscasoBEa
UOrhPIrHXrpID68kmO0sxBqgFCAmNiLzEWCsg/ob/ZLYLpAyh0AyEkP9fVRYS8NiMi0qNcTpxai/
tYwjbVP8r+hiFSNnYCibP/grAVMpgja2fOSwFgavBrtr3uaHujk3gBnhUQdyqomKMjGU2u0dfwbf
UQasAvreIs+vT/9/PyuofDdFD/N4Lvol6DoHcWsBSFYaLv36sxAcy29zCidQERujVC+M0vMSoEV9
Nc3wth7AVIkaG1tABKnPyas2gu2jUfv+kVNrAzXZ8ioiyQReXVizJSM8tJ7T7abHCwfUuc7dLzhq
tebXsqE53fJXpiw8w2s1n3Da+chZHRo3qweNUZWqVEc7ATq93zlYq5vEFTCfJdWV471HkxiBbQ5s
zU1+jkeNkK1BbgXy8/VswBTDErbKQtqWXdyWJd7YnuuXSmvrJ2RJWc6lvlwc6yAHDFRAEARjYdlG
ireJXaDXehDFBF+3Hla4P64vB2OmbMzicO1w2UwMxrhOGVl6xny9E713g3sRiNFXu5EnZ79kEP+t
MJ4meshFVeDdBxv7z5IlJzJiea9KzzVrI9bQ/UxUr+E/nWQYdbUjMO/+PCmewURRhYzZE4/R0Dj0
4EPCDMHUev0rUaH4kJf9+v+NYtrJtDIlxPneH3sygFzYaW4B+2kltIBHk18LXMZLILPY9nseGrvi
MuFPuRtufoxawdKUWRGUTMKtePIRkPdaAPGrFD3XIxvjnzjrsVRo/3GSWVlTIYT2rpFmgZ0ygJ+t
HGR+wX0JLsLc4f1s4LimH1pb16BhV/rtqrmPpPFn0jHUI9a2qbbDegqdm65b5rsDcwIEv/zy3Z1B
9sfpOaHsKci4iptv5/MVrBN7A8powhQlmtcn9LyQJSs0hr+SuSFMyJ5RTuTOOqmhli31UM+2vsFI
nE2PtqwQt5HDJt4SCp3Rfuf8mU7hZhkWULuKAyiQyXmQ7VUzB5KHZWBRmmxjGfQePoMMimFtQUh3
hP91B3NZMSizf6BV8dEREwbSBf3XL+1ICNjTvJUPkRmjwlicaBZSegyUPIX3vZy/gZ2rpoLdtSUb
PA0/qQOq+Lv2cdyJMsxw/yjvMz6p3xLvbsy/iaKaY4YY4cOtkpRbL8bZ//l+0ZZCVv8glSmvAcUD
lpbAyes2DnQxioef2eG7kYu78VcQiJ8mdzpgby1r+lQNcl07gA2wPQbBP4N/xnoTCluCGyHXXwkV
AGVKDzZ8sW7+3RanuLAJQBh12Ym7AvwlbQSfN+SH+4eSmsx2JnyFKxsOn0HoBgRjFluzZ89XBPgg
7N8QwaByep8HI6es1QHQuAVYjQpiUSoHlVhGrPBhlf+MIWnJm9JHtekL2izNgn1/UPws8ML9z6kq
JM2zTzrmHv0503b7tzh9NwbWD3vcm6BtVp1fsUZFPfYSJ3FilM3si4N/nbfi6KhdcGE7ykfPkjGe
iKUCdBf431VC4qQM+y7UXhRjF2FQ6EosCtC3Ea8zzZPDtNQsKSrLMU42gftaZhlhM4/FSDKXVmFz
hoz6lZZ4UfJygiCCkQEyyc5eWEuvvHpeVho5TXVM9GsuUaxy7QD13avt46rlgz7a60i9uvrpinRM
RZFQXZxOLny5iHpErjQI96WpjLMSKzA5qoJrIFN9M73VY1INZZFhMLHIllQWJ62tBARD/1uObzZH
O4HN5pEx2/5TGGz4x2ZRH49spFUVYMinic0gNz5B12EWQvmjA4grRvf3wEPWqanUOaev9vk6YZgs
ZYBz/sAukAbGC9CPP3Mp3Zi+ZnmLLyaLMywEfyaXiJQbFZ6QiMgAhgQKWWdChZqiREj909PLcMMp
GJqqR/F9NkrOpmJAvfoQ9u7bS8vs+OnWSDBgZaMa4/MpwzhHzbKhxEgzL2hbCW4gbBeXa3iCvIsv
5uSLdtwiu2poBAy6YfEZlCV2MTcQOqJbHw72APTCW6P/a9GOnOgd7fK8czVABSbJUoeWBWmGv1ty
Ka/anNyWSC1LxJ9ZeO/IxUEVGnjWS/d9ADz1CGW3/LKQKoPy0MhYrOSIZY54/Uqm3OVpYHqApb3t
ra4Bw/mwZTUtWlG8bIDdxPpwPphEBvKl+rG3i1dhX2VIFSPIhWEAB0hnb1o0f6/evheJyW6WygD/
7QkybIt/T1K1YA8mr899PKlwHGrXgk4OuPGl6e/OxYPcfGmhRWaMGmzhgEm8NLQXEkdbFVetZhjM
6mRS95Q9AFJp8qmCk1qJrXtBjUEJ1xT3ysf26NRqDljFiQB+8Yljdq/5zh5j2h6sE1zcy3OZYh39
5XxtVOqnukiFIO4JNoPwjk+5JfgnGJax1u7edlwJ9GRfefXv90+i1isbwFvhr4W4K2bfQaHFdSlP
rzJ/vTqtiK1D3j6CiA7FJ0jW79NoW92ZD29PwvNQ7KRkKqL31qCH+pxAIlTCp3A70UJ9nC+MHxSx
y+5V6Y6MLvJlyM8fT/Iuqt4AIsK/cG6Or8/kw4861SU96jUb3l+6ocseT8gIHCQ8A+BCCNU4ycBe
KY+eXfe3k3xj4oeIT5018IcGGy5nstCrLKJK7Eh1D4y2H6oHjAjrAb6DR7sE8vXAhUNVhkmtM/Dl
Lgf7df4Wr+gFxerilq4TE3HAPC7cXPEyLETX+lnzn1Ued1R+ZhYF+bbZMw5etJgPILEwiDhqkFPB
xjCpnux+5GIehly/JC0KdFfemSxHDqMZmGqz3/dz1D8KUjgHWskmhrNKqHRMCVo69H3W5eRWL8fy
vfkrA3KqEgEo01eQwBk0D02Eo96vWsOr5b/VIr9g8KtgfU+TMljqdBMYyZswCEd83mywQqSn2Pxh
+ul5Xp4dgb6jTC8v8TBVySaHzxF7f4k2npmlh5TGCgWoiBT02YQf3Y9f5Jx2jnhp8pTI0P0beQBA
yuO5eJxhEtBJb9hRfIrM2E1gb+x31XJby0jiaOP52Bx2wjDh5HEmplpbK8xHZ+M0yfJd8dB8AogV
RboVKYXXhifiIW1xSzA6d7dw9oXdaVLJEDsV9UeFtRH6KnkHmI799wrvGqMitSwu1hdGkNIjT/+g
/Yp29SnatSGJ2mHNIfZOIDJo4FxjWr5g4Agey06ZwqxoIZjjKGJUI0Zi5QQRqWrRfRuMxtAbywl8
CxrTDIooBAtQYPKwHwOZ90HS+J3BKbNS8LEzYTBlBbUuXXStWrTES5MdXU4uB8yxHnTQMk5wNUJN
TerD9gFX35wGDdpmarmjWhdj4YZLxzKjtAEqpYadsa2MZSrtfxcwPmJnPtTmn9r/QJ68nEEi0CID
V99KdR64JHnZ35FcJVNB/9zfWqjmggUynfreCo8m9Wm1K4KarlG/QEZTnr/UE1ofF4gQGTKDO/Nv
gk8Xg2Vy7EEMBolju73uR16o3lkFaeQpD0Uv226UgJtm3JTIwnL7h25FahsBtwk1dWvJY0feF778
66WhdyS+Nypw+vgTx9Ybtm0DdTCl9MvibJ4NRMVcqEF2EF4krZjNmQPW8T9GLEF426wNZPWyMu2z
HGUGcSr28HBUHgavFQHT/QJP9SbQWiLfjDyzbH+fbMoEqQYOccXXjtsNm8rLWidcIJtk3uvBUmXK
WXBEjjhKENOeueRgOrQFowsBR+P25cmAeu6VDOA7MZltsE4ZtsgN2UvoQzyKZKIiOommGV2F8bCY
sj2qFUA8OhlPyoo2uysrR3bF6VH9YzDPf1aRQdPYEOkaamrhqrl5erhurkWujFwAA+VNM/d2/Qeg
zhLu+//PClWNopKZPqNmeriBy/2UhRAr/FAllr28801VXprxiue0xhCQBVfpOI1GUNs2GjhVHB+S
eqEfalu5PFIbiaewD4mIuAH3t1psLeooKgYhrWEAsKjQIlo7yu0Lzruxh66NrdFyyN2UDnYa4A+9
4tVweqfojToa88l11n5aHuDX2jQndazRxydgaj9gEzrGh9whrAzxOXX6x3Oe7BQtoiZ7UlI0wKb/
nG9ImGhCQk5xSGVZUcM6c6h/0l2RPBhmysoX5JUYjgqhssQKThtVrJH3iOaPrdVl4tv8nJDzlyVy
d+yPuKn6kPTIKWJ7dK+aoozHb5QCbPN70QnXAYgjnNVjniBSoW0FA1tGLkpegTCXICk03J+uhqK9
nybtIzfZTaVPhK6AGLs3NGhBxxOReJxB4RienO7U70KWCWSHGpOQFulS5uNzyiFugIzXX1DH+KE9
UevrKckQTbIr1W+eDMT+VYwbpHd3HPB//S4RH4P9Fi1N6oJu36l+FeNng8BlRXsBWaJyjhSs7wwu
JmXh/uwl70vV0fo5HTiHSMshboURZ2hABR4eN0Wv8wWBgNDvqFhNkKaR5TRxAkz5MY9jS9umKxhD
l4p9TjWVMCUofnwlhKloufCv7ItGNsynMvovelruxc1sUdTUdn71VtHWO6fxnJlBK2fiEPMxFdMS
batKLiQxyeAZrVejn3G+tXfdMlVTYzA8TJKUnKRbftYBhEgDAjiumy824QnYq9G4j/FFmqNHzB4t
J82Eufx8nljfQQzuzd6vwZAf74pkgQ3oFOmjBu74J5MuuQiiaTsBChpOPZjyQSuKJhWR9kMOsxIA
uXRFQl0yRgxAM4ETFTnJXYd4weQCypVXnvgqM7w4GB6f8L5DB6gbNAF2mqizVi4tk5CvVQCAiNOc
XivGSydEWEZR0/bG8O1lDZrIGTn5kor71obXa1FAylsipgiTjDWkyD+EeFNVFEkbXAp9OKvMNMU/
9j6+wVA6FWB+Cqu40ObIe+MLMbhObER/Uv5ddJ/LlHD4lh2GZbuIyG2kNVWlMSq4ncNEfoOPsbqh
KwZmRwVr5SyKXzvTu+vx9h7RrAHpWDfofKlX7bUXAMUJ3N2UIiNpUcLuNjvuMx8ACHi45tLZgy8k
yvSRqWeROjTBCfSQhdvhmzrCD7AHM7psUcutqht0n0O5IY9d4QnutYC7NSznZfygBY9L1ul3ejJu
FxVlHk6YiaQ5mmkyEhtbMtg7zdET6u6Q93bgPoKfkwGPaWStMWH/fcsF141nYNzZ9/MHmoQsOhwq
nX0AhA9rP+zVxqvvFYehXLF8JI2BHCp0UkiP69AftR2JVFbwDhpI8Tg2Y5yRM3b4s4xpQLvvXW/L
/ef+PNzC4RTUbGMaG5mogmnEqrfqbhHtgJKS5zH04FVclNjuZWwS/0tAM0CbxKJ+v4TSW6+7mHK2
fl5l0jUgNIEPE1iqusjNT0URkT5r+ghmfaNmKz9F0t60ZSN90jcXfrtOVJUHVBsP/2ikeSQ0AJoN
ncp1sHeP9PM1y7coNPhTGL2j1+r22DDDlDXj+nG5xDl4RvDopLEGaUYkq0gfmfg/puHkGQVcgCEr
hrCHTmegcQ1pfIV3OYwnkaeMcyCulMJGqm9yC0K8OS7Oy96e2lNjnN+UpZBd2auPVHy2H9sty9d2
nJdEx8iZ5HX7xwDXNLyf5pIBXh/6VSvbEZW8CNA6XNx8sV99vgrBZScfTO3t2nAYAsO6LflqPec0
uML9aA8QtzM4Z7wfgFeX1QWq7GZ+Frc3mEUlFpzBel34KMq0zSZQ61HeBzdsVASU0gn9Zky50BLH
6JN7rjCyFTbFWqautWTmvWkr88H1wA3QNcDLHmfcpZuVYJBp/7dBRo64yNR242qCOxRVUJtdFzzB
puuraCK6FRCYaJK/oCl6ewwJaNBYeUcK+5KfUUFls4oSFYSgsmoL8JSuiLkXbJ7Qm7/wHS2P0t1g
GcXI808YbNCCuyR92q+4tseaqZMLbe3GxwCPppMbh5NKZhgGPmAKsoCsRFByN3KvYUtwjtObOynz
KsxUFqaqhJ2HBpredhM5B373q/rhF/e3zfP+XX1Ksx3ROEvaaH2KNx6XAQGOZKa+yBrvFtxO6U39
EKNmOOFXTVjWitZqqdA9/ydaJX+QHc4Ro1t6R1EOCFT9D1qwPDxG6cpb2XAF3WCNZoiIOMJhtbKM
h0KaMD27WMFgGZBKF0paIkrmcxzc3EjV+eicU+qoSdjUUMMFcSuDTCPFNbM0o8StOH/3gs5xjDVN
H5OUOikwIPI2LovexhWiVfv30FxRNO+6RjirxAjPv8gyknammID7dbhgcINQbkvlUA2tNPV+QzKT
jZpIYnWxniL6fsl/K0ILw6HAYZHMdOKRbX2gg+d78U35Ld1dqcLJHiW+W+17q7v7mFUGVRbDHnoO
WEg+vhv2GS2FkGMgkaT4o8Wtv9ba4CiPO2WAfo2nr9NrYHXN/wTW34kmzjuZj6CeS0+FvAPhs8K5
AMjWjE4hVOaRqTlkgJcsVspe4IdVfXS3ooyYvPOLT3mMczYltT+v/jkqCrXBzYqqd3xF3iivm1CV
sVBrI1XCYoBo/JgRUVIbdcbWfFKeQiGZnhABHPzFCYM1Q7WAyVumidL/x15aAsBrueu0/KhisTOM
EYHmo+y8WuxqUo6fgaRvaVFHmLVQMJehED9n/7LghUasXohhboGEF2YU2kmcetN29+IKWjBJSQ7+
SzYxf+mU4qcoXyRqASiZwugM1A2aMXWG9L8iZPnazu3iM1qRdJgYOyY7MI6Dk7Jdp1Gf41VcuKOZ
+bYrvaKraibvk4DkqJwK0Ox7EkNFGno+8ED8AiAE/EJ5ib5cYSbI3/8wkXigPBpWEJLRqINUCssP
kXlF7bxHfYYJNkMA4nmFibyQ2Coc9wfJf3W3ocleYljPpz1oWXIjRaBCm6jPFqx3fd5aS8wynb3u
XUl6D/C+bBlfV2bdtuZ/AuTE5xqqTeo5xF09Zl44D+QeaYVlfjFDIGxoBh+uZ7YwJm5xiAXd3xPq
XPx9wOeOdyU7YHyJ1aNlHy30jYMyEnePeJqOQ2ACQOZ88+i+6Yofoe9MuMoC5ASOGyA/MYUSBlNI
Wj6ar7KzanT2HsO6hVtZ5tFUMzEgs4Miiyybnj/qPk3J/61oPyozP+pRHuqlrnyCfOPLgGPP5+bq
oddZo6mb3XiJiUl7ApLCuIvOdssZvoqvLgsxt81O3GD4jMG0XYVWzZmDSnWEGGVN8aPbGu/qEi5s
zsAw9cnCVApDa25fJXtvuO3lRB0xA1UDngl/C0+odPIfFrih0vfJlvAGyG8hrBRhYSXaEYy8ZWq0
BU0IVVv1pL+GFMqbxePxnHk4wOMH+PqkojR/tvBE5fBx+QiFT2DfGU+WdIZK1NvE00C1IEJ72j00
FSKS+R0eNkAmiae1DChlxtaSIAgpaG/HFC0YHCcvL1IM/CkL8onrPmW1dKBKeHmY+ft8Qo98TGHq
PpkHkfXHcbYc0CUMiuHIuR1hQ7qNs9Vm84FzqkTPP97Lc2wU7lfpbk4oj2rPRECNSiccAZFJNgKd
QXtkjSRwMuQcIDQdqUN1ZP4we832X25XcMdKsKo7OirqtT62PWrjQxhIdSGY9pe5OW70opFi92FU
KnIeOtlIdNQ2+0Oz4rOGTIZvgu3EFYtXDCNWFZL7QzlPnKX2KcetMKc3KohTgwIrp7wPqypzmRdx
4WMV6ABLtvDks05rX9/bfNA21FDHJ0K+4+uWmL8CvvE0r9kFF4AnD72rEg947tUkb3ZVHSYYyv4D
/Ng88Wxp2QI+Q1E0Nxvp9zBMwr6OOaW1Lm3JlmH8uQ/SvYrcLFlqP1q5kR00URXdnjeRoCWEF1S5
OOte9dDocRGBvsIIcSSwMrov72wvWqG5MSLpodLHI3EStrlfB86JT/XxVIK2VjSbosVQkFk0QKQH
3Kzi6otLLVxyeI2oN15OXIGe3ev+i+q2R8biohGWr7Oe102PfjY7vEM4AmNfHZ/m55+zDaD5QNcg
m5hGAfbAcQhWDbgR8ZF7AT3iN1uH9n7mfmTxS05Qoj01zURnBMsbDa7KO0nB3MBByU9lwMl0h4zh
8duZNEMYjvtrg8h3kn5as6TdJuzP3xGb3YU/+cwRcijtStWEtfqfJDkpBSCncVu0lCrX3aihgJrV
wa2ivIFcp/0nZKRJ60ElMdjKEPXMKItFcV9/KBK9PDpzT6/0KayYpCOj0c1ijkdMFMVph+FNFZy1
fot9LICW60z4TdS5aJugKe5j5eH3lsLRggVQTsCZNSjlUjHIFWpSyCfhxLyb37gYkkIPYLZkNzgm
PyhnGqe3Cbhbln4gPPztPeNLIrgenIYmgv0byiFULvzBg2/VIUWF6i8YR/TpPka2Z8u/w+mkCrhD
FMgdNLqIc0Gj67yya0LTPnBFiVK0PLVuP/QKZVxiVMDaFWz9bss4ld5x+cO0eWt4+c2rhcd5QToF
EaZuS4kFcbC4gziFuEoYDKC1kRjbv6CPPG+bjFk7R28fhUA23TFZ4Eqhq7OF1AI49sc+NIoji7ub
uWUUu2+PhRtYoDI0FLvKC8hdJN7fe7AF9hAwJh0Y5ncjFiRYrOsTZuzp5pnLwwPaZQk31+un8mGQ
omSoVCnBFhxAI3NTcrdrhAGpdPby8Gi40mMYDYuV2eiX+yd1EoVHI0AjdjDsfX6j+HfF5AP4A46G
b4/FuvJp+SrUBRxb0sm7PSC0gCK0jpU8NbWUBVMKf/ieht9WTomGKJ2xv0/xW42+i3DKyyJWliAW
sMqS4ATiPK5NaJp7vWU/aPqmLnS6ZDOhE5gGz8WSvqgc1ivMJzlGBurWXM6MOd1lLkbJKoLsk5UM
Pi+XQXqEfQFoJTims3wsNAcxcanejTTUAPJUtj5FMHy5s29xUVy0GpC/AmTa0SZ+K4ZWvyDvFQDB
Av24Id+gLEE6owdY0IKxAvuXvOrQDidxqgsYO08IbeDD4CdjDZ+fR40hjTdmaEXfnJlJEUobGDir
TdkqfwWOeGqrqhkXsyI49zYQL+LG7LRgIgDPB29TQvdbJzZooTMFp/0QgLz0WX/NpS7cqbkp7laE
q4cAD61Mrj859EOivPr01Gz7fJABIFicxDn/WjK1k3zjQtMyJ1i8kk4nmpji6GJf0C/KuTEPvipP
/sx/cEOzILUxzoBqILf8lTVriQNdA3ascLo2+4hdU73qZj9LlTFZRzA+rTCNazUSxkLxyge2M5Mj
AVyZBK2PpFbqotZ15h0E9IR5VvNqRc00og8IE0x2rmwnYUrOkv+NMX9zlocQiV1E6q0Ndca6HZ3P
XVM2LrIouVNikxZ0XSLQmZp7pEMGLkGxyp3Pih4vWI5wVa4JGZznLBn0zpwvPEhR4rw+3BAy9OlL
bdvWCfEIR0CXvm4XDclGyILl0fuLxYhkSYO+FLVoLMFbAuov0Iyxi09baF53X+PS9H4ufhHsEb+L
ICKW1wMWQ7sfFD2uZFMWzu9dkMgggnpmdKEOyQO1PtkbqH/kDP3hevGsk8pFX/7tVxPH9CPWev7v
Y5T3mAt5S0QO5eWhy61VsqKBP9+VPTjrfu87sInydmwcm/1DmqcONIajb3/gr4ZC9bOzI0blm5yZ
pKuJz9TvfvYs9kHl2LSQp9xmzAzyp9e+2O3GPocaLjigd6ZktjI8/Aep1JEh+eGz8kfXC9iw2MqA
mQhSVIlbWCg2szZyvbp689/HY1Y1++c9p//Xuo1FEfT9938WRKYe62acSXzFN4JCaQX5m0si1gci
RLA/j+0LjVFQSpVlxJ7S0rTRG8uzBvFlTcZ8+JxZz8To/4BiE5JHZqNSifWq1OaUdvVa5rvkmMr+
NVNMlZTsR8VxrJY9F/rj0mbpXI9m+WVreE1FoeG025CVWmmZTaVR9uRp0+3FIbgn00OSynvmIiMJ
kVdVtQrQ9O/XIOZ3FzGso2/Y+IHiHGBkuKw05CMn1SgGOvAuKryDT0AOF/ySmU1i4/0yQeFDDzmP
fuu/qH7ld5zlcWGJANxyj33S/MMIrCfEYY1l9co7dwdxr5AwcK4bSSMQ4w/+LVcy88fK49uElQOA
dy94x7x67z3wCiauH2aXNjrpIBetRFc2v71AN5Oe8uT//RYE397a+4yJr0Q0WB/kz9CpkUUH6IPv
XgElA90sLRfP9gr+NjIquWA4ISy2ifemMoKQMxca1cz7gUK2btXOYkaUJk3eUUaxkvB2Fop8g871
i9PPU8NurzJ1Z8Yzy64JLGT8QXW5LWHpWH+kKuod9vLozJAS4ybsMVefZ4iDwEcrOSTMH9Ipl1/l
KnEbjvYoFWyaBQDkbIRvbP1WCkLbwKupDO6ajWRuKDCAGiEmb9pseQUUH0uq18ohO4KQycZ7ke53
ySDT2ygvP8h7RzjEKu/zmVDXvkb9PT4UvEVWkh4gmSiamHa+OEBoiHSDrHPlptmShfYmjbEkyzj2
iqVTUE4eBFZrtG1ZPZs/E0rgzfjMGy46yccXPjkMsQ5BKxU0eg4K9ZZyX/URX+fA5IDr3t9pyNxr
uu0ZdbFrIlvMKbs/0NzWFCuuT5bmPXrjbpnykfDZLf/IxVVPbh0JSY+M52OiDlvj9jIxOLVviRSV
QRRStzOVKo+WCKsFa8UhYQRe5/Pfjn8iQbCsx5pjhpnDTLlsdXhkExdr1XO9/YAlG7nXWfEid0Px
pA9RVZXudJT9qnCumLLWAvXwsMyGZ3JTR5XZxB+lQQlnMRakk9yxzt+6i6Avc0DpIOXnDFNE5Blx
RENrIZc90lc85G7eVS5j0zgNK5vRcAGILpjZs6sL5z1QUKmfCxm0hbBdGw2oRsisSdBq1EkgpV2q
SvN3YFuk3lJyKWHPvN72sIBrTR/B4deXNP2f6CYb4Qo8TF82CSXYxLDJkHwqh1BhpXnrMIz2AyeH
sok7sufRUEEIrK+z48JP9KHXIymmq27pGeRpfdhB7ESlfOhGL209LD/vbEnkAdoLjDUQIGwomrti
oRw8FnHlD3qrEJX4cWC8OSoWZvN2m+zgsJ9MDwk3GXPxICZH4lAnAsMvLjD6M8U7gPX0PhhrIsqn
YqFB/8EJ8l4mv5daAg/uZxOsise5sOPmAxoOPL95g6Yq266IHpZJvGRe6NTf5yqMWUCJqIMzoFMq
VKGt5MsKaNkV9OF1+P1T6k+xyQNyd5LvMVU/xswr/r+Z/Xok/vBWV23/Sss4E6LXWKE++nOhMYTy
nxtPCv0QyW7amCfZlMChgA4BJ9bhnZr9gHbEwZcVww+uQKVUIsF1M2jDDfXy2cFZjUtBHSG406/F
b4E8S1ZZER5Z6QXOz0HUA4jEOWCi2loyMPNG76/SY6fwzAULWUfNb9bFaiL11fJb2b6c066w12Ly
57va/nnWkYiD1nsHdzM0xscmP/xWp0i0Zk96aOwZgEKYrRawDTA/qlXPvZ8u9YEAnUWa8TwRqF5B
YtdYq5040vkRfiCLo3jdEQgf9U7HnZh22rOJ4fLzuqRntDPXG09P994FIvg5CXZPVZINCX8s1sNa
KlnpBSMgpUTixecmzzTzczE4xF1x31fcP8W940b1d5T450Nt2ViFdni55/GxhGpY2A+cl8pH4J3i
h9iEMmleQ6lptp4RtX/hvvDLCcaLBVYvR118m5h6T06ZQDK0KbxFiF8LXpPJx5Kzc8jcsAlM3u7F
Nd/ny7++75kuR53SOo5GzpWSveDgXY0c3uG5MzpCxRo46zU7Sr3bmD7k9W0KJluCSaHOhSQBWaQR
aVjgyhMlRUFPyjguE3TG4Qdvuopzi3kPE2cAN67m4S6TPTPffmXMx1px3zOKGzfDPGtNtE3Gald5
+FTiC5molajSQgbElAy89nH8zC2hN5N2/6AmCDdDStjscbwb11bUDoMmXAoeabtTjhPCEcqmoU6+
+dSF6Uz5xNgrU6azy4bC9GIQY5289yF5Ey4QQ4p/Sv61K5KfzE1AVR1iOMWLO7E/A8EGLX9uxJgo
tCt8vNjUlcTf0VH2EBD27G7nA3CD8al4Ct5o6RntiX/9pkQObq1/WEKhZQf5x7uK4ncGzyspvuC9
hnMahQnMM4bf0sDSU6Vef8PS3phr2LxSjxGGzN41E/LcQxuKpzGNgv7PN4MZ5rH4MdBUJsvuR0T6
WDaW1/SUPAdMQbVwr7wQBTi5cQkEACYlOnTNw8n0vCfPPw9H8I0g9UKPBt/Yrkvh4S682Zs6+MWM
4r/QMS3OeWq6Amdsdly37Qt1iLd87g8C7zZaOHzlygpLJ4r8QHe3Mk2SLJZGJxEKnbjmV8SRNrxu
UDfcSGepOpT+5tk8qbWhaJyqqurIslUVkQPpt/URl3qnBub7TjXoWbUCqHH+RFSTWdyloo9jSzpf
oCASjueolBbc1/sQ1MzS90Ss32mtpbR8XoBHJ9p1ohh9gt0bDxzb0TsKp4JAOOHHj+45kOO6JDVL
4l7FMYdUvVYOgvvBSj0/H/bGlQoxnrhc2i2YnGJuGdAZPDWTWtoxUv0hikvkLa6vnVufMANenO4A
hHHD/4Hz6qnv2Tuseduuj8FNN5FDnuCsam5cp7MkgkDLs3MXpnACed8eOTKAlTR6q0S6yYr/32rz
8MfJC4X6YU8mn9f3j1fR9K6Qqxg9VCRjmd0qhSxEaboDo/4THIk59ZBP6fOOlINmYQ4FsmOvecg4
M4Lw9kwjeX2FxTJvilJijE10SXaUTFZr5P+RXtnU23q19vCn5RNwkZ0vj4Mo1udnXxbRrcHsx7bM
r+Uvj+3tY6ob4aFs1wlYaKjso/vQ0yftrfGBAbKxjLZvfsZdERwmhhuLu0hQk/Kd3/qYR5hICxhW
7IeoiFK0ObMDuRQ5+FPCRj93YY5Ww+u4AejPAX69mqzzlrnEfOS/xuyQpgUxM+juW/psPV+GOdlm
bL9TRr0JtCxZLJh8EODJEnjsPycn5FTXfkQApINKrt91ttLeuJsJlc4O8OOwKX9urlhyIZt7BBUt
f1SRElbO7NbXiZ7vul/WdAm93b6Ff+zrmfFlHHs7PaLDmHjMvLa79mDisczFQu6vJaJkBUr4o386
miH8/FWSoPDtPWZoZpELegt5kEAf7aTHF8HIv0t1bn8C8g4zVpkI2EDrWwilc/muOy1KWYZlrkLX
eZno3EbA7wlQjR/f/jwoMt3p8uXZHkKYBkJbqLlVw27D6ktHg7UJ/SohJ9p5nXW8s5GP6aIzNQQ8
Q3RqgjltujYVGjnwmL8eTt3aybFvmTMs80aaisxtUxl55bLzpKCxSYHEphUzHQYYNhh9JIDVIH7K
GIJpxcJaCGUQdiKeVW6rl86IAcwHvg2sSRca1KtnpGg5I4GJsH3ttBf2kPnUhozRyCUQWgLmdN7E
ATTa8l0GzmMBmg6wreH1CB57doamN6vzx0BXLAy+5jJAzv4+dbOAHqwfHEMOoQJgCKABXgK2j/ET
wDZtoisXnzptgY8wEokE6U2GZmbt+JuVtD2oIKvf+2MFKIUoUzqpCN6eBWKkD7cAgI07cxYBNUrx
6/fLydRO6bU2YF3NtWLo+CspUsm5TJ+g1ruQuAkcIL8CjLlPX/bSo719t+TOx6Lzo8OMtNvbui1M
cnUly5yOi2kJGX9AhSw9weUUm87YW4RMd+gakqtXHGEYSrAzP0ZUWzLU4Jq+SuNf4/h89ZA3W2dD
1cpi4auq8VpK2CLkYy6vTuPgUPKB+57DNSEAl4PqYeyzTj5KtBC32e7rg1wWH8d9EXE4bZoEY8hk
WH8fVerFTF3VeOf16VtYSsAegaFFocihzk4yqYRHtc6CJravubzVI73+ZEtlxlx5A0X/6bnLjgmw
c6bhIU38j2i6Gq3t8gpMUHynCh9W/mck+GnHS/H6720TlZ1caWnqWtAAauaffQtPvJFHZzUriw7s
wdK2VcwhGM9pzKZqYV0fMxN538il37nQ1533mM9eQ957ymeGn5b4FNjPqz4nYte2HKGdVOYQLrzi
zV453QKLZTuMfyO5n3Hg53SauxHnwH2Lvh9B4YnGSwHh2nlHvnwPklGubfF2sz2hezAHjmoiHy5P
0eTk3qhL+kaP4F07+FbbM/5ws8WDYiUNoNoC37twsV+Z18hDqxUq1yE0LCegrF3bid+KGIgGgOhG
/sabQv/mdUOt/8dWI1Yy5OgZ0gtl5yBZ78tcvchvwMy4OUVSAjW/IkNg7147mgRJTo8DZ89sgK81
sDPYMCs0dfVAv411pYzV/YuFT/8Gyr9KCFQKYJWTZ30kfMiDKReTp1nPmNozMVkn7q1zGMQSooEo
2JelugAAKJsh8Dp6pPiFLVc+KqJ7EPOIZAP/aE3PJEEu+It6WH4PTU777dMV+3jNEH3Z7oRG2B8I
yC4Bny0kV2/5Lm8JP2B1N+/hgrmqBtJ4fk2U0rfMh2h6CdUIiuNJlc3gf67GK+9lQ8u7xeIzz+vY
YRhtsQKXeO9jVS5tzCqMHbcNFtL+eO7lOzNgAMHgdPaWNaCK2o9DzhYGVU9OdbVOrIiKro+xYbOq
bJPvBpBhqfmSz59JbDcIizaaNpMC+/GjriYK5xiPi1YvPqC4vKqySiaytn6fvWPzePIOly2xaGiz
5CrP45VreS8BrIC5GnWGu+E1p3xYwvjFo2/kDzssezBPXKnJhHHUa1tJs2m0GE0cCYsHDJUNQV/0
e//hzDOG+OkIWIwgNKJSHP+qAi41qWelSKZEVZyN7/rDgRTw1TzNPZ480q9k9VH4CZ1oiqAkODAD
4GsOUkgR/Q7TcOmXmB9slEm5/oaqMirQUlWGZUpzFclkw+MuzU30XUjh7xfTICldykB+JTAIlFGi
+BSGuYu0IiHmLc6AfEzb4W9UUjrd3RfZBjkK6WBhUvYCiMpIX20SeOg9DVj1EvqAq25tpmxWAQsl
KbLAUqaucDrG6su3HTDFcFhdfXhh6fIGsL81wrhzNOjlWIJ3k6ZCrqDi379a/wukAtsaMEqHYFxL
mLdBWUIr7Adk/EKDuNsa/lDcKCjKgVm/6m6BRHNvHpcZxg5sxnA3ccsC419827rQcrJkG/E8NNfN
mJXHfQhDXmhhl0ajYeC3ccash98pCJ3PLo9LQOkJ2KaHtBzUfNRFZzO3iBDw0uSB/s+iN6Bybmxh
GNxTA1FtZXLANdIHLA8nho6VSqFgJJYh9dpC0mBCQPrJ2QxJToiADejEe0bc9FVtwnsCdF9a+z5/
pTq64wSx6diAZIF0RkNcC5BzOZhwMTnkYPXDvFF0M3Mh7X10bdLVdIOo9xIUMlZ6n8sAQgJ+2wRI
9VXAUn3b0R4TyFtyF3v4NRwbeKcKt8EYRvRYTkPB0q6qhcoUWjpDv2fCM29jjyDGkZpvgwSs6PZC
bHOywpSXPK0BPOq9GAIImtTwsU/8120z2FRGi78C66vLbHk19wPFeQmCUiWu2iR8o+aw1+Ao/HFL
Hd+V+oU9De12kjoyLvM0hByLe1tdrn4GkAV3N0Z5merp5VS4+rBJva2Z83RoJ2QUeJJbxaHUPn+0
jVJM2CWGPjw5brkxCpkJ+DzvXcxit/G+VJTtBmphwEo1uSxp0AOxfgwrHqH0oEbP28zU9v6huG2D
5FqVNRkQ8IIa1Nnl/jg0lK0LH2ZPLFm9GrzYhfE76ryAI/xSaqiAIAsBdxowUJUtBCRNIwQ9UIIg
L+kgP5VOm2+LVLtUthENV2e3eZUoqeUJxUm5Lqaw0PVbTakrJ/thctS9hgAQ5XD/FDMiOBQst4aJ
AXXKDBD/dFUIIkrwlUM8lJ6MlSI2k335pRRVJoaPUAxb/RQkV7docB2TnHp5/unHh0F6liZylKEf
+xfC94bXxePL3TKDQOI8PJpKjBqF8dlkm0aCBHyud1LtisBsX1qjsQBQ6x4jzaaMuWWduh91Tzbg
KqjCZp9t61bA9R+/vgtrmQtv8tnhMZ3KDM50IkNCyjQvmVRvGX0X4cUfum3pBTxRGlHSPkuhI0gu
cfIponD0H1Qml8ZTR7JRQp5J13v8h00fFpnqVgMVPm6PlxQXli2Ry3Vm+jjfzjTMQ1VSna98hVHL
HUDbqAQa6UMqIlZyr+PV+f9fTv7M8+cAj9AxlBBJrtbSoRTklNzc0zu2AtYymPPygiKRPsugjn8T
lXTxj0B8De1p3AUnFSJclqF/BGX2mtox9xFo2EoYjk33/4Gc7vlppdI2UYxX7XhxUbjM5kuMmuQE
CywRfrs39n2PBWavZkKqCA22BahPVlQvP5u7RFUn3yP+9BvSrTO7EtjAUQrVATHeideNaCpVhqU4
GQ7ezxlde59mOLBCm466BK/g5UFpQA5hvZR5KwIp1aR08WmPcNMSylm/1rQkyZHqZzPsZ9qEc7bz
sa996x0kc0wu3ZUwa9fp5/6wccUaSTuIgOo8muXqralrZmjTleRTU0ukDkxA6JbQt7dY6tsgIAkB
4FrroskFr7qql3G1lZrXstlqZc0dR5K9+VVx9bPZsU/z54htpJ4dBlE/e6FJ5yGgPsjUwj+1U7k7
COKuUNy4l6mBfa0tjOjSX+J9dYBmc5xNcwzNHG2l/0kqpX4mA3HMmN+diB98Uf6D6opLeRQHbat0
7CD1SWnOEBkEsQqtB+89GoVcBztecmiw7S2y/OVgCCzljbTgHoWHZpqcFE2Y7l4TEqRNybXfgHKc
frC0cUuTVHu/TNZ0psQtiRnp0XltYU7V49P7TseYKuhYffTONnThh/AKO0vn4JCmtIDGYQljNGOD
CplzJLCNIJwyYM5rWF8qV8KZt7kNIc0rlKGp4TsdsPF/X3rayw8gwfuazuBJhNF1HPZjkdsL3OkX
Dp7S4WgzmksBjdfNypeXIgGg3dKUpkOupOygfMDEnh7iPJZghz7D9v6EXKvgwqG3y3E6NADXPrfg
X7aeLOnrUMLgGofLIdw3aYDS3LUzeze3Rk+LuUdESGTav48ufkzVCiH9BNUrrwb6+eLy5V3/baH4
90tP3i+AJ3ADhVPcx2W4UAn624BF/DJS04gt0+lUw9XTO/k5UihTOblJ1ontKpqr2Grg2RM547AK
dl6KBZ9hQQMhkgtRrJU7G13oYVDOndWlcdPqM+ppQUGsGqeXeZKL3A8u9HaGWrXA0vbK9LbiCikE
9xoMkz1CxQHhXfDRbDjCzBu8Cv6xnE5h8C0U/73OGh7vz1smpfpwPJvTpPmzan6qpZEgMj1chJfy
4ygjoOt4Hw/CROZuBkzpxfwv5W4Vgn11WEVnPiFPO0GIb2Uf0WqOI3a408xVvZkX6MCgRl0xYnVm
4Vj0cV2X7lpyhQfmgFcrhTZYLXXY/CkAtcnPlo/H/O7prq1yetAK6d/HoFLtEi3y+KQ4wMSWK9qX
JObQy+eyrQIa9qeVd83aCwaihdbUYfALfKDmu4qWIHTm/A9Uupl/FemPRsKeZQkCe3MTcCX6q/Kz
P0A4wUh9FVICzpfENpZ4OFC3F/y6143p3ERp+9AespMFmljZgxlQaXS9biGejmVFv5VBkJJsaH9W
ThgZkV2y5UMp2zcWo066W2WRmK997VlVJ3CCt13YxG1fwyP2T2xXIfJF+6zOCQumDUBjV3eWfCc7
sYAHcoL35ytESlADJeMs+ShA8jIM6aAbzrtjUmoGtzLXnynXbm5EbqmY1Xl4dgajiqOOugPusKyq
WgovNbp99u5X2bAvg/t0ouRAJK7rJZmOH2MXk/7JbenDwhHTgD6FjC4Ocnh4GoJetqNRjG23NeAJ
xnOY/iv/kFWdDI7HFTeAUq+6Mc9soLVzw1wa/2j3XRd0jzQvq+zkB5S4Fw/vDHqN1Myj1wl+5wDY
FsfAf6n3mKtlld1d8lc1cVHEzyR/jITk21odvbR2r+x2qR1UaAtqlVsrWvmsxPL0EuL3/yGVNx7g
y+Ey5Ht1xdSmD25pXLvrCygALqsoTFWDg9ay3LYMQgv6LpXPK1QD6lujCxvoev8oVPvN3Dt+TZnl
mlbs80jmSxZP/DnWY5lh5hUGDdbx0JLP+c5sqHM38cZ5u8GTRHqwuCTjmDvJSIMyADU8uzXPoVCD
782GT9iG1wLHYdbnqCwEhOxe9JNeEhhBIFKRNz/IZnnsetuzYd9X8Tcg1pROvEYKifMpQxmMThRU
Rxp2S+2twPCNcFgcfJmGYSv/Fuv0mP/1J99nPjEj21Flp42sPhRVzPRB4EWJj3U0iSfBK9pOIwQv
3GfmcJiEAMkoeY0B0t2oTMvJpAEK9oEYZrbtPchfvTMuNM/lhuLdbbCnqmjxXe2lOGg03TyrGsp9
7lJ3uEV+Azk945KjoEFRj78iLqmpuhm2wz97Zg94ChUQEQMWb080nt6VfM2QTrI3jwnnOqZPtbwl
joW60aYNHfVCFTBCFJnUg+YNe9AsvYD/D6Z43X5dU1++Ufsrvu3YhnzcnwruxW2sm4vGc9InXGkA
7+TV7j1wXFDwW6nAr07EqrEkio+SEulN6heJOyf0cnJA8ZwIfU4vlqSGKEx7PBGTje7oLmlQgqxR
9GVsbHbDN+TUmErDTI2/T1HCbOk+TjBJLs5GgpyKnbqoRvutyMxfRR2QTP+g5/Zlxfh1p3qJL9al
EyWPGXW41ArsikvcX1taCxTeJy0pafE7w5JwFVV6P5ML5xRKcuhIqixNOkYAVXZEergj1oEpAo/C
nfT7nEz7kSertlLK5bGEfMKBw63PzHPskP28Jqs3jkzQ2Uq7F3pllgYQk4g4a0IUqe+u4coBUweH
ISM+UwuXe02tqv2bthyZrY7/XDyhPIR0znGVm0GnCElbToEYBWjD0rY67jdJndiE5DgyvBrhtrin
FdOJFx3Bosq8t03uhli0uRJHMFtdjz0reZPFJ8J9W8wBmCxXyf6YYD7B8BCD253UgEv3nD/E/BvG
b/7dURB/l6OfshFrahUOsJZkqk1XwKSoFvzfFB+mHtFBtUWGNht8f11p2R2lGc4Lam97qZ/6ZF3z
rABNy0eJ1PVyazdNgINf26AD6dI20nA4jHWeCSkT7gRRCCThGyevKGhjSCyf4HykBvd0IFuHB1X7
O9KvcbURetIZy+AqsD6etO21NGi5NRpr+zknkhv9CJlMdhKbEPnCKOYvQ++pxbRSlEC/QJ3E8QuE
q4ItwPb0J56geBOkLsTKqO7YsCfEKNlUX0BYtwHl1dUmggd1lhmVzRBLNO9FZHwp5lmnTsJyueAT
1zDKimHkxfRNe4JDYnBoGaOk9Vz0nTFwWSRNpbPUPPlKoOJa0HyHXw6GpaKMZ7EnwXoYKnJaoclz
7+pIv4XieqgsCZEnSWR1yd77dWxkbAFVWPFJBwO63iTkrNhdn/NC5LInQnkK9CLGE02JHZ3ESUWL
ShI6iREeEZBJ6dpMEUMfphfYf94QiQhfuodyjRcmfRgW/n6i/I3ZpNiNT9Qb9DJ8fkC5eiouxZib
cOyZ3aTOjSL+Td6UydczJIZ//MtkxDxEGDUQjPNyKGVEBjSw5oMbJBskKsByC0Xqp/kap3zYyMLD
8drMOIEoPGA8debzh4BIGzpjo/3i0bVUCvnJ/GHW8mixT0XMPiFF9zrKR7Pffni04S/1xLEL+X7f
nemamcI//byimVCkYp1mpNx0g9a44h247baHl/YpTyTK3waTsxGKha9h4FU2rTpa/KfA2q8N5uDe
baqJ7KB3lFU+wPd7wP+EYw4o9ezZQHLLn7Ea3k4lI5FwItNQ6nm5E6oPw+7Ngper8/Ejlmo3tPJM
n3a0dN0VW2IzU4EWmU04KgRHvV/HgatlCvpZYDJWP7fnc0abEUrjpnprH3QgHyaR90jzeSEJCoL0
Kjjs0bEb4Glscf+easXqV5oezRepht2r6jaDvhP8fxqvSZI4gdSTvt34Ik/K5cLVBfcVlb3R6dBF
JGxd6g8nUKkv9O2N2apqYiCUJA7+b5LHdXTovfnaYaERQVlv3n/tDhKAAvG1f13ZgUxhdAvOp6s6
aCJwd8dNlPmTOKAZPP1nKrlsrlTzETsUbK077Hj+Q9peGj4vkmr+P/qX5uHBRlkUgfIwobUfQxDa
12qlvWHaDgXEgf8m93o9FaqHqf30zo+qO71W0UIxnv1+2xol5jkRzz60LNbsBfdGqF/4XZDq56pP
YYHAtE016IiiUUyFa4F/hWR/McVreNF4BitpZubE2And4SqEwisNya84y+Iph8/DBjsTVDJCyCir
nQGPpi5ZWavvfE6WF5Vc1jfJYJq8fa7NFuptzD6mFzwTv4tmn423XiDwEhn0expejgmTqTIWyUm2
mLRZSabBhKRCz8PAFgAU5iYG5S59Ap1656fH9OpHh1gcEIj5eS73uFepg8e1MKDmHaS1khH1K1G/
fCLJil8WCpkXHzT02beV5WLjwI5EOUZ1ToQ0fazxslZ9BmQxj/mt5114S8lXgbOWGYwytySzXj/k
9q99JM+s6s3pujTB8fKVVVzEr/QQfqZ+mvGsr1bSHSIESCJ8sqCNpE+qqZMKSWb+XNs0vFo6JC2z
pF8IZAohuehUK6JxQ22SxxRkg1sKaF49PsF4Wtht5qlxGMjbwy71PezqetK5mtYLrLZAjmu+frb6
9z8IbTq8jacnWZvlwQ/XBAToKrwBed1l/29a8qlWwA9bYxAAgUIlj6mrIUHASepGQV3T1QGVCHKT
PaDqMvG1StXc7tMtYDm5Ju/rh4fPV66DONoRjdMyWPV4f7+3OcjS14e2/rInXvGMAZh3YhJvwXMC
mTUkag9c6KAfhQGQHFSxPEjpAnZuidiTDQyby1plVQB+D/BAUtg8aPqHNNAv6DZ59fB5Tq7aN+gc
0ImxV35mIe6uBE+yJBa9+Jn4dfsK5CxJaLtA3L70v9zZxRqEhf8gQyZjMnnGhoU5pv7erY3dQoU2
APv387SvKEUByc0F9SWb4CdOfQCENH7muT3i/YDkNM00q0OQJGNX+daVg58GKgn0CnUR4ToV6eK+
4u6K61tlMQHNkPaGH1eazjgQrNk8iaJJkrVq11sowT9ji+Zp5LXzCLYMVfB/zgs+PbB42cSW868T
VRdkg4migsErjbOGWc3Fk9YmElHMbSZWV00VieARIcZSeOvoWVYSK9DSOb7afDJk6ihSoq++jXlV
IGLgDavXlkkpYHhPi1nfFMbzcDqbIVHxUoWrbBbLnR3wgS73HIFbCKFYl8tWaVMTN0MLYa+1OHyc
tJ6ZMzKPiczQ+34WHYula8+loAXsrBByKOv0JvIzfk6MLZwxPO/8L7qjQzw2+ih9YKDxoPIZ8xxV
DNlJX3GEi4hHurxs81zL9I36bR0902tMBgimjTv8MnTwQ06mfbtIYRi9h5RmIyyJ/PDtt+N6zbGH
mjobuzLN15oyyEZgtfULrZZwzsqDK4dhulhWNxgGQjtEL1b+lJIxOh7wRvroMDJiDSPpH5DLImoH
+K3k2FkdTW1GWr0um4qN+ns/qUsd+lgV5IaPU0HZyUK2LHiuclF7yf/1++c6RGSxqxTOEhnT1k99
MtHijMxJ/ejGVLW/UveXXmVoNcTNWqqFwNzgQ85qtb5HwF6TbBucGnm9NV0IhI4TjU6zdPRAlqSR
hDTM/UEM45wntCKD5lAEbXMWKCKSEzFwUsqkAMHjReqFpBn17+SwlqlTi82GLlcIdZs3J0SgjouQ
BGGqsKIxaj3DPIbW1F48DGnzWJDIh2PKxYr849WEF1msgdX1QoZt0E3V2S9ElIBW5ZqTtqOBM49Q
g50jffay8DKaS8drM8FDXdGp33CAB/FYEHiNponXyTbejCLjI1f5MbT/mvqhkxaGfoiLTySp0I+H
nOQGZbd8vVeIDuqUakXOePILKno3RhSXfgHOIZIVJ03xob5Il9EM1k6fUqFY3TZ0gogd3B2EYK2B
uZwwQru9cPGe9LoWrsSAo+t8hn1NYLHRd2qYXnCi4yTH0kD39NnHHmSRNVLlXCbFuTC4G2g6LYz5
4oHR8mpdTEpOe3S/3WDuv2FjYQQOSejpMCXfc9I0pmrAaTBrfP2UIzLb1ZnO/pXZb0QMI+d18Fon
EdrKATK/vRcleqbX3qz2rnhUtVInb/0s+eCw+fllUnbhATaKsKNKUFHfjYsWcoJvBl8GsHutwrbw
dueRrzvPxqUsOhSpe9FZ99L/KjvNajEwaN35rtBAXI4/KsIRxFR6ORCQsnEGaBJ/o3NwDO/bPBkk
fGd9N7/CTkOt26W6pkTiSoltGmNFvEbjk2w+4DdW++tVbCz3fgggG2t6uhfK1QyBtrZa91ecDot7
Ca3Ommmq8fGjIQkIDdX07o1NOpWz+pMloNwP9jk80XYMfaysqA3vs/r1edE01wB1tS9uWm6+9wfj
M3ba1f5swktUvPFXAWCxwikVKzyVNNvA0+R1IqvcD25XyfIp1TmOaJzdpMWauYaREt13ISNj/rbO
f7yor3UkoMFWEkWl6iwlZsKAIgL1Ol25OPaUUjiWlqtN+ovvBiV9Ksa5/q67wVuw7rwz0q8xrAI3
twEAnSdvf73oiW9a0Afpc6Qe0qeqU1y4E4rZJqOJdaDncQZkoIeJvCg2Z67COdNvdh4i3ptmNe4I
Vyz+/ujDIFHZ62M04HVoqQIsC90kwT03QODMQU/zGdywFe+xckbOyEOPGVQu+x2paift4LM5UMb2
ww6UdMbGlmurfgvNcE8HZ7EcOpkOKpnEAeBmuzsb482vx9XvOEV2PXyD9ml3yBS4/HpWI/xOkywT
c81pxQNYPhuzpgV1Jj4e1t6V7DKe+mEAnuMgFBasMUXbesElwXH2Zvy2InMx1GYbQOKVgkxnvNlH
yq2bhv7qS0R/thcE0vTF9IJ5MBHpwMDsiDe3MDkRv2AsBLJUaWeTazSnHGv2BxtGEn34V/S5x8/7
3yTm5ty/0RGoETPkB2Z+zVlGtFUktNJTmxoZxalq3h7G6KC11XrwfhPupt5a9/7fYI4AaQfLu7aD
9PhRbajTaZurIodEK8oxgtzwy8zRCVHxOPZyIwv2LMvXj19POldxcVh869u4ZsQH1nmFxeEe7WKI
VlELJDmGHMZ6PM1k9lK05x0Xyujrv03AvGDrU/1Tzdm4TrsZLbhRv40bY0A322Okl7dtI9T6c+ud
GLm/mQGWb8okVFOZGXaRMipyUPBf+MxHbzBByCP8z9eRrGnyhT6wtH03nW00KR/LM09hAly0e9MU
mITkrfrNht/lWht/wkrCd4A5vjzEVKbOWHOOXRYFiUEdP1j9TKT0KAhm1BQrOQRKGXrf/CPNQFrP
yTw5+Ltv3UdBa4rTQOQgncKXLxJlIxwvy0k3GOD7YSkLfpK9X0sDCmCKX7f6bsyGWqQPf0RBsfx5
ObTiJF1WI/xDmj16e+hE2YbxlQibyyLqwoheKaaBJQiLohOPqfOheT9VjLeVLp3Numdt+/4Cr65Z
7O77qxue+SOv+cP0eZAvXMTw5MkmDGPleP+r5A7mN5pJR1KE8U9xpX9Tun/qQqD9fLklo644gHL+
02qGbkVTJFAMhT9f/5fULUeZo34+UVZ8qGvr2vOF8/Zq/gcnguTf2qWLzBHh/wGN0Q4mtiTWiWW1
h8COXn2wD9jwI7DuEjQFInM6aW2GzbxWpJS9WvaLAsZIEZ7pmpQ86ylFUaWgV049GuD623jCl9W6
FNU5U8KTjDkvKFKfntdzv1o1UaBbU7n7XlmH4ap1C4UchIY51lDJdGEEobe+qVRr2BMAy1FMtSKh
D1BEcHfuRo4wZeOh4uaJlT34+Ogn09pTTuCDEQgycnuix/nqRvGDuuBjEUhCaS7senMEqDd4Zp4e
fz66pBtTqzMvE6Fpbo87r4/84y0rPDzc5mP8UlhGbEdV1Z/jQsKJWaRWI47ILqZjL7N8VDs89r4n
FFS2SIJ6dNxj+3J65GsZdNxhVgbzLQREbXHcoPRxlgfqwSKIg+nTjvRoTjumm8MWCbG1uXhgZHer
b9OaO+9ZKRxQ3/40+QP3W6BgRvHwqQFlurbBC/F7zNVXL9J9p0QYeicmrxFtbbJSDEwH8K/O41lj
/0ua3GloA5c40GbZ7cjtPoGGFwC0bX8cHyt8pBp2gQichgJVottWeyN0tFMGyAnCVoQpiCejYqKF
UstGAWSJI11yORvAT7UrOOTbxwPx+4J0oswYusSaHQJA+uxIDsaxTnwPuIDF7uvNIMU0FCyxcjra
LOi7hGGQfjQZClzVRWCL6jhFyWr6Uprh3crm0xbAF92VCdDI/1Fu6CcecdE7RhXztm0pAhy6g9VP
Nb47ICey+gTdAC7I+SdSsTC24E3pnMele3ncNvszia6vEteasxhyE0JINRnOexVVK4+QbsXOz6er
kWEVlt2KUB2Eev2RDuFNJUFWUnTNj5+9UU+nKcul4jw6W6l1i2swKVNo87lmSKQ7dLzMrZi4eN3S
9TDTUABNzh4CaCip0pdD4tueRX88ZvcHfddgGNtCaVEGMM8Ecyu5GzagCb4HHSDIpe1130BopKnT
dgIatHl98beTWHgnyzJYTk4eMybyGxnPyPRLnjvFsqkRaf/fTHwvWcgwdvT+U1qG8HCPtGJxfUOm
brkeQjRfPE4BXFjBWQ1yLaXpkWTrMq1rprC895eKaw3RixplwmIyIvkYQbAX1KoG4SAfCgJKT7RG
B0kbzmFrepuLHE9GNztpnpPNJBfo2tMqRaqu3lGnf2zZepIyOoyQotP6RC6MhISwLgOxziNzldXd
qikV2Pq+yGzCZ4hxSg38I5K7jpRuYyeF8ZPBeFWLwhcWZE9e5k989y9pMSJHjcOP44yjmI31M2CZ
vXdCFfkmOx7cuX2uRlek/yCDSJLe5yFJnaxzNAXLsdHZzP+k6f205kWHZ847lxC1Bond3nCQr13V
FqdvPUljqTdw7pZyV9zhatP5Z13XJ75krONJrR8/osHx5q5ShyFkQPDdbJWafk7p+Hpi9uLs7+4U
S7jfiWax5uZAxZ6RuNHe0w65XxyecpWOZ0/FKeuZdFUF/RCq1mOuwrCMZiCJFm2TdP/z2JYUU1ef
oy95vinvIxgt8CWelzefTJzMiJZqrJS6L7u/U24tcZj5u2lbIYXf92B5cs0Yel3JP7DTz0KWjnCh
JC4wOePdqLxC9PuNnGyM9chxz9CgLStNeM+WNX5lN1SB/d1V6fBGvmgjzDTC6XGQftJPzuEaW1AF
PyvuQkf5qiCD6ckrFBb+McRsb2nsLcVSL232oFeIoqRhkO98B9cRksV+pNpBRhGkaeENTbnPv1YA
KzgBjzupBXJPhaooUTdxv6yB/bCBWHNKmgfcph7t3LdvjmuJhH/5I4YmE32DVC58lJayMCa1LiVa
e+HaZ2LDNOZjljw8NiLV9O9bxP++/0RxjdlV/zqycjP+RRRNfDtC0Japd9YnPmTthFv/bf4OCMDM
YHdTu46yloDgNGxlOKEaC66j2BsRpH93wjLIG25IeUN3toOCMAj+Z4vKL7b/+yViwU3f6+zD2BlE
z+/o0P1EgVvBnLERHSbpldpET81H4lTvWBGHLrSJSQh6rHaVePlh++raMqZclxM9o0TY6evhiWeh
uGwCAIeLtc9Pw5Ltj2gcJSvmzzDtNr5AGh1DzhP6G4JMqybyQ6z2So+0CQ/C3r8Ia/E2KI4HO2h9
2lDIcYV5BVyJY+/ZAf8kvOniyT9ePafVEaWWhXFzudDH1mwniDAShUFh2FJBzCAA0EpZp5dFKMLv
F4HbZ31Rc0lMyAJpfhXJ1wV3B3QeLJtVGedpQdDUdoqsCdu1Vqx91/LBnNLooX/ncjFk/+juqusC
S1ybxoKHNEmG+W66+DYMfSu+0Z7CG0rECidAnnPnMBopxjwIOsmVpvQ4s/NHNBl7EElDP++AXLdW
9AE9RctG3zFptdeVe26CcIvKM5iJW/VDozIAogP7riC7Oun0GEZB4NHcGlqzdkUblOzufjwmbLfm
q2qQsByqRAUtW54ZX/988jGd6CKayN/vxGXrbD6g8Hyn5s+fmUpu/vij4UxGL9U/9MJSGbfnnuhy
EyyM7X/m9wiUudDyMrha5HAin07K4jItG7RLY5APZoEjq4rOrCH30M909bTQ56hVfZU3Sk8YH0BA
eY/OpcyB+nfNEfBDGBtezewAQ8tElHD0o+MjW5oLIeWotjMZpwxPIz2VVHPWb91BYwAVmfnEtV6H
OqMNSdLnHbtcKMHqXfWQacfBrbLXm4zsPXEeMIN4ObbOQJhrJTSZS7MOFXBeelLI2cj+qXyHJNaG
mB3wFr1GKwP7WKnHk4EEXxI3r4E7x0SdVjJfk3Q/vvmF/lG0zQ8pT9aXD1uyC8WfnxZl/aFZTIHl
LaCnK8nxeNLHcsb2F9fk4GeyYvw7b+yo1SJGcok+TFooCfsEwyqwXeUdFcDLSXUWF0c1cDlxtYox
TX+ai/T7eQxhT92/SVPTlipTfuRraS2RBlXjy0LFuxpa/kHkpmz3kKtPJ65uMNIQYud2grnk/ejq
fDHixDVAEfvynC4QYLneY7i95oajTE69oReTyevBta2gQMtNWDH7Db3dVzb5EH2Y5NbFKLN86iK8
dftuzEnEES9d2vrmO/+kPOnduTItG5MFhxNkU6aDh0f62hFJC9xEDCAl0Vx3Jo+ZZTJbo1xcNEP7
oPMrrvdhfl83iZLkvdqnMj0U3R4EsRARtPCP+4OXyjaoBaf4qyFRF4JQxt5HJyOfVH0QRPvRxzMS
dSu01j8YsynH7hSJTAeDtwe2Fp4r0/vL+UaKU1eAFuT6E/lhAGrpM58A35pB4js6too4/e/bt5QG
CfxgugMYbdHORC/HYSGZiLFzZxJEa32GeOywVwZ/63tBvi/wJh3QlaH5NLuybzoK76PVU4fznmtx
JvZ/0D8nfKqCM2aekeacswdbH4er2DX1z0b9mmD/3IKppJT/u/igkT8ChAXcSCPe3Vd5xICau01M
2msy2vj1+E1vdIm5N3iYuP2cfkaeAZphDR2aJ7/1Ob8b4lWTOjP3jWP8HKRyeeFKao9038LJEpaG
/on/1WBFP4XvQzNNV6xiO3ZnNKeQd70AGs+52fq55Yej5Q87xHClijWhApPC2g1r254GEi2+eGII
zLMYEW4h6xUvj2MEkpJFESXyh6ZIuKgTvoDXfi4MPyoAIiOP/tr29nZgdK3pRsoWMy1mGX5OQx+y
Qn8Obwsl37RqcdbQXd14t7PBDeeUvEktzaTsLygq8pPZcJBIQbR0EXYTlEJzdnj4N3xWyZcKwotn
xDvci1w0LuhjlXRCVwUqJOa9YAALRtCtKkmFreaEETBMgAdCx5fOXYzr8PRsP78kvJMgrjCouESx
q38ojdT9fbKcZI5DDl7l4oWBr6JBO/I50t8+6Zbo7heJmc3yLCFiOxcFnZJ1FhyCuI+6NlvGDkdW
SwOSd7UGSl6Dwo+VWttgu6ncJHPdqQ2DJr0PTYWP23obEB6Ql/jwfCzFG53zj4ehxdvbXoVCqJfs
mgtmrjiaXdh88OtQHEuQhOYTHIYCxCilrZiB9v13w8owjbNHvZpoDteCqwKcBU2Gxo8ExIvuWElD
23uHu1+5zTTkIadzF+/0ZJdPzwCDB1fkKtUr3oedVW/ETz2580W/iESwvhLnJGJrnjVrMApoxysV
21AIjj3UKNT1Z/Ehz+obuw9qG4RPqJjAPka/DV+AHUYFNOZcOXb7YIrjLLAhOtUEVH3NIdRPaW7K
3M5ED0ybI9YulBOVQvE594G8tC/gc4vgB5xpansBtvqXcKNExwjaODQpnk9xcPwybT9g9qvOVKz9
yyCbHtRiI+0qhLQjwvDrnu5fRjfMGGNv0sMmXkUp+F2B7XvYIFyoeQBlzUpALtao3WRqx+vCptxZ
CX9h6hW4qbSeJ00kSkB6e6SMcGQRkiBXDB3TAxZJegDMtbfcYbvAdCZ7YOx0i8vt/4F7OAlbKoJ6
4LtqMnzsNJ2k8vUbF+JXSKACwWEMJvARn+LIb4aDDKuwx9WtPBIGWFvg9iNM883b5Qh64BWpvoPN
rXAppMFWgq3NM+4hocD7ikOgyrJDe8HmjbqFgWSFVpbsuK9bIe2y1hnK7M21jqkQSGSkJbfVtgzc
iAORDL1ySu2WfftfiJJkOhmgOrZwZvCqhXlBLr7XnIcK3tz/Q9lZC7CyLuZGGlBpOr7lAfpin9JO
34JJ2G/rRzk6mREniJz9lkZMZut8Lv+j9Y922eayQj+SfGW6bG9p1fRFMLw7778Mgm6mmZ/JRhRL
+i44/ZogyqBvLFaF/QnGL8AzloSHfbL1t/YAnwsSpuHrsMZd8iNjaAm7oymKObi1hQk0Ez/vHWZT
79vMFebPlnYaAy5mCfEttS1bwbhB/KNFDfp0M74KD/p3wQje7xfSQ/WgHgSXGraIvRRGZ5BKgOxJ
v1EtGMYVpkh9ix29VU/dfyxewH8XuNAnDf6Z1RQFWRD75NdLJzRm9kqAqLfLptrYGzuXikaV5zJq
gtnSakyiJgWWw8kysI9ZBQyeGIJHoWIFSSkju4q9Sza/G/OxJaEhFjRi1gvM9OaMhCLZiJP3K1Nd
Rhztz4bxL3DE8Cpv5DBS48UpKcN/84+pThN3EvlHmzQ5FbOnWpoTnz9eGl0668feRxN4pnXHsaqU
UJrRf2IMT9I6n2TGWBns1ZbfgzAEJvWF19pvrXONvbBWJJHiShfFlixdBeZJx7FeczQ4V+LoMaXF
XQXjdhZEUfjFirqLrfJL2sOlitOf/glt7oqmAinQi4zofKLlESEGTcOIHDgD2fNEOufxR2YOMRRt
1hcm/vjeT9S7DPcHtR9sRIuMCVdUbSbDIeCw5r6bd2EtZjjXb/D/IGpodgEeJfgZXQd10Nh2Gqd6
iRp2fNUr1hTxMfH8SUZsW2zDwc2+Jx7rRNNRv09HqeToFVry/qGRd3bFWckahcof6+cfx5uiuxNN
5Bdd/TeWMw1u6sec3b8nsr3FGMEx4k8502lTUly6snmcaiv3cCBmgxNIw67Dm/mP+6dplgFXyz45
230SqKmcHm6cr7a7FUYpeGltt4FccujOpeD0fEnqhnshg7imu0PGs+KohbmRsSFdFQ7mkdM/+mdD
1tDHzWaaiIl2h5UN9cTVXYJUNinBA/jd9ayQ/bXo7NjDriygbec+1ajebEh/J3uZGKVOmfG9gI7V
+TFr24fOyAYMal+9e5S9B8Rr6YrKLHNtdyjeaNCWsjg68GE/JG/yTfUYsrui0KWAywo6bdeowmrK
YIV4qR4lW41sr7x5aTj5u9CenD/SEL2QyaPB+d4GTvEM1gHiT1z6vnBT3OnwNFNYFrn6VtX7fDI0
KbE0xQzDvy8vU5KkewPCFwgq5zpf0M8XT3VqDotkrFOYH4N45VsbH9UOKu+4I7nJp0Z1l90w6x9K
ZW+EwAYXgUA5V0ezOh7wlf16Kmxj7Mks9Orx2nJt2gxZVYgWpeBQISM3b/EMyqX24fM3jwFXk0Xl
yNDzp5P+Wz9kBSp2S3NQPV5b/9KNT1blJA5lAWnrZVgQmz64jNKIf8bzvA6SHUCLIwN3vb/c76rV
gOcOjsFk4oUDwfFDPA171cMSOi/nLa4TsFTyZN3N00ndC15MjFc0yfScssygGVzRTgAg11ltRV/L
N2QEKnMvYy7q4TTONaFNFypfyAjq+bCj5r6nw72Oln6BM12sT9NKiTN49U+lzWZD/BC4XNjm/vnX
kaTOLA82VpAlrwaEiSqu9gWziyBifLbk4iP9J8DQR53+Cgw6abBAdL0MhlwNVRPndxKIqMxKJyYS
ElIm4qItEAPbwg7o6BYQoRqE3nIN3T5wSmlfMyKXX8MPI5NRxjeNsYvpJBfBPAf5QfroRglPsiv3
JPrfB2xY0UigiJhAegtgJGyivlcXRcScO5Q09iAycAh0b9qC27CdE2eNe2gJWIRdtcUFjJK2TEoQ
Y5BZ+WAZvzhkBIyEvXuSNedmGUVChuK11rpjapRzEspk8HtBUvTwsKCwOAW7m5cChz/906wi0EmN
1FiF2iJMdNssRXp9BqNXoyn3OjEcy5pzsIm9fTPAu1SepuVmEqaPoPljPqMtX/YZB/alTod5jtFn
JXNA09MHV0WwCxm0LGAE39wxa9v907jVVBOPq1CkoMM++g5zVPbUzg3Caf8h7UWRkv7xENZt7o1W
D8umhcZPoQ1i9P6lcU5M+GlOhi45r2UlwM2sc9F+E2+0DyGBEC1VWyPcAcX2M9U6Cb8BlHHlwW1B
tZEW+VKGGYUsmHGlBsVCTWj9Fr8JaW6fMKpfK7Abgd3711Nbgp8J+Oiryzydpqe2zlCDIweG6YPL
n6PPzkTr3oyvX9daqnOG93G7dqeDwfceL90+jLNV50SASGhn+1rG7T3JuKA8PucZKhPVS3CZlhLs
+ksGQaEmmUy9jUZkONFtZrfLN3HA9HUglabggulnJ+StGOI63qiZs/XIZ/kcfLN3EkdtJtUytSB/
PBQs3Gqw0c3tCz0klMW/E+uw2HM+H0AXtDBJK1jtg/tkedJJkdKWsieJ35dL19UjlCks7kG5z9h9
dwH7Lu+Zbh/jNAEpOE3/5mX6rHL7lmlw2rLnmG6t1PD2m5Xl0eACHFivI+059iEDyvHUk+Qnj95c
POg4/IWD5P6xVwm5OiSrib3Jhuxn7aSX5h2yu/hnPxb2gDeHpVxnvL3y9dMUIoDhVaiL+QuxHE9R
I6Ebdzw3ut1+GhcLLKgBJJhLYcYmD1jcD4ehb3ThKFJwSK7EK7bKnUDcKXUHal5BeGx0ZUmnMF4d
WdTf0In2TO9wTh1YulwkWJtKSKoxYi6tsieumiSDPEdbA8elVC2dmhFANvqOQMtjWzRQBSJSMzoM
Jwlce5gS2jJSgpZn5HyExN88Z2dCJTc8iNHtHj/YRdqf7YyRu+TQi9WJ64w7h3ytK8FPnAyjIPHt
08H/iLjJCq5JCeN8ah9GgOjRdKgg+jloORnXrZfzV5saieQhWprUhi7mtWU55E5mveFYLzz12b8q
h8uAy/KzKNrTnbte1CJ3SRY62EovzhNiW8SifOFVWQTuxoerANy5RGT34gQO1+gQ8N2v4oixEfnp
X7LEMzb1aVuYaU31jiWsSC/hsF7dtwbZZSbGkU1BzoLehWv4CUePMJQoaI9FOx2aVC+Az5CXYQKb
x20qWFmO+H9iGW0CRSsIcvRFWjwGO0iL78Ke0ezogzvFYasS9Mp3GjXhztU6qhNIl7KZn4ngSlpB
YPsVj56Vzu5e5atb6gRN60wWpKDwU2PcJdk5KPZA916cJ31m60CjUYldIdOit4m2upyuVZIAJuoX
Moi1Ia+pJ5o6zkZAjfwhnp4aWJ8rEVC3PdXyBkimLihfIo173A8pn35Pq0OCo6wMACMdGKpPBvzT
IrR6QD/8wvpoMo5wwPr1grW9yIkefUBxbsjJvaumLTwLoe598wF7KSr935oZXBdOt/Ry3nodT9pD
y7BeklwqjtbtfrIXz6vfq4XjsG5Zqqd6KWrnR9B8j3dCQzRHMW8BehwgQxcu0rXT8aXnfXTaSefh
MyispwlBBBywZYowpUOaY75PWg7Ofe93FwaSy0IaQMoPRMrLqUBsfAETiKkRebE5oI+7EchVDbqd
45UkGWNbndoV1YwJ2C+Yn4IZhG16JWz5Bk45DjCGrRiX0RkX4cZoqmIffb/y/1lrAJzYbkvdn9wq
Dsul2ZiPj7Yqk1AOwWRc8+hZOiqIpym/AaEsOL43X3RTthGWkMJmePD9jHhlskq/OCp87RMb2oiy
Cj9xg8ExbQ7cXRq2DgnitGRqgdTUXhK5gSvZV5oklemLyiHMx4BiizpWYCGYFDuz2Er4di/1/t8O
KRvlkK6xab8PANy53TZ+hQoUDmIm1RdpDbLlTXD64fW/Own8vde/LfRAGvEvwdKOKKVgSZMTS9+w
LTCmKz+djCrKC9/4uzUN1G3Q4/L0xdsWfpRDq6+cp19Ddl+3QzNP6VYqPnWRB8ZifzZu3EcSf3FC
RZPBcoYkVmsx1skHDvU03kjBZ29uxIPxw1KDPp44FtuiuTnmt1ND53vbMnDIMsr7Xnyfw/gEy67q
NlSH3gdTMQYmqg4at50qVqloGv4RfjWY2r5+3sfmoNe3DCOnALCG+K1CzhTcuka8rWE7HWAI0vO/
1hNYFv1HLDbXbo6YaC8y3fSSVwdP/qbi4CPs2/RwejDrFNOfCPG2u2wwiS1nufVR6qHVrV0SmyFo
HvKws2NazmqCpVF1WsgmoayE1UCzMRLYgtw/UEwO5TijogBJ+idhE8tL5k32u6akfYuENoa2bX37
9x/PYdM+yN6iCjTtEQct3o+B3gJujS9ropNb3BfwdY0mkMO4RecRVlV91GBLhP4EL19r4yC2edvx
AeB40E1tOBdm4x4UXT3cVOklf90P7tFXWryLplEVJfQu5Dxmv3uRW9xDSK55f9ul6cKMQt8Z8BX0
WS/lDrV6pW5UIgjlE65vWeXJM8KIpYbDOLVdplk2sgPlXboSRG5ivL3jIOA6iOXDpke17jEi+ymC
MTi25XZ13TBXWXY4rcwe0w1j9HOI1uZzaQsyeEE5LhLlLDW14sEWT5m0sCJf5qGIElkt9oXVgRsR
n2WWmOLSJuQCtnX0mjzEAJr54BrQYsxOt4Eu0TfZipk7jq6tjblKWg4On6cTvfYyzYT1dz9k7hKo
B+p2unAH4xvSdkBbN3nMWIiv2EUoQZDB7ZKEqOlTbmna1gfh9HTxvZrqdDbgwRkY/H4U1/HF/PE5
PrnFRxnlHLFBh7f8/N10EYogkB96Cjg9RMfVNpB98fx4b13zsxRgOPSAIScRPZRxRmwHHCbs3tRK
9Y/cWp8LhJHtGBy7F1oeN/hm314gIu7LgQOpdG9G3d6Z9sZWvMtO0Imbi4pOqr6zi0wgrlxXXD7f
TKMWVjQ4obGqsG9pcQh9YRiS9IB1uPSwvvmVpBAHHV1RsyYLxuqWefHAWz+P4mvPgcUUgUzPZ0sa
xCW6UXnABZDhz9c+2Wy2PfUOlS4GHeOY7xolAOTXLYiiPVdxk6RP+xvBvlU5/H0MZRcoSgPSc8xD
ioJrS3yCms3DVLJbxZYegDtc+0Y4S2S0EnfY2KVVqJC9ygfd8nfjtxoTu5s0kjDdzMWiB/yinr16
MA8wXOWkxxGQUdXKRFwJGUey0moAU3Yiti59zWPELO1GY/vSvqJZOYiZeEd9XfcnHMDM4MLxm9I1
6gH/VT+hLB1gp+WlH0GWQGQ3F2xapYAAdhcgdCyCzh+35RBK4mDkxVnWCplYT2IvxnHyWoHWlhP1
MXMdOjEVSLIouaB6cYP3Uhzj0UghHuJese38hE+ai9J22yNi9jfFChlY3iX3GRgzW6yfgav8TrZI
0TA5DEP7GhuE244R9dFsPcTwmkcierfkEKXGPicVO6FuVzRSwLHV9F6ZPa25loTFWh5TncsSbjER
Fe2AVB5koA39qPHQe5n91ZD938pXSAEri5fOTdzPsG3Ib5rAGzPVJ3OGfdW40bNKLYqr+beyEjBk
0pGkzczUd4MJDTxEfa1P14vOcB6hUvEUHccwhjzYs5BksqRZhcqCmNuo3uyccJQ3tRPYsrtOd+HD
ZOoFawx8ftNB4SnrLtnFLUvJDDXwFyE9MX4pxgFAU5cf9doW+qGxBGWFmUF19QhefJsSLexjf1UI
bV53c1anprgudNPpwBXt7ikHl1AEJvp0vON4YU8KzW8iYe2sdvYs0PADWAbd1SSuG4j5uEzwJZPX
HLD964LTRy/csenRKgaEFZriaGJ8fEKvKvyGRRlbrRf/ON0d73dOzVH6KWekY/6cOJflsEy+GAMC
tywdhXLOOnaNbDsW8hwtOTtMQfNOhUg4zBNJOZwYA7txLWitD9BT4r7YoZb7h20noP0TsD+A7xvY
CYoWczj4XwZhhyAEqotKA3Ywa2apfttO0oVFLuAx6V/CholiqRK44xdF95x8zoXGgg+1exmVIj+1
uJqILQ0NzbnTsELdvpSco+zdo2jqGlOJsCSYlvm3dAt2c6fgBVdyITCd273VBKLsDNmmwyXdqGik
Pza41kOPQO9+/urJMCttdyshuSO/UTNKA4DPAgr07K9LViKddqr3hswsUzX3/KzupIW5eyxzmeYW
UwIMHBHOWBV/GsSq+fT2Cm3mHMWn2wdvM3hQzxYSH2ewbQKghzS4LoGQy+Ce7UpUMt0CjD3o6fNA
d1IC6prQTv5DdgtIYHFWWfPS9RSCQtK6NJpf0vFkXrzRyxm01mcMJ9N/VIaNKyV66LN8oDnJkyUw
1lDYI1YJmTdF5Zyu3Jf4znU5HJ2IeXT7drBWSv3XJjXpdKZeyXbQugi9rMTxd7ynMEkLR+SdLVU1
Z6p0penBW74XJeUkTJ7pr4dbZF/2ACDXzlHmO4uivkj5xakt6HGuYA9l997cOQSOBefEm1QRiRNe
YTqQCgSG2jtxyg8b0uFeOavO6IxmeWAVbO3Af11r1SH9JzyeH/dTYKnqV0Suk9HCLoXMrjHFFAF2
LFddgS+SoSaP104IWnGba0Ds6KsTeuW+ucyg9MgkWaHotfx1qbeCNT7w14cZAZ3ZsIS+Kv0+90+T
zLXl9mAucb9FQElUEPSwiP9Zgz8j7HWNAN16lhFpbMM4oLiKA9oVrIZh85EcuMPNwvCsFF4ktfLo
y/mXTpmP+b+TyFv5Ysimm716HF2UQ/BVVjWmVcgOZsR6iSS9qgUoaB4/DnBf30YmoUSxsDz2jVgY
gYN98nIdgdDNrhKYwHyXlcFjmle++8OUb8bFZWKcWjmqF2z1RRdxPabJpIB4zR79h8ZMYY2+7opQ
/V1pxQ9RWksMBcV/p7OcdKu0rqTP+crIsCD2xd0+bohOEae7LmAVBDb+fapDq1mioPkiTshV4rVq
fjaEDzF1WHrxi5TfCujLUHudJkp4DGprLekzZedacN1n1OLCdQmxFhW4032D252G0ED0amS4cfWJ
4V9wXba0je16t6fP9SgK7tNUwfMY5uFtPPPu7lQTmwzHK+2pWj7VK2u7rY188zbalJn+ucfnQ/9L
91WloXLA/HYB+9+v80WfIsQHXRz8c5tTSFm/sz2b89ZMET1OvpAQIDXWSLzm5IVdCmZfkPTY9xm+
9wKKcFjiaW873E37meWqTh7CgP9MFP0fmUNzKi3b7B/sGs93dcPJWh/mPYE1UWDjaX4AnQnd/8d5
sfey0bI47ZoxvScx2wVnzteql3NwHrcHG9OTlcezDSNkfoBBWU7aPg0tz6+CCpSmMUEhb2HfazQ0
3epGWk8gChlvY7h1BiBClqMAEs0aMWyUMH+0YkvPrRpp9VWUxMHyJkEl8olAwN2b4fGy2Usa1/0B
pIdFMF/vvxhyySj7jQxW1Qqsz2ad1uyjPdQTngRGwurOYgHgiDCcf25QPNEZfjyiuPzHq+NOvVoN
UOW1NMdQHUFCoasJdeBvG4IoujprkAaMCZDMjdDcs8SmUzGyUgV2V7c4QJ4aYxpbR2dl4u2aISNQ
KdqBl5lAmOU0Fjfg4YhBup82HwXHBTFXF3dNYrinjjb267cGfK/qgJdT6usR0CKn2c8BCYJq0QQ1
yndr1y4+dqkn7QfMA1OQgA1iBNfbyNFcf7mRc11pWI16elzGDjAzZWavTnWIbvykAkyFSt2rsuD0
f8UoZqqAgjXs3xqMROhrfYycDGrCS7bp7OQW+hl3wsGE44blqrDdny58NF83dRkabarmEV/HMPBS
hpZ6JqdoGU+hvgXf086ywALGjXJsL7zb4EpWVbidaLeC2SVLqIQ8ZZsCJWPn7Qk1ItZD8bjnNAwb
e9mGOH7tMiv9/gZAFJ2I//FWCDIa9Fe9aYnvtgAzAZzUwFM/rmfyarzIF6xbnEC/nx6v5ylq8riL
K/z0xwWnk+6yU4b11qYrN/dI7cgrLEUBioHuO3J/DHIZ6x4r3o66Y0fKoaep7QNgbqDuSW52jpFe
5wROTsFzQzxaVKUKruYX7NOjpoVkcjLiZlx0ejEsvn0gLuiqKEfdLliLT2J5wdYJRElvD5ZZgveH
slczkmP6baGucZlA2rzrABDi4vxmTjVC40k9kjHff648AEz988GeywPeWJdEbjQo+1NcTyz/DcCE
q/9847daQjOzkbA5Kfif0MTNXto5rXZGFBHiJahsrG88wAFmPPtjSYcQRCJ/CoQ6bF2twmtlTLF1
hGt1QvmTkzd2mcAtAhnZ2E7IP1ToPUTKomONFUlTuBrjSftJr1UAqKUwMtNTf8J/+Qvjur4bDvln
2Zhnlrmsf2TTcwg1yR34e0mHfGhpHIrbuYKj9ywtNhK12BB30SdhcrEwdg52OjPGh4pi6mu2eZeE
pg0hYFRA7EM39UoAjnkcDfhne8vqta4wy1hjPTunOtACoAXK2HU45xRmqM0PMDL9QCxXpAbCeM9E
axEVqolB4i5yG8NezzwkuTdsd4e9hk3003EDb9KfZ/DpHq1fasEUrj7i6Z6Rt3FRuo0Img0yQ16I
OMEgCB2dfLvD/WQILvDepTwCA5jOS8b0HW+ktz4xngJi8l4iC2hxUYgzq7dvDSPP5/0MLi84hoDH
+iA3VNJRfRKm87dTKHu3sfBM+zeoI6qzv4KUcJckGkVpP++WRANgHE5fQTVOtQFJiQIrSV58SpYT
/jk5ZxJYmvC9r9aJgvOm8ob+fW48/L/JtIEVnDzRw4MQOpjWNsec9KmuyRz1iQFvhY4e/kbzkd/A
PDECu6OsSK0CYdAksdi9OeRBKaweqybYCcec8yVMcCO4Ey08AaWFDeLrEN22JvF5d/Mo7r0LCyTO
+WQWxttBbYO4PqlGrfnPPTmjeMChADKo06737HlUd4/9t6Ypa3HeV+c5kUw84cWWh8LKIi3czEEe
q8zeo2KPHZxR184bFHjA0qOXRatg4QSHnowWgeU4g4F3I0vR18KWYH3JIEJnwLrCgi1ABwZoe+po
dVVaClo7n+Cq3tjXVgOujMnLoJC/Adq8zRHzvUh4JmoroyEcGRAfxJsI2ivz7PJp2ZSuwcVMkOB5
lQosB97fPoMYVhYEgyHXZUHux42W/Jnis+00HCysF1qJliPFfnNKGGeHV9va4frDMRt6dDMqFN9C
EDIxmpJPeIMrCx8RcaJ+9qifdD5lf18jWjRsf2+u8FWxtdPQ0jP32k+jk3Tlv73lWcrWprBA9JEL
+ucq6wHuK22iMqoCT5s79goHFLl/HUzfmqcBlsYiekLRF9dfB1ErgJ7Sci54YUZM4jj/WWwvMxcW
DRI33BiL3UN4SXzNq4dHyJjpq2DklNqVBH3eAULuyMQd8dnNljsFas6gV18ruYS/yJut95ZtK/M3
WtJIGYKujIZgrNcq9TlWL1qty0BVpxyevEEYChCrPgtu3jtszcIYzV8LRj7DwITp7TGLJPzqtiBJ
/WSj9oHmd64XwD0IRK5e4wc6nQcvRA+xChw2wiANM9Oo6jh1GkC3YSZJ8zNvwyzHal5VtVYFkBd8
1R5DYGWqhNIf5futQLs7JVDLp3334rOEF/l7eRl9LSLkAejYHvl9r4kBNa/s9VJKvwjrDYQ2Z6Fu
9Kl56yxnBvbbjQfSgih/SR2CFraEZeoo1O7TnMopqCLsvgoHpzW8EQVASBXTgDpjJn3EZAeLzss5
2h8M5Vmk1JRs5/D8KmEEuSpt/XV/f+S/UwBaGQ91K4GwomWjD+kWjuzsOsbqKwp8w5XpXtfSgD+c
z7nB/8kiYbVqDIN51f8zAKuoW8CBYm4NzWjCUKePKHTjoOmN5G9u1i+JpPUaufyhGY7RDr0SFo2z
MGt7R2hGqVRLeVo0OKAPFd4fvi3g0UhlOOfQurw40YHFlsMVGh3paSZBonZpQjuwYAhMfrBjyMGB
Ek8mbfrKpymEBmI5q9kS783WMEAcNPBfN6jc+27qtxf8kS1Fvqq+dGkjQm4mm2C3Hy/6fgGcsYgY
uttR7taPcAq/asIKpfRbSVcfPStRaJmWybWu9/zydE7sIjcMpfcG37f6cHpL1/uyy8EqU2RFzUe4
m6ixiQ7FP57eKPIcuD2Hg8y6nivHNGum30ngDPdfdz3Gh3WBYY6eGhLeHtIdxbRKeNQllX+/iISt
ef0cDOVwz+9k8nvcRWzcEBRgStFi4TM3L+enunnen+pTEgJWtSVK2m2gKLM6l1hduXOHVv3Ocfda
N25fHWd2nJbNvtHHJsoYn7mNWOKzyn5NssoQx4y4Bg/mgYXvl4FNwrHCtDzH//c/VYXvluudsTNY
G/+St1wyX+jyZ1WwLCHC1Vr1K9btWZ4gUqnMQJYYo+liPyiS61EzB7RUE1+m8wsuJ8PryGSSd/M0
xnagPAaIffZRb2t12RhUZe5dUb3w+r2C4zAFbrNvBVVDjEFunJVG5LJh11I0N4qVXxhsJNUiGkK9
k7/llHTSIoK1OfVwXAyWhESwPJhQLjr2vbm/Qwz0uymualDutI4bWIln4ZVFg+v335nidIr+aeMv
o751HStdVFQC83BOX1i+u2UnoS0aWyOaXORrK81QQfyDCVhVOadfA71x2iuOYLXNGvm1m0il8bFJ
f75miq2ZoFOHEtynz0gJlGARhD09eRp9G4sxZabTRF9BFpKc4HnTMs9+FDDKBBdAFDlPlHCocsMa
eeCw1DmNER0/YFY4oaBSJOK1V2hXcfVKDoWLdDAHkBg349BoB+Iz7VLPjzBRwxdOsirW7IZoGkea
puwCfwdV6oSz2gWme5H0CGmdOTjRNxVfL8A7Ht24m/PBqRSLuZq1POL9GI1uGO3LdpC7gQ2DijNp
IsKm5OZqc/2E4YsvtyRg8suijFcLkUwG/CK8d2Mr4msHgeJdJ9TaEs1Jv0GIZUBTRKONkQk9cPjK
MG3OpUc4uTBOSOBJ5G4ezAASL3NJgaH6mhT1WlCucAS+7OhqbzXjNXOcNoh+WFbTL0CrVN0IgC65
aTiXp8ARGBOeNLlmwmEkN+qVoFZsdd20puvj63Ri84dbyxD+nBVKn0MWFGMSXja+Q5nJSofnVtls
jzp+wUZ854FBlJsIPbysSDILIF9R8B/eOuwg+V2j2fLgb+fAMBoyoPbw8rzZ8D90DZkNR6um9Zrq
niFhFC18BOHbul0w0dEIoMez5qF0ahiVnzDUxXpzxH4aImzlUZpGOtkHS0BC4y5IEECjRNIf0dJi
V5u2YDzEjBEIB+lg1sMi/bVlJD6eAEdQSl101ND4Qr1B77mwI2FX/H1id0HMewzlGp+bDb0S05Ee
CvlvwIiRgyM7kED80y9652I3g39pWCLY2u9Bfss3czhXISudCfAfN0vbEBg1Tse4hr4BYNwk14NG
JiWbOxFIrxv3qkHN9nLxaj0CcbSV1hj4IrQ5bN3G/8L1VmX+6X8jzwnV1dYGbaksoUV1S+Shwg2t
gAAMaAPeaNm+I/pTgHHqFOqgpD4k1AIx+ym9WO9DY3ixGq0qQfqMAenu5g8WXYy79Xaibdq9GjY+
KjNQQ7wqh6eokD+Eu+4SqIBQxesQms6gGG96Ilpv/P6wKPVaYduS5ufdz+X0Ghq/dbMZcpl6AlEw
fV1S3KKAyQ/airMeipdqZ6hIRBA8xg3CMrnqYz0BtDGC4xGoJ4jQWSf8pBxt/EA+wo+sIIa5Mkpl
QQaRTVzcjMX/CaY4OZ2EDp5yj09vVZQaXjTq11lXGVp4O+d0issPsUPxCN01LdVnyt55H49XCE1p
vQm+OzpA2LmdYAFi0RrfqVyBZzszz3MUpVyl/uTIPbhHPkq/O+9tdmdRXl899p7BHkC/aEqgSBSf
t5ddu6xzk2jSDmcfEdGhjbRAAHQbbgJ5WrsoiScoXuhbVJGlK3TRrL/rOJWobbkK2WcL85QvVTRs
G3O+TB/QtAkTKzwf0QMWEDus6DSCr45c4rdK1gFROEc+UqHt3ddrVovtCq5CgfKrIboPw9vpe9te
nBf7888T5V+gc02fR0if0QHDWyBuw996zFaXc6B4IoFOV00d3RNBrMAFpWRpPlZyCh11cjB5LEO7
oY8Fav8AqoekF6vLVofK7GvvSoyK8Tg2UdzDLRNkWYqrN8asEdGsev0iXprsChk1xqtDErp2uEf7
NlfBmvLnDboZv3XFTGFpinrmZzJwtmJKnRzP3lvDYWKz2DLHctzCYbe7nDRQE5HLmZBrp9ZYfxPf
v6OTDPYBR6xTCoVkhFUYbDJKQYjWbhzSmsB2fAdzv5dFo1vibXGDeSyIxDWjiHFz4sPRKiwUmS9Z
nN12lywFT9Lc1GXX0IXu3YaEX7V0hwNC065zT58YsishAV1dn+jPgTHjkUEK+5FKZXFO7RR6JAEj
sdU5ZVpAzG3NYBo4++P9XRxHODgumiMmn8LmBRFFs4Lj0Ocotd3Y0YPVq4boyDQSjYEahnRFc9Rv
AZpxG7K3o6VkNNCSUSxOnwr3biH4OpI0jbenPul0w/gISbrK0xJWHrnLSSVdvywTbJDtCEhYErVF
rUqdOU7d8UYVX6SgJsAIAyba9TVs2E2l1MuPk4ANMYpDrvCRvS8pDTAQAwVsfgSZJhb1K1l+SoH+
7r85PNdgRgGIHA4HuGPtJmZHdTP93yH/Uwo21iCMWJiNIjw4lCtU3e4pq6so4OF7OJJ3YdFpo4Id
+0FCJH39+LvDRKLWVhsE+34ltDyBX8ZyMHUVp/ic0FTLVZPTw/4+n5+oQWyFlAc2pQktXvBA+uPw
LS2pAD9ZNDbjsApcx0P0/++dNCp0tx1IA9pzs7mJI2JjZSYFROu5Hf/mo36PhbjMerVXo98bwKZf
VE1S9CsU2x8Xe6FK7xvmhszxy4DGbTpT1d+c/YfXgrihxDuaRoFwSdDSx6LSXUXTFw7F3t2M4kGl
GALrx7ReS9ql6eQaoTJtH465mDo7VxUjXDj7n2b8gbspi2MaOq3qdPr/HFyC6SSJr8ojy3zxicYR
WgBFT7bwMSBQFDHjl3Vf102FZe9fiBt4AHEocHmFJdfXuOX/J91X/rZ0TMpzLXAH318vEhM2kT2F
dHgxZWYEM8U5R68mxiVLN2xONH6h4xL5ids3QWCRqhPGylc8GV61xfeOtR0E1JSjAER6Do04kZhq
eP8L38i3SoqqFI+AE/BrtdOM+Y6zKeyjkDoeUdllmfO1KRtO5DhxK4l4Lmwt+dPpAsyVUDEnYO7Q
t5sEnggc8quK6RCK663zjBQ2lP1qQJxnxQGt3AiOmd+h1nAIVLLbuqOpL8T2CuzYjS4j5o8zCxZx
IIyoD5qlg6ioNFJ949JrLsHB5LkA/FFoyuq246NEb1tKzLJfZG/8BqLrSEyAwr9j5ttPiCPp3F16
2Z5Oj58F9DqoITuBArEAPYsepJ8BPx06IJn3swXoJo1Kg1c/HbTnXYYihL0B6niCeNzXe+nz6tVZ
Nj5ii/Ee/fP/TLHe4s26pZ/7/p9ayMfN4Z9jwguU5ZIdfGUacyFS2bpN5/VoHpoPS3/fgsKV8N+D
JR8QhDK458/SKRb2fOZxx+whoC7U25vdoRYkEVjPT1jljcKSLb1m3Fqfr4PuP1SiSa92HJv/aE1X
FdqQb2jQk3aH/GqvlW7U+1lK4cI8e8dHXXiR2IF04Nfqxl17o+Fjc+TTbeOx7u4Q9jyQGi/OTEa0
YPnZWFWTK/Q5j9N1ZDwmg+1wktLWgNJEYtX89wFN4zjc28S54Iq08rzYNboaRezePGEnQ2g4ChtA
Z5m9mIvkY1SEyE+WcWk1dKAyec2vIJpQaB07kvd/G3i+j6t8ypz7OVKsqocO0HIDocbVCwQkkjCO
18OrD/LEKDvT4niItHscePSuQznMnZN67Yvn0/1f/N9JwFrYF3wWKxiVuQqfZ6V1Ot2qFPxvQqEw
lmFmkQpRHKkLcnWtcYd+vsl3j791ara/scfgkOAbC+3cviUBPEForxaPZWEGR11vlhKBZDsvz5M5
1hT/wr5eyTSITSAfMRkCM0J0rVudzE6jt//J+d0Qj6Ih+C3EFbOT7yUS1deqSs+osrxSp9IZYWwR
SUHocJQD9iHSc5+WskqRIAcbeBfMp8ZNRc9Uk1HPb6SuJmSDJ2OQ8ndpxsL8M9UB7GtHZRgW+Ll9
RarYU17i9LxHEruRWnggwhgmgt0MmSIJ2gEme/vXqDGmcg1gjiWju59s8HXXsf2ivap4VkokHKbQ
wQOmOw2WiIgaAjNuMRPZjhHiDUBMla9VXLeS7T6lx/7kgAS3+yEymD/yJQOT/j9clSwjSRA3ekrs
nj2XH3mpbZpJdag5Ah//IYKB/jYVT5Xdy7IlgT0bIIbvBlGg9EadwxmQ6ku7OH2D4ICgATMSFLs8
CNWpvYjSs6jPjPvO/PqPTqmu3U5zE7OBqt9sPCtWkEOsexQbM8bO39LrwLOPpqOFlUoS5k/UDwg+
6jfI1PoLbDwX8sd8l+BGjXZphQehu1TtM9Bu17h8t01banYbRN3Ttq3PFVGqV+ouPX2tCqFrSPph
TAQUw3TQS8vLPNJXCdSreeTghpSY3oN+wSbRw7tJ603xKcAF8oJNxGS50SRKR3TLPleFSqKp4nd6
CyX7fYDpYHQCj4M/CRMAF2TswdFdqzVcQtvKWha8OydDrKmK8hO6YAD/524CAAC4JWNs/n6pl6DO
ZYNbho/96czPMs4VhRRHFcKYvwzTXOeZ1bFx+PfVhOMsjb4pzdHLV0ZscKy0td7MF3gsAAKMbaxh
OVxUbkIrmnxDAv16MIVNbPIkce72x62tQONJgIKQOfB6YPoEiS0REmNTobqR9ckS1H5EProkpeEr
k9f+8f0zwUk+2S1kvgW224rOWxlP6/CKMkBeD7jPkiC8qQ2Oq+0lqwJt94bn6Ly6fcs1b+wBnRG4
SomuDAqyWsTgDieSm+t+uaDjZPG+v0UhThwaX4+FWLTcvmHlf6zpdD0I/GWN0ufElIsbaFCTltsV
57+QKonzTvuT8W5Avo1GfJuWqDWD1+vnDDvD+zPF13BU4iTaMCoNT/hFPHpUR349Bn6P60Wf+ZeB
23xMhugjf4cKs7TtGfXotDPMLqCb4vBU61zMIjzAy/AxkuN0Jurif0jSnMr7C+fEbpwosQdT0dRA
dt2+0XIhPKQSiw97FHpA9LCG+TYPF6kf5ztSAZ9fps/3kfRNZsK0PzKlx7jenrDS4bIz9B+mLnbD
SxIr77+YWW9ZNHjHC4Shb1urgMQSixN2z7UwGUvCTeu7U0klQNz0hEHT6FFgTYEFLa+beaZzVxQ5
/V2kDjvw23LolOCT9DokSod1woDxhOWYlnymr7ggO++hz/ktxsovztXq9YiYm5uFf+ZE62jWNClY
v5OC/NzzfmBPD88WOIrh1yJovamaSBiJN+iDAaHjh1lLGyfJuGwr0zkj7VbmtuBEm3fl8Y1w6IBW
IMlNfw4gR05KaK7t9DQBSaeF0aQksIIU6vSqL+rOQuRc3kEAZrx9w4q5bixfRpfCay94+6240PKl
LNdjPkIqqrA271AdLsRuoS9EH8263k2OE1D1lOJIrSnPKUyeVyRWhJAvaIF+QStDuu2VoVc0KURx
lsEWOIkCOJnEyMkAIjHhmiDoqK4LWOIq7sTIpcmEyJzAxoaDMkhAq4RHXLj8GF8SngEnqcKi3aoy
JHNYzZmoGIAn6HXHBiUKbFvaww6ZNtgip3N+yC5paSW1sx+4p/zIYWo2xlkAvZGvPRPUpSG8Ysbw
MfZ7iKEnWme2LfE8Zs0TLTJelf+08ujXAr9toUr1HSD3hq1nfSCnEA2/OZMQZpj+y4yu3slxK0i/
SxhCanRiS9pfppzt3nxiERcBPjGvNIa0F9wHc3QRfEbx2dFiFsT+d1EIe16y/tWcTIugM3ai9qNW
s5amhfAZT3OBzFEf7lkbU3aU+WRVRZo2QF1B3txluOI3uMkm3+rqGZnNYe2eU1ktRuXPlBcEHMN9
QySBzfY0Ppa+aIWoOgEV+3BOntwoG/HE0O4VR3P8iHcUhuQoHJiwN5CL70rrBMEG9SE7LAWxsyTg
NRSK/r9TFOxs3ftXQLdJfqx8VroWqdpyFR6UQXm+s5JCP65Jhx1qmaI2SleopxUjo6sHVz6apU7w
KIXF4fhsSxp26Ah/JlFFadmzWBT0RVuU5XKv6kkwFzVlLOT+FHVgZJ7emtR5ZWmF4uhQHTb5Qh8/
RqsihijUnoIYxBzqZfwlhtxgy4E2ZWs4EV5gHfpU8wbMWBsKk2le+sjzBogoFHDqeF6NXTw8UmeB
9ti6bVi4IDGzRoOXYkQH/Q8c7C1QqGNgGsodynlrGTlJQQCBAtbfW2DOOLfAeV0coqWY+TwrYhZ1
TbEMapQHs3yJZNPTRykF3NGmjGkNZDdD7O8GpUxwXIMcm4YqduBN93Wq7/+Jbhx16nFRnw0+l2Hr
y1K69PW9dxRSBIa82K9shWWrAtOLcP2C70mgyNeq72pQrDI8Xao6mKj4MFqGlWdpv/wlV/ZlPvxC
CojZHOXCn5CBZgyUarIOyThZrsf1jK+6S9MROg1M78fDtYrSL3tWDpgYuN8C6SM32QHhle4bq8ju
cFHNpUW48JDHISu8rzVGAIghveHDoUJNOcrqjsIZOt9JjUxZWY6CrWpOCk2ZaJmgwCTaz15lK4Mr
fsnABXDh2RJE4AW6wK4/mZa/DnL+L7ex/co/skk7pqPNsxZ0lmetYj/n1qe6IhUKzPjjaIyLaqQd
RZeFzJZlEn7hmVmnJhtQewYX9kFuWyd5saE9HKnrDfoSH3t8MyVJa0eazZ2GGaNPjyHtwjXy/eyY
EXevFN+CrrEQ36Sz5wQh+Gh1L/tUZa+mB/TXm8IPQ3R0dceR4v71F6JIjF6arm6C3wpGfKcvYwoG
+oB+mlO6B1gWme/wZgCqk5FMm6/HvkxiY+urFTlWjE1ZSR1mkk3Ec0KYV2czWozQ9PoRQuPwZN62
GwNUtKrSToQpO+qVzkd5Ht6looSC456+MIOpobMRILfQGk8ty7paMCbiuF4bfJ/m68MGlzc7397w
H/q5uk6/WwpyKzGYUZ4My6sPyCZwzv/+OaKS/iR+maFXOCcwBF6shk5tUWKmYRUHeCTQ6KzfIZjJ
02dTPnX0nCnMNApZpkskBo8TA5e4OUi2raEoY90o2KwteasKIz7x2WfuqfPsV/OxRyfHKgzhEDqA
+5dvpJz7Vbi3iVbobTIu97evEERiKEEdgkllD+axGF0qP1xS0gHh8CSBdmn8y7tbRjcVw7Ox7LNC
cNg90/Wvf2BOpupO7BwtKfoTbVyEayUW/u6L05FmcwMa8bplqOXXoLFwgd6rYh5oGmpypJZAB2QB
Z5LSdCuTD5c8zag83whGjMFeUWE9fIZpyxo5J22DqgPAiNNpdfc3FKRQCLVLeScHMQy0osbVL6XT
ztBaXqAYlTPymzXxQsHGJBVOFeInn8Oeqkkr94n9DA/NwXrgOveGJJJAblFzf9YY0HZ41N0cqePW
ElvbX0nB5CVEhC4BdhjOPX2rFe9HPGbGrKyIVVFkUzfZHZRBFhgksnhcUyghN0ePwX5aUHOF+82N
YRGdsmbNRQiIFUDGDOGfqflFNFFoVeiEYi355LB0N6ljV35lwA97Jqy9N6nNkecScotPsdc67paG
imjw+M1t5Oq5+SXUvosPd/aq86oMFyn5cgHiSgdBKVnvqrM4004bGujM+eGGI6MW4F7RLMsNhKzh
x89P0pMwodXyCtWt5hOew8xStPgLk4fthNkT2HHxgbpnRrQh6Dki7d/lBpvfJj3Mb6nSEIQnEjRi
t1+PwxdHmBjekw2KFlVj1u5FyfpuJ8G6pRhKyMwF+zRO1+9ofdB9GpD2Ne/XOWfphalM/CiiXQnr
F6+b6IKOG69LERCRiB4ezV7o1QjwQUdGHNRGy8iHhUB8Hc9gtNTmHzeFswg6IXswczCFIXmkPYnY
AypdVvxtc/gvpWp62fH+IMfGPfCYnFtbDK0Ipq5+vQsSzgA1VCn8MRvdwd7ZJPQ+kngGSArb+EPA
v+1pz6fjIuxGHTcrS5Btou1Ns/zAVrLs1okgk2hbufy3bLtRwI1BARjsCKIlqWvoI4lNEErTN2MY
O9TNaS8xhFIbecfQLXt1mIPQmmTB+bBYz+zflxE1mqsB688yCQi6NVrheGW77udPlNThhyw2DwPi
O3Ui2O8epRfzsG/SKpim5CyqrPx9LrXw2zn57SR3ztxpoj205nORPR3LbLfFSEjg24m9iJ1Ylj/l
M9DSMFUjL02wYBfO+Sb0jZSnVPWQc7C0oOqKuk2K3WXuMiMPB5km6oh3WHYFLL654fQphrh6tKgc
KmFCJzPfn37INOX5ULYxHNkXd4/ETJR/0IysMCKk9bky8leN4+xbtnO//Y4D5yA7h8ZbU6LJUpuT
NBqVs2ZYJ6MjY+dCUu4rbyVoN9mW/FsHmfH9+pHUWSX8NGkyjzKtc7FEClUAtc/3UCsbh/VIinDb
HLi6t1RhOH4+R//3tpHgHq0xFGJOK851DlM34ZyNvz4WlVl11AZwCU/+1x5vO/1o6ySjiUAUF9CC
nOnW9ujRaauoLsUixmpFAsPJGobRP9n7SNvumHZB8HCX5ZYzH9hwUy09DjyVCsvyAvVyJaWukHLL
LLw44DWHO7Tj19K2zA1DvE3M1kU5R9Ml7D/94lnyTPKiTXChbo0Cj3q3nKzwqSrge3155k6TqHFr
v4FZIBZyyxUZXPd2IE/+s1oCSWjHFIFpUHHDfkczIB1dWACH4WmGszTUm7KvymymIxiH7ESuihYP
9I05PWYWp47W4mbHbJ1wtphclanprVhGujunRhZKof28ZlFp0WtCyi+ZrCpizmJGzAhH8J6Xw7OB
iFDbPQIJbgoexuXGnvsYUnjArT87b6N+/PY5jIPdTt7CAYVhfXnxEzr5+S4Z0HKK03Er6nTodu7Z
yjZKsGZZvm6lMj9JzKZfjy1DtrEebnowZb2Pppx76q6HkdUuU5x3b4skWoe75RngX6YsUZKxPRNQ
Arsp5svki/wVEtDDT/JolajGXV97uvqaVG9TQ2zEf5yxYSlKN3Y+sNNnrnKrnKeG8SuKN7S2RyZ4
XSgiRPBNBf97SAPE1TEJop0s2IkMnwPsQbYqRs0KH2VZ58y3TgDIn7OF4enkeqhi9k6fz8tn/e9y
Q80OkyeUNrxRRxVJpo9N/V28xIm9Ur7zkqumfrUTJ+iNJgPY4Epk1TzO3nsJkQEDu6qp0YvM72Gl
Mb5cFR5KaU8oFyfU3PCCgMYM7gU/mwlpSvK0D4vDkFb28s1ZyLTfiFmwZ2YoN2jLFsOsSO6rPx1K
03lHtYGHgl3ryeSkDekM47EHAvGNGT6uYJRB/mkrzG50uAJypXJqV4LjRq0fMGcZX05L78f5BcU6
UgYy38FSuyrZHXqEhhLmmS+SRz4Pn4YTWEy/9Q9bItRwBCHqtWdkmvWHag0jw7E7Vt1VOIjCdnjK
Z6+fzxJvkfM6eqCr+JrP1SZt0phGEPsKT7OC6br+DL5bZXGxCne41qcX2noRW0TBLwOhEqt4LwJi
36VwkfJUwCN/UMtrJKf/F9TnY0WEcT1maI+jWjnImSNy/B2/pDixBl3LkolfjXESCK6gWTyPCZMC
yGsIloBDu85zKZFnzDT7Svgqi43gUrzBiNpVJwYCn6K5+4urlDfk89be94mJbjmTqAAJ4uzuyS0y
KEtyFP6PnEuJlzvdywhsf186U/dn2Ps270O0BV2KhHBDcrtjYNAK+HWSxa8RemCaGhdJksdPcyrE
iAXwniHUZrwj7yfT+ydZT9RNRn6aKHYhgNXT7flHFoCdtScZUpl2yL6Bjnxa3sqMSgecfr/vtaPQ
rT65ytVKZAa/9UqQmFqcEiyWO8U6uVCJeIv5UMicnjzhYOzYcxj5OOe3jnoNcaB5XRTjhaS8fGL9
pPKhV9+7nRq9aacWUFRh8C9cQXx6bPFXSjUQ5ewB0aNBn7pUsmLM1sEtkZd9UVpBLmtWMObI3U+f
cVpV5vh7WueU6L14DHQfscydwlazsdN5B1ujjQpxAeWi+yxfiYcrdqvLP3I+4slnJvukH1wTbXfR
a9dYLD8bOS8mEgwaUn/WMZofetE5v0YRjjBsoaeIOlsFY5G+952mC3dUODHZ2XNjw5Um75AD60PI
nts/IV3Cg4gJqMPPw2EeqSyI2r/3SgovDCJBo+lTMkJUqr98Utj0RXQrSnMyP4uW9p4yDKn7UzNo
WvHUHHq6UwiJst0ue9rt/319z2N2idR4bap29m2/w8Q8FEnw2lbNUmNel2f2UQgB6N/wQOUwn4SA
6TEcZ/Q+cqEAIcaBu3+0UF4z+6tTTulDaBQirOJQfcJ3FIwhbw69Mc0bOT3yAgGwvg9b6hp++26v
kUYK/9NK5gl7CLg4In488cL0ngOEoD3I9ADzcp9jUeXiqFFjMDYhTU5Z2O1ueZvIlq7lze9IkFNO
KySDACSQAlHqF87dKZOk91grNsWIwDOjcaZ1NJy7NXANWEFAfrt9TYzIBGRS9BvuEneIX6F/h7AG
GlOtpAPOqg5NxinMnXvNcqIHV7bn+aaDG5NDLIvAlquvzEm744Cm4rIqgvWwjd5ps3L//ihoHE/f
Zn3yTAfTJbTZ4Fbxv5cHYuXaI89tQxkFQ5DlmIWNeAKlWGSWW/r9Jw3fe6+1Gr8C+wcnP9A3aV4T
7721FcbFSv/EF+1FJoZqw8+K9tDi8R0IESkq1jU53FigKzRbLLVetF1kVsgFEWb1rU2hw3rESYwi
rCZ6HUcYA13r8kjFK6Wx4ZOfrJNX7SrOGEK10hZJzm5q86D8OE7XFfSUONCO4yKKwd+nLWLesfjW
Ax1a0zVdptagpjxUvZgwRIr2zYpxOpBTckMSi1AGoADCa8IabzF9FYygIMTIIgEQTrC7r4W4Avev
6CmeJRwZumnF4im5XUrwuOL1BTF9kOhVHocCGCayhFTIrggBbFnadsOucLQEbRaqG9EThrlDSvPy
HSwEixV2GJamizvPu0kdz/yz5SgLGgvRIObOYGA9vxaO4hI/+DHGuJL65B7mJbdKnv8Avwcreodi
4EIJdOCK+FfdQS3m0VxNuRBXAcZeMlshwgei/zKfieUxIBJic0rTRxlNH/FCrJ89zZD/MywWWuoc
iPUobF+OSfyG9IIMlyR1ktmOjNhLIUHg06ziE85lQ646pMogerZheNff+BUa7/twSxBDbvap8LTE
6HF3dG3HQeU8YSPgCbO8ojBOAeJaza8oQRNFdmcHgMhBUDZ8NR9h3JvsVPjSfc03ZCFhnQ88Qk3v
R2jbUZj+BjRo1vjxgtBPWm9DpEpbe0ojFnnIPhQdTFVrA6RpOO/iSA9rqjIqVfpDOwcZdjae1WvH
wpnFH3knBEfOnSUX6Up6Cegqikmh/TBaNpCOUBiuJaFc0EMYZ0xIGk7BAJ8LczqRDhH5BzjNc2kn
dw+13s5KRVAwweffOt1xvQSgmgrzFQLahynxAfYWUeSzFwS5vDg/d+HZZJzq2QfrjIdJ6xmJbeeO
0EdPoX8/LatK66dHEUgj5jiydOMfE57wvFvdpl79o0l3C2kAxbLSrwZU+RvZZLIQfThOMWb6SkC0
iBbuczJoX288/bA/dS6PrLNOwZBOoqHgDwB7xqhAu5/DitBQj4YpNRG0E+8xvlNMGf0eX6PbQbCN
Bab0qILBUjrixFffkfmrBpkgUCpwsfyHjAyRMDgNSa4HR6oVSpjZNL61EE2qTgOGoqdvKmQMAriO
KYDxJwsyjOdL0upmTbrv41K/k+DE5Q2bpJlYgY1CBUVp9r7fmYJtIKfIHKoS4J2/+Y6BOeTX+Mr1
ZoJUNptSLBJ3vMOvIy0iM8lnsAPkM8XpjP3nsMrUKdW/USJ9FiIi6znKuS5LGE1Y9BiwVa2WBi3t
tHtNCz4ToohOtsrWF3zq/E3kTpj2+g+fcREG7bJ8XDIAKNk2IkjtlCBn1R9d8RgjGV0IcsGfH4L8
l4g6TSfdgcZns7hwc0WtQV7BrCdwff+d8pS+eMlOL9FrevA6xgv5hcHVIVoJfDhg1Mm4HQ7dve2V
HWdM39BQlJXhy7ANAEPrZI/z+vvJmj62dWEi/jhQedqf+UhoT7HAuXBIJefEkZD6U71rudCvinm4
pa/GrEZ1WAlbsqryGx+AG7Yel3QMTimB5MaSNaF1E0RapnOuUTY8kZXrMM/CSH6sAhBkGOcGHcBa
JI+wF4ZPRWtCGwTBG/wX/TX7ZxaH0BD4fbzEA+sd928gwfHtWBHlCeuAxZEyTZYDPND6mijuHWLd
97G1rFBI0XgNe79bkOI5y46jwBbwtTpi1ns8WSDthxASCjbfOrIwqAw78Cj4DWD39/kcWXHfKR2u
UjCAzLEnD+LoJSNZSE5TTEXti77N8YqcSkHga+XtZwas/FHMQyDnfghEzp9fZi2dJOfTqJwgQQWB
/TLlaS5114UP2+j6pFNuJGXwqZEMGiqS6IorSdEBXj93kZ9EQ7CQPap9BU5ErNvo+XaBOrrfRHML
Ql3qFBrUdyP3M12lTJPPRVF1pgmd/0mrSq/QA/tk34yWqC1K9Bmcv/tP1ijbkWT6Scq0Wm+hbOHS
nn0BysE9efNkxGZ6Fq9ncZ9djdvWH5VIIAoTHzwBSvTiLG6NELG/vWZChxeBA8spOBzmqTASfeMC
SgcaPLEL8CK0zR7Z9juaLHuy7HkwP43qimCuUgoNFLJHgtVi+Rl+EuxJ5oh5d28EZ9TkVwmUZA6M
fnE/u/D+Swp+6wkO8RTeowVUWL/HVMXe6yPx/Zdt5Ga1MNpDu0N33z9+ut08upa6fG+t9R8Kh7Wp
eTYNm+PoQksbhaE9s+pEqSKJmT79DERNHiHU3mg0HQVaCOWSkYezWUT1X0YFb+IMvJWTfwWj9CTs
Gto3VyAmRpIDzKPznzHvHfMXWVANLvDsvjvUzsnJ55BCPQBaErLuOSzdI4xLR//rSxzcOYS+b22G
pu8gsJQLULkVQwe4pbkpUIhPyn5cdAnoxlKQRyWHgur98hXeidDwLw6TE4p8leJ9uL/o4EEN7CGs
xlnwqBSV6tVRTy9R613Iv6vmncgdTovvUXISl/b2MZmAdghV0FaVHylzm4meD7Y2L+rRG2xveRce
xTy+Xllb6Go0J8IooN2mVQXIJws6P50VAxU0teHEnFQXNtQAu7Gm83mEav8654RH10JofCcZ6/LH
JCVXKEW7OVoRSIzJWrrtBEGEWjErDJGFhcdOvN3dP2oJk0RjQB9onBIZq4UIK7ByCC/uTG98yl/N
ZYDYkHpLeGOQoZFOmh/Gi/obgEifiYSkxbHnT/1Ig4RsEhoBYQkHFz9lrRmL1N9gMOl8CGJqgCB/
K6Dg//V3i2fi8dVhbcrpIBUI6wqqcEyJKjYIiuZR+Bp8J16Ji6ZV+714mHbIZgWKbj8iUBkRPnfu
MQblFp0DYvIEKdYkq7hfBVAZhtTUe9yvIt8xO3D88BJPkErB/Cr5+PFJTHzQWRYGtVlRQzxxZPv/
m9GwZCm1PWjE2Pu+lFnVfV9nPgLakB4hPDTT7tsRHcOlGTdSwAaJnIbHhV/7ZtOp8rf+Rc3LiC/n
hd/rX39Oo+yr+jdE0mMMTNEEbBNNd35GeYF4f+v3RUDnFS9Tds7P8ko5yG84TXgG7PJ2M8HU70Zf
lJ35ktVp4hFl4U3OiYvytU99aZ+gcj0VmmOgAKQh7Buqjyo6qWVjyCev5s5IJIzQgWff3ZtLw2yV
7ejxsRkdvJZko42OnWirLTl8xtb4RWzFHYGgtZLwtC1AnkbmM245c6ZR54kQViDl76RtcgLCqgLK
E5+wAlT5D5dGPm1AKMu33+IhuKICi6DsZkqCp+ta7wHV4Hky2tbn/6ZS7OEuiRjeEUOYko4UDYAL
xle0bfRJa3TAfwWoei8uHqwzXIUyYRJqtKQfEzIR9/DBx2GjlX7HCipgEiCTqH06R4ftImW3NDaI
i78mBXFgL1VWyytwj5HcxCnH/aA5rzg1anUD+Pomu9s9j6y7A5Y1EyPJ1Mv/iRHbrjDJs6SUHQpc
GssFYNYQeKWNPWh8bRVouzQpHI1HC+mw6Rn6woB6ThmylBMy7gt09gE3dJyccCZxh9cvrR/HrBoL
5bZs6Mc7XNMMss+BW67e5Hau4y2f3GTCOrj9z3jFIS52flxFf+5TNjGNngzyap8ParB7tFJHKjQp
OQ5TEEUKIYgbu06Ur11grVGJZAwr83Ecys8MOe886lFbNF41GQnk3unmDvEbTQPfbt2DR7sCqXVu
qVFBNPrqsJFjH6UoQ1Haq7XVSlkL/WtEorLGOiIWWHd5eiUvvXB58sGFfPFgLUsjn1UXf/7irq0Z
KDnR7HyGH18OGYwT2R+CWfRxQWs3Pvk2KDgx6jG9CJlWxD1XcCOjfQK7EDYh0BABsBjBTgo75GD/
BOiPKossj1/esv+OJOqiqw9lY025CaDu6Hv6zETEpDX16l9yy0GiaPp1jOqIQDVE+BNK9zLK+Wc/
PZEtcHORAZ0TIMYpdSxv88UBbLE0AqnO21J4Eann5JNKCC8S0rez4dJrdRNeEWToMnIS55yp0SGN
/HZPEoQi/W1k65gp1NLAuFIqJm9eZkZgMcZ3s59UoQ0Y1qq8lIjdM+KFkZnOwwG4UcddrgK4r0VS
xJqKk1ZYg9u9kdAeIMavJO2HgHBdd5e4fpl3RhXmFHpURiXgq13kihwdmVKyjD0hBTsCvTZ10w7y
QRinZxYwNDhysyvxWnqLsQxspzsNtScjd1FODijWUe1MhXA7XrO1FqBbqvdMv0HKEp9+1BxqmfJJ
fMHWfzE8iRGaJSNtmKlCW+uBNV3+V9nKe6dnoGYzJoz1oKHyOgIDBgYWKYaw9PBbuIh9M6GRD3Qf
iPOkHi69Lp+kQkMNHKCKffHmKVe71i0NEv5qoGVqTdFBQ4YYhYQ07QWK6TqGEyTYdWf9kerKzmXW
SWazYWhCipLq/afxeAMgRqnCU7LDUs0+5tIYzJUJg95yE9kKl/nv9t005WMxCsdS01Aa5l36PU0C
pFMMdt3UQpNNT2BIAPxpg6jA+J38FzQJ2pa6nR94zP4T132VnTbRg3hdBv/rYsIXwJAD7h7R7ofO
372prE/X+EKdg3TgZXD6DKJa5Ynlag5usmoFtNrdddV3RSiNP8lfxeodfnV9tGjZx/egCCRqnxp9
dkJFjfk9bcPhT3iwEdCrhhXA5vb4eSbHuDK3wlaNCPPLBMldplxUsNLOla9PeNJOIbHrsdD2PkIP
xt4+yM37+atvfEd/Ve44JDtFvLydymJXdFBnAHuN5WRroh/kUHkRjsBbuQ32GA7qDzWOEwT7bvf3
HrnMUX6xtJM8NHNusUyFJhj7LVYrBaGTlfD2OTzgjXmKvVEKA9nkcr04ZI/j5nLo+B7hWKZlTDD3
m4fpuipvS75vARgCZtsROoaKHlmL/smS2DwcpWsJkjL1PygQWwmdvP78Fs4A2Pg2Y+ePlV1Rv8e+
Ro/ZiEy4b0aU4R1krpdysHJP+A0u7yHaBoj9msOrOsXoQ+wFOM2dMDeCqiYnttgwQzi4qhshxJk7
0X9JDC7zMARY8jZThNildejj1vPWsCZcbQVOvd+llbitQw+O1G22lKpFPgefX7PYZnOWw9lOpjTr
G60meX/T0kE0xwbUu20xIHKzGns7R8o0gjid8Xa/5LIUSDbRISr4Qj+edOIW8wu/bkEXoUDo1Bh6
ZbQEaWS7+lIMFpOBFwkqjHGcFUzRD2P219q2X54Xt232gfohFCUGKSUciYFVZAvxD8jpiGnPfScc
WK/gR/de7qgPL8+PjYvLpmMrd1t9uGOIXcB2jjsyWTH0vfBDlxxoIYe/QKg56Mb/oPyeJojR5lHd
ILd/mk2r+EMZIprFAjrxP/3Lgr9/QBeIQJhkbdbVPi53hsIDncdOWXFchbbmVo7lT596HPSgLznl
jI1Z66j1qy14TDR/FEPp7wrg1WvNkfbRnl3019xceciisj86Er78HQwpoxVr5ymRav4bsNim6zZV
i7KdkIbEgynB4nKYNoLyY3pl8EWHqscjbsjaonHW4iI3NwqOL1S94jm6kDGW7+9LZvcIxzWpTugL
iQQh9ia6sCzZ2CX0omKDBbg5QrepJOAXAGxxee2If0w6pNbfZY09nWUmwHES2Ltg5Pb2ro9G0J6d
BJ5AjKlei7puMMQ2KzBph7rCNGZyE6vg9lOAIZgZ8/PBDWjE7jISU6o/tIKChDoah/nrzi8aS3rh
LMCaj3S/CEkIEl6F2UxJVWLqccgBJJJ6o8+jSbd2XlMjgBeFLi6zyUI6y9mnBFrSVrvDhnRHxYEK
S2wyWKccBBjHqEyAPcCGWMcBxTqqX2hrXi5DIWyTMP+FgM5BK5cuM2FHDmNfg+qA9jci2SWaMnhL
BcEZCyYPrrQvpUot/SRcfKX6voAXhT2Yp6HYNy3LMqLcqCT0WLj8ZZEZqs5P1PywHr8adASLLk8P
X0veDeyVVLSweBMlAuODIdGgJ37V5qPi20oqKeAYxIBogyuOjzJKIWuGgEFTrT9mhTpM6pgDzP1I
q/31qQ3ctqmg+jeiOPWJOzTmfbHTeOmb5LF5TNMXheugpCgpPE1uwjH2zVHhAfsmkPz0RIHM2L7D
I+PziM5efl114auLcx2xImK70+XSTHCVUJWS5EKd91FmIADotSbEhBKe11TC915MEJ0Wet+ns8rH
0kdRFpY0RGFS/lC+vGxbSdXJOT/h5pzTh+nZaz/L2CahUfuX2h6Kkl20ESTUpCrKIw5VhYnJO0xn
0sEK8TSeBJ9AyxDEubbQdhObkx8m581Ilpk0l+e0wz3BfycDxy8e9oJ7dkMY4Ia+U3Wzxhcu9D1d
W+aqwmc2irufeEI61lSX+bVDl/pJERVGHnLwPLcS6QpD/6oRykkk7zVUSZBprTiTh/39MvO61Hja
Z6hHqSJCl8WRtOR9Wlx+6SzVUW+ZOOBuoOonwWw0gmoLaNuhePFsQSDth/DObX+yrpa9MiXG9XEX
1c2pc8edbdHcYzad5d/IIQo4hoqpn1Pg7QmF1lqAzqAnjI65/7z4aG1nnBQ0RmreXrfvq3dUk4YR
qCpZ9wgrddkIzya9WOKNhVaisAErBpCy5UlTFVRr4Q3cclElHMILiTWxu+mS7mYtloQNlkz0knba
7HciVwX1DHH793a1nDBk4uLyf6iV0e/nDGaER1ebcmhf34htOSALy/+xViVScTzEJkfxE96gy1O1
E3FZpDAvLABoFN9wNTiJ1nCp6tUhtj4V4Y1PH6m7k9AnaRrVsWl63LFsWg/GfhcujNwP5muHPIRq
1nOjv5weN0D0b7665HCEvNVnVEZ3aFDQ1/WIfaoSAGMhKEY6N4gpx4qez1I3wbbkrkWZODHcv5ao
Vcy/OP8YD75xdrbs2jNIo6PftE4DGTz+oXUmiGLVW1aFoWWpdoJU2oweMsj5+5MqP0qYeN05dJF5
NQIr4CziZN4jyAQEEkzjuhoPNQW12Ct9xHUVAwcmywnNt3brjFYIE+OJtktlxMNASocTw/G+5HF8
7GGpdargvN/n0tRfo+qUEFAa/k/YRqiONFORnhGAB4DGRNbBwfkXCQxXQea6wrZy8GGVKxzgcKsR
WBMLUtJgLilq6ClwFRz9ms3E73yIGW1DSy8K2m+Nfz2Iz0cgTAICqM7Q6yw/zGJmiQl/D2k8f07g
IF93SLVB8QQdFD/DFz6uW1b9Z0Rs2+FiSpEDY7WgUdoZcBsw1CQnaaUKERD4toeTcC1a6HgRiK5Z
qSD+kSnP3OIvsz6QrjSLhaISaIMjF9tiusIw5jGBGfSdKcZLxbBZPdSNBX/IX44bHFiSolK4TgDO
NsXzZ5j7TbFiFkN2TjpIiFkhs/xim1ZQABMmT7YEKRPJRKWukLMwdGuyYVCxLxSwpSVcslBZej9N
9rWRuGZv9gEw0peJalnYY/tX3GXvBtvkb6zakgAicwLhUhxZjfLMsjSank2Rl4CIejDv95Y6oAd3
GM0oe1kVIw9ffuIK1ovFEk/GBjJIakv0y/7qlasvdSPD3ykQalJxwt04UEZzXKsLAk290EDXETKj
k+8vkKa7e2Z1mARQGgrf2mJihdZ4ok5nlZJe4F+nly3KBgdvcR+DwtAbMlQ8TtfYF9jJpmejAlbn
t+3Vp1XYZvsbtQYSIZ4oARMMtXvpsgZ65XX+8v+lzfZhSmzlEdiBbWy5z6Ps2ueRf1qaVn/vRZbR
unjN/AJNskXhuijBolbukvdBZGBvgTpwkqNEcE6Mom1zDAndLVcny4V0AZJPJSc319i7eI/iyvNk
bpwfrQpZ7Uyv9VRkrxZ728+AlwhkWi8GWCB8+38A+JxcEEePeMqqk/kBu/j0VdmgtrXIsoqeg6IN
JIUDnScqypxDpd/hnap/CYCoLKbooVcg86Nuy0W/OuKxApfqJVqaqc1xo5cVHCI5uNMzGzXxafMN
AdDHIpLbmF9CzGxL6CN6WwdBnx31ZbEgAGDDIIngwJxk/ufe5WkHpHtoLOfDMQkj1HC6mxEvIEN8
6sY0M4kapFxg2sP2h5r9iGR8Hdn32VhUx0q6aMm1HOrWtlJYX/Pi12ise2+4f1gPuhW+we7+fUfh
fkvlbG3CS6XmUyySIEALaZ2Rr4acG7VDGda6AGkX+6h3yfRdAUibB3hhFst29QJc+ebaz130E95d
tINvZKnAtCqkTn9w2fbYqyHhqs0Q+FpNycNfEt6VLP2bwGt0SGFQzPvXt71NNK1ZfA7CvsS5GrPj
CRMHGmfjsLXfO4xfQ45H2juQHf94no4e8Bst/srPYA/9mdCnklCj+ImjVBZg7LARQKYRWW0j2ANA
M6WCWOTNx4x0FvoYHZtKE/K+sh9psR/7wBanyYMeC5+3b482sZXE+EY10Z2J7U2n1AJPMsbpqK1R
S+ofZooINbfqP8kTP0EsUdv7Xv/KwYdz3yeJvmBGoF/iyx8qKmWDn5yD6AzPsWmF4N2Vm9l+xkpb
lPUGuEKKUjYY0eXUPWyZY8a/pzEyXYNidqwh8Zyib/boCOA3pC+pxx4i1P3S+EJpNqmvwQ8iYwFC
VOozh3BSyHcmxn8kzdGknWu8u7zqChYkfx4c1XxPG25Nk0RKWrn3Hw7n/WnzLRh9XdY9qm7JXu5c
qGE/8FvNso7LHEBCC4nC3DSmtslDXPsfFg5GqYtNVbpf1Tum9LI0rpyt8YNOXXSO0ZRHUCZKap/t
4w23Cb8bWfAAMVEUiBryklFyPrEWDo1FD0M610We+iKa98akqTVPYjz6OZwwQWI1rC2F+yCUJ5uG
2gL1xATqBfjJDllqk6qtrebprg6YqyMGX5kq5PiwCO0bdaeZoPxz5TL46YUhtcLlpaGKVQkfsVeN
rCdHofAlRx/B6VI1I1hgyDEKiHB0p2gjVjTXKV0uT+otwy+FrremnNeNEjFya/1ekUdMu1FOg1er
JBsZULFxB9EmYvseKjKihAQyld4sOX2PI2WDlISORmRE5uGp7QL1efgsSbhDrsgE98uDhB1nZWZV
x9tp7DWwXpPWmMl7RQmg7ign56yr/Ep6kF+fGGJTXcwrO5xY9vPOlN7chvehpJ3SoweKvJJ0ZaFy
NbRZYiISaKK5vSz6r5D3WuEMjHrw2djENcrMur6cDMQPXWMtxXm8BKGJLEHjw3X0ez3L13GiwUNv
GUTUrKPDqwEdZoq9RwyAwmXKR42WHQdnhtjFj+9Fw1iKuPKUd45Gt+ExCDao9da8GKlqbvYzaJnW
GrB6uJ1RzrsIMk4pxMA8LocwHPWFHrGxdi57ZJVXu1zqrmlBN62hyBWzTGEJGovJdRNCoS1I28Sr
BOIcsvs3rEXNVz83JrGSfK1dJF9foLGGEYEtlli6Pz8+OfQH2hhS4IdcyNG40amKtY38lpM5U4ji
pFQJr6jqocCj7PX9X2d+oGVUrJ8znO5EXO43O79oIC/kq1NT6oLvtoq9UF/gKFvoe1P7ZodYIaXS
vR/sEpCSYl2ltpgka8D+Ua5LhBHxX1CX/ySEkVmnr0XP9RXjSIV53aRuq4PC8up/7zHszOJKOmyl
ioUJPgGr9GrhfNNkLym2DFguzK+D89gwKiX6uDATe2gln/e7AGwvLcs9PyBRpQywpocb7Ql8fA66
0n5aQhnS5zHTj4hRtYfAhV7thHgscumpolQGtV3WMBcxrQj0mvoz/KC2ymI2LJVgcyekDHLlIUOq
/Lmg8D78uppI308FZvWWRIDjszpGUZGq4p6CEZ90UZQX5ZfRyC+PDz53beerLY+zGHyV5LePgXIM
+KlSwWQXhbtedajs11oMVVAGu+PPEy8tvyHqBeuTSi6xirgPFEUNsPtq69r3hGd+UUDQeCrDKCkc
IhjSJ55ChRZRAIpo/oTMj390TmNUqhociiLkfYxFMEyE30+ixkt3HLUB40MX0gjalViDLpwY/wrD
Y2qyhhkWfKW0268KtMJF7Y1m049Yt0T67HWgmSk+LrwUG3kPZKGWg8EQprzaCSvKmYdoAj3xMWBR
OFER4jit+wHC7H+SIHgwiakYBDmyDeydpeMksPWT7toQLcy6MrX7TTSSF/l0FR6zzN9P9HpWef3n
RryAX3e0sMz1klLBAujKNxM1UoWOE2qx0T8V6tVvlDt4aov8m9hTTHIxWUWLI/3FLs6H0/S9kyFt
fYIF/OVsZPpeqn/ZxDVRO8ZXMv9uMBT1ONcesHrcyaaUuKbttkBbSqepn4w/NC+5KX/8PIDGQP/V
g7sJ2mjurrgP9ddYWj2wSYsDj3J8x7mzQD6XrCd3VlgWEs0B4n7DIxpgrB94KWVePzsA39oFni3b
YU13yMHCR+jczGCtWNUGJVyXCUCB+3Msn+FRodOhciqF9+zTtxyn6X1ds/lWtkTeIYQ+RvxG+2PI
kskKIsfj7PB6h2QxlIsxYKiIOtYB6zGm8YG4ko6lDXrta4XNULTZLDlTwkqs0RxvBpgDcIx1Vj94
5XYIwx5uXe1SXX3kXarDcohfOTwHeMeOYGChJsKqN9EV+pPsVo3irbi6nE1oqNnT1VBAq4vY6AX4
DFP8AwW6gPri5s4msmwrNeMnQYZiAL5m4fU6Rfjy3xGcryEHMOaLYZ5wJy8A0tNNvH8DoGEnjI+o
RT377ReA9/3GcfuT0H8y5krP9DeJUrYX8WtxfhDcrXXYB5pXescXYlxSKYn5cUWpJI/jLXglcHMU
wuEBF4SAdYU2tAsGrB428yxhASCsdO1D14CDi3czCzV9Aik/qmi6jJRXRs949ELa2ylK3I9UgEeM
f+b6NXbkKEsN6qcbz5+OV0XIz0VLuWTN8OPxEqm7OeHid1BCitL47iumzUGn5eZ0X0Lz3TDtToY5
F+x8z8TeALM1JvXV1Wpa9w+BogPy/IXQXb64ZCgBWQp+qsX6v2iKKUtI33Ptdk9EWRfOvOYDzxnY
LUdUgo3sRTxoY5rEziktb2Sw9yC/laRvgrh4JZvZCfS/Gl48U55fC8M34LEVOu+jmh8eIvH0oMUN
uORWPZq6jN+LFTwrRW4QzO7ww9yqhg8L1obvuRVhPrTVcODDo4Ry85veGrBOWq4o86D3QPlACyNH
jr9jwQge8LFkjnU3qq0lsNj+QL81cMnlhdcK/7cm9v2rF++2eQ15mQ4xMBwHDl34Oazy+Z4Fln+C
EHJaJemCMR55X1LQZYqkiEWsz6Caa/HgIfY+wQUAWbjsIAuScyP59HH/QEpd7D+cRvnYKtgtbI4i
wcsJKM8l8eufLlzmhs0XIgBRu7cPd7tC3+t3HakCLH5UUZfiKZ4L4is6Ekg5/TFL/LxFt187L4dh
eXJ9PrbSwrXikDCg4ikkAKtSxfKKGjk29FANfveyKWwC+nn15i2vqgsp0j2OcF5Szig8BLPq8wrW
DlPoy/2o6AzoCLN8eIegNEZMAmX/XB09fH1xo86plGqGf+qW5HlmjqecQRvovLGcX05ayx1ho618
1xp5vSrXOtCQKAIPgj8vGCHXeSCJ6UUYhyjW1D9kVPXIvgWu2/ssZhcP2JM9TvarR3qx4BjvRZjt
ZoIglKabLRUhEMCHz30iDVI2iW4oi1BFe36egacbJWyUiSKl00MxGR6ILvrM+WpOSHvrCVsBOtDW
IAvMB0MAPzb/ZNipfbmQuObIt58oYQ9EbwB0zt+U6qPW34YYUkEgg9g1C4xizjqTUwIqvy1+i/zs
8rPD1JjmNbuybwxxP9Yx5OdnelBK5kILdS5PY+9U1JdKRbxO2Ylx9i5d/uQQmE47EYrBWkyC6OhE
97gUVSykVb6iBI8FH5DA2s8vBFNk4vT9jhls3TtB2ZKTrp2pXtwvWEA19UGEyCl0VQg14WJqO8+3
ZPS5LIrWYsIbtjQIScfmgyrvepYYh5rC9Vv8pmrS07qhTHy5eh7Dmv4AZc0zkyYTKRHU0H6jbjFh
B0R1QOb9xiXdEfB4a/lqfuDz68UmOBC9F3XLmdidqjHyJCapuM+qEz5EJu2ChjodscXOm59IS4cS
SUJFNVv11NtLH/jkhzGaCv3pPtKLN4aik44cXNpxWYRGqr2b0yb176LuYR85nLzIdWfUdUTf0zjv
qROqgBTsY4JJCmubcvBLDX4Vkzw/pNQ5P49WqanLor+gC0fLJifQWZGgNEEH9po46OXwe2GskoQj
5ZXlIKXDWm/GGHmeBQeeUnDlYag5RxWFe7JFGc8BKpFuITvqvCDIG5uZLQyiRWwTaPy0iifTbpIo
CWF/oHmuytoc5uHR9CF+QUKHRGJxw4l3lbBL6rgT+x/RO4cjHewkKkJMO6v7avsnyTfXkzeUEtaH
AndxRSx+cm2fs7CNJu2MMLBU2UDqLmKEyJcvxD38txECA77iwgs6Z9z+YhjQE7fMEvDGdk4lgTE4
SKhVXBNyotqUklj/DmNJnDZTHNdvZNpTCic9TFT/uqjxsn7tsUy5UStFTt2q9ngvac1UcDr5YHMx
bETXjsBah4s9vW/PnP9h+tByCwNAyP1HCYn/ot7Lo83EAgLLAR3FBqD/qlr9fjrAp8p49FYqaWYF
vPaF+N5PJnja9RvISa3i51OHXx41Qu93A0bbR5zJWU1KwBp+806+bYa6yqeMIiwAAEb3bQfR4bwa
9SuXUsuXc4lSYa+1O2BzPi9N5dOSHAgzNMwnNd1vNwfsIX2h4+SnQOxZ708CC/HqW85gMhNslbF/
ABpbVvZau/46dEyHOVsPpnvSJIZ4nMBGEmXF2zWD3IhIvCNn2rYUJA0rWg5TJjNJUUPPk5519KJX
3sD5cYHZ8TfPyAA7mVw7PbbG+UD99NmovYbGOidCGICiGGnfH0SWsKXL9XXTjgYq2I3GHpi6reOc
VwoO6B8Gu+CSRnJJfc0JIFyDskNh+Q65eEIr/Yc/KibcevjsMRMfo/Y1saOyRoxZMPxxDOGbg59D
Khdo9BAa+Sls2vZX41krBqQFKfrrP+wpC9fJrPW/8MEE3YfjgsMxFkcUFdgS5m9UyRSno2WbryNN
J2fGX5Y7cwPxAkrPkpoIO5jRftjBH1ShsUZtDs5193FGmkhjfLrHJggf/jObhqSMoACc9ZoxFnzk
LWHQtFJIaMKJstRsPsvp6B4u3aikuf2uzh3wKrNDOKAv5g8JRfmyDuwb07Ow89y6qtXIMMrXOjqv
rE0AbQ8ZWQojnprUmxXauS+v0UTm9yr+DfKItPf9WwNfTHdZN+5ZtEjNmpZZLzhkdxr51HIdf73t
yMKLVF3mmJP1O1JgMtWOSyPkPfYpVOc9cS+qHGAB9+QvM4bvHSvJsmRrwIpytJnL6tfBSF5F7c9m
Ra+6XFph1n8WAEKAcsLLK3CDxtQqbTXAR3V2s6sS2sCEPsLSCEVeql/yFxMzBp+DD5LYi/RxPbkb
4U+/DD3x8i6lYDAQG2vr4brwS3CcNXH4t4SdzsIwk0vcEihhDfqZ5gijJHfjFhGMdkbVVLHdnnMj
7wEXmL9RZzMyuf78JnxTqFMDIlLaMzLjCSrNrA+auuzFXEnVl70KJRj/eRDRpL6EdD8xvQ4/+NCN
THpX4a55sRQr/FHzm2emR3ZufK8/Hj0OP6GjBNWad2TnwMrglEQKPTSsNHZrtjdi5yq4NWs4EwRW
cv77Dq5ylKljZeaaoq8hkW04REKkeE+V0rKOJx8nYrgBMcWAT5FnLQdoGKF2gwxLV553fMAvlbgI
qNLYlFTlRkZyJ8K/8NXGC0Qjv5TrrChPO4ll3bdJzB74VTLsR/MrwZNTfUrm+XwYqcP0/ZWg6hdz
Ogn0PD27Jvyy0W6LBl1e8m3gfoBkAiVG93JRSxX0MdGDuSprQ9jttnmxIuHP4jzxHMPODJ2yOm77
XAerXOoZXIEcm0tlXokpJyVxKNPougwijRQMNsAOGpiylwaEwi4rKkvasm1QT4wCBbSXMY3pLX6U
zDGBkraE4UtlhY4i/mhPd8QEQNaLCvWazF6spAVNubbWBFfRVexkfvbY5TfLWyKgJuurD9NNXuld
yUmjS2iWLFr5juhhJ5TepDyG+K1de5ljDigmOPqBmFLHn2ejyvrovyOUJdFJ3nkUvppbhGkovs3I
vBEsczETsPUPDAbSnwKNbflhV/nknT60OpIqj2IEPWCyVC5cgcriHP86qb6ivMZyvy+Wub4NtMYg
e3MEAHKO7RqHI6LwyZ18nRQOoe54nwtlblRRYhhj6y+IvoFVvMdKaGU//3LGe/9nH1HOdPhPhzWd
0yDItxOKCGwSAH0Vqv8KrogmMJ2Z32BSriexUqHG19NId/xH1eJJGOWtiMHST0iBdg9WksBSy41S
LDdD3DDkC6ZXkT4zWvfPgMguHOT3xdPL+B/hRnGWl+qh+4itBi97ZUnssFRc1vuqNInQiCT8dbys
wPNkWKU/+z2y7TV57qq8izK2bPtMCPIzhGQGnNBvDF8qDFd+Zxlae5gwXZk9yuYGMtmhBI25jY82
1dtXEyIsUFE3RyK+GgYYIH5/DcURzUt6WYOXAbK0+Sjgdfw5nRlk7RtXpgNpNuwsnQBm7uM8PSeI
GdUqoWvJZ/c6/LClL/cwVfj22my5N3/Lb2vU1aomjR/PdSP4oUkByTRenGjzibtHzbT58bonPpLV
E3nYBXNTCM9mjofOyoGMi2EME0EHZl5dR+CsV89e6WaEOs6a+H3TCXYnVCramBnKQxhz9Y549jXu
oOX4IkUM11R/fYs7NZD2mFCjfBnilurYNT9/sQFrhGqordw1HAgaEKtsLQUiw8XjmM2dvQrYe5Hq
3qxiia0yiy60c0CzBDSzocxbxmQ7SzZzRh2qziAreeTO4AKI4pTmftqS4cw7g8vA/EpRbwl+Qs38
IFAacCdGWb/2mqxghrZMgNFHKVEs8jFsrprOUJ5LXAgU6K5bjFUQKqj2PPDUgpn+W9bl/LHfrfBI
hYddwRw4eBp7cVR5UeHwZC+w7hRV+WWiPEllIIklzmOOnbeZHMc/PrO6ZjZXaCPviQ2VgIPH47pH
7dAPlqgZFJGioLsIgHXJ5FIMTg5S7Cgov2QDQQsSHQwGPm00a/8yfCKXGO168UUeMjzZTiEDB60O
rxLbcKr/rtQ5Hd0/pdb3zpSyc/bxkmdwYfsQ3kibssXLZ+7VSmJ867V2CSOjLfPS5QaWirQeMeIH
r071DcdFXS0C2pWQjraoDDX7oXOkxZrXJmUF7h77fkFMmN9q5FdjB98EpzFdaXMV82ilq38euRI3
f30SWj4cZgICR21eqo62JBOx/lzgQafEsCxk5wvOSs+clQu5DeP+RzioqrBXKWk3qUkDaBJG2UxI
5WwpcGk9xVyUbSxIayw1AjULBjcB4tZRH7G37TPL2rw7TleHz0dB8hGJXLmHssV3JkpiD55wFGjd
FRv42lq/PwjZzaaviBERjafp4vOEvpfYjYvrrZAPBU0ZXfK3+z8zeYhFvH0wmbQz6XpP3wCmuJwo
1Blntv2gacLLJ56zXxE6Mrpjk0EIUcM21nS6kyxb+Vm6Wo/NI//CO/inW9uSOxVAD7g17zpWk5C3
drOv0QfRECItNLnTYipvQ4on4VEvfCk7SbdIO0c3Rgu9BWTK0IXk4wz0ddSNpphVvRVnPciNAOWw
srWgx043Odj16zOcScIxDlIpGFaDWuGWNDk99fzX88jW1RhOVYdUVLcx65vn5xmccRqXOvWOp5Yl
HxZb4NbKXB0o5fVa2/PaQ1Rik1xD5XB49z+Qb0OvOD7Y5mz1E2bP/4eav6DfF9mnw65BNcBzPNX0
Xmz7QJiFir1fw1OJxgP/d1crfiLuPhgcI+7+TNslQPu2ktISl1XTMxoI1cUVEV9a1qOe1WKblKPB
wbSCUrozGXiEGMqyimELBnhIshSWRoXYTYaQkhzD2+mgbBl3cRw1uyU7ppfJjHFOr65Ex8xas7P5
AaJpOnFjFd3C7tOqiAPZumZrCc7JBAmFFG0xSL7W2etBtVzBNOGjy9jx0z5qGw52ZXf7P2H9ibwZ
tB/aap/jY/hjKS4cvtwEXiRedMLA01keXJ20sqw58Pg2DBmbVCMuRSmZ6azCp5C9HdLCJFI1VzVL
ODgUDv5D5IQ9zTdYOvMK+7kWXg5SkwI4kTWKgKpbk5TEWAEyaoCjsiADbjLHExhwbXxvtfWBsfvF
J32980gVvDnRehUzxHJPk3POm4cZ2V6L73Eky3YFeoTrUSf1dSiOPdeh48AhrDOYT+G4Y6nwevQZ
Lm/lC2e2GNcnnwLbJdIr4Lvz4m0adYF55mL6PV8nvhF5yG2E9SSN30+IIfW+52lvZhtG7AZWL1kN
wMgY6LVrV0aNgQNrdFGs6xrpI2tlvOFas17hHo1V7HxMhqq/3uYuSJgcxYoJ3w3bQT3jCvXBdV7M
8FJpujM3hknJggg6nBoscXz3Opdlq6kW7HdY4uALqNsU/MrYSI4mbVK3tAjy1jdfmZt96vQOySAG
w4oYtrtR09vXsZ3V70g7V5ArJbsxVa9oiyOjN6Jda5NOXXxectM9cpFNkABDihlAJppJLcUJSRph
t/rJ0FJbTpXX0Pra0oXw7QIGwpl9I51AxlH0uM7o2gm43lFetoMQK4UQeKouoAxTws+u1FNubljE
4zFxh7fBbJ1XHH/eH8DcRDcx3b3y5U73X9/or8zxKYtPBG+lAoOY2C8ud6v1ELSMZRobcX3DZjEg
lMNls/62Xxudwkbf1CBL6EPdQqYdz1wLIJvhdHqEhc4cOwaZdMziToGaQZvnUzdDfWxMyVPaE2Jt
xXKB+SvpghSjL4ZrdQNfHo/vTpczD7j2D1wESm/oFbMnrIsGZLCzNKyvn5Z0p8GXgHn+xCBN9mod
OFOa/SgqiSQty6dESng0naTPUAItXLERA7SBd3UaZhBrCXq3wp/0YdfAY23yblRE0BoQLM0Zlfad
EehIZIV0cM75VvoxB35V+EZM0dsP+c6QY4vwUURJZeORnFJjZrkLoQbaBZ7fJFCalH+hYSwh/ybA
UHdEkmMuUVjw/DP7LLWA5lqPcbYyFooQ3V4dxoLeYG/0nBKmJV3Q6AlONey5b0enMcApBWzytpIN
1bENk7zWGPRfZqmVW27SoBvzwNUqicPHdZgbAk61qZbij8QUc9oZcrVhsZQq87A1H6DHqCzvnXp8
EBd+NQRh9rOWSeINqqfXjen9oUydiWHHXqfGFrJqwsVFNJ0yX9Rb/1RO5FMhFECUgzyZRC4t7Xeg
PDclzLIF2w0BfPozj662rACaQ7D5eYE7rynDQY+W5WggBFvxY/PuFzYAG8+BAA7W2FQJKr5Hce0g
N2l9SbBLZfW05gtT3r3j7AUMl+WTRIzcM6h0xi8AZcXs+Z7eMLBVcJs0q6M3S1S1LTUCUmEpqVpw
34qD+zHjeJCRSk0WngZr0/nrrcs21epYtepXLH/HXs1jufWqdiF8ZI53VS7z0xqkDHNBsRwQ3IOC
qiSHOZGP6AIhSAWy70L20GRWvcy9kWykVRdVU5/0kgMBQS77tzqmuNrOhbfw9q1yyjqx5gU8JVC4
XT9GoHb0WYn42Qe/LHKwWYBLRWPh2yvimAKqHQWgbqb4btRs5DhLtND3CDnq7dyG04SgyzO2GZxK
BXt1f4uN4yXLmietYDWVqFlDqvSj4nO0UfqUylmwUD2spp2T9FCjaKkI6zMX9MPL/p6hivcBUj+f
QyYaUlqGGDfDW8si+Ce7KkDiW9dpqc7qvXTx0plSZIYyYQphnmoocOpcTU9hMf+JLE+GWKvn14ai
MFVslYDBZkPz/2qpHo6G+bcba/3BK8mpD37gs9sQZ+kge2MBT7VvgiA1YOlIFvBTn6aLK0RMs1my
8SnRuJiA88+HyeTIAY5/pQvGMN3nleNgAA38MRNDXaXQHtLcYmGGJYtq4utnxB8kVN9jV/YmdJ9W
ONS1JfQADbV7wG3vQtpldEwvfb5a/m0Run/iSuPA8lsKzg/1m4AlrhJV/QN16/UjnXmsejtSoMo4
qFly4TAj63Ra0Ov5VbMF/YO7Yp4xC0aX1HdmHUp17d8lKsGokPWBFZlzODpIhP5TWUMc1dlxQ7KC
lrDRPF+3eisAf8MYrjbJWVlEOkz+rvBo+MwRTGnLGhK9v4B72PGj/scMnf4Vbt7Z4BQTRdSROLDK
uBr1RkHdDPW31Z5VqKAGKtZAbhjA30jnuudIHFldBWc2tVotY6wUkKAADTrCYyxJ5MqjauypQIaG
TjAP+43BjfOSqJwrfF05uw9EEhEph7tvwOJRpH2bcAv1XoD/wz7C1qlwl+cL31UzOFdcSutDdZkK
TD+SwqhJHoVgqvRZsBqigJBjqIhq/0noKxzqXyN22Z1/ahY/vbuK3cQ0ehsaBZl6/jLBQMB8pr74
K3L0FVoMq03FFYkB6+9GUqPB8CnGAxXOk31d7HhmEAg34QBw34xeVZ1cvbj/cL5cgFrqqPPIlqPT
DXZ3JK9qeCsYErm1Bz2vp2unyFSiyPPF9u8I/1biaHgnBiHg0SZ+fP1KSGOPxYdbkJtH9oLTd5h4
mirMvSV8I3ezqlC+o4u0EopL6Q6XvBpW+gvNjFtaB46Mz6GyCUluxBBb25CHkcrX8b+Fn2GNn1q7
TVZoIDQB5yTcBTE//xFPQ309fgoGmkgahQQmSIrdUEikyoWPkggq37Gf25fUtCVSkO7gdlPCMLdF
+py0CoPqSI4rbz387uF+7icCagi7/x/9MK+IoPGxSb21O4eJ3wsUbut4L1j1d3v0r9qp+naECNZC
PH+tPN+cxfrIbQUiHSFhWoGmsWGxmHTG2/XfOE6PAEebybWUHVRYPn1gHQheIM372NCbOaE/EtH9
uQcy+5J/U2KtzpHVRJzPIOF0vlqflOCsOo4mE/C/RjjyN0e/lcTZm6xWOpjawXVGP/fNxmVScUIa
Ua5rr51tppJ08R9Vfhyzaeo0CsJGOKKfjVUS9sbQVfxJzwrgxwlga9ia7bZ6l3t6+QN5yyXBvjvK
GMtibD9d16+y47sSQ5Xf6noAi/l3i6XxMtgNBdLXzzJ/PqWfcq8ZVcH6C8AAEJK8jm6x1B13dr2y
MfPaR1SHIFAJe1Vvboh4pIbXgMK5Cmx+JwwIbmfk8CxGcwINCPT4wnl9X+Nves+bMVBVGWnicwEL
YchM5u4iOUB+TmSMwja0RQ9ky9TwDQmOb5IRjDdUnVFro1DHe+fLuGM2TBVkjIrJtHayux1Ng8OK
emG60myVQM/rAIgpjTizwhHKcgqXLMwPtjiKyDXR6xpGtG+v/wHcoKVSwZOXw/TpH7LrORWxBFtO
F1kF5/XegdQIVP7VmL0SKI3dc+XperisA1yBSSBOajeiB52I8M/SsNVlmzZHT10ZQVbQuWJ6P92p
NAL6IUv7pMbEtbU3lA7srxRAN+kwdy8kY3i1UvUATmVYbhxmqHGpcBLcvUhRAQtJ8GR3Jd7hGUKR
zuzSzLAj8HV6CiwZth5ujCzLx/FowWfihUrokg8E/ONT2uoSkixGYoois4wYu6GhOb4c2a6uaKgb
ca/w/w4LY9Ffm/9dWBMHxvYMoRL8keBVmp/AOfTJ13tUPSa1c6bI7kSSyovcsan8BMrdk9SI/YhZ
s6s+WzV9GUIqvTxEUXuErChu7fHJU0Eqdn0x2f6bu6l2aVrj5SQI2ahTidP0b2JysD7eztSpsLAg
ZGizijkPzgaqNGGRCC2eV7XJUqo/kK2gZzx9i0lPSjw8hk0ZlmyTelI36CYhBIYEVhNA96ujXtqW
Q9bULjTyrfZdBoZ0vadUt50vW90XsSHd7OSKaR6rrJ5cv4DBrz207+limPsQhAiZVuqKM2i/bquG
pYjEr3h2ioc/rDKHBE+q+nyPDENcU9wPmsc2cBRmwpBqQRCWD4MC7vh3NMp63PVHCRY6sUZ3Ztlt
MEwCC5BTtE1Ao7qJLz690JxYLA6sSuTl5476eB4aczum4IOJlq2Ffx4Z8QEUGTiiqjXEYzf/a+uI
hmXpviNIZFZ9cMuH6+Yocgi8R142M7LMT4Zex7XKbec3T3IT+/+eF2BLx3AtaN0ajEA94DXBsQVk
z5vdj9jx0gSd3Cfz6Rgrf2pC4S7pw/k50U5bD9wNERXoyjT6Vm6u5K60hY98LgYAP3N1wUtT0KHt
0LNxURkLwH+zdBsQiV9orxU6gR0td3F3dnOoBZCkkJSlMEHpnXpk3UfST9yg7JM3qLveFg1teR7/
l24Gixp0h9+zYoWBzT1GPKdA3fIdDH8hyQz2nLYNrFbdJWw7prlVBYZUFFExXq0XjqQLkKEsRIYe
wg66NyvizuN+FtORme2WcwHCOvYWGczArZ6ZpJdebvyfDCvSE+8oATJ4I4kZLtEBaA5Ct32DK0xU
GIGZXIAH/DoIz70UB9zjCZWqzxh5FJaihs54kJSBoahu6JyXmTQj6OZ1b9GKeX+ujQ/A0deYaURZ
OrDmbjVe31FeUSJeomzkXwPMXaxr0UNQA2wdtbmfSS4Do6lYpQSVV4p2W6EXS270EuYr15lsU4QI
jXZ83jipojwlL1CQoSvxZ8GADLPc+Yug15HK9KJAQWscB+ITRfqvCqSB0sO8OdIqh3MrOMvaPp/X
ajGX3Iq2qFWvyvaauO48lkBtpA6eqq3bHiZ6aFtZeY5+uypzYkMxza2ooYkF6EN3JMbsXufK6Sqm
eUI4r/zAoIQzqYDGqKMwbolgKRxDpCc8hZpSUmOHWLMp5Q6d+4sS8Jnf6z2APRw8oPM1gSSIO3ZK
iybOOUZ84mWG0j/himoAQOnNukI/oQB5zfzWDs0YjJSEBYfOxkus3Gro75GXtorq2CpWLYuLGVCc
zIy3bFFWvYyBCJUqYzqRX0gp5rAfnEDblf9KW+yegaA5d/uqH3Gg4AO+IseYJsJkRBf+4yhd3WWO
BA1OQiQ80n7Wz+bDYPiJSwiggyNdcWsxZdV5aa35VaxzDAq83a+Y9fzrXlIiRJC8KEAZLPnKApl7
Wih1/0jhl85d7osRBLN1VJZBSjxPmezLFiRfsQOxTVYGG7ILdVtXK3HrIkqZCyFWiab4siZd4qjn
emQKEIFuNpB02o++iIwwmR1IaNWy9mrVb9XGZiBv5fCtshqBUXO8omPn+bwWUw7j1Gk4I4tI1HQ3
XmNG9bELnD3zsSGCsx/Z8DY/tBa/gRv2Y7OCB0Av0ZakCQvU1A1Pk6A3vWOj5jYXOk3m8pNUOabm
umZ9HKqYI07lx3p3upvppAA9U8mjzAwB+DhY7K5jc6eMc7VA667c22JgndUJaNQP2RsIKDfjVjbi
FUEaLSQrOqHuUi4uV97gpHPlGSy2dtzxS+fAINL+flMLACxIE2KL+jCKPzH/4vCpzTfJ5ae4NiO7
3nlyVQIj9gOP1wZ9m9V1Lwv2He2ZNT8hcc93NcgLoIctisRQdIorCgJK7xvvyuHUBiMMTfsca9+J
I03kQ3KszfyT1hu3RW4bP434cay4FECnfUQqEqtN2MoB3vSKGLYaHDZP+TvtWklyM2XbH1qYYYnb
iwL45Kirz0txyXxLZT8HHZ5QKrgIGE27xdl16VI7dsZNFKEnr3qVDoyES6v4GsXBilQN775HHXC+
+x/hy/QIQHxRJoSyryXS//ZdO/xyPTI7OXM0ckYBZoSYkvWv3OwNcNmJG3MuBUpcafALVH1AY1KD
FuLYqdY/8TqvUYnpVU3qeonIm5Wl1XbMAvq8GwAiATOaMsKLjFTrjIGnVqOSnEMicc/nBkIln+23
T/7I2FmQvDqouKQBxggP9SDSE64kkbVbWThExMcUTFTioajy+WhiRmvXNV8n1aX6J8DD9cqPbtoG
btC8mGxFtXaDIhpxY2yVeGUObB7QZvuZ0p8P5/XAjOz0OEgmB9pnv/4wTezbcXMwPkP1BQsDlXTU
+SuTZerf5LkLwPxXpoj7njemCONJwiklVIkBD1jyUxj56f9vifC7vOGiT42ah/6O4cJ/q7K4rBzB
CUyAdhawZIeC4jd4g+AKPV6UWZH3LkrzaDpA1uo+l2pCk+7CYk4L252OXWDkAQhz2VMMvOmlO/Ak
3uK7SFqTBUPG1+hBfVB6Gypsxxq7c8yjBk3HrDBHAOMrTCxIfOtk+d2XXxbN4hkJFg1uS3UybCYz
wxXibGDKaWtxQ61GYbQ9Ha8Dl3p/7XF4KfriAp2NGNesGZuF+bbVwzo1bLIO2lhOttvnOFSxrTCk
oUnIfo8oaAgGEB8NZxJYwe4LzAbjc8QbfvlQ78ky3BRVNJ/UXRgSQFCwfaHWfsrlRqGSPZMkly36
OHAUelbUKGNrK4v2c5eq4k2v8yH8ahe7G1zK9P8jc6F9eyci7htqlzat/xdKXQ+Vc/PdeI+Ybc7r
ugxozwMv+8eEUkTqFR5CbPXqt12WRRafPNN+PyHe+5Y+Sz9Rkd8/Oi5aum/CEb/ARR/HtRKssIv3
DTEbySgyvxEyl2rGtufGsqNyEgWa7qHD2cuyPWmSxBNNYMGC5eZXw+oqaYbMfEzEzmHS/FZcgxUZ
52peVyzPsnGgJDzR+qupLTYt+bbHEB79xh9ZTcGTemrUXpdyodAqJYWq+cTEBBIgk0hFeW/7ApwU
Z34xMSbHQpDwFLDRA2Fq2hDPAHqb0tctraOf/H21e8As5M7iCRYicjz/EuNrB8a6cQRw25xEffmg
CkKU+rpUsMtDhFg9oujXn48dVuUUSk+Meg8DtgdluC70yDHaMHG8WS8qvgSozv4XVqPlaK9UR0n1
Myf+qkAqE8psNNqTTpaRIlrIxQJ8TZ88v2MAM+8zm/Ck+KcYfJB7ZJB/Z/U9tIwUeLfvbPBA6kAb
78+c7DEgLMgFs8xIajm5KetTlLcdXWSwjhKUJn6V8NnLKYWy1FzFb1NEWWyzz70NsjEmS8Khwu/1
GqWm5rHiK60xcBKYPRmB0jwefS3uCmO0tB2e6vfGcmINQd5wZEKutlYcjS3B/ZErkS6dTjPt3/Yq
V4VrYK39CBA5kF3V/UC0LH5xEgW9i7UxiKar6yzPimLB4jv+CVKKch05czw78s0OimuP0oTQpYh0
wDVDAZ6V9vvuENhur8nPG6oKOCU7boeaZ8bzdX5H/VmY5Iz96nTL2Q3MMsEyiFnKxl0mtAVe99P8
CdO0U/p7XwbjfqsvhJ8bkVjgelzOiO4Po0mc4soXDjh4Q/qDnT25j1n4UYn2c3H7VdDrFhBmdvcY
N0AbO2esercwP6WpY5I2yFKWxMo5IDeBJGapcWpwLH5F5K3g7qk3ABWH4M07jXM9guCHWmZnq+U7
S3macCJcSg5WDMiT11An5ieS9XaKvo+D6d/spSmyOMUWS8TUjVu/Rd/8W60XxznZknSqrPbeu/ms
gCwSuVBbwB+lADHH+LLUsNIwMZ0kNp9j9T0wUyV1X3AVSP7omxuCeaQCgKiAuGK/3dDG+OQg6gQS
P5n6t/+0j/s/r2AntpRxKgaGlrlvW6fb4A7JCUkdzaZoanoM+1C6SFsDAhYpFZBWAKrGe0ZI7cXC
Tx1ty74B1vxs8Vyc/7zpcJwjw7ZFFeFCJuKpNpM+m6zfE8RiVgsrFR4F20i9XTURI/JTx6lkXfa4
/9QVSw+5WXPiw436LYJ0EyO74Dc0eXj+fojiltluDxQyCDVd4zm4ItUTzB71zq6HRE8MpA+BdAjC
mSHHbl5PegVhgavr8tSpY5WjCxtJxDYqmk94x+YJOjWWcNmBQ8P+JeYe5Y9Vcrc6l2rFkiBqvo4e
uQgMvb4fxdhOTG7aBdfKdUb3wHkZSphaZErayB6uft0NZk5223hRkbsx/Lo7B5WLp8SVnEy3CpiJ
b3ZauYnFtOeWIIPMkOJ57uQxHV6fM6BeR5o/3qD0WvxYCFljgO4OCW67IZALttDkiGWKX33zuuok
fl3/U79hI8vXYPQbIm3EjKuj5kYUWGblko+/1zelinNMQkWIJJ2zqoldS00n4qLjOUuiDAzzt00N
ymE0HyruIW3c9rCrg3MMuOs+bZ+lBgLMHwwt+CKHIiMD5zsZsdtPXEcFVIrtGuGbcnBW4BbFcaBh
Z8GNDZdNNJAP5Kcj0hBv7ZAEDtAFgFZzw74sVC/9aOSr6k2hdvLijr1xhOUwKWEvKkWomP11iazN
0sBuvgzlsYh7ha4ZDp7IAqgaostjxb8rOMipmrMizzclEkKfR1tpFR5umDkgDjEvN6XYurx6+Cgc
8ND9MZaRXPodnN/3wwdy5zgGxfZQUEz2xTp/2Ark6/p6gJFwLOz6/yjjK3XIhejvZ441TRl3qMq8
R6DDAP1odiTsmYttLh7dLhvpzgV8JNrB5r2wUD9KAIYEh01NglqfTT6ByEM8Q9hvPm0RyZIRn+Xm
V6qC5Swzg4l9PvcrvBi1bcLwVZOx2O6ncYAU4G6e0n7QX7cR4uvsPt/ikoloHLGbcUIZx0uxiPjh
b7P6Ie5zsvQGQ8AkI1QmC+cYpE8xM3i+WfzIbW5WSOGIu6+a8a3bzEEiocYoMERfyZfpG+W835Dh
/XSsZ82tcFLcCcexVxxi4f4uk5aNFT719Vwk8V6mWUU2jCKao3RslFuX4WXAyxPDcVRatSIKFIZh
UN1q18ZvLBo4InZWxxAqJYjMGDcWi3yC4n9PNAl3h1M7DDK20xYMVMPpOIH1hiN8EBM5qTv1FVEu
5t7ct0/3r85aC2/w8LnHuCxCUPoNtppoBaZhBRNLtxal+OYlUbN+WuIEcAozQp5JHCg5+oHhXTTZ
+ehxej25jAK6IMoGZ13s5QaO24Ug6AhmsFl86/DoYF+O/uyqXIF4XBXUMCrcqL+KnYzN8QbSQsmC
18gyEKkYRZMVBKuH8j6TeiUzfpwbItVSZLOQcidsUggraLIBfsCilTtgVlAVfQR99UW0ajmgGMAA
mXHLDFepE6m0GDNRWNnP/MCNFtn38hPBpvpdmELkkCG6XZcMDYYUBVeGjpNmGqCQ0wYPRzdha20S
BC9csZ/SCr01q2YpRlb3J94tOulduv37wG/qjPoAVmYMh2eu3dc4/z+lqO+MgW+mTQeiBt1Q4p9Z
Qh8xyrfcbI7IwLUoBuRNxxVoWqvtjMELiQr6b7oCq7znFsF5OQgRhUPZGiwbH6Vrm1CYJp9LVuUx
okLjrFaoixELMC3k8Pkuo7t+ZR3nkF+jiHzjNVkP7Y6/fy208A/gK6tO5i7OT4mbfJqCcyOQH93/
iCbwYxEAT2p3QgR3/cD+HpXxVuS6cMiBYep4q4ugtZwg7es3d3d3+3WwvtysgVrzmIjowTbRF+1U
t3o2wxrY87gePq2t1rF18wbRyDCAnzWraY5lwa/ZmE6ZADtSHvCXvvCyZPgfwrReUKwsi9jf8ukA
z41ryHBmW8ycz5OXgyrTcKx8KqrvQOMeLv80yhTiiQQrAmib9ItEKyfIzAIZVhlhqHZUBiZtKzL/
jnlgXQ5M3FpSVWsJtehwQ+CChtXQ0pWbr5Is8kKQQzpI+HriFatIymz84vn076HdW9yX6dtunik0
eEBz31MB45E+UUhDEEj1TvN7sp+kEDAqDvb7a33+2MDrhGrMYOrkXUH8Gp5HeicJ/np10Ng9YQCN
hDhsAp6cysJ0k/FHf0x3dVTge8TA+Uq2JXD8wxF5PPOG1LFAycTtF7Yrc0ztyUQGOyjdr4I+tljL
jgcdkWhba3LOh5kpPx3KXk7wHC/oypPevPWi9+RlSdRG8G0Cl6MpDHOrpAYUyFuMMKjwyryelZh/
ZMYGjsRPqdlRrTDddk1PwN1hV3NYbYAXTIenRiQGcFywlpnSb31MfXz8wtCFIA+LjpAXcNgzFo8R
n4Crohz4MWiyAPVLVUGiRx+/W3379YrbMZ/4HAoM7ivX4PdZjodvQvz8w6FEwB0/citxmEcgqvMy
HTeEcMBdGQbld0Ar/ov2g2o9L+0nuCG6UfmnNxCBHDGnG0tgoqcTFSDfYe01DemnQcsq/ugw21sa
mUvcpxPxym/vJueTIpvhLraUUmvyPGUleWUHsxgbyAy65Xs8CdGaVxOjx8a/vOkj8C6h0zJLJOaz
ZWr/u3HEb1cA+aJ+bHJHvNzOPcIQFeKMZ8e6Bc7RqsfzrT1Amu2yvfbL+VwJynkN5HAfDwOB2/RE
SXSIPZtNtUeaiL5lDvL1+8dNl9D63hZHiqMwDeBU9csDmYPZdHI+Dz/dXs1qt60Q5bqwHuGAwVVM
SwX3xHsMjEdVieE10zX+bEy7BMQE9TFhmasSscw01S5uzVKWy23mRgYm83A41pcSSpxXpUW9PTCo
L0q7ylVJWd13fXBfmR2aLq62DDcg/38stZL9/2tF9roKQkQAPQGlOED8OWYX/9R5Byql1sx5eVpj
uY9yq37WF0+XBu0ex9CDwTItjbRE3eGfIhICp/IWRG+q4IbFzKRdZzj7rXWXMxogJAZZcLho5Oo0
CtjG3l1buQn/DWW2Oxcd62QiNzJK8VMyw14iJVlUjUbdrqYZy5ceTDXySAS/PWIEjFuwyAWdEkYd
1GXUf/qAw4m3sJjmjziL6CcOjrJXZWUEXzMk62P2OuVHruQTc/Kq99PSm//s5CiIfbrQTz9SEfsi
N9AuZnAZdb+2LowWDCVdimiaxR0Texumzwn/vnLMOtJmso/rFH96IBVbTFo1iPNLFyr1TKpuHbZ3
BK7EcEOp5kzHsoTKgLqT8z9oaYcY6rE3nYajryiprImRAbZTT4G48Ryp1NnGOnWFF1aQ9OcafmRi
ys2Ou/KhHTtt3wyay2xsYFeumdgZGx6Bc/lP2kpyEAW6LnSdNJZ+pD/yBDGAzfaHQ6/ZAtZYTka+
9B8k43V5OIfRilp0Fw/t/MKBbVD2waOpVGmeA8EzPdmWHbIYaFbOIksIP1xqUXrpKEUNuqqr65Su
HvieMf4FEVL0zotCwXtgKSgfQP5uN1YUmrd0UAt0f7lTpopyW3vjLmGqjr7TNu6l5QrjjLmsqF2q
xZz1JwWl6zKCH3EjBp5rGslMcqsMUeOkNpmZRIUXUivUVAG3XhNW0cEqLwL8GP0uSDn6dAjlsLKX
FPUEq/ANlxndalJ03NV0TwHTcvB3e9PpiTM0x3KBuVS2N8PzKGuA0WlJdVzG2DB5wVxaz5PzQs0E
7qZsOZj0ZMuXsJZ6BgxZ1a1iygBg+1HNa6AlCG6JZoeSyUagLi1yMVq77d6h1YcKXxdyiiBtbdXA
DY4bqkpOmjYV+KfRILlWVuWtUXyiJx9hQeCzHfzFDHi7hT7XECCFhocyj0jR/bVAjjKnIxrBbdfU
lw9SFPGf20pw729yA3WzYkUuCBCWodUzZPfeczTmUFvDBGwBSLuHgSWQRJi9VUR0GitituJ3fNpx
OVOyEgcoYfdc9PX8H4vQHbLQjqF1e9kppqkXIwZNpWEBxK25ZRcbUIfCejsYmzMPM1BJ5h8wc7xI
dYK61OImNfWT2tle8zlO5QypUJnxuNoBSJF5O2Lo48FeET1hapetBK9hb0IU7ZU3Pp6qvKISqFaG
yEgMTH3SkPX7qN9hsY4EbPHqJ3OsmlX7O2zImQf1oQuHJ/Lgt4dqmYnvkSGGgm/H2bqq2fROYew3
1WCocJE0c5cqnaIOyKlQ1HOxOz6DVQs8qpYk4jefD3c3j/DtXoZ2/5B0yHyi9PN9Ps0XFjznJjv/
twnltkLRSedJuMkShY7xgWHMpXNzaGuz7huRN7GenSG2+bJr0vvX8r6pYSwTNWj6TWKzpAREafPN
NLs6TiJRbuqGvky0qeNc8an4fEpExiaK+FNgsHduSKz1JXdnA/BTIu+DLwQ4V1EmGRYjZigLtlo6
pH+jPlmeyxZCzuqmOcrejN1rrI1TO1Bd0BTzeIy3VkeIFjE1fdseZq+xJeFETjwCNecEdDDrP01y
fcOnI7Ht64NDSRn3bFQCxbXcn9C4cBEAmy28E2jw70iOfr1U5offVstC8XEFunpshbGJkjWawyfj
KXjbT4drlTEwzojuJ2K3fvdDhzt6BQvfNCrN88AcATxOlGW4NP0rR2WC2qCWzTCdyf550Fv1WspE
5h3aCjOo18DgOB2ipX+bVyxh3aDkQ/Vv2edAHaUZBqdBheKNl7mSLaCN7QJVQhscM1GYBfvazbfr
fCRbiZVeYt1tqX87bkAJkNIUpNstTOfGKoY4DESpwma2cHYmIWCHAdUpFusZ8MOt4Ve3ZI2gVK0u
AkM0IlMPQgVaElPS7nfIsUwsUzUqZQr5+SMGZvIYeH5cXxdARjovDPEBvtFxBN74zOPK9FMG5EUa
lC/nCWazdh/79WGEmJM63FPeVcoHWVIC8DutwchEYnTy0ntgKWbgCy7RLFxyGkLWSF9d0M8Hh8JX
9YHte5QJxq/p/evd/95LdHba+8yF3mITBWZ1cW66/2Nv73J9Y88TRYP4xTHbkY8OxGNr+qaUXJ2C
NRjE5RXfMvljGfS//nCDyFhqvePRAR58yl62haam/ZjGidyDsAWlbEo+dTPEsPa3gBN1o7SPU3A/
TKI0MaHUPVPaU7jOx38/ogkcB6TL3tTfdeN5B1d4XJUbdn3fBucC0DxbcI6bOavly7O0Q1s2lM9P
anqa+D0H/Pw7DsNISedtlsx7Lb3Qw1SGDLtsBHUl/TJZ+H9bbRDkQu9FuoFtO0YaDWLrCQUbO5sq
oOyaBqDwfvBA3OJBZ/9p2WCgNBfIL9PflTuanDcGLn4GeTCx76KMAO1aqyCzCQsbNrQ0cq8kNNkx
jhJZAZMC2aph4DJ1JHbGzq3Hb1tS4X231GVhdVoWdKzgejxQE/Hcascx40hoqfHdaNjytibOcPw9
ORbu3EcZM3OIo1hXZ2aNbPXlclVmfzl3biZ7MJx/Bund7NwWmrLDWAsA9bxoUum1TFgrnHeZBjj2
bxBcKo3oe4HkCyLT626Yy8mTyFOybqv+LI79kBeXQ/7WaHK8/3RRCPO5sinGyUZcy8+S5uo3ZZ3m
HlgOXjw2PkW5Z4MJvbIHb/pdJXercJ9S3zw2dlnSdsACht4Af6jDCGjWkNd8usfzjW3E/GW2rwAh
B02wh5it75Pn2+uI1zs1F0Eei6KsW0ISoIMTmDWcHzm/bxQ3/nPS7K8Gdq49UCBgTXBkXbW5EjHE
2xGYzblEJbuX7WkV+CDG8ApNgr0Wlv8R9iXa7QoPwUNmylRlGXZt9dxoWjjbVAspPLJCjU1I0p4W
yZwNDC8CclBWZ53SEfSzVMHA1KnZRZEhkFCRl0TpUHU7RfEb/6aoFseaOjlb0Jk6WXY2tjvcTuxQ
/qUo/ujPssMSLUeiiVHxdBDWg7i/hbl5mWSd5r0+G75lmZlxeIxenZeipzAbbeA0rVMjaY5CFTIs
vR8XvNa8bcpI4UZmaSj5ufZS1YUtngb1rraj4wwh1T+MYbZBtEfEKP6BhphwxUXRlnrx8hJ46QhZ
31wHQZkSouhgi5JtDHMh/tZssKY8xGl1Dn1+osfHcqHyRov/jpN1s/1O3MMLchsZ0BE9NnBsX6Xh
qLBTQCFllN/EvDCTYcm+58DBSBQJOBgWUIeULCMIld3VlJBMVmFwGLKjbThAbNNM0/QVbL5r3CdU
uuM9c337TNi9BhkdG/EWkKJDHPk7vexbslg+FwvoXdG1D2ILz80ynQw3MR7LWqxA4+w+e/M5KHYB
sqsrxG7J6T3mMC/odfw6wyEVplj18p330mqLCjRxBiB7o4aD6Rv3YvH3Dgb7ibiC/QHmRiwoxJf6
RhROCC4fFeMFWdFBZyNggHR6xY4Ntpx/OlClqZ6xv8B2ZI2LZEp+vFR9/fIcb+K4iUw7wYS74AvZ
IxFD6x2fptXrSh4nt5en/qVdx1gcuM4xnbsBPL85YjV6XcLsCMj/UHuvPSurdBBykF8zyYeLWfIp
TmEB/6wiJdbhbh7VHJtcmnmn3tdjgNomlGGN319YXcjXdb0za2VdDiR3SLiiP781vEAMiluvMTNo
OQ992ot+c0KcLc8R8wdmX73K0IgLlI8IUj6s+dGthL0jWKvuBEdsJDNbRYP3PFyjWVeMVgdl0GDV
2IWxwT17xegTGscSG08Ov9gFyD8XloW8uCj4jwPLn80EvVBJqGUK/M4YIEsCJBGs/2IW8X2pyv/O
LGjtoNaN7pmYhFVmttSi2EhunaY/dDEqF1wmCIcQOvcdU7pekvcAmJ3xT9R0cwkN9uWOU+yTB8Bo
0J5ff3VCzfkakpkqVhttqRfMaJdWWnPi9lVztBSsxc7jMH1ORxkA3HnUuc+hi1f/pdz19C7+ekS9
S2qO42W6hgyLeObi2ee6HaITu3t0tAT0WEYehy/A1ImcEiYxAQoYdwJpxGHS1cpG0NaOpGmj7xko
1pUaZZqkMh+gQDgJQzoSmEcSngWieTBowHim1nbZfsOujPcDO8SeFTurd4NIhTnUBtxvFWBtjy7E
GmRo85HMh5SX8OnoWJJPUqsWJ4mZxwP5f2J9Qmihyso7aW0eK6OYESa1viYWCusX/WsTk9EL6b99
LIYmAUIjAtaWKByOu2PGc9dtNhOtl2hjInV/YPTsXuiNiSLBsuKCCHU6xZzo5+ICd9uAhPvwFimg
gxiLXwPXcbVWESqUnPUtJ/DdHugQTAPmQx30q7JIdpv2Qwk1ojpLa1YHHaMZChyIbrEVBpat4Vr4
Q/gWtvRJMYn79F6it9W4+D+xmAcmRwa0adorcXtzPtl/2emFPKln3q4OkUY8Z7nFm/AoN9tMrinM
vTarxxsq8k0JSDqdcQ/+SmpDZCekvMHaBvybV19j5NkZuoqe9SiKmR1ORuWjm75RcENR2rqAVDCG
0MfsCxFcn5yVI4fpIgvsu+9t0WbfstU+bdQEf0xMyb23RYhJnX4oqpgWYhvYCtIlEvJFc109Rwiw
W/Fblt3nVXn6xKy43LCJaMUZBu+kVl/aR9/BW/ampXUgBKiPxVX1zqiW7AVO9JjMcPQxNF2ANbOX
MbKOLXFtRuzRrrCnpC6iAq03UaAb8gknnQjZq0MBiElvAvUeZqsAnt0yLShJP4Y9pJF7uuAxgDl3
+dgg1TOV5D1kom/kfN7z+M36KAt0rC8Qt8qZmALKvJKtCSAmZzi+194G1EU2998tGnThyYBP0KGd
BHLhtMF6nWkY9Sn7vN4ysHSTIVKqZeMmVmdGUxPIqFxb1imz/wcM705J4rx6dIrkhmzNd4iFpV6i
ZXUCh1QXoAbLYBsKjtynZWl4xGNvc3SyYeOBCVx9SwzBBs5UZWwKrxab68X8NY5PsU2OVDNtV6Dn
b/oI6ex/eR5gnGZrYwvmRc3nDduBQTSGZgqFGdbLQloBWo5ud2SYAm1QwP5/qEOOngOsEagtMHXX
7po7Rz5XVyfmgFurDWK5PQqqmoiNVQ3lfVQv4QShVnw3zd1+azHDYjpkTCKw/z4KzYGC84uHwoSy
0TsHJ3WiIvtpx40xEtu03yJT6a8jx3Jat2AWL4ffIGQIGexm3J8wpNSQG+b/es546Qudx815I1O3
7XBMKiUZ9X9U7se11CL6V8EOtieq/G2laN+6xSLhF5qE/WLCi9drt0O2CwUS2zAwJe4M8jtMrkQp
Fts1cTPJfFoh1wPX1jjp1dtbPxrG4sA2TU1fKN+vp7i8/bsjn0YRxVpCRDX/WGkcwJ7ICfFW1lHW
tEKCioZAkyHXFzi2Tm67V6E9zuVSwhIvNM1DjSft93t/XjNZojnOvnZFdhWJI4agta++SJ1hmxCc
iK0vcyGpCTYb6g0NvCdLLk0bYbirgpey8seC8rWFSQayhRF8XXQ/F1uq5Z3w/CzNotzpigB42qF3
jQ8B+vd+uGeRdTGLwfKil0w5PWmBVcKW1N8fIgH/qgnZl/o0F2cjtARFk6ObkbzitW/4Kf+uK/hl
Isc1HS3SX06k6AOgh8VUWj+uN4GZRGjxdK9hQJXaG5ukB4ZdQ1SnZqGMfbO6yI8eJHnX8odvqIQa
iQX6ltGfsy7W/85FCo1YJtUwAYOHMNVGPJhilDPFBTzr9NG/D6Q15hfOaizIgFnuSv2oUHmDJnPy
dyW9/R++5VPIvBCB6IsIkD0sHQX46hPzah6++3XWO4SECYvxJfKQ2L7B1RCZ8/e00sn1TZdjDKIA
Hs27g0OT+1qG2zebe0t3/Thzkr80xMpAbWpvFAUWi00C8GAXEwgmproW/uNei7XgB8kInnK6dBsD
PMzlVapWmqNWAzm19FLrLR+n9fStV0R4tp/0ISsKAiG19FUmghjj6niUDlECjTyLPBfsUuf2o3Bs
2VyhVziYsNk58qYLuF/4jkrmlHAPpVBjUz93FXEw9u+sYJdBUytuy7YjH0JoKzzoX2ahNFdlQJMQ
adfvfiFl/wwiF9nopPr/Z9d8EvvAHtZYPfmgRwDcceWd3lsN6pfPlKhI6aZ/vhEdHPs6Z0VIqCh1
SwW2o9cq2j9rIbO7QJNNA7Lyf+IvtoUgeDrF+EldBXv5qyDm9s7cogpVVjzx8VVBvRysxsP3Gssu
yIchJWxBHmBAzR430vNjbLk7NBZBv2xY8bvJgn3z1/1IwsR2Ub4qFhVD0Z/Hdc5VlmaAZdpZORZd
SBpsC2CUqDIUJbRfphbmdG7dXRpXRjdGMcvNVdgCM+8RwHQcpVYvkkn6edM5ETh0QBM1mCyGKf1J
24VPXuOvqGAMcImUKriRNrOMLmE4RO+4ndxyVjzC0JNRPhTPogdpAzT4XV8oCSzv+oPC/9MrFFcE
RZzyDH0+vPzG3RSYPcvVcD/YCdigjH2ZWAiTmO2f8znQ3sdowwpI1mSwfd8dF8wqhIaqqvkxP2OP
3VZo3jNI5TYQlIwZCQjsuIL56ZZMkAulWZw6EZ4Yuv9IFUY4fqZoiLIGgzVwT4MDjNbIHq82Rv4U
vmsczGGF9Wv+bUQDNvIf1s8WgJjYloJCMMF3x/yWRdfmgAoQBxU1mS0I6eUTLESmEdY+vZhKSyTp
SX/nvmjRGy9eNPXi8m4iaygqhT8U/C8Vmk3uJ+x0UENfo4DSyGAiXBLasDDx9cw5rx/FJJ66LHgI
7AbqPLr1Vn3IsHusZ8PB8PXeAJgpHMgPeyi8FQx79l2mGqfzyMJy9fs3sBXIHaBrQbWsUdEb/Z6F
s80C/aweCBpEorxVwvhoHB38r3piSP4w5vYI8TwJCML0I8gvu1Dd1GjVuB5HVNfeA9uc0aRaDdzL
U4GcohoQABjhAUstX/puyRW/x/bcSBKIZIRwVxp/BBzAFOsaVw14Md6sqJp7X03a3zHJKqzWxrQX
+fz7i89M3xBLLJ04SSBbb1p5EUU+lt8Wi+1AKJxvvZ7rB5MtPtEUCqMtgh8YrRfbtthoYkOtKCQU
uHkjavM91vYjhOQGWc6YofJ684T2j0i+h5XweknWDWpBxkT0nZFwmB/ZS5OMwByHqq8mk9zGDOry
m979AbD0DN7dJp0u5wxkwFQwxSvJsAfjSas0uQVyoCsgs3EJf2TnhR3srBJNv2uuOTSkTgAFkCY0
MBFLBFQowTPGseftlEAbFA5pG9o9TbQbjPVMEP+MN62YSutiwaV3xLqE8/5T3gbgvNJvQ3ppu4Ih
KprIuUN5CkIWdeNasW3Sup89sSlDeRq73rnYFwPkDQ5/ULnrd3thPu9y1uMIWEl5L+xEoRLIcP9F
54w1iP3kmIUWjsmPxJwWf/debTCMLcpnxeNmpHAq79GrfwSyicJkdZlWllMPpTTuKaOccdmNrM2s
Ec4mpo5vk2CuouJ9lHtt9ByUh7cZxoxFm/cpyRHfhpqNLu+wvwwrHKK/HSEGZ+RL4uymP43ofadN
fNvu0ELeUrKXivbVSDp8Wn+XQ/xReLBZZl0w50A6yk/0UQ0GYFJ3fn5Nq4dSUJNmw/Nsk3IutXgi
6o7oj/x1LP1uHSSf1YLZLrH7parJuOT1nlj7Utsk4rtHaRZNKGkfdc+kHUWrp2GUcAXNZiU4NYSr
dyuBMOMc5SWgz/fN1PG/EveTzNjeCVSaVUAOsLoSfHsbEUacBwvf82t+fK3s2Lb/W/e46znVKyvT
PreAEq1GVme+PQbDXvM49+rHRslnANKBp4mEV0On6XvLqjHPNLlF8EeXsN9QDinVs+zrwwQqIU+3
0MSy2DPGP+bHKuh+PO5nNX2WUAEW675+tqDge7RVVNtb8Ft4EAY/O4cc3Ey5ovMvpjI8/1GzLQSF
Jo5mvfze1pq52n2ep77cZ7YDn8vG9kY4EXszpS7ouGvn/6bw0hVSVlKpB5TctJk6mw4NCWKRhB4N
kNHvjaWcXUjbCf5AF9k0OPe9FSUrD2qyFn7W6nXO3g/TgunEGJITGQBS/5VVekNMt3Lhd/f5FDZw
3K2P5GdcQ+CBNOPzyZI1XxdCxgG5VkepYl+tYa5FCYeadhbQ/QbIU+/z7MvG3gMPxNrQKzIcrSkT
SQOFZHfyhwxqBLBD3kmJ01i5AKgbaU3+86NePP6GxqsBexhLkJESw4sgdorEA2qwHaFVUrSYZmVz
wsrvN258bF9Rb6ELxE9VLTHe98iMklQDUKblTyaO5hs66HNqXgpqB8d90bdgEmPUqSEuRKGg70C4
sZAEYKXVMJFWY/eBzlEpFdBCN7PLhzNDLr2LwfHUJzlzsQ9MIQGGYNmJaHtYsvugGhZ+9ax2hBJH
O3RzLK8juZawH1v0vneFx2bqUt+uN5xwM/ky/Cl0NuIq7kb7+YCznlS/cdKJW8z7Rryiu3EpDJf4
sXl23TkCWwxkbAcw8qB8AwOpL4fw+DqK8LQKo2vGZicjSZBWreD35UjoqUYb8+KTwTX+KwMp1MBQ
TKmgPPI03mqM3FR8SMD5R3uoK50DuzsE2DvanjokRKeXcssGzfhFqn0FBJl5QEc54axaybL78qVL
D6x521lm3EzrOnwmpZaJnhJxrbDsUoX22aAKUHu7S8l+9cQ3UTa8hk2Akvz/uXsmr+xtXJFd8ft5
CbPbdAXCRpPbORq/zO+9SYAu1wm7zT2iRx7CjuVumOws/n7laVQelIRwg+/yyyprKJqfmEfmQKb/
yCRrX/8CtvL5t6eI2K4B4VoMpIvzHOf00X3cVQE1ra09neKBtg9R2MQpehjCX50hoyrvI0KSFLZ/
aO9gOgA/rmPEmNq9tL6H3f7c1xUtGsfRhiquQ0E3uEjsz1Op++8Wg6rTxabBoBxmqqdTtC3yMBDu
9/gfJbcxKui7u03LT6AkjcZr5R+jTcoecdHSkozUnxAeR6GLKfoBxD/Mp/Cnt+nDOTgcRzoTEbDU
WuO49tpEpa07FlwV2cHGH+hce+8f9PA1s/o/UnPV/NrGow9UsRWOkT8MI00xJsyUZgg70LbpkjGG
2bcm1Cxt/qlHJ7b72F3U26dQHNZHV3NgH+82JDqLlp7QCefuGUptHD3vmoF1csQBYZAIsR0Nr+5U
jnAwDWq8tAaJpRT3pvXrx21Uo+BmDKnRko6pH/lRCJsKA2LT/W1oVm7Cb6W/PETbZBpe252paar4
V7BfceFx0QcrKj2WRb7K9GLOBN8u+QMBKfyx3VoGwd35J+hBJbucLa8Kcl3E2x6eXYEcZnJzXa0L
12oHQQUNP93fZdcfJnvd4BiAAjrReB6Z1vBPF7HYhSlbzTZbW5MEE0ZUZ9jHO+uux0ZrRbENIhDf
zxmNoFhk0wHMa06YG1TkUkeVLcpIP+HreR7JAjurwA+NT2exjwhJmMA8Z/yxDTYruHVLDvJ7jcgb
u/aZK5nAybbcHwAEFY3TDPitRGGsY/G3mGEEuRXep1XW9zrgsuESOLHdKFETKK4nlxKWd4ZS3fqo
nooYQjnnHwd5Y/LKzdsLLrw5qSO7kcdZTd6/quTxWcVUHIYsDtFrBIv02iNG201U74nA197zh03L
68CDidLs4VOCGGItH2QqpRE5bYEWaQu7jt8DvjOi8BgDCaW8RbQJZhHURJfhrHgu35HV1g+JR6qb
Y023zg6GuGf4tjVLtaGoYYMNNNrGgYnyGqHXdBa2R8UYAeuwi/gRH+rTRZ065uthoP/nIt/j1gWP
tQJtk07y+38T6rt0KWlzNRVjjVubj09p/gTrOsWH8rQATQMcF+CrijtJYcTl56UB8XmEvT9q/F3x
zcnISzoTyoXTLsDI/2uUUVdvptUxmke0ISuj8aB1NUROmy0Fmeo6z6e7mG1Lq0wX6KeJSuIQivcf
xW1hc6HsztKGxP2/g1wGivyEpT6N/TDwfAnK2LqHJjdMwOtrFx6G0B9O+gI4IkQYIhZqFcd2i5bE
uud3PZKnKpmRNToSaD51dwaP3Z6SNkLjlKEIv3o771RhPNpfqIDfj/Vo8q9GwZLqivzjSIRiSc/i
plcv3nPIEu+/aLk6v0aXPmqluzx2DCRkUSgc+/OXE4o6lKbmnUPtEBqvFueyKIJhba2cj+D16cQH
zjdJaJzidGkkoPPgWfxAS/3ZOvbmZnOefcvq6S0MazjeUZ9Dzei+s3SX7muk+pK3AqDtjKzUfNgI
kSKfc13LyuKuu+F1dynjqV09giCPDyKOtL8Ju80d3hJv4v/frv0ile3/x6pi0S3wJXM4ZEGMefsJ
JGX5f4bs6BgxkEA8JSQteegIUgAxXLmehYf1K2ZJQ9XYrxwrx9TjahbcVJFlaK95N5dcyjJqzEzW
EC1C4+31P32nPBCxPolxH3WKOb5TsZyn8zM01xTPravmNXNrC1huvT8iR4QSs48+PQny9rmO7JD5
C3fHjL0Plrqh9dkigVTBd066W4zJHjZQQh1pAsRJCde7xGTHzNkerdTFTW5KtbPKCWUyQ54MybMi
h+QF1/y43EsShz2h7aUkzTnXqU9DDwsU0MMJR2oOVvZZa8lw1dJ78Z2VaUmSBty0SmnQ1z3RXLX3
YMjT3jBd7b+s23yAz4TLaufJ8L50/sjGVSiGrBgsv+mlE8DuA5XStklzc/1kR7/K5flR3xHPwrYV
hrETQa+qGsyW7yAJTPZvakBuwSs0RPmXQjEu1XH5wbMF9WzIIk0tmKXcYnraC6wgd0NXiSz/ab/1
alTYWk45Kg1wJkGxeGhRVa25K9hPKHE8HDcUAWoB9WtR1S+y9kc31oU4WEE5yiPH9wcDZTcKB12L
zH6liZS+zkRW96VRmW2KlvOM5zMsWVfBx4SZn7RS8XHVZXuRpgTwiS01AWyhMx2E/mVzkjQv7hH2
6h//Ec4008DbWB4hi8CjiO12P5KCA0RExIYbHeB1zIqK8GJWMYoft4H0/ecIYFJ7lWfV9idm9azD
oG4vDknRudkm0hDv+tyD3z6dbSBpTcFwSqBrQFV4YxG3+q5v+G84yfNVwLbDTcDFpMQmKnbK9s3I
FX+09fCbfylD4LSZBtErge5VKWp1B6j9W9Tswk3uP2LWLjQqzpGJoDZI6lK4nRhnW5az8AGaXOfp
cfjHhN88Dtitv88DtoToyjnuUlkVSYfwZvw2qCcSbf1K35iRSLYL1xgihgeRbtUGLTh5PIdmrLTa
NlCSioQdPS02HzwpDhr5ijojDvTr9AVUKzLmBY1GGSK9R1zGlxrkiRuRTOHTCTPxqvLCxA1iFgJX
OoWJZG5g50h6pLhReveMaQLZSRDF6/gSPAT06KSsCeVKEycqYfCpqqUWu2uORkdFuhbNQCaNI08p
m04FCN99WaYs6Uo7SMR0sVGyYEf5J1xxDQ1OH4uaPDKOMIhZRvpUVuZPADKY3bKIxsSXIDTR58al
wW7qMGJ1KiYHBftRQLv+kYctL/A/LZ56VuwcbQ81sEdABlXJFXQ6BFW3ha7ZnFqlGchoMZSr/yIu
giaeM0unZ2ooh6JeXCGs6/LaRK3mvfjehr3fugZQhZWVr3MWmpzX4oliyfc6HaPyRK0qjRjOiHEj
pWelaawLLdjztGnEN8kuQCwgVRGyMyhXDoN/g0xGh7erbhnSd1jRE4TQlOcJAPobrln9nms+5dgc
63kg4wfbMIEKpcrXBhIDzdYYDsju4qgcP+ja/mfo1af4/PkXnKACnCzolJiPTem5zDvdQdMKgArk
mq5412b0kgXNfiIEtyXDcqLVxIxCG20nJJblYiIY6FP+dsyGjvezvLcsd8SLTqNTk3WQWHCPji7f
sXL4dooXcIkK6N3sJ2VIWA/evHcSNSe6XFx8DFIneCR2If6UREhyeHAPy8MmNBJr8KBfILX6Uuw9
37JuLsk/HCbG9DY2lRcg8sP2uQLI+9iwOPpKiZrBqimhw720kLgQzIYGm9rspsai1f7S05S+9oun
YqxhF99pu7aNAd6qVpZowLMkZ9sa8uiWPfGGVE56X7HlbAgXbDT7NlkHSmskCRwmCrVYQw5Axa8M
rwyxImvQHJB417SYO7r+jH/N3ZbpWhes26WZORrdYDtSBZJSFa5ELgcqgaLWw9zaUunrUx9fYBfa
mNfYrj51J6xq0Zv8CnmKt3wyv6Vz0Y1TInQGKSVn3KhcVy2XTKtuiS0qRQ0PxquduQ8dxjdvb5ku
burNFRPKHlPhyzPCsFDt3szaokYkFXnB5nKpPqYdaMrCOfffWVyddRG+iVdsWz9TOxYneSfvUv9e
y1Q0KtYf8bFjYo7+d+dvkSfnDjWQtTMATclVN2mqHSszXRDlI3esSA0WF3I+uyOObCoYdKuI4eVy
2769WJoQshw6nQaXo7qvg7WMq6zjaDYSXtyIHh7rquo8V1VC2umkWdRgNLC5RDR+HADJpNU2R94w
calfE8MhDKPrk1hcfs1Vd6DEwiy0fq/+xrsyiWDhKucf50CVyCRvLMJFYtcHxZmUTgYHD9edVFON
dNTs57wpqSa9LBWvFUvn9JvST0gYsrhfWQmpO00w24KbkggmHpem8CAnkcLZjpEPzfC6RqF/Xcho
IWeL5DFXLA9UdPGXfNCqNbWF4ofjSu86TMzDpSR+TM60j+Af9MBE+IudyEDRNN4mXwcpQhtiqyBH
wtlqotK9s9zEVWpKFB6VsLcPJuuaXXjLiHZ4f0OfPfEEzVkKKwb9BfLvt2qtBbBXWUKuKXnNNKgn
6itumh3CBKnznJ/efnHRAMoEvBHxO6s81Xn/IHypq0TmfeeI+ACrN9kUYS8pdoWTWB6MfFCd8wfD
y09buUtAotjAgNeWy4OkZ7XGhf2riQSpWKfdx4TobDSBZ4quEoJy04h/uBbayQiKhmayO+AV5ul4
Q3t9PFJk9zNmelPjvnvGv6sNf0dzUb8dSBBpAkcXybkoBmb+z/5vyQvT3XXu1f8mBkq+20aPBs2K
JRPtdT/gs/dy+DFZhCVowG9NrVPywhtC+yosdglze8AMWZm1PhgqVv9KN/c9kkK2S30DrMBdHnPR
W6XSfbqWIx0IMCBHpUb0OWhHLbS7DqYDvjKmTgXy2ywyP9u0SX6ev2vRxi6NX6mEJbnj7qDk14kv
syrRpvFrJhOdaoMG8y3LZqFFKAHRrDdIswfUJCxWRpBhheS1s3GWZzgtG1FTTrIoMbbYZmstsY/L
jjB63znyiQNlgEqQYYhq74sRDWc8/ZLHL3Bp5LIIQfgRxm1gNFS1By7dCOqZLuENBgtsiO0EmTa7
l3VZGkjK+P/Nl1EmG7qUynKmtcW1m5KQnkMWanbwDRokV2Ovh9f5fo8n+dHOhVaJlrFQTvAtTSSn
T4AmpS4IB5s6KCMFXtSUdKJfHZarxl9p9jb6c0hHqsicVXvGHhr2wcsVt6Nwq579rC9d5SrzFQn6
2Plyiwkbn5rUGkBnwLf94SLthv6zm7/oqs8ecwP3VcgYZZLnuvDOdeGZdfGtOLn7N9x6GkM3wv0p
CgmeLHXedsUHMk0QFMPipXDb4DJnIFAmg4SVe1Zf0nrvHEPdQ3nxiGPcTwB2csCVsWvNpGETG+Xl
lLxB7WuXdyh8C1VA1AIXKfJfa/GAIe2ev16f32O9STUwcSwxmxviSZ+YDErP3ec7qZm3ACEhMTGz
AhwzufIU7ZiqwMMJPotjJ/izMOZeTJDb6QWTFKWQjyxfaSeDiQMdJFmbg2RTijTnz2HkgZYypSoH
k9Ln5kpBenHu7i5h2TjcgtsNj33kaK/xhaByTsJtQ/qf0mSSG8JuF/8UxcFUZekVFNWb6MbQn9iN
3vs3UZc9wWLZ4l+M7p99uq92FTZdwWhLS8Luz/v7xHokRRNuGPoUQNkIn25RH5ylrzKO6SFsZm0L
6cQmlHRuBzzuSi1CBzQuGJXWO2NBxp9qWDHoDozSc9LhejWFiY1GUWNwz58fMdaeBs0OyIbtUTe+
AIwrTEqjxkoBXDELSPS3KJPSITMp/iLPSIOaFlZ+fdM6i9zn7jUqQIYkZ6HJwkjLTdJP9Ef68XcI
FG2xYmb5JMC1v9Q8yMcH3cNk84zeSjfhO9MNwOIDgBl9cxIoMoOs4KaJZalmsM4QKHDy3IAIb38J
sGB55aRhs8e9xl5+SzQgYoZJwUrz7HamDs5m7lk1l4sxfbpQLvr1MiNeTXExVZKD41/uCnpvxzAd
+tC5DEg+vFSLNBkRiltSqTEiyFtW2GpmCZZ/YwA4X0EB3M5A9y0lutiVEoZ1iWLb+MKd7KYmSeDt
2QiTxwNTrSMuCLZouMeLKLahHys2YErJgE4HhR/Te/yTF+f4hCKwk+u4HdIZ0QNrK5cq19tbpuNz
ZC+QxvxhgAW7cQIWGijw8qir2w+7bFCwwRLO2Ah9Dm/SPcdho9FDNBmFxOIjOhZQm+0OjPGOJcGO
CJaDzs5JdyQAUlUxuJuPINWHfWVPUBp4DxUegQdlhmgYz7L+0j8W5ad+D82pNRu7EhIojehGqaTB
yQoZT4LC2nG2p2VL8THaLOnE0SrHKS6iJvNvIxK2vc3Gcympr4D4muqBm3HQBV+11c84qFN8G3iB
evGceMPmOGiRkDMKa2KwPz5MvBpe+kaawvdfbhOCmfLVktWBJ4vN2GoCssbH5CcMXp/lW8aoadOT
2AB7jUoiQVxDi5MuViCL8cEAqJSUdF5fJjyOpihRDtdm/iwKB6xrvmHGul4gHmdT6oko+OT7VO2i
7jBiySYoGB5Dr5w2BSWFpQvmZxdArCqqXnfAo1A/haS51sVO98JU6SC/ANwzqHk5XaRFtm8k6WfC
yR+loaouctWeju9Qb4Bgz+5NmHzUfh5Lk6+Jd/HxAYHv87+OGlgXeeCtXpZqbkZwWLJMGjTnwaRo
fMo8aT1bv1FaRvK/wXTdRASyUveMoWmKsqCSd2Z2OU3IyouNT8OjxdfzipaMx/EPZKeNB9+vk3eh
9gokfFpfEv4OUxtMoMEz/F4tZBWi7kAr2gzZajJNUWYpRaIUiPnjfD5L8G8SgUwS7qN/v9ScjTRq
KOMS8MsoB7TalFP7KXQUj94qzyn8/iOclyKQUZv0eu41S8jZ8xeDzW54AjrQofPKGfVOYm7gQyH/
gjkYMdil7WYe1yoRPz5rWSTpumgqj4yPuIEYdw/5YyCo0AZXfonHNR7oODKl+J8lVHHiy9ycWyE6
9rKu1kQyQUUhxlWdM4XtKIyyU4gYuWvlQS718Aq1LYOE1tZuv2vsncRK4zmYKClEkxgXiJjr3ua1
axPChqJrdJy0XfcgDz0KWusqulygBMB/R/W3gU/mCwuzcWeaYymdnGBI8mGNEH0AMqPmu5h4NFZE
OW6qowCqO8VVBocf36szOsRXfLgB/idVsQ4sjPW6e7CvNQTYBajTpVJQkfqbzx+Dn40iphhtXZho
S05Wj6GrdFnlNbohPB3BjGa77DPRHM20dKGrZkPpE1QOxOpAAmxYIYzLt6QH7kFnU3byDG18ziLd
g3omZV4bYCHdr1+pwJVplNbwRT4iHF0gLhT71JnTWocM0dHmGdi/GifJprUGV/jz2oJM575k3cVV
Od7iY1ptQopOn+mafVttsdqlztOvgu3RtIGAMPbk7zQ8hiJ4wxClhVg2Kra9Qk2JysshkmTPW16p
8wAKltwpkgWP4/WGuyBVyxHm9Kb9WMR3NSfLr4Wmq8Dz0Ab1ZZwj2Nm8UD8+t6/uHosP7r2zEpZt
VnbRKcv6mNoMTD4B0z9mb9gqbhjy+PGbMncq46LBxizpKUylfHw97hjGFmm2ZecOhvi01dWiVWwd
96TU53NXsJhxwz6TbGON8ULUjeCHNrimRnuBQZUMLZ2IQFc8OMzzBlK5rkklrij9YZ+hAvtXzfTJ
aIU2uh+pJFkC5RWDbnGD32S/S84PRjkDro09AaGxenGWZgUrPyE4eoHJrZHaS+7sVROAZ8mxH56e
pSzuuYIAp1ina6yQ2UlA5Omzgg2ZV1sGxZuDCHVg0Pb0W7IcXhbbbykXVYBXB6T9pAc3nQPyTW+G
K/F+I9OftIuwyRXTOTY1/LYspQpDMxbp2JatLGYAPpBqyQJBPYzQiiHvGwetLT0D55j9+1yuCWHl
pVagfiF8eiR/OhZz0c1uS4hz9PUxBnAxB6GAfUkwJ783nIKWXHR3wpkIFaWCmU/cLNsVqBOGGrT0
g4XT+ZtnpgUomd/LMYvb5MzbtwkogoBkKf8lI52AE9ugn58e7AhcpR05HSOEW6DQiS6qmo5U02EA
XM9La+avuW+QNjlQgR2qZoCToGeDBSUYWABSP4o1GPmldbNCEL/s8JA6+DJt/YRcgzG1AIRjYXVq
w0EdOyPjMk4ZhBSMNnTNvYImwfyeJvugw1Ee9nXR7ZIqUsft2NyxjnZdDHB8JERadHGdKeugQu6N
fH8Pm0Zjv6LT0vqtAngn6Zm/yrU9JhhsAZ7Vv7CjyDC/2ovQeo3PMnJ8tOG1GkEg0kyT3HsZT+LD
m+61nEzpU/Lmei63q2lnhs0+CgHcS8ukCtjqolhCRzlDi/bFIE4Wit0FVQjP/tTZ6+JOb9LDRq0Y
Y1YNj0uGt2qmccrO+I0Iic49laKs9+g6omMYKvP4ZSP6UP7b61d2Man39YIHRPzNbe43Fy6YoPom
uzFNAUhT9isi45Kw/WQfC7V78CafHD4egc/xbKMNZ1CxCQ8n/YJ7MQVqM4ZAPyfLHtlpIpAc/olE
cxkdYSwRVXHg7gE/MujNjMZSdnj+cylkWz2Tb1JBfEIbBHu0Id1JDdIbCMZddCqJUGz5b1d83PQd
nLqPefCHd9eFnxQGRONZy2TAUxO3pcLtlFoSLkPMc0R8wwjjXCGrItZdb5J4Eu/YZLxZuGKR4rlh
7NyWmPidamQRmLuppNT9Y2CoEfaS1g4/PX91CuboAvrWoQA5XUzlwjEtvN3ml60N3D98cvstDk5C
XqDH0auGxqElcxqcYEbNpmji0qjvwgS5zZ6LJQSiwEY5HHcqRXh+xF4x5t1piKUCPorco6qESoK8
Vc3pcs0Owr/L9CcfL0bbjJc/wTnkT3FNMraSDl1TN2XX06AquufXD+akLeil+8WShvxVqrNoU4X2
O3rkoxC9tBhIjBWOpInvlK+mYUTdXieSy7mDHF33hywWcCGt8zdADCCscss4uhKLVEfQB5OpAoNV
m8oIyRzlbEchMWW4o3M81itD/WlL49AhNAIQNylirDvnr0JxzoEhybzhXES1X/0x8qPN/DRfiVYy
WI16y9DZxwPSVX2+AjjLIlD7RARvLtGEL5x9zyPXQ2jYIhkvC1fqpgV3w9uffnRd13Xc+0ENMCyj
yLs7N5lD1LOhSetNzV1hgVDX5h82BxhLmBUAYa4muNs9GxEXrm22fgwlxJtNgezkIXsJ7C0kjDSz
3Yh2IBNS4Zgt2tOkOSGHobYXVvtP+U2nVQDe3oUTw2ViRtBf3KAbT5ikhZly9UCEstJvlG+Hd+IN
IsBv6dvLtCMGevGWYzRhA8OXaBfQKysF6Ykoo7P82vyC79V3J9NR/0c2ldjG6h2IeCDXnBT68Z4b
hDtzzy5FX7NkMUrSggorMz3S+q3kZy+RYLCXOhPeandm7Ed8RxYLy00wi7L77xBJ8HCDgVzo3czK
o3hpXYfoj7ELDfODUSsRiWeCAiVInF7YPY+siUo2oZ5COqz0IXRcSzymHBtQpNS9G+kdYTN0ekJx
ANFNlAct3OlxNJba2eKDNw41hGcqeQugDqtOaokkgM4wCD33N3OmdelXjObSdZv7FX+lLmsrVSd3
NC0LKl5nO6y3g1dANqVWqLM/f2yCL/PSDHdz6Zd6A1eGDMAIEv6dwVdJUb4saxgjNCVQJhabp/ti
MspnY13KDreC7wm91N2pKIzcOIXvk7DH1Bhxze3+TIxK+xABavBv6Y5Q2Ls7QAn4Dh4Mi46Aa1BJ
TV7Cbv+T0EqEqq561BInEq4IN5bbACS4S4gPpTmOXFF4gT1rj0JtkaI6hAf+ayClj5jF14N7rKQ9
jVX6nnYRsNYAtdTx/5dXLHR+sJGR6/TF/Vq4FWWokDIwCTBEPs/TwOf7ZbKgZtdi/HD41PzESBAC
nixAhm4FusFwv6vevsiy3vRUA0gVXWtovCgWIcDzPSKvQSq6D20EFwB8W2kduyc14I1UiyxnQXl6
DHdLn9jkCjS0fgobKvisA8wrs1itcU9z9te3II5qyvJfdwBOLrfAyzbs2PrI3V2ZB60Z0Sc/3F2K
tZtGJzE8gpCahrR2LIDMmIDXiqUDb3JppksIROv+cjRH4wL1KRDvrBmg6R9ZoATglUYg11eIuWZ0
wBSQwM94fOM9rk3ESwc9vbvLXnw0gKjc791iTRbkHjqXWocI9I9PFQN6c7cFvlnnf+rCzmAPmg7Z
G5F7kVFadcZdEgpDgWED0D8R1uQcixNpRE2j0yL8t5rHxwXyGC5dSmzi50vRzxwq6jsFh/BWlzw8
8Drm0GbCA9mqS6LDApwRzSQjYJa4ycqD8A6i073mzhyxy3zbkPHkdq5XHE55M00k8a34T3KP4BUD
/HedLbwIwEkB0vxmPdtZOhcr0voSTP4m1f6nshA/hUpfkA8gRShifA6w/gBhmKEgT4Q2sun30Y9y
5ZdYTtVpquFzDctNFVr0ORzaN95FivOq6vDbdoMvBcx0wt/PAVy6jilFqsCkU8oD5BArqGwHtHqV
PtcWwPPpk8/SlsKOGnJPZQSwKOwWQ0JzXI5/WJhCibdnLGeqjF74EZePvRQwvDQrMkfyc7JC6Xef
L8TbJ/Ia39Otcqde+BafM9uOUh9JT8FVm0y4GvdbeIbSa3VFqiwF3okkeFVC4eg5WeVRKjG6ssH3
wr577xjfFowQrWTpfCf6qEU4x0hwedCTRbQfD+TnoCqESPjQ3iqBN8I3wT1SS5u2vUa2L/CcJKK9
tJbSSGKfZjOmTi+nlTaq1xvP1iejJ5bPjNp2VRId1c+s6pVu3ioxozREz2WKPmWGykuf18Cox8jB
lCJ1t9IM5j5zrvMUJTtXycFh3H1U6IaEuQbyS7XnMjSlY0QWebK+7xD2S1vbdkdFEK5wXb8xPqYk
u1L9FCNYggXrvUp2JBGYRelcu2A1K31XWky18CQzkdo7sIJqXqY77MLu2PQBhgojdS73wQMAxhSz
2HSjWVVnjUonifE8/2yVxduRdfJObVR5rsZazNtI1PqjdafD87gzGYMBdynf5VP6EVF6TXQ2uJDC
ezwfevq9A7nkrCOCD/wrT07hj31etWewCIDBi93vC3RsRy5OCIOBQX6AcIEYx9AFmKWe/h/KuWbY
wgLUG/kfFaXSIMojnjRrTmMKFdPbikkyFOBrYuRY0vops2W90MvR2ZVtuWYDhPyethqTya7rZosi
/yfEjCt1riWPI9jfeRgojJXPCYn8HkeukJKp/i1JZ6BKtEiNszYRfZDgXS95jPaY9GJ/fxo6sPoo
OQXf+HBHqgCLdiwJbRc8hk8BYVo8c9F6iJlFygQqJI0IcxPaebrP09ErFKsGhb3zZ+BsZJ3OhQgI
JlLkyYN6H2sRIFG8Jpnj4frhBUp9a4sB2W1C36bvOBvdikSXzRz9RkVu0HQDbaD50uBOPtjmYWHN
hrSGKpdZY7VQTGbDKbwg2ijrF2aTu33Pj33VVYtX8sy884ffsTPBJPEQhxoABmWtCZlQp4BdLyaP
B+R6y6s+wpFgGBJkJPtbrFB+T6U2HB98qp2NAc8e0TJ+XTHWmxe4JUAdeiyqQTvbG2Kp/aDw4bmo
wu4Ch07jWa9S9HZS/tH7NhRGEd1ihjpJsAJbotF+YPCU2ImzZVZROwNTJW3Z9lpvMyxuugSGcsRT
2OASFTsIS3V78lMP87s8KdMtr9sx6rtm0XqBZub41jurL8Mr+VqlegNs5uVv5aBAC/H9qdl17Kfz
EwtjLw5+EcBbk9u+OOj3Wxyze9osMGufVMEzqqJmdyAUrmZ9cUBEZpuuVf+G/x3na6p1Pia3xZjD
U8gr4ahY8qLVaCdRP81P2UgxwPPBXY7muJGwNEiRGm5LTJoNk0lwD5YveSaHNAHsyaIbJejqgztJ
TZRtiYvQuNHB4lbGPImeqfW+p6iaYOyT44hpgc6VgJ2X7cELEbnAMPpTEZPjQOqxB2N8e/rToBu3
CrGPurMlUJoTs3JD1Y3krD9vGxl7/4gztjoE3cDkDVwRhg4kvhpgeeMdDEVCJikVHIr/kJWPH6M3
BoYzsqbNMDepkYKs8SJ/4FCkGkYxe3lywCVDu+IkspvUotU1A/dQTLpQFW9XkPwzaZz5kwpiT9Le
d74WjTlBHH8lSfyeE8jo8m/JfCJOs3tHCf+4tLYhCNrZmb5C0cpR0NwF9MzWAKwKojJDnOOXkkie
barkSjqmzHjDu5+xnzfrD6IqDd3gOPboFs6H3u3pIf86lLfYfbmY/EBm7H9x2rN3YJ3dXKa1fqzl
X2vSuLQgZBxxUnMpnb5Bp7z/ZmIassJKW9VE0qA4AI+jyTbB4KmmPK1kAEl4aIYAlme/YjAp5bw3
7/VSdWQOiYVlDkK2LMtSwLtfFyShSWGJ2I9/PJrWNrOFiIyLd+2+jfalx1fUvZMFHtKY1AkK/+zu
k8YQSjB7m5xHvSKjJitDk4HCxoDbAMehqnqpeo6ht+oXsri1dp91ULI0NoV54sQYOgwZJ2P31wXp
+NqR0Vm6dTS/ms08nAM1Ghwu9N8HmjWs6g11UWM2X+fVCrR9mJYxMf3H/ispiTfUKIVSV+4SWqFi
QhMPAPOk1m0J0b0eeykOiqSfCeUV8C+PrPu6Ee053Km5BAs5uhC9rKpCZPdfXWbmBzj+QRLi3LhM
SiB7HobfgyBnuAw5grFJ5G6Zwo6bXeGqWZShDIZ8SMj8iUBz4gWykaBy6/wqv8TgqpIOEb12vxtr
o1rgqGcHBKO3IXmCaHFAEKybLuAxWe2A5SUIHx4Wql5TohlSp564JeidHIbHjNwtv6ao9Qs9Tso5
nYEMRYr64Armo10/HVcPxIL/Jutv284EuMdUaIQT5ryhdtYUKMY2hmf9VsYSrDxj7HbonAEH8GaG
St1ZkydOglyilG5A0AvWHQ3tquBWtfO0sXbK73sWlOAnUKtJ7f1ALplw+XsN8WAeXbzWr+S89rE8
kazdydj63LGf9bmeZjlFYXkhUYK1l+Wk7kFIOCX/nUCystnutFq45McOohru0xcUU9gMd890Joqw
VLAzSaxvhM4CGVuPkebEKnhFVepZdXSUiMB8Bv+REcLbMCy5jE9ivqW4DSIcgffdUypM0cjpuLir
8DAwUaEV1wiqhiFNf+hSD9OTFHT0EF7SS4+aH2ax6iWH9Y/vGsO7nGTQTUTOUu6Mw4Svzb5gZ86q
pcAYNwHtMJxmaP0dZ19yAC89rkRWByt5Yv3U7C4t3lhpDxyMTRZjcPYLHFU6TRIejUMfbPLsV2m6
Nt53cYTuFYqSHSxyOqlIAwnnLppt2lOLlaoAyXIduA6q4gwB3rTuaOmngmfU3XzyahM6o9fJ1oGf
Q6jeMYZVVweP+DYbq6mlEGjz+K9FATQckZGY7EcBNNf6rG3DQUDiBOEcmYSO92Mrjo7FYFlM3rUB
Tsf3EIWKuszWzRTRx4BKh8SZSeFiBqlASvihZlu0tDilIWL2bMovHDlrSzJTVWQF6RA0TrowI4Q2
d8JkxQscpYZ8K38rEp5N9hu1MnW4QWepAGfwEYhqop+iMFKCTCeto6PBZ5C40p5i826E/SQWliRO
yKDY9lMDZyiZ7/yKpOcqAVUNXwHA6A8ZNF1oAyXjC75ou3D0z4Hi15vENlI59aGiXrZAaopsjbjs
BMozj7HxdvlEuFpEz3RV0frFhc60moYt+FT/PiLudkPj+Nv9b0ZQrG4q4f0Fhf+3TN4N6zYGrOdf
PfQu988PoqoTwCNl46T6TQjJnSUr2HaZ/lvy4J384oMRW4CmyP34PWE74JROyVLt7sx36Fg7I/fX
FCzEqeMKXxEFMxG3Yke6BPa6e8Q6lCljemhSI68q5HNsCGn2l3GPDl6ylxdm0q4eSAaa24h8lRb9
ufKFssXGvE8hn/EaUvxc4WHRapFXvj5CkeBVm1nrNyUW+QSWohS0uvT5QGNM7DvVnB+4VP19gxFx
Ul4M60gQ43uapoy/h0zNkTjlSJnG5GU5eIjZmQGG+pxWQ+P89+4sMy5Oi0PDauCHx1PU2lLpIp/Q
k9+4BuMMdWvlrxpLiBqdEyORVtIWpSZ6eGXvOz1lzpcwHd8HmGnhjV4FCOi3lB6ugIQ2IkgfRg03
JTevunl0sZvsFdl6T57LElVMgzPie0+TnkT/gYBiDzy4YluDYbV/nDKX2aCI7FAw2PRUfq8fpboR
3X01Gu1vbQANTlyT9FiTcnttGiUbC3KbtI9gcnDK8iSnQS+oelAmKjzwatSxxyKtEkz4fCIWOi7X
Fe1wydPeuagWfFy9QM6hUsfyiGYHncoSQVyS5ok+PaosBQLn5xaBkDkULRERINMpsZLzGRrX1zL3
fmGpy3znpjbFUsaf4BNgolNuOiOb70EuC1iOwZycBkwkD+HHTrTo9L2wuVRU+iMI8aW+7v7jn4IL
0YG3R20Ckix7vR+VIN473LwcuW8PX3zZ87FXZkbT9tRhwHykyNQ8W9EAZn4yws0IH2T9x1CT46zW
tYbyWgKS4DRtTBd50nJojzfWEaSUw0STOgurYw/oUQNGztYEJin4DOt8zU08qGnBVWR+vyYAQXb/
aSbPNQBBdlg7mZB+bYsptroioACBJLf528g5XMlf9UpAFU2HBSkTV812NH8DKpsx5/k7Y0P5gM+G
8QCbHga7RO/jMza1jAf5oPLbrTtIoenPCZU/ovQ1N4BCNbtjowXu3mjv3keq+g5iVL4VJeoaoU3m
je5yrfX/Y6qAlDLsxQIqlEKheITcPeJ/HBSBmvurgOr9JvxUqMibyjbhs0htMpQeHgMuTTkCkfrZ
h2b3zl7bYdnjaxEgyZMeztB8KNFWduah2iwjWRIqMU/arc+9nkH7wf6KTZB5riT2Fhs5nXG3wIFW
eKdLdbQWBenEPonWejbyo17ZwMRudCqGtd6PSmoaM5GWHeQ10jGoo2Ova1TbcFOAYYdY6ohoxtXf
L0mO2zeU4h2i7QzJAhjHziSIwREHW88hSMVYxvhed3LcMQYz5A+jD6piSSMH29envpIch5kHDhzs
zn1MvjDvUdg/HhfeDYjt5AOFNcq/B2yt/lumIXoa1L13+Z1XD/ItKSvHCaTBravC0GJPwBpRLltJ
Gb0wgc+bqpQVrXk+nyA+znCxk06go850oHptEXs7HthUIX9u0H9XoF4oOueMrRf6bPU6X/93njWC
jqieKorPg06DiAo2aogasObCVNxAIm943x1UIWt5f35t2D0531gZO4SngH1IbctcDGasVJQiHsDg
uyA1/2og7sjUse4a/xB58oTtKZEVGspYqvoXtjTuDzM2CBqieDGLeK5JQc8liKAjsJ8xv0811G8n
QgmhDahC++pklP2C+Dtp5kKIqmmeXa2q0CxbBQiwo7q6p/IZajJ2KtIqkCrHkw01uJPMK24iNKmN
dMkOZxgMJh6UX3v7WWGcrfHMK6m1NqvT6QcQEUxXjdjxBAtyYSBBMUHyQ/KlTyCBzLQfGUMw9Isx
9ffH9+iViAPbuCLjvormrckQV3vhBohJDyvIAw5DinzcTKYBf/SLw5Yg9Hf9cwYjYt+l5PzXOga2
P2XpcFqqpjSbA4QeAesGLXye72onRiMw+0FTaXOxTuNM5F67SDLmEPRxhFPsaPccV7iYl0ldOQts
yr41/uo0jDaro8i+fI4cj7Ne8uIEaSgTxwwsIBc1MAcoo5ZfZZwXOc9PmdVaaXKw9hLkkJhPcCSY
bZnlfTJXEbgKNh8QBTGh0gv1ji3HS82jCwZGsdKq2fwGVX8Tl+7KIMN4jSD6G14WF1NWUFkbARdh
dN3v0J1qhNBh9UGGfPhpfdePFJzGUOFrLHJFiuBRDgqorBNtW8gSy2pl7EkG/kLdb1CuuPZWCST9
HvnS7vn2JdiutW4+rIDW/R+/8Q10zCHzfua9Z7n22kJEJwDDF5ILYPydEWqcLCUiEKLsWehkAh0i
f2+XUOQbjbxRDl9KZshj0CyKBOcOE5HgHjeJefQgQcTdpLAnO3eyFYTV/3KJq6BFNZ9k4l4m6Xm8
4tgo/9DJ5xbj/MD3hwkxT7Ou/vqxauhj1K6J2RnSA9v1w5SzinSRfSBdjzBtYuLcKb1l9Zx+XUwl
t53LKtnRb6P8nUMNm15jfCHBGLa2357u8LenkOxotvOhzNtLTwhySKerKN2p9dXviW/KRNltTgTs
ZRNOz1azWXoRmioXW66Jcd7sr81Gfc/lqrdX2y3cGaE4av6mG9xs+p7HKUReGXylluoi6I/YzVPM
5EBm8JOCOLEeqjiFUpXIEXbkAjFHSfj9hKSweShzhnSBvJjtMMPHmAJQX9AJBkr9cPQv5t+p5GeA
7Yo1mUN0zWfow+d2c4FloPCl7X7CPhBWahm4VFGjvbQYPojsrwg5TRyFzqc8AwiVaqE17ykzg6LJ
lPOjLuwc3p0wXHRhP+wnbqLfaCwjrg73t8RuipA4J/hePccRPGxJlVZl85H7uB6Bq3N7A90EsTu7
EjKQoZykKdYCY5DLxXap1Afd5waulstxpN1ESqXm++3y9H5gBIccLDlWCqvzTzGuyb/kfQODs41h
UJH1vf8xfWOBNMKLxX3uRINWLvyJWW48zUCdFlf9mNmueyYkySb4KJgsCfObdxY+dZeKD6csv3KA
t/W6nM6d7V5v+1/lQZ3iwkf6rUd6n3uNp3MghU1ZsBk+S3oSke323lRtHKcDCbq3NCSDdvIWq935
Aa0/qcxvgN4r0YSPfqhWI7lgvfADL5oRmZqb4mHsWBns0a+HHPedNm2ZM4s5GrYon4hbfoeQiBUi
iTCR220+GnCYWM3WpPJESYad8nQ4GdxTXHOfcvFy928CrlLOF5nsFKi2DZd9Q5JuR98/6RgWmwBj
TPxStGgtdxhkT5qqD0CknWKwxCN+KBd2Wbupxlys+IIbRLOb24vcnnWc5wpxCqh0RBc+wTYStyFN
wquZCFCX1YjUlA+whsxg/uTu/MkQy8H5d/dPnOXqMxIpiVqNsRDzPcfzGFA5GGrx5eJvbFFBdRt0
R6/uXygcj6ntItwq5WWM0NbtarFgD8Wac7YKjpwLjmQtRy4MGzagMQZH4Ai2eFmGoA+M7EPhs8Hq
Hg5MKbxjov1zx00DKgtIHjc1/xgpInDO/2MCUh4W+JgwDaKXkANEkBPQPUtrk1MT59cCwHat/luh
lRg958OdH2icSmEp3DA16IhD4OJnPH/ZPx+gwBPmT7vS0onzBQsOf9kpDpONeCnc4mLApsdrSV9a
BG53gISs1y1RjOqx6nZHHjZdos+murGwMki7YrJZh5HYUreLe7EI8mFqHqq3mcrS9xjSVs+1ifGG
EJLOzFZZm4aAmi6u+n1ZoaScWKniSDrxe8cXZstPiKZbV7F726PgXm+ryj436M7bcougNRktkt7y
/Fn1kyxKTczw42yRAZEFXJ7jMY48yyfhmnuL2Z0zXk5rNYkq7cY3X91g38WCNntEKT54IkwAXR7t
k4bnQq5oPUeCvvINUGZrfCD+21lNbmTjkl1BHqQN/0jhirxWl+eU9IIM/4ckYbgMsYnsFwvcZdD5
SaBjN6NNPSZqOt/qheLTuu5BxBu10SKFY77Ziv4rYdZ60qe8DVhZVDfbOSf5PwIxDQ5hBtrD6qqA
gvsFxaJL2VKiKM6huIBKCyh7eJ8NUCPYLnvYUYjOSe8qoUAOHhg5vDEY7WcWAEbRJjBSOfo3GzKR
iP+RQKa08SVUl+waopTI/HPYRs4ug+t8p/l0BsPVOOBROnbdCKTSScQBnAEILH+HLRHPTqEvoRTD
GwSIb8bxauIOquYhBD/+jhrq/mV2q34mz1Wy2voLbGfwP3vzfswBge5M30j1p397oHHylcobMvMO
2iNBoRsUxRhdgMhbrabVTtSgCOWanXk8ALqTc4NXnRuypaNyOFDQSibRulvT2q/feOotYLhTICXr
ttpKuBidBS87B1/W8qjRvzZvwdfj70KnQrJ2v5hInMmWGE1wdalhxUhq8h6CNKgGsVKShuzR6nOq
guqBaNnZwBWNtK7FNVaW1rcc5Vodj4hmSbOhMRhAEpnzlbK/Sq1lnKMmyoPJFwMVKWD9nER7P3py
VYc3pPMVaov4+gJXja2eoEFBU7UCEQDvq/4oZJ1OzSA2SEzAdqURQAtItlZgmct0iXdLSqMXDtZL
NrpTZqrcp3xGQ3Svj8i0MkFuVpTXezr09zXFKZf7rkIaDtt/dg6GMmaQKuEe0OGDBA6CeSIeAHnp
1Q+rcLcVlRQlzLUc+lC9ZgQ0LFMFwJL78375jhKVXpNN/jfh6sm4Gl2FWd6yotN8g5DDUKcaMKeB
auI+1/cjyRfUcTZbQS3h19eSf0B56OFxSduUkOSX8NFoMMzWu5am9Cvs0HcdrWovWr6lp4XuDVyo
3b18IjC/WVF/FXQGqS74cRk4mmZb9nqIplC4+YTRCvzZH+yyV7yHxnuV2oPlk8kDtOP4qJHjsp0P
NYFHHKMowfgtfh+D2lFhTBjCScHuGvOSR6uCydHhYFNM60fhxQwrxf+/wSk3FOUNoxXU1156pSa1
8IYnT68xNR2HrSwuWPwzciELrnRUKsFx5AkVWzPYpzGPz/RyojxXG6zSCoYuTAJTVoGKHNG1qUyJ
6rhr7MR1WtJjhu7TV4pAsg6FQ/+bOYMi3ybi9ddJeYAwBrTz1ovcJxwpFuUPSrq9ySjK1QPFyvEr
Ll7oOma9+0RTMhsLYr7bGlc7rFFrwtNrjA3EhgBYvPpXYEKDEs8H0XHCsxWZESN43QOGtb11gMZS
1RXDSislN6JCAwevWN2D6eFs7hS4tKrh5+KV6aef1NvvF3XkkAAjaZGejU04HxPWYcqBgxdg35pG
36m/vOahIarZ74dcOB2HBlhphAnVs9bKkzvDHvRXk0FBEsYuLWfkN/oYZXx/Ov1F4Ildo5Wp2a0I
x1Msrn87PdcQmjnpPhfVw8QMBlM/46htGx09z/h3+83MAcZLb6JpTwXTLJ5nZRgP+IpfyaBEMqnG
7HEj62jkPe4TJca7ca47SfVUpIUEheOjIfEsz961lmjWcSVxCmI+O2W1j1yng8HilRPNoMNZX8M0
+OwHE5i7HbVw4HM837E3Xxc9Q258GAg0s/IUsSuDvqJE+Nu0YFoQQdIsJCNk2gaTX6OQ6q7AWgig
UwJGYTpRcb9Nr6gB4sfqmalgfmoasFHb4o9ZcH+TTpu9+H99pq25iByXcXwJMtmUrUE3XWrolMQw
LStBTqUm3tAMYC5PzibCf0br0ZnhXx3wjJeE8YmmdSHqAvPzMvL9Bzg5pEzM+sofgNDrAQdluj2R
A7Jsbv9KAfHdmDh1B4hBDou5vkrHNoZl6DNFYzXc0mEaGswRPS5Qvt21+faFlWFnVhEiy+r+FHfe
I8gWjlk1O4i3UF9b8Zw7B2cZ1p3aaAejbcjbEqCKZ1EvmDR2Op6c3ORfaBc/25vQu++OWX6KvuMR
aW8++VI0vttu9bXudCshvk9HLuVjLINGst1cmHj8OP20wnMU9/pXdgYKa3vXRDPG1//jqBt6aOMv
AgpyFx3Er/KKBxhwhQC10RibJzP6SqqeTYIcIBwXY/h2kNenUXsLzOhv1b/fKK6sBL/F3PD8rGtJ
k3txS8RJ1EXFPj6OsFmwK93FJ6x+uYqmkITv0xqrxxrtvLEAIscg3nbGAWqqq77JwqOyHydmm0ua
EPmt07IV9zlHK2s87YP/6wxayDuFI2IxZIyjbrxSF7SZ51by9hWUgN6OdJCEXqzrVBw1HucoGU4G
spUrIUfl4kDPmMv/Ds4MdnmGDwoS8MmvAiBOAD5Qzc3anASiwDSON1DNaWML37yqAS6QbSJr69tv
WoE7RhDDqM3OJkUNbkxa0qILfA3cCM0zQHch1deOKqJHX0HRB17n9ak7UH5KW3U6jDBcoph5Jjn6
hAbki30ZWoywAPbZIV1Ib+9avG/Xx4ziWJUiQhKnk8tS6EfpN0H3/PBwqQawl6b/Oiz8onALY7hd
9A5R94UZDY36WUX1PKnWfV6M+utfXTURyzocWf+InCHQlsRhJf+xGfjJ7GBpSkYhmZ7nddxUDJGE
x4/NNEKjBNi7wB2BUwh8paXruZbtj8tGwYtc/YkZWBCANb8Rgf1X6Lw5sBk9bkqI4Fc2xgB0Gksb
xHD8lEga5O3d/M/pXQAssvEh7dVeEGX9nkNsVMJ+KLnKj71jeRJ+eIXRM1Q7Ssa0R4uGdZ2tjdaX
PlEOQgcW0RzOMYjaY6ROME7UzaP9Nc+b/xz0Knkqu7+yG9MP8DhYtitZMow7vz6GYs8uHkyu8Hc7
9wp92qecaxd1IoghL+hzFdr8gEjaBaQY/ahNpp0hh35glfuAIsd8Is4Mr6VS9awfzd67bfkn9lbf
YH2SVF9jtRFc2oKlwDf0glW6gCTfKaqXhHrms8H5MDJdZ4TIBJctoQmPXVDr7I3x/EX3Z4bpW5Ox
5wukS0jPzlPORPC1cUcZbUcCxwVUHtytXoBnWp728HuutrdausUFl3yvgjNNhn3auPMNenPCKE8Y
ADZd3CSoNTCinfbWd3LczHeOQ7S88phu26EWpcdZeBOITzhnkltotMP6DHHBcv65icMMtPO3z2d7
pjKGCOWSJ5ypYlqp46fZeRRQhcUQVAHbJc0TF8EzVw9VNJ1O/73LiEFYxd0L0UFxEoa4N28uZvdY
TWPkt8EXXNPPokMj7/fUtq4KUoyHvu/toi0E4awQFKpp0AFPlZPlYgB5sk1Q3rlXxnqn8OiwrNWY
cdJbKKP/ARNhL6mCT6977XMlZ1rOtIQASaRQS2YIxWOsGO43GwnkPhZb3LgQRoUIku6JP0yLQVb+
xXIK1jad7v7LHEz1FxFUTWwu9NF1pgE6GSppIF+PXl0QHA3RqpSQ3O+zO79qyt6VsakNhTYDAQ55
KhmVXKzXC0o1FzWHcaQJFwF8+bhCqx+v6AoNzNLmzjnqohePugb42ccAXhrN2xhFel/Fa9sbkbCZ
hFLXQ8Uy9mCqz2TY591XHN853ZSbxJf9WvDC5PaEIxR+6sKwRMkU2bSW/w446n9yoo8/J1SpUBKI
n8ppGHMYCvcrjt/tLK1Pm9/1/V21UEEXw6zvrnVJozEtOUGyFff7kbjfz9hG3CA+FgxI77pPG8bl
cyYTO2eojzy2VKncTmaiuwM1Dy0wnD6r2+9FbPlwBShVAgFWr+zi4SCtDtf10QkNqNmZUNhXt0n0
xxKMDvX+sW8UVuMJ/BMSO8vDeBpenmNb8URoaSvmVzlJVKTdea4sBivRMp5G0RRUQGtiRMz08Fes
+wp/zzzFmhljSnUZuAMGLMeHLogP49ExP1+xTERWKEzvWQmiTDZjyv2xUl/hzZO8FIvBS3fKxQlr
azlH9bOFFYxBhTUpor5kBb/5NBAbYhlGkphU0hFlwlECAh80q2q/IRGmxZWENb0sgJFPpMXAlrIb
MKhJFwj/grXmM8Ap4ChH+xnaGi9vOGQayio+7X2ryVgD0mbviKY3/gvRCbQDw0ylLBWLfo9nJfHr
opYSLWaXlZnTGY65fVsKEHBGeidTytmHQgrNc492CaT3OpjbKkcr3umvqkj17x+Hgo4QBkxp7Vvb
junIoaWsvTMqlc8V9PhXUrzpSTnfT8S/guRRSrmF9Db3IMgFyB+VPiUR6IbToLr1HwmqdpQ96cRE
/pCn8B7PKGOuGYcIqV+983a4+rXVH4mwVoBM1KYQJw0jrzSBnBTQci8lnl79WKXdxGzJQcQpXbmh
v3Imhxko5eS49QYrYCkYRylESQ3x/AWib6PxM4CcbOQM/PT0W5xgGHxtqV3Ln8itloWltMYyDyGw
fMGv2UX8qRIqGqbidhJYPlaXLJ3Qpalew96mcWbNVIf2N8suyLDYRvBSuERYvaWdb1P65+9WiP6q
pFEt4zpNWU5xIKgCMdtfU8r3263vMDE/pma6WEvTUvKiFlTgoEmJ0329tg/8UOIuPF43aA3BvoFW
OZD9BB8qXQgPrAlLxNxG+hbeWHygabDYTvx5Ri24Wvl0NmH0TUaZLUT5XnTuC/Um+PxqO8vDENW9
sKKPEFuniRy+C/p2jTwCXtNtmu5EsFYbrn93hS4wOel1TVa+zui+yVOAunM833BNXNFXuBv0qw2W
XUW4W8XUyoFoe92hCqK3ur2ejI9PJv3pooi5XW41E/Ag9IazQ+9Q24iLYhbzVENdwj22DcpLjAQ/
NRoAXbXL6hiG4Hf656v9NqKouwKPKQt9diTTp1IUm0qAYZWyDzOU41OVIDXG7jH5JCiAHgYR287t
BjoMUElLTxIzOLkYuNMjM5GVnuFRQcqxt8gxjejj4POf7/XTYopkcNoNhovwVdQLUkDPo4HlLC8/
RXTpMba/gDI4wImYuLyLB8kqi4vNz1rdNFcpo8UdLzJ/T/oeDRqRiN+mVbhzJfC27psabygypOmM
aW1sVmdqLNdWJMzI/zyoHLEFSKzmpr3CunImSoNeDAmjJuDvBQzTxSCp2mE4MI0Q5MgxnVyRouvE
+BHBvOJYoaF6B7KogOUDnpCmlQipDJfk0ss4Z/q9TNYnwDXoMNpPd43aLLKqQ7MI1r6sarafboC8
JvDOK4pSq1XzHAXTWluo33EmkTFOtZPMqVnYT5CyrJmq7W3oogNRqMoxDqRwM+loZj5uc8YPX3rr
50WHCU0LrEy5HqrWk791dRhOD1hsUmauwlYZVjMpVmxcoKbqx1c4Do3D1tPW49gY+AR2FJK3VMTv
z60ZPxHhx0s8lV+Iewqe1zyO63zd4NOz87h+hT5+SLip6DIx+0nSuM0rDFb38qN8aXtGm//ikp84
gwnLriGYh/lx55x89lAVsqWMfAEKfWBf5/BBDoYTsIMKxa+RWQuklTUJV3K9P2+kOO6u75vLDCR6
kdkKRRexPF10ABjIX4pzHNHUHnxz7pzyQp6lKaTFoe/Dk3bl0buZcvd7VWR+TsHg2RpLJwBN7uU3
4Bq1FwQEYL1P6aiU7QbIJ+1yvKuZiFDEUpVUeV4tNLnc7WPZnOn0ZcZorcMcyvAjYzLNXD1FQ/pM
jAnyVGBbECX1eCzugzDcoQnUCIuP/JWSP/zFkMcXsKGwYfPeCgFBt3BVxP7vGmFEpsHvfhj195QP
meWMxPSgMM65etzmTOTqyEwrZkR3wz0jo+RI3W048VfTecEuEF0FuodVXiRmmAYxjCLe7wNxT1oK
svtg1/BvWH3TshsGRcYCHUXXt0TioBvMgTzRB8X8ydLxKzbPDfhs68bXS1aP3vyd8UUOJc7TZVMO
y3oiYc7lKPnPIq7aeWITub6FZbTWDTlf8zoEX7cZEy8yNnEZLpYZfIA5/Se2T+8efo2Jyhe9UatO
lR6tQ1AbrOBXkI/i0dl/ae6xI2N7RqfU3KM0J+QPt7mqWFLG9kF6oRrEUOAsMFfSU8wc1AV1GMyu
w3mXjBFqEdbC6UHMYvL6AVqVJeADoppefjGTtbC+JTKt9ljPb4IiU3NTIJ6p9AhC+KxRaSydcepf
SsXawfSo+G/vc0JJ9gMqeXBsYQ/zJLgbrV7sZLGUQg7jJ3Cdep5FpGHGSfy9Od/qZ6YBocO9xVmn
SJykE7KkfdLP7hKUWhr+bKmECex3PwJ7vF/481QY/3VDytePD/fcFwzaHF4yz1TVLK6VP0Ey8xN+
sZgfU9ZnviFWk3hCewxrdwC5FQ7n8KdO8yFuftViFv83/gyyO8NvmDyYawYW5JcknOzCS5Cllbz9
e8ADBk8Ygl5YSzhc+dGKJGSSp3FCZYXLLtts1ZBwMcTA5MOG+g3EfYHPo6FzxPfNBKBBNfXGi4Lt
7ZOtB/ujI4eWs64PfiZnlkkvrER3luwfHDf76oRLUMl7QHo45TITqyluolXQKvaeJUR1Toos1RjV
q39CWc8S3NFQs5xokeklZ3+2Gl3x5upRLU9hatxdYfnaTxsJeVATGPmvieXaaQIxQ5iEn2rdQQUz
5LuRHU9iz1J1PGPfLFBgtH2IZKXMHRJ9Ym2MC4FWfyGgnS51E4i2hyGJProm/CGRtu/KWgmsx/GY
7cjTdNYw+nbrNmCJiS2qiHAtqU1diWvR/o6lUsGmXbl+AHQaLjwd5A4UyVl8U2BnqlLDdzaNpGaV
0PX4BPsN5fjQ5x/lquvCuQ45bKn3hjdnrb8uCAiaMluSJvg6z6QPn2rFvuugYkp4bHrSZqigrs6V
QhrTvMAZdVZyMpf8HI2h79dUeD3AKOBqk+m4gQ5QL88oo6L6mrUdBXyml0OPA0JfmyDgLEsRezHX
c0cAF3TfNRQxga/VBbsWP0MMx+V7Jl1yoqe/1NKIL83/C0XnyV8wSeHnb0rMeXjRrrtaTcTAYahb
k03MstHaZip5+WZlTEsMsDbWJMoUr75nmMbvJhcsy6jYrDvWhwc8Sc4TeiwRs0aYNxvwrGGazoXf
rGy0wSMUdUSc4dmnjY60oi5z1XzZD/fm4iHsNxCaUKuzD8aMcT9UxlI4ElOMM1Jk8cjoIAqhvQ+T
DUgvDGm1iqV7Sv4Wr6cZKbPSPpvQ3hK7iZIvBtD61dpR/9/1dj4ujEuMWLV9hzs0mLI53Bb4tDIv
/1W4lmVAIqFlNRNScukzd9dKV0CB/Emf2KAvKKRnIRpXMTPYHaseRj2d/DdXsljd8fbG95H5X+pc
yd1cT+9Ecl4HLqHl/X8Oz8kZ90ByLXEjEJ3S3+yI+iU0WKdaunrDtTR8DL0d/kBTh6g2nnUlS409
zqFjkzah0HI6zy7Ko0OZYtShLzV+KB4K/U/zyB4stO1c77w5UzrE1qxZmWoGJdSSpupbL02EW8IM
u1rDVPJADDqlEBAx1AvIsheXC/ReMXlL+YPnJbvKkI+2AHSwcDDv+X0bhsi2mLrIOLUAxeKDfciU
w+tuCfCsqyqsGPySq/az4tUguC+Qwd04YX5wuKpaxAb6TEOsRWUMS1Je4A0xiTckc6zkN9lfSutE
ZrtH4ThfbeFIpnLEEqDwWBIGwQLm/KAbDfEEpT7snAqPk3PTkLyGBnAzSZBo2fqVlmUqfEr47ZiJ
FHyyp5wX88mZp8BnCNd0bASZp97r1v/iQ3qnyJ0Bn967thtEriAayl6Ba9BUWawVJOlbbECOciEZ
DnsAaw6UTlhV5wVPeUEa29bhhpQnAu2KnlbRCSZ+yqV/D1OOagJe3jiK3xmZwzyMphznTGMR2Ml7
021KO4FSG8LlUPt8VpvOjXMcH01+cqFE/1RB0CtkX75QkMfPNyu0rwpp/za3+a9zv1g6TGIrMZqc
yQiKcAt/zQBYH8vLoJx8ejAhrauYdkXBXt+gvzCF7btNsBOcbmmk9U8THZcdTDLiezD02tYECJFu
NTDTkysewKjL3FiE8fDllDa88GGTErhn66VzT3m/50U1MBXiQJ1+3Yci7F6MP5BLUxzJphkKkkpP
1GcallBzrpu7F3pWMfCOZptB2PCMLxHfwu7mxEKkEF/v2iEdn7T/mQPQxWo8qrX2Ajj6ZUtF+g58
8rndEwH/lkCjCA6KNGe+G3ddeEbJNTRiudskiFRqFuU0awqbVl2dViaqsEmyXVKBK+lxgkwperVK
TSUCnF4nkGdatlZLu04NE8irKKFRzacnla/VbsWISmKsxMu0zgF1xX2vn07xnH79XZ9hNMJTnEem
WANLZclAtu8ijz1vhkirFv3iBX+H9228veuC53Rr2W0mbZBLZ3mAOA/Ls1YLhxonzRmDj3N2OLok
hfKv4kh3CRrUJqO0voMn3Va1FYys15FKV+WlKfJ2u1eELcuu052u/k0uLknXCM1AtAI1u1VKgBis
2b5B56EacBFd/R0vMN/WT3qfedtR4X6byJCp8KSp7yn4U2+81/oHLC5MkfeH2rZhRTkN+qs9MJ8f
gBJbkgFB9NiBkJfaMCj/ABVrM5qMpO8qyZOWQi644JFjC9FlTXUdQv5KdoW321k4i+VnpipmyOQi
/SWdPwNQwCfLvwR4GVn2brIH3xDT7/K5KJuaoSahZHX8EIxL10zHH+eMY5X+QxuLtGcvN8t+0/ax
GP8T9lwPduuuncT1GSDKSb9FjMQWzP2vLfjsBhTFIU0zaX1GwbdviyzSQTSabJDOqHUwYmUHiKTn
audQGmUNQpKclw+l/NwBxWw+bmAReNr+UQmTabYOLuaFMuj6vsHl0/4H003uF7sq6TMRqZylOIlf
hgaXD3LTh7usxeEEl7/Ld33YEXlHVrK5bUIJwYNYB3dAS9plty7Dx3k1P558RaaoJ0WKTAWPu6CR
k6KWBCfMjOMN0FapjqCKJMgvBsQXnE2u7MLzmjAyDLMnq4+VORKFWzyV+dmVSVSYvDJFrh3FZYZS
AlEwkaI1z1PgkXyRfOHR4txhCSk7Wbrb1yQ8wgZnEDrRQ0LQyvXyEWySFpyWWL4FlFhjGicnqb+T
wHLGbE+3fCNtkJwaxfT+nBDaPVzpKiGeOZb6r7gBCJp27kD4uUBPl9WaCSg9BBOtvlwD4KitpwCh
e9L0/VTxiLiRgsQNarXC+f1SGfE/kVCrczLFPekVwsjSVYvorHJeBh7KYnAnQV/GdVz92AHdzD3B
mpIqNfK6q6NJ8KpxP4xTA+u/lzFjRupLDNxI6Kber+3RGpShoYyOJeBA8bNrLs4s1oaeyTPsjgBI
N1iNl0eGOQS7bfGV9ami/8S1t0z3lziQ73sFYL033fzsP6ZzTbbZZ5PChYGntm8pdhL4bXURulrn
Y4N/Fi5vGxBNPKKsWzZeadjW6maaaFixUVSduY8GnvvqzSUI+Q822cEB9hcYVnJd8Jwt5J9QbaNm
FOHIM+KX0bEbR5tF2cHEjvEey098cxy0J4vB3ehFNMPXm8BUt1e3d6z+dkYjxjALbPniWItTt7ee
sNIc5ynAFogEfOgOUIao+D0JfMV/MTff772MQLhwdN67OBhct+3DnYYhHWW4IQvRAirhzZD5d8qf
G1qHNfbLVuYCPLhTGD4MY4EXiBPorZDEFBZTy+TIjijSTz4g+OsPJHClvqJYjvqpYwafVZAeMWmT
FD4PmPMBOhgfqKi3mSXyjf8PwVqUOsomajZP/k6pj9QdA7cln7QDBj1dMesJZqFSOVk/tgCMSICB
n5r061WroNg9U7S8/jCV4zFrDeA8aM2aa/WPRIsHCOWvAwP0zmw7RzQPjXwzhjZuwCOTTkBvwyHy
ydJ3x8uMufXlbWVwajz8kX2V7hn+v3OsMysvKI8Ee59Eav+6VBQh/zdbtjcq/LPSHUfoTMwJtYaz
kY1088aAuUQxbgvloEAg70INWuC+C7H1VgqqeP+tPuUn4aTVfkRLuT3EmIYzTsvCNOaLRORyGO0P
6WIYBZjB58ttU5rjGR+IxX+NxjvfDnxCswuy9TjAoMdk365WGSlx2a2YAuAJ2VNohOCYT1kB3duz
WkrkyG/I57cxXrF4hnNhu8/W/pbqwjIZtlZYJHoOjDvrembg3l2IHrJTcmP0V7TsUDr19j9kp0T8
jKQO/jP0G3Y3RJGJW/M5d6dGHRumw/gfpnsnfkOiVsyGS8QfFdM/d5ou7dfjkL1bNQZpj45lm7i8
v1UaLFAL/PTpm7JphjQ2wRtidwr6AWY1ObDkrkgYgqsqUzbZkrqyYhOSmr/NMeg83rynTBKIKgvn
DJkDEvLPkiffEVY2KuibTNlx8ZJ+L/eN0LKPovLj3VOaz87rb1m5BXSTczBJSq+grxgeizP+oOBq
r4kZ0taqLV0QrkNx3is5wr1XfPvaISzEJeIVBYyvgBYAr1ZKVwz6YMAeXF8zxt20hv1TF7XHFKQL
sxLN7bUKbT9l0k/hOK/ZdL101QRxVgBHiCIecCPE5X1lKiKkFN4wf2dn+nmuWuvQvu9jchOV1gxx
dG+3a5pPFor0pofDMWnviH494tFV3C5MOdyySnnE0+3Dprk/xQJ8Mvoqq6RantOGtHRM274ucnyw
L50hSUni/5jwv+0e9ZrjtvJjLzcq+90KiVx94/27aKjGoZwXikYqbHxYwxZDJ/9bz8tWfSB00f3s
TyYb2GKbFrcr3Q643KNADmqFVYnuoPBhjCg4eSp9MVuPeugprZiYca+0Z0oRn/VoCUaQTkAY2uu+
Oo/LhWrdvg5q/ojMiVDtvHjqY3sYdvYizcrjwDX03sINcSJYFYxqjgbP1UyZIil0xcuiIgoVDaC4
uZ0oBVpphQziqCzgDvXkZCz7E88S06tnEjZ6F/yKiyNj90uvqO+ZXpWtvucwRtM3W0rjsJ5+ISYE
hbGMTGJPO0cTjf0TMrbh5e/UkGX8ynXxz5Pb84hJcSek7LPFt/pPa8qEjzznpTdQkCUvuo/p2fwE
TEyFml3PMh32cyaKh/FqV5Kw3jvf30ZKCxvWfKs9ul159vg+UWOq2X0R96I5wGYvjlTGxmOUJ0YE
6RKy6k97IDJl10v53VKHPMDxcCXe6j3NNWmMtsrJzXULbIxzHXRY7qkVgh7kaSqKuaJRgLMq+QGf
TzRoyAOu/u05G5AyvOnBccswfJJYMJjD9gVaSQV311Htq3oJb6q/duHAyQDNegQS42hs15WPnoik
/hZvviK6oXwxIg63rPXgEyfwdgZSVw/sDDhNYcD/CtRqiTrlvI3O3bhCql+AOonndEVJQUfIfCFa
91dKWwhMT5xnFq43YdNul8mYh2FLopAUKZYrcVC/XRzMaJcQjlyemKlaeGfZdnGS41vLJhlDbp8q
eDpBIIKwKqwn9VLXA6EPmNKOfQlLMteRaHFU69ktnf8rm9TVAwtqcNB6LPZcfYI3+zFtQ5BzN41N
2iB3kV1DIw35lcrLyYZJ9VrHFqv7rACFUyotxWKbBrcd3X/Wnduu3M/ONu9ggRkJtDwxi/cjeoBU
3bvauCKimOPkWmygwv9R2u9zo5m/seaI0dnsJoFHsBu5IDG9piz6yEOAwmNFBO4e5ulySTYJUUyO
Xp8bHMcHvw3tFvvrNfqVyCnEsYrKdrsI06b1HoXdXRHxueXE43Pfgqs8GvDl8tw84uLRfBMhgIie
wmQ3d+5Fp3pgrCOso/0W8qECtje6NnkcGK6lX4dYOZrcnWIrdY7tj3a53/VQ4fXR0Ppfc2w1sBLJ
k3VMPALQVX5w9yWzhB0AvPZAbRjAZX4WfWqVmKnaXywQ/17SMBo25CGIY/Xu33Lo6Xe8cDnKIJJl
5IynjVPQ5m/tH6fMDh3iwLuYKDh3sJ8203UKyzt+Ay4ue+7P+jSW6pE3RjkcgLTn0QRg4T9hD14W
PLwFD/GN1ZR1+FSshO6a4qrXDZGFrDiZRCJrtPJItM6/EV70VAJ0CH9zZZ1/9u/qrxV6Ytai0skm
fkNTstoyWNybsth/tuqRB+P8IhYN/anBHPixb+KRSJYV2R1xPugHSU28GmGf1/PRf/tuCZEQJP+r
QMtbhS6Nvki564oPn9Z7IKted+bi9ZTr2PTmSOjQ9iRva3veBz3su6pjMnvJv8BF4ZkLFIkBzKLI
9wNlTElusUNbawODQFAV8dgoWDRWs/NC6706YdDnN6Z7yix7rvdngedKPkJEKos5QsZN3KlIzHql
g4oi0AZjLFN4BUDFJ/XUbjrrYhqqqeLhU/qZuByq5IR5y10DUTDZOwKK8sZwNKabw9CTxcQ0i1op
iJfnbdkbGjTXo9WbxoOAPoURBm6y1jYLDKCxWZbO9TR6UPXe8wShY8A/dXYuylWiLgpSTTFbDiLJ
L/o8Gu6gkqdp0rdeZASl0Y0Iq8kCCPofzq1MFWKPWQtqBwVmCM9kJeDYLNkN4DGWjmUhEZUwOinJ
5jF8oIUjyG44lHVguoxObAO2x5SAfNPgFT0a2xicyLTQ4//OXVEmYSWFZywn29qb2QHQlogRZuNJ
pQ8O38ryi645sCBieDl5EVNRf+RABjCP/o6RGHr8bJkYOwkX9BlGAwnunpjoUDfna/p3K6xY/1z3
CqGyEPI9Jhy6yegneAqbdywdYy7SbaYUYn+9bqrnAa7gK2RZzBxDmCWFY+P9b6gjnO1meS/s/y+0
SFA2jpA/WENRfZMO64398SclLe/PEfmymXv8Mp1LzGXPn41t0HY0JKU8y3dMohv/zZkNcbqFQveE
D1HQnKj5ojJJ+IGB0MVbJtYqwlAjJCsxMLESHMXL45kZM3/zJaOoGP9TzmQxix7J7ET4Dh4ch35a
G+rk/T8WRo/czpAxMY2ag9CO2lCKkMr+gQ1Qya9bA/D3s9i4gKCVXfziSBjksiO/qsXubT0Eovj4
TJchYSlPRM5VlBsrDK5PpByczOLrFd/N3SD87Kw1jpmvnDQ8z1dyxlSZIwpTJ+ELE13a/iLrvGZz
XoJqeHzwkpIyf7q549MbS3zGKUbfRrRahi1DxdZbWeOOrk6TyigNfGJz3OG6akEwKpwmFHaUu/O/
VqWnwldDzVBtqHVolGXPxopTb8knOD+ARsT0w4t8lojtI01xUjK2tHFgTJMuAuV7hGCbhKmQXInc
dtG7ZwWxWejweSqpbaL1cxUFy+Dmig3p03J9B0mBpdxxc0l6uSzascbllYWj0U/dlWPhq6jdnpzF
f9iSZLmJBU+HtoTfXNeSRyw0PImpT9fA1QI1b5MLajG6aF7Iy5ymfZIhQH8CYETYrR5lyWvqiTCE
/txbtk6m+pfWeTRfWYL04H6B79GFJwHJpR5eguReRArlAIcPIPKInzao4JN9SfsAo36pBAUMyE5M
Z/Mg/2VhIs/iHRzDNNGOK0GrKcFkDKK1A8jwDEcuxT608I0NxHIz+vK2rDMCZxuiDkj6u9VA95tT
PTdq9cau1V8qUKitjT6zRCX9H4UoNtlTDdDE1DrYbMFS0qtqMCLshysQ3hUyKYdsjJnA7lbz4FJj
w3QIjv5Id/7YU+Gv9ysPickLBQ67/pJeUjJNWbSQLWThj7xC23d2qI5l/ly1ZMsVVlSDefKUw6C7
WmICZvCCJ44dFwjjxFu+wzEbs+eMQdbXrVoGD26CksFn6dTDCqQ+AyiDqSX4GIDJSYXKPFF6XfIw
zj2ifPoGdGdSYnBFnv7dCTIcrO5d2KU0wNiRY2Pcw3sWooajhWHa70XMZx1ySoG/JMiMObWL4Hc3
qJbz2w4MkHqaGMPlfZwakbZLyELYOqNb/96iOagiNJ4dpO/VSPg4Ya6nhdMKNQ9Wpoqj1UOVCXgO
P4g/A0mAaDn/jF6Fc4EWOKu1qFJMX5Ti02nFv6r8awhQzgUIkfg/70+JkhRGqC1AOEpi1ZXQD1w2
JiIQPgzVtJA/ODmQkJ1heGzfH49VTLM0oZzy1W+vxybRZpm/9yQ6zBBeU4TywS69tZ3VyUj3Yg4n
xmRfzklZP3s3JiQaCN2QgDdvpwaRr15iIds5ni9+yXrJOCgzYQIqUOS6Eq6hiFmhuo7qcoBTAXBU
mNrgZ14gBFz7AWml5kSLlgukC9hJvz0RU+zBd1i0dj5kQzsfCOZB9GLac+Y85OdNtUBpU4JyjbvF
QWVSr6yIq/ZLXMS9PC0pTaXLPNdIwfpsGng/4fh/nP+H+GXSCpvOXtvQ+zvoaJ6oYB53IufQiU4O
R7fVnqQnBpbHP8bPWdPEDgE7re/ldwzos6MImXezHD1Vd40ln4heZ2laN7prihhg18D2C08PrwoQ
t0997+LcOtmkgStIComGynta1ihc0Rus2ajfYiQynzWUrNzFmH6oiFNQUXhv80V3OcQTMmWuTOWR
GUbt3ROchURKsb68HzmvaWsSYbnkM2CPqic893808GJOMktdNC7wQORvTuiwiibK3w2qivL1fhrR
jLLpshLqe+e5UuftkfuN9W80D6M3VN3ogxVvb3XslIBQiQuUtJTB4YsI4jer7hk9Fqq0eiWmGVBV
3qvPjPdGJC+TPg6TJFjg+QbfjmDC4X715+hREU58rlcUwWR8jEgF0BA0uEhyqoGkRMdISZuZ8idx
9YgxknWeInIIk0b9pzNwJAidfi+Cm0Eql8QiWyhaKLHJA9lqdy1rdAOCG7u/xOwpDUiAiwZ6CFkU
vjE4IDb5FQFU8i4iMsLpfLZzElZYCfwBjoobDCMwZX+u+fNBqG/QzfNTSgmZ/c6BF19Mc1aV0OGk
EBt1IFt5z+9b+ywru4Y7gJL6c5le0TpdI0AkMnnDzHHO1IPBvMRRhlFmZPwOdWvbn0qQ56tAaswn
7NygSRfVHBoqUIgX6ijhL8GhCPYJFH7T3oJB6d4+vVgkj4++vLUPRL/bYGNtXCLet34OaMrpbGPu
stwMEDZY194fgBP4XOCQu3f5m/6u7TDABT8+Y7RaziIB003t+JdloyYaXnfAGcZUvuCvNqTVcq6n
YNnSM8i0N2m6kyok2XgYEU4noC7tU4sJdXqQSLH5VvpjpVg/rsoRMZbxfuNNvbhywAQ7nwLX//Jl
kNM6Igd8ltR6SpHVw0hsTa/AeVo2hpN/PxgR94buV34fV3DJYosby5ESibgDs5xOVpL1fgI8FuMW
VNgFQembGy6/cvqHc7JIQvjQKMQOCOeFAcfBI3jXYhJVXXMndu9jwI2aY60FIggDWJY/FAu4F20f
hJX9rK4RCaGd1jloEBBoWKheiXSB59mdH14a6pLl/LrSdOEBgycymgIpvdI8cPWcmcuZc1BzcqdB
5+aDMmec3gWzvFyLM086F3ZMxLTCL8JVz0hfqWkks03hAAVHPfepoQW/canH+53L6NF5xzDEkBtx
Mwa7Z+40wndkG7Gg9HByhS3VFT1NhJ9FzNTc81Md1jyz+IBij/FU/bTGYa4HLNNL2y4QK4Nc6YO3
VYA0BKDXI/fkM/birLLn1aM8MUWg63nbmA1HuCuu29lbnhKl7mP90uIc3zTtKHskz3j7uatYOFB4
6NpHWikIjjsM5NV9UW7CbdtWms/P+jfCl1by/I8WqOjsbr3zUQJbJJt7avDUjGzI5l6sSovcC8ZC
r74oltz/X+3BM0zPJiQ+6bBOHptJz7w7FxrOM3f+1ktrQ/wRPnCIGCaOoD6YHYZAZ9y+qakPM6Qx
arVSB2cEJFviMJZhA2wTdL8W2spT24DnKNuromepPrOTWGouhBuz336NhV/mwM6ZDvPOwCC+jNWr
ryl6jbnXaNxtFndN0a4TFhx62AzzBdOej/8KMhASR02vf/i9i7M8giVLAGUiqaBIleXJg9Zv8T4C
2duIIwnoeK7yKsGJjbSAQgem5rDFI1sFqVbvXeZzELQGZxm2sEyg9M+7AypBytvggXzrALY8ZgMj
rMvYjzz1/xF4/EBmGGyc+0rEm8JWduz7rxigMEXyH6chOJlMxqAGDCxs7B14bQEK0JaJLxVcCi3H
kCXeqzBMCtA1ai84NMW4QQMnSOkFWWPpfGkE0S2aG5YlDKUyYLlFlvsxapBkMxRh6/VeEbt9YLVL
iEogwWurZNbHZjh0s1jbrHFVzmcPjdgroDNpy59jZlcRMCsFpkNGaBedCyt9zxoIBVoH/4baQTof
s2nVW0PT8bsCTVfj+cJ3XRi6XubTtHCtvc9zPTo4gwg22+S/e5qGpEmAkywnh7o8TK/d9Ho6Uopd
L+vhn5GCu5DCBZwiVy7qLqPv1pQ+ffSNQydhiOAwaXuW96mJe5z3ZN+d1c7i43jQT4AeIdGEAYqd
z3Dd9/dwnUR01qVEmX6LzUbGdPSjXfM8IpmzPaf+9ifD1DezA5VZlsdlD0Mnpgx8ZY97SD++jB/5
1MPPBXL9irTflIIoNmZZ+wNfBbqty/j2/OvrpolgUcBBP0MXy+WsdNFqn2d8R3FypVN2GjxuJjQM
9N5YPPMnbRxn27paT0OB9UQ7+tnFDd219FiSv4Mz45f/fRJc/5d4ADr9LPE5yMG0zHgJokPwqdGU
dK5nNASnrb54Wf+/I8YPQPGP9Yel0OcSVhwEg8Pkl3ffhsuV75nKXFiRfyW7/ijwdKCS0E1O0uRd
eapSqCMBMIZtykeI++2MoDGoTalbsaE8ahegDHue1TuA9qtR9TrVmKO6VuQDnsoIsH1SdxxFdomg
1iu6+gM4r6dV82FI8+K5htZgCq0VH9VcYQzLoJfBHNgQpf5+W57gVihVj7qKQFHYoo7IkpUHEaw2
SHoUaZlooTLsbplrtUKYAYQ6fN+VVd/Kw39t4B13G6OJgiiBHMWil69rn7Tb276oRDxcS8I3M+zm
L1HFPLL2T5fSyn0yGfQpbONwZOS5yOn093fKkURH0fpn1MxGe8Rg/DLGI8WHdkLfljWgiSpzYVo3
60vFJQtYRgDBgen0u4TSw8U2TN5KJiMe2TrelYTMRpenn6T9tkd4t1Zc+1f3CTUUMlsATVz5H/Ln
6P385UcSEXa5IWlZGV3F2Y+DN9Z0xbhtyjLRG23LDjj7CHz506zxbhBNb32Mbi0idsEGOrOoYQ7B
o/knSi3XhyIN8ajChrq1RI2hGbtecGB0Y2as5EUSi74swFCZ2mEJ2S6LYZuINBxtWQfMYz5pIqBF
gcv0063UTv72+ABVHcuI7TVE8akvWXpqHaI0zSLyO1lNBzZ/ixvsXRE38C9Ubdk+aCxiULUujN1F
Y5w9sMzaFvnJeNMKQ/cF0+At4MGVqDsQbtsUzHxX/6pQ3EijdH5Cd7N/cVwCSB0w1oTUPQ6E6mb9
UKI0+3iVG+5gXiKDZJgEEVDWihUyNdj+unuY7sLNEb1c0P/eZmK6wsp/EUy7sbZZjBABhA2rvlig
saZBxXll5iybqmt6X7BFKmuebE5XULRw60JlYfV0aS7xA6X167Q4O6aJl49L/RODgkTHV8oaCScb
rdNPCfpmOHd3tNlqUcT/T/mopfM3j5ikav7c0046yHvlqmJTApxYvOMAyXdUf+r7zLu1n0OvAllb
olxrd7+Co2NxVgPKnv+UpUX/vfIysvrJRILqVgyEE6+u17PcJTeRebdD+AdyZqetrecPfDCkjQZd
u7dUvUCtBPGHbmX6+QjcjY3mLFW4EYhrs1aSFgUafn2AiqQk7FS4vWmY+XbTgTZeDw2rQdlKxGlk
+caSzKrLKOhyFTHFWqhDx0b1XQ+x09RaZDSIs+Bl6oV8WqCjkkgW8w8g8QzwsI+/GbVzd954I3Xk
zrcehX/enjBfSRtME5fWo8WrQ2/0R78cnwjgQev7gKD33TPbsTMuPiJSZ3dxS9vnLQ1mr7GNcYbI
Nz8dCeEFiDjMkgTsXNUUwtdbpfsdH68CW3e+8iH3iAHHlZZPukolqUXrvYOvsVZXmPrTxLLTCRai
2Kc/Wg+0RRBS9yaY+EqzyhRm6OBnzJ4g+/HO5te3ZmTyrtrDalHoB/NY2OlKr1fITJqJ512licsB
PvonqYY3/TIA6cKFwW98IqjLJ1HGkSdSasM4AyDs5G0GCg6y7v2Ot+2PipgdTSfeB9I8yM/mp3QW
RoWgwAq9bkyZghdCCI90EhuKERjYOMD6u494XR0bE4EigZTZirRTlH3pGcU1QQ6r4IOGDgvs3GKD
B/TaJb2ziXIladU+i+APxBu+VKvoJaPI24dkb0oGOvSr+x2t/cpd0BqSHMvRExRncl07z7JZoi7y
rz0Ech33bbpEm6jaHc6Mn8U6NnLhh/xyHQ6B6V63waa/S3FqjH9yvmdaFhLJUQRPNgIyQ4ZRKfe6
lGWcyiTzP/TbLO8g2vmXSjRopg1h0wmcPpVjoyvwcOTtKxmqUdcrV1M8zSL3JfeVRDXJZDd4pErI
jDXq59/szveEYw+6hnFoGUeXXKzCJU2wnGdywF+XhGmMugzU2NFcAJsyvcPLq6v2WNAxwaCybcG0
j47eDVVyACABscDGJkw+mICpFDMslTmWpikKLFp9kqkLverYY8gO0pMrtZKWkisN3tTfaGaHHtwE
vh/ZDJbY4TNtJgoE9GNPdzszEy1p8LErHF7P9MHLjnn+iH4oc9PYduvIqn2zsD9hZzF/eJl0lmL5
KL4PEgUxTnwZD5DMm+MsPiVzCak9JV69hVBQrD/D+i9abv4HOgVO5mpGK+gqYo15R/mTtvXuWR9T
lQgB7EwHFkUQrUn8/1ptuph0wLC5k3nKCn3F73CAzRJg97db7qVZCGKze4o12oOm55pfWbv/Ouzj
SThhFacCFc9uLy1C6Vxr0ifGDqt6ajATf1E08RXqpLgELHe9keBGns3Tewr8PeY3RGmF5vUfRFGF
5CUO8VLQQfXPNUoP2hqHOi0Rb8SEutQpmmGUbO6ryH8nFsjga/NvRukxIk9W9XB+Ivll2xFLU1ny
1yliAj8/FcD3KXS5kLU+DhRZwqTZGtJlNY4CyILEo5RBWrfMcccqn4Ej1KnuC/5L7eBZFNYY4amN
GI7raKGR490cLEoARrRBP6wFsZsCFkkq9fl0uf+IONZAZZWYhq31luZDdwaPHq0FfhBULIoBB0UM
169PLd99hYAFsEF2fQ2Z/OH/m5e8mQQx+Nr7YWT/121D5ztkxNWxIwESqCyKNN6Awm6C5GfF7J7J
9CojSWS7mVetHPw2PnJ0RwESxG4JCJ7BIKPkYKfJLq8W7ZHXjddzA4WMxQNsCxtqf/ouSRzjU918
E2Bca/n+TXH6FnN6NarBIj0PMSF2avnEpditsniDTNtcXgdjWo3zoUNNxNE+dz8Sbn+uVNrPhhkc
kq55KtoxnVXTdNNIolG+f7ntjXcn+nMjZeAMgeVRmY17wg/BuQHGGSWExu7aZmnlZQ9htqiCReOd
mpriv0lUCW/PDtgXkpVNnnUHauxxfeJqSMwiXOD6eOILy7yrcr+RNfYN9vQiliky8tWzdgjc5dQ1
zbb+3pE1a1YwCnSOVm8PDWAV4wkThJdlN5alKsD6UjjIQYgpZek/9/FvTsxUKKFitbrtA1kN9SOj
hYL9DJy1TtdA/lq7Go6BxdsDHrRYI3yWO1JH0rCNpsC98UEY4gVoBiTLKJaI5MwVC7TouTQGX7fb
hB5HI6Gm9wrMnSt+/MEpgveR1yhfE+6ne72vEAIDhnWMYY5WElLJcjM05WqeCOJUqCChnDsr/ym3
8xlfojySJRHMxCdDEHxVFfgJ6iGKd4pIRXhetErxz86JWRCClfJAQZPVVLMwVDp4EH7Qw9bU2BNV
+SRBhCqK2+llZcR6Ld3PjgJ1boU7EVD/g5EAdCTWk4oDqEFwocHzZj1H6Va8wyzf314USi/6aZmw
65LrgrAYSZlmpgy9gso3lPyljCRyeywAGZ0DS3y+PEso1339vGVTy7aSbSlb2KCEJs5Tj7qh2FjJ
U/Bg5AjkSA8cVITdFZI6Rz+JgOv9rcGQtDptwX+yzNQCiuaz5Oc8U4aEiDHnRJ93HUIOWjzE8aQy
ZLaJkkPyFuPoSdnjOazSWtNjo+Vo7oULFq9h6j0EBweALcXLIQs3LOEuFScVhIQaHD21Et9Kn1zd
02vjON2eJ5eQ0MUg4nyg4Ofw2Zk/AZV48Rh/ldudQ/xAoTwOxPXQk5CO6I4Ulu70AvWK1scXZPQQ
gwzkmbe7STmmzclyTez3wP3erlOO9Jl3UHsPUzKmnov5hJaBuTdv/w8wtOG//3EjxyD1IBtXWHHw
xTKfnolwaoIOcNidXKGyHkKZRX7l2awvcrPvBFkbWRtcOAx8H0OWo2BFNPV8tdgcYOUd7FMEqDBQ
xsy3CUiReshZjXPwqgr8Fxg8QbV0hT3jIL5gdghOe6qqcRjDe1CPaOZh4Wf3pwb9PVnMOJTeDukc
VsXnN/zaOrOb7VmCzi4GSHEAglpMwKxxZz2ZPIOSkEZsb2j1zfG432w8g9KNyvS0+rYe2vYJgfhI
ZCChUlzlu1grJirZzNiPEAkFALwfSFZHmkgbnM+xhzJ4bQRItOXHry1cr3OqsIb5+zcSKhaWucDG
UnXa+0FkgLLCAGKyrkjAiG8bGsdVn5lNvWbrP+mAD3wLEzVydFpTnRD/wsr37nIoGKEUBJui8Z/r
2J8mJ077zsJ3KM29O95OqlLLslPagX59BG6qfxKuCBpVLTAWVOxWGMj27bXGgpBTTRR4QUKwkzTe
DOvAnMEl5UjVyi8nAL0RxQvh2CaXs9/owklIStxVHGdCf5Fj7qztbA09qJKAyXSGVGcWQo2Zrlnd
3l1RtuZjYt+d4WSED3ZxDMe38V00dt+1anMTcg3MuZep/wVEwPj0l5QtwPlrbDSnEuJ1nKUfbCkv
hq020ABuwfqayP2122QOSut0i5eqN7w3aI+7qqTgMeWlWUyzoQfni3RBFkinI/9eZkwPt6pHdSp4
3eFE7Fp43+gXRJlvqaqB4Gt4nQjAyaQ5W5GV88zPnjxQsD8ad8od9ugqf2ID2xsASF396Hck38id
0O18q1LeRP14u6wQAR1YxSskZuSRtDpcbeZRexykAsjYUWiiMJ1Y+c0BxdFd0MVphRQlM7El1rv1
NbPRS0j2A9eZvUm44URne/KAYnn6iUgkEjDGMT2hfyi3PO0V5YluIZP8bm/n7VmN4iqgRBNbfa3m
7uVUkogIBCKOTDlCWlWcdUWA4ZCuLx+HU3Thbky2CX0Clwm7jRSxHbfizl0gZW0E5OG7qGjB8TAS
W62q36ZYoA0S/GuLIdiTCyrcSpRevsR6BARg7dTBxPAxs0RSkfrwYl/x7jS8OE4Lsl4YjCmlTRvD
DU1vJ29MJXot8sSzMYtgQ1z+OfRjXzI1soxzyE/Hxlo2PMDyqJ/TKqs9eiQXIecv+xpL93ZKA+uw
00LHpJUAGxF1FvbgIbaQMeiXKQXO8BYqy29rd1wFVpjhQvP3zUQk8CIkiN76YT8IUFYmDCO+Tsc4
eUYPI+83qCG443bZfct2ub1sSValrHuSo5r2Sw09DEGO/m4MvLXhQOKzQKsoTJzyTjGnsAHP5nxL
BrxJ21HqcOxYBvSdiMNIGAGxAcb8g4FcKzv9H0CApJZub5Hev987rxMXAxIxJIPOz3BWd1HVpXCw
C/edlcpNXexUqT154yjihatiITv0LsyOfwTuzpcQSt8J8DcyGirAaMfX3CUY0hDZKsmvwPdlQ0An
FIuv6OMMotOPXqLSXyITlUeRqCA4WVY3ggF99nKkWWVJxl4lFD1/S1DEOuwipRIOUBJYY0ukskkq
JirmmlyeE86VBU653db8f9RsqRW32FZ2ZNS78w4EwwUZAqKE8hPfxIOvUowO0rEoDO8dhuWPLaL8
Lhy+XON44xZetPJjJD7ohrUFvG4SRXVKW/zFDNERW9e7ZIQXwTPI09TvRe0wvjRsjt5vE0pX7mNG
28go98yv+4fOdMtO7OuTtXyGHZSyUQABUbMC7E6T0HVl0YRmcM+fgl//wSJOlGG9Pq2Afo/fxeKU
Ywk7nlE+k++1VPOztx8LnC++urwbbdMj8iWWMlWRfcgCbsowGGs6T+n0VvYSDXQ8Ld1XqhNli14Q
ol/GRh4f2rYzSCcOk2am+ErQXMDvTDnCWX7yaww7r4ixPFSbPD/T8pGwliaPng4Dss1v/T4ojnyJ
hXaOfl3kzixxphxvnMeiwZMKNpeBiwyPTwf8A1zZSykbCXYYLBcqtIBZUf0A5yDqVzx+azlUc1Us
Nz5vXfg0S7ilTlSiiU9hvoNuegks3m/0xbNTTEu7KaDVcBmLbUSK/FHlqFEG8tdqROabN0LFPARE
L/wJECoa0YmfejHJRVj6qHohFsTRQ8iBMwhkJdEwNjbP5kVtIKRF63gxRykRdBgRwsUNmUuKQ5M0
t88Wnu0bXCKimNJmBgtBlr1gio8TzVxfi6JvWErf/3SbB9pp29LvmMylKYmZNe1Xw1hkDNiZoznj
WFgdzr8rf4R2IEXZnOWs64TfVe0LNYD2QgI+AuK4jefhdbbYKsNHOWT1E1ZtArhltP7L+PWzu7GS
w+/gPwYg5MeeYEQelHeCneGlYFwqaL7NO8I/nTDqrD3ZmKd8WjzwfOCe6KlDw2QJP2/RAICHsNgv
/tawyq/l6GkB9rYSZLmfExmW1tWh4ktzq815eVzmtJ/IoJZ/XOA8DFQArWB5mkIiMGG3yXjDqj4L
6u/bf3Jgc6DgzUCU2keR2rLBR/4bTGukQh9SK/vs76Dkk5BxO1g+LLSgTu76FVAieeDnXRS4Byz3
Chd5IhlxNRWQFs1gM/0WSD1rqbC7sBelMvGQDj6+D+MJh+zSNMX4nMMFRps5yS+bLsbirXJmrAtP
PyzdIqIXNK0y6kVQXtbe09Pf73+/qQAsAXy8uMRexanEO0XoSKm2JdutoPf0yEPmW3Jp7tPXy57R
D0DO7n7XAOz0wSpNnkGq4nioeYeCHfCa/POEZ5i9dqz041ByKvSI/PfktL2Cw2mHd058VNTzTdN1
GdqeeeXuE09pCkjPY1w3Xtbi5Pc/pjufFCm3KhbatoUGV5NIpNeJy1ucTVDInQbPl187w3mVK7q5
PiD28kYpqYhOXFfExZ75b+D24u9GL2jQ19jJW2cQ/+HYlf9ed0RwSTnRm1MEhOYXgOEdmSx6RgoG
TsW6/VHjx3OIbJgfHdj8TyNL8/ucT1bFxoNQnORi7HfUbhF17btm5n5n53kdGIMhJ2DzDJelnHV7
GR0lBut1BBOLb8XYCPsxC8UTlvAc8tAftH4xJTfppscZhe5pv8Vxsnm0FXa9fY6vmQh7agXEPIEt
p1Y1YzwZj+8xxIE3jTXv8FtUu3Mo6G3/UJvItVE0a/tP6Gn4MBsx+WEM+Kxr0AvR9XFZ+qxWat23
6fHZCf8S5pNhTYoWktn9ACzFAc6Z7ZLeB9s0laR7iF+y7FkI6/Ahp8WhircChgx0x+6UU/9WQb0R
jHorTEAWXg1/ES/yH1/5sMYMy5I5X3NklifKwQ/yUWLZNiOf0L6AL2XICpLZT4KOoZWVl9MiZwaY
ZWxBuCeDqyZeANYSl0kd9ka2gRVjbWvdcc4O1kEJinjIhIeb8gypA+YP3QcKd04nOhp3QKQqvEg7
VkXf3UwYPYPBPmwwoxmWV1hE6cxtwy8x1T297wir5SwlFSi/5D1QyCfPeDpy4lS/7YR24rpQ0ask
ma+b0NRR/0Y3y8032TZZ6R5tO16t8jyBTeU3CHa2/7vftCHbQ8mTpfBA2zrpDpxYwhUODExuKBjm
cDXjqAWpx4A6771Cbyc1rxny2rn2CTi1Nb9Yg0ETbnr0S8JsnY+jxShBUNwfspX44tJGNgCdh2vF
u1Td5DYv0kNgEvS6v4FJEAWI4o7b8UQJ+VNkX9kIk762a8pJj/HPtGz7ijrNUnhpfZpePvCukoRV
yGkMajvp0Sj53Gzo+vVdptM2cEwBxaCjLtIrrK/RZfhZW5PGDH7Gj1SpnNfOuhziwY9ICqZ2XaQb
awWXTu1ECU640V+S3+pcqMSfPan/ffHRTJxsShvCauukF9yD0306FeiBmACcS5nLRPn6kZ0xEQwf
JsTGQABDr/uYe0U1WFCo9AmfRTxZ1IFaH/tK3hdn1XiLLLDjJVouX8y22WtlNfwrwG2R+nCZTwDx
7rZtRpLmvCyS4dtsOoUewW2vDC+9dHxoGeO3tNyOyhX6D1kIie5Bw879glaH25xQDgQfukU58O/N
60mdcj0LiNsw0vMMPvInH5bpbgl2z5zZZW4yp48Z83h9UZWISsRP6qFej/sg3Rvz9BPx11Zz24en
/SOxiC1ajNZaPDMbt5pcSeuvLOkdcrEEC3q/nrUMnYpa+Zjkvz0gxzuVhO/7uXkFGBZcliA8m4Cf
QxKC7OrKW+lKu9MRdFU0TvbCf/38Hr9KMt/pJJFeNyfnmgqK6ACxy8dnINiHjuexDEerAab0fNNK
XmY8b3i5MTsJvDWUHWMpj0AKx+MfYiS8LRDyoF0jx2iIr9zJl7FulAyxt8FyxuLBHYtkCVZEIilV
U0BdivwE30yOmqQjTxmjLxKvGXuibrVEWUaMaBehAIF/S4SJkMVeBpAa+ygitDggCOGBqWQgKnba
9EOqgsdCfi73hCWCb5TyVhc+cG5CfsN9fbZh8k3PzPIjh6KH1bvPcsLWGCTOImLfM4M0zVQDUjWL
9bQVbn1GwFWpu1SKM8AKwgyyUh9eUFK29qkSaZwiS7+AU2MkRw99ur67tzAg8VWY+DRxGChUExOq
SKNrJxxAZEsBB8NKhC1sXyYsAdFG87G5yBX+f+V1UctxtA3kKF8xomQvlN5HCZcWtkDafMbJLiLB
F0bRacKYR16bHnUahl95YHlAm9na3kHrFLngFImjwZ5SStgVxle+RIjtCOEvVkP4K8xFzaeV9lf5
ctpyLKVV+b71cPg74hw525EJC3w384OCcjq1egoivQK077EeJ1S8dP7cHNNrBku68RDoNUQ+fvW0
SA30M+2D4OahHiGGtR/pNy8pThUQJCsRUUL3iS2/nWLpta0G2//rp4QmAXr/8FC6lkbcC6IIlbXk
Phfy0aoLIdM2mKtp177nVvMZ9P/zK0AOU2PsJwm8hhHhozAsbO7Bsz5omq7y/agM6Pz7ihEjdEjB
qZD768bmSG8yzFm0yR4tjSL06pjPcj6ZwzQPTx4rePGNEr2rMDiCQLl3+P1jGz0Vd5ex5/J9me18
icJIyrcffsm94tSqkC6BD/qOBUTi+2m6z9Os5A5rQjClCUMao6JRHA+tmAJfTV6oui0o0vuCLveM
In6/P8QLeYpmGaqDe8aPfjDVR6zhVHiWWmlcUgFucWD9tlksfC3c6hKpbMKqQ9EwvC4oGRjvke09
gm8rY+FcdWq+eJauRcUKZEvpWTjX1nD8zGK2PPjy+TrbzgW3mBwAAWTY9I4Ck2y81B9rk3ONjJpd
F1s5Fatn582uwRGj/XUJ4DKZ6c5RWtepWvpLWB5bDMM3Gdx/1xu5urGPu/tESwt7BcyoM8NzElAu
yoBC3gE1Wh3ibiHnhL2cnI0AU9SDU+V7dq/M2ruO93hrKchEOcfzoEWpYWH169Nt6LdVdi+/3iNJ
M3Q1Jcd/cMaCUzK8Csxv9jNMX0bzccygpZW8dzHtWrtBL5+hCcsl30kj/xXfzKe1aF6YxPaXVm59
44rRSpRdXCC6ufVG1JlVPKYfR6T9UmTkFCARWjbrUzQu3F2Y2uFONfVs4w+DnsOLMBZaLng/s2i8
b3uWTBT6iZip0BDfwCL0AkG44NDfYVIXiNGKDaL74Vx06yvSMlJ+xUsg2VuBeF0J8OEMUSbjEsnC
UW/fe1bujYlCPtLbfTeeHDLuxPO7iB1UpMAIqI+WvOtSd9Ph27XZhC5zeY8POpoGD1zTv3QL2jg+
2ZUUdOlG34F7gqoPoG+2sVltJBBy3B0+vN4y4fKdiHSeoeC6t1SDkjwqBZ0H0MenfEC1raQg5CB1
UhptbkV+HaCWJvlLxA/jVh8Oil65YjJXS2zOCXlyOmDAW0YSMP2VkBAKHxsWgTnJqNGhJiQBmxft
+ErksZavfRdqlo1KuYdLxmlR+p1Dv8aL/XvEhMT/umRpp8bMidGq/BbaclO+K2ZdbnO2FVf1rwWw
i9t6tUcZc67zCTTY4bX45UMZ+TDS4/tFncxNLx6y5d3g5HWCNfYYZgyHBt6FCrEb08eioyVec6Wn
BHZjl7U7J+OReRf0zbV+LVL1yJOu5pM2J7Cp6mxtZduRT5w+EkwB9xFlf/EUksZWjRRGQrPU4yfI
uGcYwXfKEFwo25dIt0PwL8XJ+JqA5Lk5iZINAkIesmZP+5U+l/YsUc7DA9GOS2hGw079FsRy+zot
YZzlNem15wRlI/lgdTB+eosx5RH/NjmdFRpAezmKFL2wA5q/+takRI9J7TtSweiwyP3t0Wz6diPw
hyVWfJQgCTLoXWNSF5gaAYmrQxdq1dyeYvI8FCGb2EIMIsnhBqviec+RE2GEDiHC1LAh7gr+vW1G
yIqmG+4YGRwT/K3M1+sMREM9GGilQsj9HSrMtSe69qdybImYb0I/LisOpX85ke4vcwYkHEwkJfl7
Uo1MV3ii4kW5yoTWBZj+UMg4mUKPT+5ghjNDFIXAstBzANXVMx0CaqR6E2Eadz/TFuCsuzW7ZPha
oJ8wOGJrelfvjTRftNIhke7sHLeYN8BPLnMlSzYu04sHEFW/WgusOY8ER4Vk/e43StVhaRseHqbk
ZB/sMktBQZEm0dOvbvjYtqg431GPM7Z8qFc35KidnK97KGr9bmwAgi6WwyLNeXR18pXG/F0jZo+U
C8B0vd/SQqm5RxryeoG4XbbO5+UMrBQGmxEvGKsgJyLT+6Ju2xdTNKWRpyoz5kM+FzJN2ElANZIc
ysSsp6XR8boWx8d3FAvezeHNTlobgQEveUcU4EikHMECJsniXiZBVOglYfzehyeHNJ4eEbx+gYgJ
6BPIKlqW1dT7FRr5fc1+5jJkvzqaLNgiGMlBbbUC2av2D/Yq6RCwihdA8/6GqBxKU3dwLUXm2Ljj
gbbAgKUHku82KolA9l/VbdIa+flkBhzQkZ7HeLLEhrSTxmyd+cs1R4gbMI3Jhp2oXesrXjZn1xCL
p3XbT+YhZ0BF83Hh1hbT+jhuPH+a93AVdCrKYHoHIBVRK/KOWzcEr0Fdw2Bh8XUXjdHGdRFbaGdx
STeoalZVicW/NA1P71in456bNicp40penKH/RRFqPPdIA7BtLXivsX5+xdo+rzPOeMPNbLQVxlFD
PgXXxBtPCDBe0Z6ttcN4J+dPJfojDufVA3w2W7sqeMg66PBRICPGOHAYGjFfaql3xIw1ZxSs2Ejy
ms2kaMqGglvVvGJWx6hcE3/OhM6qEs6jYRBHm0/2KFWgLhHbg6wCwNhEEv/wAEKWMnXnNFAL9nLV
Ly3uZtuBgbcaxdd+pDgyXNUvwIW8p+c0VQ8O2iRYI5L1WMMQFFZZIEjms1miSBaNZelq7WqRmFXO
EdwSnbtkd6zOBh8X6XnusFcI9+Sq9xBbxuJ9qzzDjqozfyZIgwn6IP3JsO5j57cN+I19ulSx1kln
kBKzGofYjolPoa16kU+dUx3x61xy+deDLxLXmrD4+FkGpdcrAmn9uF2AD1EqAoQPlD5Z/FClYeW4
iWuTRnaKvQdYMeEK66Frm1vswIbE/XAgK3Sy/su8loEYbg/7uzwzhaVe6XAB4Weib4Xq3K/giftg
bzilIjEQW+RcUgLawtAHeTEUku7n6d078mamnQGDyQM7GIy6vAr09RTzoIpcmS1GFn+n7PcLcios
EjhPadUr1JLwMMlIHMs45KxvYtORYFL8ueleB/pL5IAVvXI+A/VlnroY3t7KqsGcBafz0Ehduvtv
sKga9dCXBtgxq9hRaRtvMljepSHuCnvwLgGohJOs3mgFu9jdDz42T5uGlj3myEn7KxcSXmkUe9dp
ma1hSug7iI7UpcMiP79M1G3aKdrN/1L7SwAurb2/sHH8IGJKjGPhZgYLagF/GtM6ZpoTduGTt0JD
Zi++s7Pqkc1BC92UoI2OV3Zuo+5j791p/xcRUY7JNKfB2DFNFZEzxrXal3it0Syv5MPK4CIqHIQS
zw3/sk3Pr+4zoT70+EXd3FZ+swjZ/ekAX1X8vi8OhhodIeNo4U7FDSVwiDSk4DcM5Y2ChqEQ8zl6
FV5vPssPQwgZi4U01c8PvXIhvvyR3AdMBUB5xecKOo0bcrbcFWPmaymn7NqcIvQeXww7g0617uyd
PR22/YyRJ5LrXCv4GQxMpu22R/hHQheUb4HD+xvCqsXv7LFRrRfNZW8eWjfJugGOPtl1Lr9kbt8n
GzRUsISrPR+T54M2+t7CHj+NE8k5zFF3BySMj/hpN7edEXoCwK0RPx+e4yj8mS8YI+TVo3ZLvjDZ
zP6eGXae/LDMreKBy8wTKIrCQYnTZ2cQOsqUrUg7xWUrN1jEtQcmCZulO+Ae7r+F74C69tY64jQm
UKkuvZ0/S+okYQBF6+cfzzRcQfXR1U6qGX4Ttm9xNnAqfdgbHJIHIUr3YwlNlgZu3KFpg0lV3BnJ
pNLPKnPidnfiTsEEAbUmHGm0LfVnwLqqx8yQ1aNYK7+sYyl1lBl2EKQOP1/d1jgpHik+YPv6yM4k
MuCqY0mj0pvLqC5soqIbTU9PgEb7JM3FGF32nUbQgmcI2iKXCQqqGo2CGzYIrNE2KHC8NOhciUBk
6YvJlAxixGQlwIx4vR1TvY2meaHa+jfOvaHD8q3+IJZ/dbLOH5zFHzzQOn4Kqb4JdeIXDKn2uQYz
8Pt2I7H01RFRKowyeaBGJkmdWGno5Xt5r9Po7KqwdttqvFGm7NTp5/aHJUFW8pQ2f4XcQDlg/zxf
ETMx4dp9Vj5tuwMRng5U1Pfz3CkSHGjeMIAR2IQbuyjdY0rhTxJt5y1BZtDzLRvCwPaOzm3piDNN
gKOApkQ/goQuWn72cG3415SfdDro7HcUfInupreCjCs6AvLC/PjDMuMOnzTidn7QYRrd1ulzzD/6
HlCMo5EDgpum6bq58g5MsH08AR9Uov7q5taXqk5w0hOrgZgZaSjzb5HTGMF5SDhKq2IqZwL/tjPq
XVyYU7oZ9E7lZRUxfekpad/SRLkkrIlKlSltdCZdxQAsEJS+RGvaxVwJ0tRuO3yApxiv3SllwFAj
a8DbL087ad4IzB7RCqmkZFMvJeqlhks0nvj0YD7bCE7x6o9zwapw3KsCUHANkHudF7l47ZDpilKa
M19n2qST+g6yCPjDObd3MAs7fKf77vT9TrKfbwQVD8F7sREi5NHa6nG52qrO2jTQ9EYq5KCjtt4o
hTDULZvxKjMw0QH49lz8mAAHEuRJ5cBcc3ridYlIh7eYzL9VHcFRnhQ0yijZh65va0w/44F5kXvt
3FbhMfWBbOCM1Xm8PIxBxAx1o+jci1/kS8ZUr9+Od51KErin3Uw/YhmhNd2uei3eoSdQTWdb0AAj
G/lZfFF/gCyaZpMy3vGaHLCO6z9ogVSjAGVOhDFicPipr9crFgSiXmUgGapsoY2qZfUOl7PpB2jJ
btHTh5FnkMIXYCBighlrYFinvHa6tOiWHs7piIfHc7u3p0BZorlJcbi6qIed0M0MTb8vTARkQx6+
0ApkapSDLFOpR5Z4EnVyOvx2sStlZFgUsZPW3NBnbZUsISgm1VPlGLTpIregQsx53g5az6X/wKYf
3NlRGI/dhCIoEoUGIInvKKPqM0zUdFoL2DJ7ypZM55c/0eN+pcSnCmJKXsuyGfVUybxwraiA2Bbt
4WLWO/BQU7c2uNMc8VKGbWrhql2be/O+dmLcjDzkUJrObd0WLVkP4eQDUZIe30w6joaQzGmJJHJJ
+4zPVylKTZETA60daVLQyZk/gMoNfD2rgVcHfWMMOxGCzNwXj94gknrSEBycCpUmzwKIw9xZpEE4
njRh2ALv96upxbzKHtO896GQ2pCM61morhmGo6gJNW11eQsbXilfv2UM8LUcfi6c0OSvZ60SRLTL
PGPiYJtdnrvZKBjXdt46vFKdXchJPx9bSLUFhghjYbB7E/KZ3MdIBdlvDEOmMsNXFdizZFiYqhIU
hWSJj20OBaEQeQkFS5wOWhm2KQ0B8dEUVX7YodaoySstDHiv0YhVNfmsLZ3HUaJIUC99GHAfpUBB
pvHyFV5paVeuIvf3puaELCCfbRFCE+gzFDSsoyl5mqJPN21WJKuDS0iujUCUjbCmgZSKclUp7AVI
Y/xzAxopSgD5xr4fJRO4NnqGiYHpHOL8x0eek1+AUe1JPmW7fHp0j4M4lf1iTA51K3zwwgCCK2hJ
+Ibp05ZKVhZIxeofHUs+Mz2NdROFtWrcNH3EZ+qeqNiwAlihDRGAjno4gDvbuHpVV1ZtbX4yH7hX
YdKuq/WM7V1AixbMTvhyxsc3t8y7BUJ1Qf313JiG9ifoumQwZxQinOLgtteqoDRtcc0NYO68q6aB
JgxXdrKGX3bmdl7FGKNTsEwL7248heZe0BWoKphl4ljc8UIREdvTymJl4JdpuQHJW2WyD4cfpokR
NNp8/5UISrcuJRucKAvicjIoU5hnU+9ldFGjbGC3D4q6tPmTCnXqHMOFzWqUJjlShrzRS8C7zAxz
RALDF5hZfu3cg32ayraD4447hXgXIKgyNpJiDTmFRXjgIqSBMJVddFMJWn6WEDcI/g7I77elCxnb
xvYU2uMR5UHqw9ueWv4RwlTTQKkbQTnwfshBzGFsxCJgp6pY+9Q/xcR2a9d2FUGgjvIeHEjc4hpv
MPHZMDi+mxwaOrnHrUoA5Y34wtCTxPFXuaGSVOhlb6/2nG3iTE+D2stULQIVXCwzxicAxEAnDhVR
VilVSY1lGfVw9Ju5ViOQGsZwNzjOc4uV7sPeHgTeFvcDdV34T0OYchhr4zlPNueBKA627yJ32F6m
FSRY9TwB0/tKQF+lCOc2L+lUIt0JXDN7kynT1PuuZQnHB0A5SlkdDgHlsxu0QHnZHw4s0tKqEgbS
NlzFiQqukncG7JLxHphFCb7jmqKPdj7/NwOcqcwATtU9CnyGy0ZAKaYmbzOWXkIJWkhTSRFIGB0J
2hK817qLNw6oXqjO8F9BWybVaS5tyZCfi3n0SzU9KDdWtOwfoFXw2Y6NrzKKhBmi1g0QgOd/1irJ
2FfofmKj1YpBnu+Q2b/sqxmmBy8hWPcbK0nxwpmADPK/+P06wvfVuJgKUyLe54PYZmc0izrdG7an
h5jiPBA68hiNMt2cJq51+q4V916M6eVI13mudO71fN/GtWcHdBOdG3JjBa91XMABV3qOreHe2kAv
oT9j52hpA63FGD1n/4mDTzkHsetTXY9oskNSc7fB620FlvaDr7dB2alBaz1lbiJnyKWlS5P1vXD0
4Zmh19WXitmiuh5IuUI2Vhrah9OjrvRgH6qu/1Xy8Sr0cOC9S77KtPQAyukqPlYpokWoNuCxeaLL
1JzP0SMZNjGeiNXBTJPCNMSUmqf/WC/81BcG5YzW5dr7tBYNcNZQHWi9j0HT8AGr8JGoM6kCrIEj
YCikeZpRl/P9f29bQ0FOc7iuwMeIjcR6k8xcge/MNGW/zt56urXOr+3E7A7K+Iqy+yuj8D8Zodow
3q3mUhQkia6n2u7PPytw/Vhz9ex4T2lbrlrPq8udoC9RZPaQEw8bvixQoJF+H007c5lnB+2SfVCr
sZO8Zo2lh+gkJDHEn/sk3qUJbhF98H295WgyqpVZT2qas/FUVL/TpHldgixiYb8rbPbEWy3ZrNUY
E3xtnzkXXCplUG0h26RBkhd6EcaSzBXW037NOT4ocS9/DnIXEi16wwVI7PuMv3b/63bLHLKP2SSj
ORNSgKf6w2dJHfcP6kLhNUeb3mNiPer8yoWhFPPdJm5a3K/fbzrCWKwuEy78tITHEhQj1UkkcLY6
WpaXIx078SE6RwztTivlwcQxXPIT66CxN1cKG3o+iE4H48fwBHBDdJ34EaL23BVgn9WcnJu9tmgM
sRuVHvNkQuuzEQu0uOL95rd6zE2ai36rcBpx5iFCoRLTGSpJGseyreURMa1EPg6tnR1Qe3D6i5hB
luBJzScO5DYPE0sHjqyH0aXNsFP5ScL9GA8IeNFp9iFxw2kJ1YLjop2l3gRN6p/GCIZ9zpp/oKbv
ZH++hDlunFDCbWvG1Yu8qAYn+YdcmrcluVoE/MXmwaMas9BKvGdwj0sMr0Fr2+uLQOusdiPvV/CI
gHaJolk7fEnzYDLiibb8B2W0V+iknCZVIvwd3e3hL1LmUEutwOWL2Ctn/lp+IIc8hGcHq2YxyNdS
okmmMshbF6EXSShIY0MUW0beYWg1+CWxLTiAGE9/vechnhoDO+SkaxceGFBJzRV2dFJxiPKDrumR
0Wjrk5aa5sU1mfcTZGPCbaj/fFT+ZBv0rWaLvTmRDsQZhDywznqLgFJddECcDEswIXoJ51RmbC4I
OgSPA8nZ0eGq7P+r++iC9KA4kPT/mlIGTGpxqPKYLdXS44ul1/J4PcvH3SJzgHX8h10JQchH4Y2F
/BFy6vhVElyKPijMMmPgABG6SCBYMLbrSnjzi1TeludfqCHDDWd0elr9P9QAjyPCDGZItJf3iWsA
a2j3dQ5HkaTNQJoVr2S1GPJcKuo7j35AQrlK5SNzhkkVYcEBS/EmREqw1oMDdkZS8SFSe1aLXaXH
4vgTyd7YFz4jseCp/mIP0QcarzIuAIrS/LMM3McuksCyBHZ32aUiE2R1Q6kIMCDUQimkZdSXDZpf
CXJ1BPkFgNectPm2Lmcx0rx3obQh56i8Nv3e7ffP8kuC48ESsNfQ5t/XJxXRcJIXh93bjAvMMw8o
ehWL1LwNldIyQc3IjfC8Nu2nNOnaV2A8IVuclN9ldhwgr18/hZKGW6Dywe9/YFPvF+xuySY1Ix7B
WHbhLy8aV34f+8ATrDB45lQqxAMzkP3MhEV+MDSOncD9qh3glnGPUc/9cTOvtM/UJ3PFAbiClrJ1
616tJAnWa3jf4J4/go9ssZcxpVup3TgWNP8lUtU9zNQIiPffjuy3yge4Kg6Unuil1aQLpcdVIZIm
YYnDR6yt035dk69bkAujicJlXiufay0H9m3mgzmEFO8k+n/t7cQiVHno4SICDI7K7IDV83D00lpp
zkciOps4IrWeU5RHWQW71mAN6BCiNY+xddbXW5i+J5QZQG4kDSvfSDx6WIG7HrfJlsM2nASLUR4G
4l3BaLftBd3rjqGibEyVrI00NTnPn8Z22TR2zdLWfZ1mUG2YHUKKH2HYkM1NaLTE2pXnG2/nRPGt
sAvPN3yDRCi9PoqK6P1OoYT7C3dVcNmu5y4xfLuCJMHifFBydiTM//RazfTz0bGuG3MJPjK1uBKP
Om/DJjFGmMB/e5Szo5HgaskHDr824sRP5sd51AyD6VSJdrVZitmx/X+0Ibp8/5N951HxUOjGksg3
IcJNESr1zNxBjrXtEFf8+Z0yhUE0+gfJw+24oP6z5armLgQ/dnpUYHyOW2lHnCvgwaOzGjtin8f8
pNGBEQA1VY3RqQAvhBLNrtxddeLbUQPhraTS/bYe3JgHJJtXRTy+idML/MexJcaCqy6iFfEOztGF
2Ch8GO9iVthlMNKyiGaOMfO4mG5Sxv4TG2E2XBl0blsnX6lt0Zkdu32ZzVsCkGghCRh1kEPSbacX
cPv3v+hxWz2C1IIiVQ5VFY2aQrSid2qG++JXntTSMYWYJevkMFjOgNtKBhiqWsvTLFbZJoeYo4Mi
V1vEotPNnnL5FkpavIBSbLk/aabPI6/LESFDP2Q58J6ut5xmOcEqQG2Vj2KXFeUg/NM7XyxLKmeI
eht96OAdOmWEdRzGJr8fS585QUakc2teWjg8A6FuxhvP9ceNmPP/Aq6wi1jUO6XFR0a+UnVaSpgN
qYda2sLMyvP5mCsqtL0nnDkPjL4wg04tbkcfgOq/9G4Gq2fUx2+pERcE0D765ywm0lpcoiMYOtwQ
+GcFve4oZU9ohSY9MXV8rHw63Nks0jDTUhauXdcyN0mNHCFbAhA0syyjdzqSwBb/cduBrUXwPBG4
9zLj01okHnvyD0D4Z7vqbXq2ZQH1IgLwAarGaHDWcDrdk9+p/dEq84MeE43daW9BKAHY0WEbIpkm
zXQ/G6JsJwTmGpAXC0dNJOPYxAGLkz7udYymAVeLlwn7ArBOYSCQKL3U2lVKtmZCUSWjHr8A1xSm
hRSX75MGb76sALU24ftpZ9feUbWzAaIitXS4VvzMv5gwu4edSdnu6SvR/aj+eB3TQIwZ1YL5U1Dw
z6G5DiNi5LBjD+6yVmFlY83Op9JbUehYwNLm7M6mE4y3+nFhj/i/O1+1+oRdwJxqDanlFeOYSLbs
zee6L4LsuJqcC/LVtns4DYg60sepxlFwdjgVHhGnr5JtsGj7TW+srglrqKZSs3LyUw6cR2BoGEK4
yfeTIFiwQhVnyhwSYg/FuKi6waSL15UnOUok/lSjxf/XyPqksA9QUf65AosdSomnPtdjKU89+U3v
YeFjTf231/GGZbSLSXw7M/JCJ3oN5EQ02G+zySr96OKB36KAvEnt8ri9reK50YX6Iz9lEHX5iEKu
AEERBOvExOVElUlvqdgYt9TJ1o7g/WYC+RnNkATrP3ndHR+8nKTfETj4g9SS+jvJE+ufqChooa0k
765uvSfZjxE8Hz0dwJ+iJGbVyfBPgE/SAHUqA3ApxH+bNs+BpqLgKNS44kuIGABvuHFb9hwkVYRL
dLrCoq5BYvDS4Zuw0A+9xeaooV+43FANPm8uGhAnIa6qV/KvfVWPJkL5OwcW3/vNOzIT/b/kwkR0
cXzfo5FIxrBYLQ5XSHE/ZGmufIhQpmEicOUEVcGp0qMBaRolMv5hImohUhtvWqc0wccxTDY+tAi4
NxeBBA91E4Tw7mRLERyxreiTm0fI1B4LiRGx/v8a5whed669E1OJ0rw4+6ODQVY1sJKo41yPh7/d
GGjX+euTJBUAdvV1kWaXuQiz43CSk9/LGfd4jmgTeh+mO7IQCTy3x6A3F3n9asaCssp1Y+n4b5Pf
0LYiCafvapYJ6EjzaSXCh+Xy/8898Rn6LU6ojumhtNv1FN58ynQsC3QXpLTOKhgJaAHJCavkASwg
VzIkyPY38eT+Nry7/OG1cBhEInZF3ofYR/FkF6QsyaHQ0XWcf2Uf1gDYmuHxIGs0cXi8Ys+yO2d/
eDf01QaWu0zv3LZl3mkKEUtq2fn8LjpAvIj7eLFmmTTp5r+QMZ94UJyvU0hwgK9Y9G5vj5mthLF9
ZKPLZMfQQa3pMo0QvU2bRs0ei2n4SqekXZAvez80vYvjuRRiA+XR2NMxlJFCuAZ8iC22BWF7alY0
W3h6zsW4JpoYukGV3NAiGG5nbqZ/4AB2axntzCSJvYkZ5yrOodwjEz2UVXZi3DoqLQuC/zXD/zSs
T7Ta17+t5qZ72iDQd2Io2aa0DZuXfg3PmdnSkuMXKx0cPQP8q5CnvJDAzl4dDpB7b1TUnSi1xtdR
EU7FDklRbT3qsuuW1UkoH57QKHC6+6fKyzKKHun5QZrXioo8OHhvBtcU6dpxDUi7bt8iMR8mCVuf
aWHJWtXkOO/MZI+PpoC7ky8IcsyoQv2YMmm/2HIJXdAE+Q3U8cguKQXzOtxJFcmMBRLy4H2OWhFo
H1tkPur0QWPDZenU6WI6vr5lc+yWDqpV62iTCH+sKTIKYStrD9ewqwhfkcggYYU8QCOhjUnTwHuS
a3/s9SnlmDUWSo1aEMZMDQU5sb6cho7bgoGZynS2N0bfpCMo/BSVwvSx5qC9WnKxMSAmIfKnHHNq
qBlf918e2Js7SveYLIEyFImCYh6uh4Q4ItD/6nfM7GSwyaV8ZDXMiWseuUUUkqdbFE9XoVwH8IeG
Rlnw2YAMOzU/XK8PyKzl8UvFGXyEQ1va80dL0bZU4EeyExki8pERI2epZzVxVkfc+mHWWGrDZu5k
DoUWisEP9EuBoDowXW7MrPJyd8lvh0PvlLvAoyOQsYJQaxdgcQokkN19Zqz9vHBLXdYdbOHkeNxY
s7VwIRZbIIVnY2RohGQGAWj5Sb9w46eHoTwgNP2Ob/eagl7elDKNoqWvjEye9t1be2dSWzd4j0AO
eYEBqedEq6YF+GmR/IMGnlKBuTazHCF8yL69RVyjhQvbGMq+86suRL6LYi7eiyACxWLwvVdUsf+x
IgSQGHF1h61DwAClubA3GFco8fdZdqPJs2u14sXy1XQ75toKaP57h3avGBD0latuGbF0rQ1NsnqE
epkYEiYEYScWfp7bgUNYo3m0twUlsgH2G2/2i3rOCcbSf5r4sFVrjbRuKsQvRYoolBByOzo5Of3T
WN5mZNO3WxyVKKq9OzYq1DN0LEpLalI0MiWCFsarAUlAacMMtFFYMJgqoGBPVxGy/PMFKGmWlVbe
ssmZG1tnicpaiw8uY5p1+LEvYwXOlZHrb/qK5F/EaTZlkSXF+wXBO3od6qRe9Dfqv434J4zXkVBC
0TOiuT3a0zuXRY7niW3kN/aUGRQrdYGKPex5/Lvj+E13NRQpTXCB4UwMFpTkwmxSJXiLblSfdGq9
3AcX+PH487ni+FqXrhKAx2zKiKBW62dfTNQL86wykZEhKV264l4+aD7sYhhxAdae5LIfmQLFIY8r
Pjg3p70ox/z0P232g1mPimDyIGoGpkJQzYg7QNvWCBTh/aruOczG+kZ2WBpjJXh59zXHKWcSuNT1
IKlGUyOOFqK9qP8WCwBOdGEwLGFI3Geq2P9HHz7hFM635pE1z6iwjg2xwzTPa28xJDh5wyB4pIHR
CTbc/et7VeL3+rdOumrumgcm1P3c/DmhKp9Wsd3AWQt/bOzIXOKRU98wa7TwnlUSio8NFzWjFY5T
CUAwySZ9OO7K6wFCKUb3mVwrL+pTZH4VGXksRNzWx4Aeo7n6zG0m92gOITWrZCEzAVQgY8Ew9G7s
W7CrX7QtBIU9wjKtJdmwtoXMjH8dDjZnsHXheLpI89FdGRpigdsNqsUhooaECbuxHKOOVeHSoIYR
yWIyG4XDiHbzqY0ixiuAbTNibDBiAlMkSPd0cCn5Qkknt5UGstYNUwZ7KOXPGFjqr4TNQ2uQtmYp
5t4kTCRbt6muONZXvxVOVw7TbUURgoc6pb8jKaKijvtC1xoEB79TdCwPJePR0qXXFrlNaz0zLAcC
bp2Fna0VBw8DrZl92XRKf3x73gCC62FFe+uD7GkSsdN6rIAKrNkscCJDYveFXdEb9lx/B5oAaXlj
SoKmIFofwmS2FWTtvj1yYJSvE4108SD4RyyZ895LEnV57uQ/NU9xfxxkCad/uPTevbGWRODR9X7W
Ft62h5qftwm6VPeqB8mvouTWhxx84InRAX6UeDDybj5UN8fvFnLgfktLfq5uO0W45cBrpYBpfTj+
HHOwbvCe7XeKhF6LqEhQXDEZfnUDKYdnRU3q1KQozF58ntRhkpyaSBr+PN/qbF1AnsTUpghb8CMu
i0fUfOhMsYukfwONWAH3vsknhV78LTxaVCEPjthJGy5V6y1WfPFNmB3FPso/C/SFJpFAv+h32TUN
SkGKSQ02nM5Z5RL45OBT2HMDjMWE+ZMy+CYDuSLCOnBGrk2t6Y2FrPMEAPO5WO+dXUgb1HGt0Huu
Vgb4AYmjYtZ6/wKmiwsWp5y1qpIiYMcdbUfuL+lkv0u9qDEVvfQcg+mgm48wy+Ajp5ZOqcXd1a4j
rGU3Si3X3ltvkJQ0HrRE6zuYkCOwQMKAOUPY0fQDo01jsqp/LZHUIYwV9Vy1tDbFEIjvmputFc6S
LGVYnyR5bM3yN4nXAB3JwfmOz4dIIh1TJ+20Ix1IFjUNyfHRgyZIDmKX+xo7fcPFICJcmngz+Ur8
CCwYrlpYXvxEzfCtGHcWBsglRjQatwvNsVFGqxVoovi025q4B9oEZ7L78yaoU35890btOzZcjFZ4
SGflGQAUTOTu+7tChpMpxyM7SojrK50/6Gx+TjHQXzeikTFae66tctixDXzl0fjusQnlvQC46I1p
6X0hfdoQOjIsLIh2/pfUwqFKbJCnzHCO2i7w35B8yALCPi6YWom53CpTuUMTGCjXKwS4AK2b3kZf
V7wXjf2Lm8JKPv9GJszaTSxOmRoTNRp4xKgVvnOhhguXmguXJYfmb1/WsFMRzdKGaevLFHgaWScX
3/pdj1kWL6gc2PhBtf4iWY0m17lijofGNBjVWgL3A2gwCl5v9ORxVorsIkUlRMTapBLnQfG8mfsg
UqIbwcYDhiW6NTFD9pvzsuCJFlsQsXRKf9u8ldeN1DmiP1EO5zpNRb2SuF6F3Ueufd0wGtpZ4b37
JySLz9GI/9aF97ClKirbDfe8CYOdqe0JC8U+yC03gm01FpH0L60Y4EHqx6kKuNseFfvVNn9zJ/mC
RuHUOh3TIEQEZa3BUKNbhvdjxjMN7HAbmaPlIdqPRFYnernUWnp8qhhLbE+yNJhJvtkDRjCBMeww
Xz3hQg8TG8v4SOvB9QP9MLuO2AdYo2FFQczzj1LphWeg6tzHyTKoHlMwu102KLZ8nfnS3aklq5iL
boI4rVx9avEPDG7CxNNuYuz7xxIQLp5LNr3d3MOOILMvots+n0E0qk17qtMINz6IP4yi5sCYBFOv
oGtWfWoIFVRN554dYHihDFsPCKfwZTNur5FPisFVc56gpiJFPyZPwlWiqw4WYWuEM5cycWbok5pu
nc4Pm1bcq0mIH23k+yUh9F4RCCiBj9ir6GmR+N/j7alRFqTus+ft2L+3W9sgw3kKZUFI6GLYTARK
1FFFeGW9Qaou2rpmAEjnC+wPgkP7ALJLY7yT6722kG7MM5fpC+XsM8cb3WEb6wh6Qd0qbFyEdAnm
UJeRT1oebilq3ViwC5NPtJl3DLM+gS98r5+JwYFhVx6t4jIeE9geh7y5yY3xeF6LE3HxgVpLvj0u
p5I6dHEAZxMJ6RnOGFoQLAQQuZ+e3U496HjxQIFkQSlNZ1EnZWW4eRSH6hwJ/EsUA9v34Gd9qT2k
CtcaXeVPg9OOmZXwn5P17LGnfhBb42QCPzO/iHG1OoVtrmgcXJnB02l+Mo2je/S6++yokLgBtBYD
8RK+sxTqFWAl/ILKaLkMwop+mxAW3ymqZUZkMFT0HyrenD4y3zJ56bgiGPNOobfqxiyzNFHEDiHH
9mlG5fVM6RcOLrE3IgwwupMMo6rvqo45tEoTaDJsX7ZwyLCLDKDcW1H1utcg8NQv3sQkYQ31uACN
KHEI/2rznPhnojYciTmDuurRBzVQ0bEwnGTR2IdlmSf+7Ok1acxUYRI8ZHo2HG36z6BWP4RMFshl
6ZcAe296/odLa2H3gTB8LFL1Xj1qZdNHsEAWftr23L57KLIF3YxAubuli6AxJIZJmaeetBQE3pnD
O8CLPul7sDOFpxHLwEe5/spMjxWpKT6f9G5aUJx4ekqpBPipvlfgs5w8sBjlTXJVp2qjRp7n/deb
jpuNxW0OuX9ByD+L4Wkw6rfRCDq6OMz42S+IGVd48xra2r0wt3D2QnHypcndovkxh+dU5iepDl/N
qO7KM3KcjuMsGLRYpgcvuiIP9nuEQaILF22G6z/3ZoIxDvcAmEtWguJoPaynkRgXOTqhkzifksgn
+qYQT6gSsxrdk34t934fg0TAH4CqSSlGbWVwxPqGgCYMJ4hI43QWn0KqoUJ7NYO5tjTItC2jEdoq
Fyr9Q2ttYNAKZTBzIeGJyFl/d91lIf2NnvVZQB07I5mNMisborhHnYK4bpI/qOHmVvNuVNpzvIzk
5mgHEvhNmpHF0yXNqJWwxRayIgyx2X7RI9FmLWnQQq6+u1H58RYrU1gW0dMauHLJjuIaZoTN7S7n
8ETuKh6Ev0G5Krx2hNPnt5LcAsmgCuImG6rvZVbDVnB3lJwGy7V/OTsIMXI4q4MC7zSKNTJR8DLW
X/9nARD/zHuxTtagAP2eJGw2ZlzwFcWpmafahLm6CGAGE59ujtW2RgWpybQ004cd0voBBfft7B7G
gcOHJZsFt0AaVkdCbdYy7q4PqwL7ev6zp2in3E/IhiXqrQFEBk5CrioR1AvU2Ic3APnI4mN5f5EA
/O84VahsoE/osldb0Wn3EaNRCuLP2pac2Iq9cfhuI25USPd2sJlA3Cjwx8vBjJrg9i0AXPGsqGyT
1Lu+IbffXB6+48k8uEq6DaoWy7zratoidsHTNlVar77YPQMe9iA68vkAzyYD5jnltTh1V4C7q+BX
BebkeW8fp86aUmnNYJ+hzwyqf8sX7iQif/YmbkXOIT+I8141slxd3ftvuQnVB6hXPYZ5BrY6/f9+
9RnHPRHZj555Il3Sqdv0ae4RZ3Cuuw/3UFYBZhLOlAzRMBHS6N9wE8Z6lXiIhkLW3MS+pF2jeNWO
aIUgVCjQhcUh+Deq/DGIptmN0UzlXFSbjdUc8JAD+vpQ3foNTtnV5sLE8Vg74+VbwXtIHoLcRNTZ
+ZOZEaqDntI4yzCAmkvl65H1RVu/UwFrqC7nJvIawFrZLBb08BLgD9vgtva6T5njqolwDheu0ubm
Fyi3/yn1U5tJe04+JQ7UXWWkH/Dg5gH+obAdkm6CbAvQ0c1KjOsC6BqSUmHdbDgzEKo+c9UuQvWr
ubpSYSceSSthH74uideb8EERCcUJ4P7q5cEAxP4NWJIf9kDu+6C5zWrT/2USSxx6UY4lnKJPRshh
9tL48NyHGBU1qDA4rxZqK14Akk6SU0fZRraxyVcUFiyap4GE2SGrVajktm7A6p/tJ6KPTptere6m
i98GcqJhEZlJyFPCGWRn7W3vfhCxJg4w0KnMzlBiZk1EL5b74081cgik1O9IEa5uvmfK21DtBMQd
k5ad8HDQEqkIl/ZOoYAqfKTwsipEiOJcQRU9CfeId+3A5tnDF0evdWxKLr7GEuI3rPGrUuWQFjjZ
3BquTgVFxNgBGHouqENK4lOW3D9AayB7/gVTk4UYmBVdK2f3NpamnWwpzZJ6F1OsVyVKHyA02QZ0
2dW023NASqlNo/8IHpABToHCEeNO10+erIjNBNJjO65j3Svwto2BTXVs2QUW4sD3JqVziWPdibKD
Q6qA4IyLw/Ot/trfO51J3z4lzc5k2HG6RFEpCEKhcWMO34rtiOvpBhQB8rN2UlotKcAj1xxX1ZiZ
RL+VyqIvVIEaRWUwIvsxJ925wu9t2v2epqWwPDuhzN8v/DyaD2//AwLaSmb1Po8Aanm/saKmEzwD
JLtWbpSRX85sQtYbHPgCK9VuCf2Iut6YcueMf+/cPArDDI3KheE8eVQ14tQxmuZAxfW44jft94BE
2HNsw4VR3ASSZvKNo6HhuwnhllxIKBjzTxzMtrpy+ULx7Ow5XOUZo9EJwbx5DRib/e5leuB/jBXr
ytABDbv2JMQeUM6uUaPuuU21xeevDJ3elszO/ZdAdz8dJRZA746CjUpxBEHa71TXrbrLlkV6ifxA
JVab9bSDcBS8K5ag3Qv7wjYXG6Tl+bXoaxVvc2kDD3+ePgVnRhr2PDWubnIgDL+Nk3nbQB89I/HQ
WJiyDVvDkc5zuvWfJOK/B9GKiKoE7TecBDdoixMZHhKpSEDkkMasHhmT4aGAetKoQN9ExxJTtOin
bbpM//YigbtJenQPPARs2gSsBTjhqAo7qdTXY7sA41l7qc/baisV5gjT+4jJZ96rAe0Qn/7vcdU4
apb2XRfFASiMMYeZOis2wO8yPkTMaysDwfOmlEOOwwHj1WjJk31/sWNNPtCt7okkqXp4A8wcMbpG
rm3Qg8IzItS0jDeNGZAa66V37ovH+DGg0/rj9z+Wjn8dWfhrPRfKoy8Tn4pgbvuChHy3zTMuzBtj
xaN4TqO3HRjG9FfEze5jiYFENZhR0OFxQkhSsgFnb5MhWWlfn/K8BuMeHNhuKJUSFBRYWQmEAhC2
AJ9c215m8Rcnum6TuJcY/nDKVtwYNK0p2GLDU+Rd+UTaNXaLzqekX6iXVAyYAsxfnPf3kxc+ZoGt
azUo7BYaTs9VU7+Evjl/f/PfnLBSGMjNvl2xMA89g5YSp1w6wjnlqga+HJ/adenlXFzDh2jXaq2G
iyacK59oxT7ud4XLx8h6rRDR0ybBsvzsglPGxmrjAZruiiAeNNe41ZjRdpOk5peui8b6Lta2Wg3p
r3b+FSZul/2duyJkXx2u97oH/Ylg7VOvZ+IYDmz3V81rNPBbXc/3jouxEQn3YCElnz3ULpYeL5Wd
yu3WucHRMJjIbgiatHik/K04h5Vt6YDho3eLt3jq/TrczplJWcs8fO/EnWa9tj435IQ20NI+RpmY
BHJHEfVDSTLM0Caqy49ARsaR7PVoB2C1wZwYnWdXT4NwKonh8+6PWIWOAJYRcXYOCFE3ddqgJeE/
TjWaVRYweDFZCYTid5p2IFp8ezu2ailqEhQXEqWjoasPPq0kGwqLmqqEx0HFj9CqR8YwQfrfC6o6
bGBlwSFFYdVHSSlIYxH0kIUJFYcuDyXm6hcoeKNn3PwBWnBz2YHEgBcy4wAGpHqyF01GyDBvpaVz
YYD/RP9gWn0vBYik3crfvbVqqVmhUPnKZ8AD80DkenWiRQineW8vIUMSnTfJWKud9LLmReKvTqgY
g8evnjrZFGk1NnX4uaKHQz4xS5GV53yc66l2dtMULaGTNvHbR/3lfHbJDUrRVeXLRl+pBL+oEeWe
0XiTP/Pvv7HpWXUH/JviYftK+drPGAlkSGmrg6pkp4jqeptPyH/DvT8DspVun8d1PDwOn8Vl0e7c
Z94B5GhxdGB1YKBBjnsLdg3KUC/gGg3G5DYNR7m166whBGNuGuOi6iE9ydMyk3DzMYN4CGhkSzTX
b2Rp/PtHPrkaEus7uzHByrlsSjslMISXUyWmWlhDrqxNhMWJrTaGXh7ESZPw5KRLkPB7UGOZjM3P
Ms9ft9GnEWtXAsGqhdc1J0amLXjrAPcHhpFnPOG6RwCDq9Qu17Yk0HveLJ8YVerMqvOB/S4m87nd
ghEsPhPLjwzS7zaEk++mSIpTbL0XztiPL0orDX/ti/XMw19rTYhe4Kb2Rz3M0JcA2wNi9ERq895w
3JLqTc2MIA98hQMdOo25BotYi8KxHAOBPP9Oekw1m+ZeswHV7AmAqI+RXVH0/7BYDGTybKdHMCJY
5bLRcLwfxqCEhgEpS4FzcShMy1jVG0vq5bSQ/Y5nZ7w2f5OTE7Ndx5zI/Ww3lE968/2Peeu3hxIa
bww74DIVNi8W+kPLtRr70APz3FTVPv+i5YetlVN8DQTefPTSzNpMCDuEyK0WiexoviE2iq/Zdwcq
qCXZhGeUdpiH0cs5U+0Rtb9DAUhuFSvUiKEO4zcSUYSe6WuvnKwLe78jNXZ+1+SKelCrAepDP110
ftJX1h7gUnlhCybdVX4qvEFgvaT0BtcAcjl5FYmHBJVcIjFAZfxzNtfpIFxR/+znes4p7WtVegRi
OIdeh4FDJC3tCWVtpvIhdBY7OMLAVh+nMjbWdvHSjFVrgBJ8PSN4hzUCA9BPchfhjVi90XiM1C8D
8IHKlIXpeM4/0qE5VkbOtxfZE8CZce84InCPb89p+CJvCaCeFs4n4ejTYxc61ZGczG2NXj5Vbn1Q
9xLZskMkNfp1n8thi7R/K2/ryE/UtEMj/rnUhVN2QarTd/6OQOwVNWQQboGdEADdeDO2T+5RKiYq
HkZ57f9GYsUOUMWpz5WcRBkB++ecnN2H0eK3p8wHyfVNT5aYoRwPkNS7ZJuIrKXjjxHjsYTVpIOU
+ZKrodSAJQn5SPUsUb+w326sFSddTCgKhqV3gF/uO9Oj2qk/axoKPMFHBINY4AyTZxGIOnbTH2AS
yeAuWcDb/H1g90q+jEIsWRQWgL5/LTJnAl0Y2oEJf00A34UeCw7v/xJEKFMYbV72F/DIVy3SrPhq
YqvhLH+6sbjOh8kGKXiF8LgMEhu1m7AKiWdjzYtXuIHWQ8oBd3GihFd96EB9qrN0Tbsgl4QAKF3y
DCgSrfcpoZPNC4fTqWuMZZclj3UyV2ys7cm0/uYPH0VAu5QsyizZcwuYouBNPIlz/khP3PGU9VKH
JRpeUWhwtQtW5N3GmXNqqNJ+kjZvgRTS5lDusa9h98RoIn/Go2mvlzDlNV+zmNLA91qA7jynGuJq
yRKodksLkBFm8tUMOX9DpcTLvnPKfbGCdvelp4xkUpbR+bHbgfOsNv0SsiKMbbG/IkWfNT/qj859
o67eXoY1iozRiSa1I6Evz9UUNUV92OS1ROzp2Kx4Bm+zPrFooY1Gm4Ea5FKRzeN3Y/iSbQ5kC1yg
LVRYuZqEjdrqGMTjIwtw2WDF4WlZ2LWUe08YiZvUixy7SIsmySfPWNGFN7eAwsNpV4zCIzvF6tU0
wusbVopJJu1R7vE9R5Sfh5xEjpEdnN9ZD0yBq6LVc/eraDedJQicQplOK6HH5ZB3xCD+7G8zhVtF
oUsjUk25tZH89RfNPaU5AQXdSQQsdS8VTR7QhTn9Zbd+ZpMiv6azUqeyveQVneyFsN4DwspouLGH
+0giHsMqfltz7uLzZl6tuUfBUXhE/U29XyhgbgvsyL8iiNhrKepIBxDJqL2m11/2/BhMIqOy6uQm
t+TXzxvP0HyitIEfn6ReALwUGODUGZknA4/DHijRAAwLhHKmseiW1pPTzsiUVd9WAdkWcgpjsQCS
FTsY1ZecI0vXNx+H56J0PX0r7NFvZKnRhifA0eZm2MFdscXgG5b48Qf5XH+NPzKmcl1OeBsg6hlh
YHHJt5ykyjawqqqVYbbgOFa2kei3fz+SD+0DGgm6uAh1B7Y2dcHCTa/kOlCy6q/iQDpey7O53OJq
LYp/Oki1ZpMyQ6nM3ncpN7hzmskDPjdL81lKUmfe6mVxhx5G4migg/p7cpFv6Hxgg1MVrWcKy2NY
sfp1Nhf8TFw00n0dxbGdHiMks5iof6tmjL2hcItayFKLz1rULkwp/zYemwsVwMDzTr3WSGaBTrif
zElIhjhaOD7DpSdqXHMlpS5KK1LWpkgdAbfdP9hZrZXdyjxKYcvS7zefbdIM0zvSqr5dF9tjCMw4
Be1Zn7OJvbZGgEi3AHUit3S7oyYL20nyqFs28KdCWT//yfYXwNrnJ6CNgbTtodv7wQxjIzJmyY99
4SWOT63u1826u1rxHfLppI/HMh8WpyLYc1uZsfbxnRQcABci3c5Ywm5+7LT/JRmH+6MBYoHF08jh
sy+zLWa+NnBY89fI903DyQ6MLyTrm8mgIET+P2YUOCVoQbpTSMxL2wN2UZ5Sn1pr1DHYPck7kIp8
scnvl+RhO0rz4Lv6Gug9/lvy1WyyDbZkej9rp7iIeYdcLEpUnblYIh6mKuU0+0wLGsqQ9ppE4Sjs
/LV0yTSUsfp079YtWQv/0uQHhDzvEUZxCpW3XunWsi1Dazs8Abdo7E961DFYlrod0ZYdBVqZaJSG
il4kCxL4R/gPnQ9y8L2XOXfl4Q3DLBZz9n4VT12erQlMgBhZdrG9Fj5ibUP4+ipSq8VykAsdqi38
lQxQa5kZG1x1i6UbHaO4ISK8PNGc8urYNpHFVuvo82fDgMJkiIkDTAR1lcOKrJdjIrheJCkQTP6t
lrp0dpsk4NVCnhUS9r6MliYxBMNh+seLNMFqq2k3udxNtU9d2L9jRqFhro8y7fZXuUuHCbgYw/jn
BDqIutXjgv14Qlf0vBYztNZ0LCX+Z6sfFuA3dK8cU6w+HtDRsi0bo+77bLECmt673AhaBLz82SOb
80BXj/ZGkZya/Gxnsr8BrHHQrssXAp65r42y4yYf00B5cy3vtC+Xd5Hr3okp4QUMg6AiiAB7mIOc
2dHI/UIcHo6Lh9gYnWOzqHq8a3RcY+dm55aE14KJoa3AQk/32ryroCblzqTcR3DvhMlAaSbNlPCY
fnruRHcJFs9n8c96x5vgxzaL5FcAZttvG/+UXhXSEZsIYAXav4P+oEzHRSMexM5Jx5eIi5NYUTgy
LU+Uo6UhVXn5MdGg5RGvkd2cyPrbBqdBr0a0fuugEl0y+14dcMxcsBHaxMIE/aB7LV91VdSbNv+A
RH5n/ZGqqkJwZuDYlx0X6i2YnaYFB5UwtGuqfR1GB3FG4AXXJHXXpH/dzd+tA9FwoBOakZE7bEVB
w5CvtNF2MdK5NecU3pfkYGtyvhKwnyMB7uG8BUDSZGOqQVkNH4Hr80rCKls1Wz1C8wx2As4kM9M2
qWBzcReGzU5+RjBZ1cThxTDmNnj89vCifcrPJgxT8pnNTR67MNi1DW34il4+jOmgAHpmWZ3zfHZd
Y3+/7uBq/EaH0PsLk33R1mNzDECbcyOI7OY4l2cNLq8xSnYNykGE0p92wwSAi7xXDbw1xOmqt0Ip
9IlfROaC9JzxbttYrGtJAeMOTxZA/9Mu1DE4JSnPrp4n1rtrUaDf3AbGJJHbyE9RRjLIdrvbnJX4
TbdgGZD3GqzrLj6QGs1KfqrEZRWDj9OVpE6VXdYvlxeZLh+9mjoV/Kl89KDkoa3G4j6+ImPNs+1k
ocCIl28dYO1cyzQmvepgLYs5dU+solcsWaynPJyB1hSJN4ap8hWdu05e+NR7zSFWHAFspx4BcAfb
l03PKA4n19Ofwp3/dMaHocpme+mNMWDWKmcBYhPw29gyxmcjSwsQ10fK1XkjD7kLH4F215d+WXkd
iSFWN3HJA1HOfZ5ng8VmV8g+gDA+WrN7xH5LEwWw1YpwbbfGNHFKM1Mu4BTg+AURBsH5klEpoyEB
D/Al6LN9nc5kf3EfXpFjBT6cqeqiF5IJtq3z4eVoatjnFqDZqdHQCGuNX6eQyCF56G5zmlLdhtjv
94DNssqusURqdhuVqEoMLuSWxy50JRmg48BxWc/qhs3Wqsr8XZy0AxcZjWfFAOH2dztijIHnOHso
rxC5vFZC3jaVf7vw9N1kBYl1niSAKwWeYS4WCl/GUBO7GMPsTmICdf0v3Xb7kA+L9lqPnFlQdiZa
edOT8BYUIjxrmbulW3yBlQDVtne2L+8mRnfZCTvThDlObElt4yWmlnFGed7YTVp30Xk533YsD2AN
H28OHt3CpEYRCxu4mocC4CZ4kKnpKBiVsrrUUESTk/UKeIWppksWx1+LA0/fUkb7w3mqDiw1FeOc
uX2V/tyD2wt7Jv1I7NLAMWs6bMdcEYsMwKQFTZ8IhaG2fhnsa9hkU/KfWSLXAvVWETbb5E6zPS4s
c4sEDlOG9kZvBwE6OhCD3ONfHwLNCW9z6bK1jQd5KpJnPuPN8herkWXitoswFt//m3mmxy7qFoy8
RnpPCMHtcnQMiVvPG9HxSzaiz6Fwfx/AWuo6ITgOfNxKrQ2piB+PThWISwoBmdvulDEHeC9i79tC
UHMTjz1N6RcfBnKHqZ191dCN8EoT91lLJ6x5Utvs4jj3pYLCZHnsgLz/WRDN4kCBcRuCDtNu+Tmw
v+qPYK5NfCmsG/Y47CFCVhQsZyaW9IC/IPZDjKdX2Ab4k+3/m/7exjS75EkByq9MCm7olW84XoFB
8cPWbw+mnRxIQwDwZ4QWdIe8c+CHOSQ/8Bli34CBd1HsVO1avFgWK0+YObDMya1gY6QxwHCWRnOw
3RFB10sg3OV59OZTPiirQzJ6EyOJ4luVk83TombXa4QH02xAQNJC6bAI6YcQ4JfBuGfRymCSC5bw
V/w1eLaeKIKZ25dAeNY0DMkx/rtwXsQfypSs6VvYv2DQMaemgXw/RT458YcvlIsRmz0XhXlFfbD8
q2craxzLAQcGfo8LIbh54A6sOl1l3y2D2ycwxHMlQ/oMWyqdaLfndUiCkyo4+DFNsGvndvcyrdmt
GjfJauFNN4Z6KtvFZUgKNnvx73b+M/GXpCa/IGnmtH1rHkJax989UiYZxxDI7MZuMaVGgn58EilG
c73mTY7y8z0Iy/v9CyYVnuRViTOdg/jFJxo/8hFilF9XV9qzuogh+h8AV+Xl+V7im6U6sTiudvk4
p+VaGbVQ5rT9q6PyN5maUDxNVv5CYuao9RoFjPjfZWABfIJxjtm/H/fsPRWGHTMUxi7Mhxw884+V
sFmX6iD+oCorEK3mwAtTHgub6H5MzoN6VJdKvD/TTq7OQM7pBQpP8JwYWfz/NcBALSCi3XPCI54W
U+XDQRii6kNFg5E3QpA/dOBAuovYA5/smXeDIlQ55Fep7T9RXDmXFNl5J7RjkT57y5RbjsPwGo/w
aY9fjwWOl0DV21aFRsmieP6XfVRy5c6Gqx1TOImYHK5HrL5D6C9bAoyoLroAbgrX9zquqlzo8M+d
eL4ilYxEMKvoyWXwsnQ6r/Q7Nec2kLd/Ad6RbVJ08jLrkqumK8xeVyuHBHKkGW3n7rYfQBj7nmua
zoT/ycdJMqN1EnrNBoQovUESh1IfzFLXHpKk3gWlpJp0UdCR1OGLBC0yHYLRMpmP83Q1hnJHTyH8
PDv2WyFs3XCqqYj+aooVlcSfM+843BPIcuFEdnd+z248p15DwPQofwTNeoA9KTt16lbX4Jq4uCRt
2mFxkm7BcSbOZMsvrTmTO17Sw4/ckf0NIBF1DxgcxaRdPxqNyAyZ1TDxbdK+cFJ7hSR6hfomzhy3
602wTSM6q5ODGZL9GyFuUH6pUGWMn+Uuw0nSYoX/4Z1fZChqVFm7y8khKMZeGKnPxUqXKGBzLxlO
/5ddePL84JZO0K7B4X730b4Riuf31Y0uyP7N8FnyPyPSBnasMSEqKjmTC9jKOasuOm5XaEdQVG0c
WUW3f7ojwPB6ip+uBguz7n9YSjJ/+S9XecaQooOPxYeV4ufBL7nBvcHbC+GVLjZjThgGkZdaCkza
WxWw4wwsLngXuPlJmWeFy6CdDtjZ9SRjTmhl/J3W40UFzfwV+Ph+ujM5qU8tA7zm9/0Fv5siVgw+
+Xs7zVNd3rAr2gq6ZaVQiSCYtPEBWcpkyqch1lQ6X4pCoY3ehewF5GfEMntAenNZLX+WAfmGr5Vj
FfUZHCOVd1v8+XjKKBqYBsXyYN0A80gakYlC8pwxUQJi5nJYl+CdnNirhpGCpByQZEq99CXBJEII
fo2zXH+ZTwKS7WlUO9wNEuXjhIDYWVnGpZQ7keLKV2FPHiePYrDc3G4j8A/wmyzdlaAI+fbnZOfa
D/rTgxOT0kqPHQPMB0jwz3S3TuASLRyZJfr2J3YLuAr/mbdGkvqJdqQiBMRvulXKITxxmDU0/ZV5
f0DL1XycjROnYSN3G7LCWcapMxozB9mXWvHc5M8WuEWlEYW7LgKOLmDEPQxRHmUbl5lIFkoj7IKs
kRo/2O+UrC+6F46HhNr4lTgqTUmWwyS999KAhRE0uDWmEuDzqWf7dDQH7si/5gNiRUnfdIdh+IoS
hz6zxfpYLzQClX7BpE6s9xqeNuq1YjcKL/iVrpF8bKKb2rP79p+GmUa0lzCy6h7IFuF7X/d8CimC
pNY9TWF7G3+4lNOrryPmytWbC/ZKx9qUl7RlSgH4dLtVxYQqerstndyBXxVKuWcQVENEiBXLYNst
qzEKLP21bGwfWk9ETe7k2iRSrd3pxlzUih2HWdu1U75MrnHsZ/l+kV/UCqRKzbvOeQdjdhJ6fFHg
zDmMBlp9q4p/j7iRAqTEawzwgG4h4RtvWSKdPxfnc2rm8y+biNTgODiW/m527AThySeE9SVCGbXZ
7bS3cR1BV6ilXPhdyWaBI/rbxfwydsUsg6efZHPDFBdD3TndiSFCTuPFp6cM7TnGlGnKMG6iUuTb
l/hsU+L44GnCVh3QG0jtfMDbUZhJFQ4quA/bvdHgx56ztOq2AnmOeVjTBr9qulsKqIrsS4sPM6tp
YSA6xWmirYMq8EA01h5C+J4/tC0Q52ANUltyxSVO31Exc4NNK3lSppOYxbUHC5fQewZ/4wMGPVJv
ka5Pz4a6ZMqYvv6pi7rTujw3uh7p5CTsruGmY4AQ+jNhYVURoS/1cnFFNb8Etd2dqVmVOikl72Ct
I0wwUYMKwf4IkwuvcXmSHa5bl4wXxPl1xgyMTMkbo4v5ovnn7OB8rvjtWPhiqu09FEQPgAirvWGM
NTWdooN0MzIAMQZNxoQxzQCpGQ0BTk18w5llsBdaeillV/Yerj8rd4DrO0C/gBKqEC5dHvmHu+kn
CbwLIT+TcD7JvEKa7H5Ww9yzi4R/0MywiWp1w+SNlm46+bbqcMW2Sx5Nj2QwoVsffZrVx/J7wcw0
vePdVHckhcm4elgmX6AjAy5PB/h+WSMizU6E5dhEBcrlslYqh7Mj88tsRKhHMhwn0bt+ipWFOAzo
R0G0+Vjs3DZmFXHm4BCy9jLDg4mK3iDGGVF4Ow4mwRpha0WgA89e/QmrVtLZ1qdbuCSiuwpx4lpB
r8d1q053y4ODH7zBvUHoz8MAXunrQ9Rb8SA+RcsUO3d9mm08N8fRpiGQlAMAAd4Y304+UxxQhPpY
nk3/p+RTlOHe2IekW9X6zExZ9X4wegIMKB57TAj0TYeJxP9qaEE8qF3sUscquarceXC/muhxRJhc
+WpjuQPazCzkffZchp9D76e2o8F/eaeGBMrUfj6dK8TIW9L2rjFM+cDSA8trWssnS0GTEODaO0KT
lYR+rr0nrJfEs2UzyHWVAeMgT8ixMf5kTMlnwXLrJYqytyCI6DOV6O1zg+ByGB/rN59uzQtPxOWI
FoiUV9HKs3ezBoy75+ReyyPN20cEwfS6NxhuWhkJ/Vt14c1hjTReMI7dtOfXs3jCrSDWmrjQDDhT
ZWzMWuGq1IC49E2Sj7lEsLyUNp+2goAcJTXWd0Vr3/UQfBDrMubOapbq3jZD8CsE5RpTZqM8vJaF
biuvRT+PgVDU9pd+ntpexHXuhNGgqVr9/0+Xf3GeaPSyYZxc7ptQ6qTs3mosALu5ak1zNn54e4UU
zQT2Kb4cOjmCSDBgHiubRs9qUMw7Qaz3OX/2xnnEftNjzn21wiyG+a8KxNyLExz5CzLqZ6qZas/8
7sWF6/Cq8v6fKrJXvxRoz640WrxyU+OdQLpOCIfXCduVB9FjHI4ee3VVSDZ1mnlAQs/QRfVHcctL
Y7UzZZAfxvOxC7UbrhOcNRIcf6eff1w/zXVZqSBYKCTS5Jcdxy0B+u3hLnqjFpr501CRRL1PxJsA
79FLYxXyZGPkQKP4Q/X10gamiZP4jwa/Kl/pxMX4w1E1s0y6VjVndoKnCxU1V4y9ZZdRpWFAYz+6
XC7pmAbZ7M4iHFsez7mNBngZo5lgkVavZG+r598VfRVaPpzlY/8JXXiAu+IHnu5F6Oqi4jkWx5VQ
rOFHHgQQgK6YsIjrBNMmEAve/HHW91pEjJiD/RrkAveUsy7MiHpgGFL+aGXF7EzITSP1Crc2Uxvo
JcFjw0vSDiGQ98lv75ZFAe/qEn7Wt4InnOHHYniTHn5Dz6+4kYOtEb96fGlJ3EptrJbCJ8NzA/9S
aRov1eLaOkN39JJZMgMb/FD5HkHxcUVMM/dqZ/yttC1ZqtdHSd6TLTFnzGV5sr6y2y3y/D/iUf/A
kijIq9L9uLUWjmVsU81v06mkpyXa7xNdeabf43N82ZpQyYvHFQi2BM+1iUm0VV3gV9WfhyAHiutA
0kMuiJWWygWqGfKsv3nDkQV1ek6AW39yCKyRhnDZfWMUWkr4h2Wt7s7BpZ2HL9HoeCTRzqajAqVw
hiHu/cDWW0VHYjQ5BCJU5MQ5+xsY+y9SgUYXIiECi5dx9us59DZr0ShsAeDeVD+/ajw3diBJM49t
AWYgs4FnjOcG8r1QqAjCYwQ5mnawCzfKw2HpE5mhwyZkSLhxWD7NKseA+Lb92xatlynjZaJonMKy
IWU9ZtAq2AUnWnV04ivmcpU0cZCAD3GD6+TfRTBe6Ff4VWpV0HqwkMsHFnqHUw361/6u/Bd3Ij0g
K/VofHSDxpE9byV6mBJoLshLa+qDsd+gGJRewhPVbsl3xrYTAyIxwAqffO1QiQGA8A8Jg1oXKZCL
AXehnVrqtpIN2mQd9abE4kvYPNj9QnbXzaT2HMUH1AJ/V2+L6xfyFgSsT4V6B83sezgxGgKPaEqb
MPvcCVbgf/tzlsw9cFqxcXANpHDFpEUZrbpX8J/7uh98dCHu5f+9t4TdNiPNFJUS9Eua+mCtat8E
Vc9gWTtLkPSDUTOjhE6IiLKyIlBy8bAdLy3DOpHZ1GOMZGXojDqsiU7L7u2T5rxxlrH8V0J5rg0w
SXMOAn8BH0KYrafT1cXBX9R509oQ307PChUSugL2Df1AZTWdWOuVqcBJmbkFF42/7C92IDgVg8WL
pxY67qyzKF9tm/nFWD/olDboq48NzZ3+yl1RgeeEWam2NblTEV5hrTLhD27UIEc+5d+r5+Bk/ey9
jLV6li/C2Ac/pJnkgv94TsPesTrzsjDClnUp603l7ieUuRLUtKW60+/DCxb8CnnpYqGHCvtPjt4B
HKUJhN8yiBhTJpGe7eZhdBkyvfj3s4gm+BE+P5JrwnKq/arkvh4DnbecZ9JcDqoGiXueY04sxQ+c
u6eAA/Ke4HfdQzeofzRV4CDx3DKwzvFsM0JocxAzik5CU7efrLMBIhGIIfQoKvWPkgT6y28unvkS
cvPjkv3MYK27I23pBbVbyQWh3byRuKnbdp+bSOmmBFrcgUCfoobhsaQOQ9BkXAT0J8NL8V/AZ1E6
U/r6NXOgZbMwy6tDFvnOuCUEKwaZb1d4yKdJnxb7RTeHqn4G+OV1qfOfH0aKwpbWMWt6ZuhKm0SJ
PTxHo37FX/YI9YHuUwjnx3fsddTFlawr1hPN//Hhtir5Tq9ta/2uFTq3GIxrRmTtPcSNyV8PQANV
mHFxYQtyIyi+he/hViJifTEEvkyvOnQa4AolmBL8kTm7sR1TeC944bOWCRY1iAQp2lfqOq5d3tsO
Dv8/72FEnO3zUSdVy2HtKe735YoOYIl9WVeLhH2sntfVmMFzTMoq6DnPYn/Wp/SiinU1yxFzEQSu
EHDeJuyGTkuxreaeEahtY9414oTxxUDbQgRTUnIXoLMFw6u7Qv2EJG8MQlsYOswzdOAla1XZJjF5
hT+MkbQsQIKPPWh0M+fu4RPwxAuGX8il+NAktubuZa1H8b1nruBEYheEUm8oT0kGlt69NN9Fm473
1wjR6ENea5pzk1sOTucC+axOI7pkxxAmJpxdKVwnriQKWdlvO9b6mvDR5XbTrjrBrfaDTV7oPRoU
9947CKw+W77q9bt7tAOdg8LKWk8qr08/DcK4ZWF9ev/21giHBPyX4QfJMVZbAPHaG40XjWnJYo6U
cN2PmIz6X8wNrWry+lefIfi8uh6uQbQid1tFdAUzN/vJY3d8+vDgIlKdaEbAivCoLOwG4o5He9YZ
tYF2LO2Jjr79JZLmbR3CRk0VvMXq8VbXmvTs44YSNhqn7dU377G63PWb6YXZ/+wvL1yG2B97fnjH
mmRMjH+9y+DSsfAtVuopszaH3tvqUzWAzkKmTiBmnZA0XLZXPq6HnEu/+jGKigQA8SR+/MaMmSej
dlh/Ftiru//1YmV9o5CzdpVYrUcgNX30WBmd+qTgltYXMB85e37C8Lx+HYtjSotmmWsrzgPytRTd
vYOsXGwd2BCX0uyCZZ/N6F/UXr3xUuBe4GZpljEeIWqTbUa60KqRyhpEtOX9qRNN4uwy6uhyw5Rh
IjbTXYWXsQpEMwz6/Rr8S9IxxJd2G9eNINZlwqWeEmrb/LkFD5AlNetIGJ00JRU0Jw7ncM35Tcd0
tPbg/EjFyqyf/Rti9Zu/dltfkxtjZywJNWhQHZDqKG4KxSUh7PKRF8ikJIXZlp+ocRdJzlZtq4nu
/Y+STOYh25j/NLJwm3Mn/iZRiKe3mtcxJfMtvhpDLFB20vw82aOK13LDvhQdr4d6j49B7W++km9P
XLIvHIpVwnVJNhHyVuvTjg0wRcbz1WKraRC3m/TTsSNOpYdjZJDPpKjBK7JnoTcrQZt7bFu1woYW
utenW4CXkUsZxiZIWdBxFYbVaqMUzHCcxSZVzDsL4Qu0uokm7c40BlY63JlFbdcrnSw6Hb/BdDcx
rMlqawoN3Xuduc8NKu6GvSX3cn4Z7PJJ2FjK9F/+C8ASn0gOPGcEBvr+3HKCM/6+NghAgY1DKu3I
NwZpDYFT76cfcUEsuSXaQzvKshFcilxUUGbZx9akAHO1N1jyDdPuLpzURX/Ya1R/QZUzvOdxE51M
h37PIIucnNYQz1Evo4152Adbft7CcamumbmUMHNzJEqQSJvkJPmXCN4JmJIfFf0MzwMLXQV6K1oi
w4kRWA8ZvORKMPA5t30QKV+RXATCVGQ/lsLtDUCfT6rJWwwpXqgE0ToDALkGqAo9hAWD/tznNrpR
CM9GR8qMkjMURCKutk+PbDQFnsvvP2ufVEPEl7jS+O9R6IHamdhV4LoA5RNISonl3hV+c6pGf5RU
rkeTsC0Fq8gpWfR6tMGkr5iT2P3u+/y2hkBYje8cp9OW6XvEw5gP9BytfYdlMAg58N6jgAKB323y
wF6nWDJ1eij3n8u5yx3WhsWN/WvlKR/g5Es0RgFSHdqVg/F0T4mXnZA9LRv2Sbdfp3GOkyw6ES5j
3rdUFFiec/fSYOaz6JAHYbFnZotcsG6eI1e44KEWw6PB5BRF0Fh+Z2FTd3hR6uFdTE9IdNw5d3FQ
YuHMl6zMf6RKaB+Jy3I0iuofkbPeVxsbcLDmO+V0DULzwKyKfw064UE3QrgQQRmYdyMt032Q1P7F
pRQKiW8jtJ7RCdNpVu+mk/rOxXTsP5EaSoKt293k2Osy2IiLvde3bv5MJrSWKWQkLQ9euZFjLe6P
Bg5psiM6yHZpRUYpmi7RjghSmXsogyo2oIbGrhZ/2dp4+EsSBSuaIXo24w7rAJtrFBw9H++/qBGF
Y5L9IWn5rxWU1WtItGd6+KPHiOgBoOqOu0dWMsimvqpW8/276r5t8erFsM18HqxxpuP9DNyW4oE/
ntMXkKhq5m94RC1+xQ0nHz0nSXzm05KRFrG0nZuRQukKhyEKdL2CmVQot8qo06Ob/l6ItxNqhNRc
2knBS2fLKJbPBYmOchq4NxlM/2rUdSvFvGKyVP+DMfboQzbNeSvKluEqM9i/vh/jKQRyEYKPCOxj
FbzRC5wvHlAU5NMQ5D0hRahZzBEq3AEC3/0NHDBpsxtPg9WxZQlwR8yhptZrl6kvMLkVW1JOLBQi
SfHPgB9wWOtqhlMzToaTc+8f+ySv7ClUUWmymRcbMg0LrnAAKFDNASokNjfUfAy09Pio0yfdDSRy
OP2qYWWoiOqZGCi5XwAqN8qPcoipNpmU6nrms2tfx/XC11vjxBp4JHt565+6fxfkogLfubYL5VKc
svW4dAQefxnEDlf7XWG13Cakqhr1164OPusq8PkCeHAAMvIsOQ11tUNe4YAmVpODrUC960BMNm3O
VbChh+AMQ9+JaBfPz1iSKJQXg31AHlA893NfybN7QbnLrP3cdqIT7quEGzm1ue0nhk93pLTmvEpi
Ncio59DbCBYQNPNCbVfFsbKHJc3toCuFZN4Nlj9R214SmPgKdpZjs/xAL/C2LlfDeNeNmGnCWjAs
M0lk6TdCnuUEIA5a22tx0EM/hNwenCrZcFqSGA5KoSlvzry/+ggEVYCgZb9tGeyDZPFWE34eGmZJ
wY6eJhId7cUE71MIGJVAp/r/D4J/tfIUZu45bweMn0rwAGeuJh5pf7+O6zFGA6OugZlv4E/A4t6Q
WSpZZmfV/qJCJWQpQabtglaXe5Exi+7tOVEAOZPnJmzAwn9Uui5ImqVTZg1LVruYBi/Y0enSgcvg
j7PI1roU1VM7NwNw+eyvi3zY+Y5YR05dCq9J3BNhXa7xVTLN+05oU1AHpmuW9gpD7wkfiNDrDS8b
y5BBzBJJpzJtNpfmFvEQ98Qeq6qTcg/6z7aHqOsapalPo/Ag+eOEqVrH3YWNOoRqvNO1gajbjh2s
xIzuFLPTXugNiHs1MWNHCsfTVk+tdCvkCQskMGEIrL3ffPdKtcdKdph4KA3E1aEmYax/iAdTn+aU
0XvUsFHw1KXhEhnhUbTNyS33r2tap2H1xkQHfEVks7VERphcXUaYkfr0thUCR3ktFB1c0stNrIIj
Hvk1WHu2A5d+4/UDpAuxB0YZOP6jWWldTQiQ6mP11of7xH/o4GbLkCGpYXd2ecilyPU/jO0cRWrW
Nei1x3xolMlofxwSYU3SYFp15ASw9K5SnJwGURljF7Qepn8YDiiWAAQgMfQpHD5vfYKNNrC2Num3
kWKFmmQoo5Tr+vAaO4i5cIQCtDyQPkkddeFbkvzH/y5SPZIUQyB4uxaGczWNRbnerE4i1zvUwSzz
379zVsJeNDvFLppngTRPw25ZuzSALLb90nPA+9p3o+nTLQTy/Zctke3iP0ixQf8yjLihLjMAGpnW
QPEikgulAzAJQUzxLGPQBsdeZHaJxSdjl5Dv5Kbo7zkvBSvbRwBNZ0gGajUNUua7gUkbJhy+ps9n
A2eMcoYTRNvJaFKpO9MHu4OuJOPkkSE0TJIho4fPoLLUa0LUoHfXLdziCPPIl72oVvKsEx9RNJR8
JxGcn4JlK01Z/ipGi2dbn79m1iTYHguzXx/QL4g+0PqS6LNuryoMLOrodWMf4t5lgqXBJ2NNB0I5
xop54odaMCXp8U3HfWNPJuoE5MHOIWLIArA+pvlR2iUPiTEemEsWiRDBvT1/YHOQdRByThfjSyWP
z9Z/UXEldf7sfSx1qYM9Av1itj5342B7lvhnV/E5EjKAB9YmNAnvuqVt0LDQzUl1nxvJnZnuvElV
votP2em4f5df8I/YW6KcAm7TbnSQ3iLY5jdPYH0V/1T8pT4pY01EtcV2RVPNWgSI9Ah6YMClTvpS
rC0D1DD8hdXcvp2TMaBQMw3jB8epV7tBxsAsm/0CFeDiiu9BEE4BKgreCSujghJmOC/l9DpX6GrE
uBAdXh3lBbxrHckAJFMkpMOlEm5x5IRW3lWZGxOqAVypkkmVLvdwVSAFz1cdMJo8JcWPpJc8bgMr
HjeRNQwD96NToH4P/u2Z0YmkGpu++h78p32KfY3uR/kVpInfK3kkqB/gDTcWBD1a0kWzeJhV6ckZ
U8hPq4lyllJZdU95IxIFfFdVXei2qP4csbolHKv4tedj/jHEbzhIKfpEK0mjwT9ZH4xgYZR3NC0U
+GO1jdZaY8uOCxpSyMQc9j7H7N27IyTtvD6KeSSYhp60G6SdHOQXvo95pDOMaOSv8G+EEFz3/psV
FjbBNREJndt+f5bqZqRXdozCXnIbQQygNanuznudlVNMCXMsWCiGHYt5PSsLfDe7m+1vBLm3iVju
xbRavwlCqioCuLR8HA9qXY0yhvw+6RPkPs0OTCVer3b19eoDIlSzP1gfAnQMuAesmp9e98zckeaJ
P1LXjXvaqeUzWalRLzRV8HT/LDgo9EoTfACND3ydDoH6y9Mva4aml+GHc7dV6bnVTqW+16I2fxac
maSjdjwJtlOgsn0/bXe+eVU0ZfUE3p1IMr+ZEi5ObKilNLoidYqQRNm/aouZ6tbRWozJ1yo/mJKY
2Za4zKZGW3nPwqdVJsfvVREwNYKVm8+kV1VUJGAyYPwaFyhroTd3jjGSzYjynfmrOtuQpKVD3HZu
kd0K4nFJybTMY9yVFp51eUkiHbx0sg8nDgpLPE+VbJyrwONaRCc92Ya5MDD21B7fRNNyGHWLmDWs
7hc69USGYp2Che0SjuhhaxCoshazDuXRrmorvILtIpzW/8Uue2kMYvQS8UL6SA517LUP4SxbZUJl
KoYhPwjvwhT06Svcu7hr4mNQL6LnDW3TzFRLajC2VAgOb1SCO1M+9sSzPRmfHhV4ed5h/m09v1OM
Lm5o1ZiFRWXb4m1BnBEXQ8cBF+jej0LLB+BBc9LSS7Gk98tuhiWjLrJyhKmIoyuxjYt4OXdNwLxL
INh+dsqBx4fBEvXPZu0q2ihidsotvbUQJLVsISWf1g9sjqKuQQ3gh+ySa/eipIGG4aYIcrmp5rTs
qS0QN9Ez6g+BIGuVian+cGHqZUPamn+drF2IbqoTIRolqiuSgZoIhNzZ4GbfHdYckXwLeVpoI87L
DvI8mo0Uy6zDa07RqKJyHl3yCROSz+t50n+kthE82k+9jitHFlkvEQNKjHvGjC3cs9EAN6iHVf5x
o1b2Mbq/bkP6VfqZQabqjxWdm2JGqwdPNrhMO4/FrnkVlUE5tGhUo+4hmPt+4BMSjpvm9cVAv4gM
ttpjtZzpE3YdpHvxd120YRksl5KTZRYm4L892w/3xtbOzxEI5KJxXfaeNJagKjXh9W/Vmg77FAMP
zTiz/7ol32veTsQ8PWcLK0viEB4kJ+u417Fj3YZM6yzYzjNxbK/0TiDMgFXvCqrtf9mYk3h4V51v
ze/Fc9rfVFUTsdD7zrPAaKxWH8XkMTLzEg1lkuWnXnP1QtUxOWL49Bm2KEPRbDZgeUPWBYWmYVBQ
ExBufMB6DqRNkc87kbm8jjaI43UqnW6CbB889IytW0LMjgOZPEvX3e6PXofTLjxctcoeH1otVAfs
rDF3ceOtWvG34OIEe5qefJdjbjkgbCAxfkzabZrYlGz9kpevBKDcGf/GkP64YEyuuQKLpk6jnZmP
mmrnNze6sRRyXNOGSJ/PCBJa4uYVQGfZwnyiSS/jPAs3zSDejc8jzvRzoB/5tiVBeHsvNYp3IDgc
ppmRLfo5vOBY8uh7z026hQtr28O8EV0VVwZYXCs0jDFqRjAnrCf4QmBgcm+kCq0X9WIu8gp8Fmx4
nqmd7MtbNXXnkTLd/aTr8fPVVAzPUsiCAg3zpVboRroF36ggar8xmJP1HoMimNlOJXAQ63oYLcP1
4dZm4x9igRCg6EKLTU11Q73mXJYuaA0IjuiNZXR7Lr5OnbLRItih3f62Ygo4X8+m7E0CLjXb+BjN
Gejhmjqv0DcB75I9+4+M6uHNDPpY7KbyL7VdkTIdY+eWa24BAnFzj3VIBdJ+T/O9gOnNoJRLW/8Q
H0rU2NdhylhLe3JAosixzDFSOTsEJNYBcAbAkPSKXU2Gu7HvxUedIM/VY4kp/tWh59yKPz7gxLuA
GntfP4gyKmW0iFMx3vqe92OKjU+71AtXutoCAe32c45MnNbbm/ufcDR/2xe+xv5sDjEZ9+IJreMA
CWkaamS/mG1rM/T/6IHaAamao/5j3rvKsUsy+iaFapv6JxnWZsV6yg7PaSKt+WFgoaHX91LqcSed
X+u74frPHg7n/uPL7mljhdIbB0PZApFMp/poI+55PNsYb9OuemMCaneOZiPWni4DuSjshunsWDxu
mucHJMEWZPLwvCtODapoiUhrI8K9eH/5Yd/wB8tm2DpG1gbDUhZuzTG/ezC0suA/Oq+AhlHr+H5V
I6Gi1fYVqeNJy+uYysK2bZ4VjEyRRkxJdS4K8lLHpFH5jNOR7CrWVbkyG4WBnAG656vxVx3SwiL4
YnJtezcl3vX/ibXr3RwQ4QwzewfhMYtyx9/d8SeEeLMbl7G0XgeI9MI/l9hvX6TGYBwUeE3G0t5h
8vZhSR3XOj110ihEh2txv0Y4oKJQh0gZWf9FhT+IC0uplmAp51voSCDd2jNFe8Rt0YmIjVQAyzgr
ndupAoynIdJLma1ABbqLiWnx4ElxD9a1zPgBhUKc72ebSyyZ2kAXOI5TP0Au4BbhRyaapZHPZtTb
ZK4tYNIoKcY7MljVJpcajhXPcWOgDzAUCO2G8kF4TV1eMbmQLFeTeGwMOp8yV/0+Fnj1NA28UGVR
GQLP0hwWY4SUHS9sI+j6nCe0Yul1+yQzP/wiefmGUjOVoj6sNZ1U5+7s8YlxX6cemZbgtlqe7KkS
QmrM6PKneRI3BZU4PrQS7mX3cG7MAFJqqy29v3FGnzsnMDWMQjELurUVtoN82NA1OuChFECYSQCP
BLeG2oPOgBlguDnLtCt1NyRL06q+BSZKpX8w7Ei01lifEt/PEHvvWjdGULAk7hYpCKHPpEvqKeF1
7Cdtv7sNzT8UVsQLqiZNXtj/L5tsEBQ66KUstDo+s5Cz4uxr3Qih1ujq1WAGj2PM+724fBygnSmh
LARFLacTmnVhGJyBf5OEQ8at5aKveNJDUPchyo47I5NYVSqO6lwEp0xuMlL6XhG72NzLKVKP79kZ
s4lG9Uq+DCyX+w+7NAoRqe7Buqw59wjH59KanhE1VbCLWgEZUkKfVDF4UxH0YiBxPlSsb5BuMYxs
HnTuo4e5Q5Ntf6N9kkzyqlw/p0+gohAPi0TBYzrVR3wqGx9iZeIIiPrpY3QRBfM5ozYbYOT4cisU
y8eES2pp6q4FxWIF1B1wlGh46gVs9hMP2m5vFiAH1z5hqDcci5NaS7XtWxGzOtWMr0igARkaklnu
YkXmWZaRCgDdJMOPIFJO9YfT/kyBarWAbRAUL9NoG/9gm998FayQKWUJQK9HsVOGAa6PZ2CRBb90
yExB96rtrbcidv0VWaTmAGKqKis4GDw8smLBKhQj/PnKVh79XjUZO2j9B/rJftZLVtIGIW+H+y0H
DMh4chS8QAN5GqGOvhcX7WP6tRNYVcZmrR8wf6R2k0zRFaDdeNmBrqhdLtf29jt+rZBoNFJHWnx2
19wyTG7fydaxph2X4sO4bAEae2ZQYvN1uaVgWLZBpqiktXz2JnJMjceRFqWK3zfnR6zqeJPVHLjN
Zh4OeEMIEAyrZv5BhEb5fxD/XoAHSrcg2/mTiwCllHIpiRDD3ePHbXgJTl5M5ON8L6Lpb2r0nKQr
0kkPQZc2V9ThdQ2KEy93q+LHyuCMzbePlPjZ89UCfbAFTwg4HCKqQZ8zGmlKI5gwuGmEmbNCC+iN
Wkc2k3GRcXEGd/RMcIN8/hDQe4P40TPFAYgGTmT8Zzk2Gsnq255jyYmcjPzgYm2Nd95wLOif3Ua+
tr4x7xQcr9+ppLeFG9+03MjJwOeOrKbN1nIleFs1KLE1zvyJGTZOhhrmKeehITGGasZIKGlzykkC
jag6pQVSmnv7GGJvEMank5KwITyxjMeMDFinD2Upzt27OnNAFr5iZabeq4CPlLqR+pLN5p4eWf9A
KfNOk9phuqISJYruG1fEOaL3m6AkOf1vmBtYM0+S/B9TAeodAcMKdRr9Wl/hM2HB3gvHNKvU2B7p
nvODhhP+/MLnvuAVQHU77u4LbfY+bqIiF3Ywa+6nf5KC0e1QVb/gqAtvzplA27AKnkz45scX5fDH
upQGE5+XARfvhIcwamZwIlUbS/g9dQfjsSP3mBB2VXAkGLu5VV5PFwijv9fuQF2ROc4N+F3Ka/0j
30kTFR58D4BclfyWK6bETBaXvTJ6gdi9y2Y/IJkf+0ZJEmLfCmr7A/V0fsd25SWiiho+stAtwP9M
tVhzhJHHfHq1qdO9s8/olPVzoDFZoaEgniKMrgTFu1NE/kmhyh1AMRctyLkck9UxClYYuWA+b1il
VFovoTGe4QCdPYLOjs4wT/3Pw9Icz3vgAFLuqMCzLjpSsxLi5POkh7/hS9Qjt4wDuE+4EzjKG0Qe
bUsRan2nIoE6eXelITrj/UcHKEhxcwRp+q7i9cgcv521IZQaB6y8nkoYXpYsBEW7HmZJPE9YM7W0
uVUQFdTR+9i9TWkytVTR6JQ6IC4A8nuE1i0ZxdrhL0A6l26rybdSXYJPk8HXkC2s3CaEGDL0nuPW
KoP9lzU/gpaYgnk+6uELL6Fx5xQM7SvL2+zIq270eXk8PGaOPwrw7C60VI2liTgPRKVdRz9NY437
9h/JNhKsjH1wI/AE1E2QZ+bJjyn+P3Za2OjtQbxonKvqwzmwchw7U3UiRR3bwo429nC/dI8cTOBR
QsuJDY1wysqXaEwL4IyHYnCHBDZxoOWTEQXnNt5Osg17ft+3VYmetplJtPQbwgjmDiTr8UcLiL8f
eHufOh1xeekDicgHUZ4otCXFkt6OQgw7mXGAmBHkmpRiAZMWFCNysbU5g2HBXZXYscR0yreMVpph
jLP69rnuoE1wtQOb2rDZIF6jcLCPIyRnhfDcH8KX5gg1Ohsn+rT19eIA44AUMYLFSOXMTY1Tzxfd
sJ+uST0Jy1Iju9iPd2+/mx1SI99TJSf8E6/fUVv26qlCLq5yX5elGKU7fUhc5dbtd2N9Bqlg/UZ2
fNCYoH3Q32NGGgWMb5DNwLn4GMT5+EQdZMpe8IG/mT0RSI9EGOZr9myBuspfkaSJ1aDuu2DenknN
WcTQsHuXj1FgxdHWCnIZ8LAGe8lwaTtnXtCaES0CBTZovFaHzmka+KEd0r0FkM2fPBvrZzVeMg9x
37/63mg3PeCXQxtGTlkc9ErwPIPYZecynbE5gx3WHrxrh0jd4rKWmYV982imCT4/qkzbFhfc03ab
VU+EpsTvvVUlIeohPeMuq4GiV2PrqKuHNx4PaPZSXhnbp8W2MZNpJtjSva0B9l9PPlfhlp206ZBj
oPKbJ4Yl23NT+65DT8MwwIRZB+LdpJrIUNgeadupbPMfsfv5Ir0ockjIXRRr5V3KlGaLXpinP+7p
zJGkbNKrows+cEcHmwE/VrBhVYlSZytoGBxiBf6CXBUKp70tr/ueQMT4Q4j1RmuNh9RTBzQWAzaV
Iy8k3lO48tQxj1X3aCpnN1kTrMhpGZ9T+3+9xMoYMrBD3hwRtiDKdjR4GfaXZ2qQRnMQm+od8XO7
iTyswsD5NF10uO9zLogkqJDFreppGAKlIoinJPHXD4pDUbDIL4HB+kD/K7Fh5z7q2E2XJh0T1vDG
v82OHmqmIP/x1feqO4KHVmn3ZZKopZ4AcWkP1SX2FtoiOvEmeKbWZ77ZQIGNNJ9Ik+YlC66n9ed8
U7lPI6WvF6WEi0sQUxV/l22tb83dDrSrDbjGdU3lgW+2uljurr2pfTGrGwHjnk34/WHXr28xycBM
jgxZsrWk2R3ZyX7bG73J4g1O4Rhs5MmH8YYpGkc8AH5cNz0HrT2gGt8Ls5J83cpy6GjNyZyZmDBj
LJNJASlfUy8qrPz9GY1KD9wNfwGZhitptQXhcCkMhwSwpcXGgPDV+oSIlzo4eQ3ameX3FuoGf6zo
vfuRi0XiQ15MXdx1piwV1zIf9cA3aH+1WleezlEuv9nVJwSoOAgWNQ7NsLm8nP3l7QxKgUfe1kmC
AGf1hnJze3t8omn+YSoMcwnFccFkQwdmNbijDNp3Cj6s7br2pFEt/m7Epp7zNZv0SGzeiHJq5+2+
mbsXHsFDOfE5AYB70WSSVlvtWBcus8rbMcbYhSELuIQoxhC6+pfWUk8DD4HPOD1PTPchJtd7803u
iIhs7PKnJCKjAsZRo9K7hIOLlfEEmc5hlU1/wi7A2Hq6hZ5KDxeHNNUeD894FCyIVFCVLEoOwebC
oFq3YW7698P0zJlTK1+DSHSOXeqYDo7Ypxuy84Wb8mnMStafP9mWhSeeCZT9OVgZVlLYF+lKbmku
eBuGQgScK3EJPbFaaQJrjEuYtT/Vp/zdfAh2lx2M7XLgJjPhS+zOgNj/8JA9vVEAtPmhTP4Jgfrs
aK+q7DFUMVPSrjo2/atA1d/tQyiwpIz9RZibVOsoln/hz3p/g2+8QIYgF4Lb1m3WbuohwMZ9Jmr3
hR05Ib7Q6I36woBR6cYI69oVyVm68uyIN287Kkiia19pxSS2tkgh/i8zsG8xlTxro3qNx4q8r3tT
vXsB++P3lddw/JA6FSJN4NHvis5mkEK/so24yKLI5Axi5BUI0BMsthV2j4hlIWR+NKYWwmFX3dDn
Meeu/U+rkN+ImwlqU+iDQnof1urMk1ztdbx+3qRW2jED+gBQGnsvKu48AAxYq3lFPkTtOfX/G0IA
eSJg4qlgu674TwjDcU7Gs8atv7xpjAjgfVW7U96EbwfoKyMYypht0oseStSIpZA9crUW4ja6cmia
L9bAxAmO1X2ckOo1tCRIv6RQr4CD1g0bauuNJsE+UbSp5VsimsnKYTw5GiGkkXDc6SC/13BA/1cy
rr8nEEPAXHAV1151W1S4d3AUFxswT2gr3tnQw58lcFs04iZWLmfunyImfiV57UbI6n+9HdKzUlYP
FfPrCDzFT71p03q+pXHGxojpSc2lzjkVth8d249dLW4hd8o0UBnjuIfls5CgDwnaD3qQFPB1XGhz
9FmUbIJhcuS8JI2thjeqBWYRJAW+FKIJqGB6OjnIblN3FSaKIUOtUpasLC7F9xlgv57VVZ91S0kU
XXBaIna9OY4ssMAXDRPL+Ee+0GkW3Jlsr9xaAdg+oo0BODxafBWQjAObwinGrOQj+ltkdE9Al4d5
TmD9VEXp+9mL45JhC38NaLKgeRF3n/i9mD6/94+ty0vQ9cYdRmZ4c1/lkD+BYgYijB+hUp2MfUcs
9pPHvE9cWEGrOEWd+cufZjXwvM6x4I1+PRnhhILBSEBOjXe/eKaFj4iqtflR/dyPCiPNLG6hG2uB
43oHbwddv33AoytHfKMasAiWXTTQUggEqArgpay5ayJjS9luOWmwuc/pjT6SMm+1RP1nH89Vzdam
cZhMKgWpVmYiDfQcLC08bAT5LMkKVeywtqFT1m51WScY2Eg4k18G3kBfEHDlSeL1I/IdPsIIhUJK
O4YHkP4YwMh2+8t9Ubsn9IJOisXSTPfnai8W8m9U8E+RVduZP/4soPn/khpOhcKz+UXcN7UNFJ32
GNQimrUjCUNBIq4+vtP3LV/vBApj40TW4rzYn7G8h+ZxUWPQHmeuyJ77TfVmnhW3SuggqcHgcZmJ
CbKj87g5/hfkUj0jeE0PZkXZgD8Bh60BibX4EExm+Tc15j7X5hSovl7hEBST1VqJRlzN/0tpJ/ol
EsjVfRTqkjEFCD4W4O+Zi0Ynco5s/axy0JCUY51N8u6drpBprg2vKIyLfJoAi58qsLq7+GmEBLMZ
CVYS5+5kwqNrWdUAS6NgLmXuSPLqnBJW/3rd1wDKvpuoHm+JFpLsXs2C8M41hLaANBRSSWkaupED
al978vt2QIkXaThtzKXgJPabh7u/4dOTocxLbSFfipcXz7K6oKDjkQQmMNqcknApcjzKvST0HvL1
tsdrGhWutjuLd1pXZFR2Xr113GasBZzggmWJysS+6IZ8GKwLMA3L+vM0TkDqDfPU2Oj4R47QjQQv
9CJwTLI9MRLCGb13Acu2904o+VPhxsL0IwvakeKodYuLYZf3jCeFp7mNw+ft0tOtw0e1/jQelPJ9
mBp9fhxrSALgd2RXkxiiIKhlNvQHwiHxt22A8EWSbib5/V+cIhYRXSmwS7BtPUex/nPyGVXlDhlW
xes5q7h+bB4mLi2Hx7QRzRRFmDd2GJvD3tfk/EuC6T+ehmEfvOqq2XlbfiWE6OxyWotR9spZw7nW
2YDqY6w7vISL5xZ5XoRzMpHGZ8FaDumoUld5DglOY2Yr8Gd2J2eGHLBkVUj9g+ZDYbTRb3iUrK86
QUBF1QYVoW3ZCECY4vPFPswUx+FpIa1hdE032CSh4HQ0zzN0OaHEAOD4gL61GCjiJx4PN5o6zYmw
2+W3i40CsLdOZnG3oIDXXDWLqcFfG9jjXkFOZp8D3+UPnvoLgkuOK8UdnOzeSFl/YTyzdJQunAox
TKCX5xjKvY4ZbyDYh50V2thEuMfFIhr7L6g+1YIKiQZYPi50dnbvmIR1oR0ZZegLwbBl03NavPjF
kU/CMVoHsFD54JmH8S206kaAOOmj/bA8XGtEg7mkQNuZK0Q63EPPQx/DBjNY+T38CAGhwFYVrIlc
t5eiLtHurbV0kZWOel4RB2BIT6SW1j2+QawiWDYaeEBS/OzgirXsFJaJzoQK2neiRjTzQUiMFcfc
ZWuF4XCNgvN9I5Ofem4Q+XTYfpg0BCu+dQnemj/Cu1BejBfClqMECrMv19GcWQ14F6sQm8xczhTl
ulS1xx0WsVif9TPew7kOtXH9v0hDaVOHTVXk/wqB5uH8kNpuE09aIlxa4nczzwJaLfF5MnDrZaBf
TmxoVCvWvVRNX9L6y0SaEvKu69iCZGH+mWa9mGuwa6sR04suvFLEHFsMrI6JYF4E9g//h9RPQtAO
xIjJ93KnTP6ZWWdN9f/YvdMLa01Be4GVfA+oDr3SUzE6Kn1Qn7B+46LIkuDJcef8g1Poh4lNs8nQ
6M0FKufDHty1YYtfQ5Rl+yPwN5OEncEL7QKIVr5nWIz3vCRR87Nc50UAnd/PqoIYy65JhjZn4E6Z
URrU86Q9d58/koLk1NOqIDBJCxRUUrveE3rVCMgz0L9VZV7rmwqzD1nD3f13avlT8hpUAkpjDBV+
sizW0CS84HiBc77kJwtKFg42mdMuLLpOQTxnAu/eBBW5wiA4Pdv38dedpdlDyLqu4n3oKKS0ACN8
Dy40yllbg3xsIXE1Ft1CLtWKSTuQPQCQhtDsVOSOLmJStDzlvf5cwTERDlHTvfbGx6o2c4wvvR/6
y38Rt/uTt0T6wWksT0Mn2F50IIn8H5oi436gzoGZxuEPyKY+1SLE66JCTIOyNJTQ05T4do8D2z/s
ipj/mIDAIkjD1b5FNsKWPfT/k/UFNRPcOJaENqxcB4xdOYpNRheDhnVJ3ZVZLhaFM4TDIldVtwim
ShGNK4oYq0MoNStgleEsBvBv1Mbj9ykk/yfe1H6FQjGrXGOQujJbRa1L+L1Qfz9g38iJaJF5Kb4W
g5RN75UgLQz/lM5Bks/sJ1l88eB72Tj/+FYSak/XNSEB6j0UQ7z22HGx4oZXw9t28pFvhz5BUjzE
zJkE7ojyIOiAqa2v7aR540cMBRDtxXIsMlKJAhyfVOklG58h6yi+SEVIWle/FmknQeHs2JK3nGKR
WrsFVQ9/fkRSg8jBZbDgnmGa9YwzpLapbNqjSjj2ECoMSCaK7HGAF9qseFk3UmjTEn6DBCsdnvkT
1/UiiNaVS6yVm9YXI5rEVx+y2lHWMlLAa1cs0BKxRJPIBfJsNqzF31m0Ce28JSezqlcGaQVJ7dAF
5Mw9wDtV01EIRdMOVrtLry2Ex0XCfLZlb4WAJu4vXDzrfhdWlUn9GTibRznH34xzalcCtrRxSBOR
cAK6Kzyhi9w6Qffi/VwMxte86RRGOykPGLHyuruq1p5im0rn7NekNDO7okfzJjFxt7SBP+kTF7tF
xHrbrAJh06VkatueZJgQTVKl8XbBzwWWfs1oacF16XQ5A0razQN0DT2OGVRaPGCCAOB3iMgdhYb7
WfW43JanCQgkakjKjZ068q3M1X5HHA1k6BFeta8daxU4czu9CgoFIWNRtxLjFpQiENOOSr3IUWh2
1+tZBP76yl+0110ba3wLaldGZrKFNaX9tXjYjWqI86Zww9wWFQ7XP2OWTqyv7Sh4xHQq92pW785d
pHsfVEZVquS3bX9Fi8xwBTv8eh4YJffQOFcgtua1iUbmO5jbj1g8OqMMtKu7poXUXVVmDkpfWJIE
mW+RQPvSMLWkqviz13FqmThRp28ijgRY7uUikyHuifJWGwwme/qPN3oVFW0D0Q9h/IClzxpwURSq
9yw50bdxKO27sFivERgT5pAWmb/5AMzIvboik6ODdQc6TWaJRinNWHGakWV6R8ccoz+jpwBXSoAW
QpQ8h4YYigUPEUexp58hQbNVtVeQmqU/E8m7LIIbs7RcXNGVFi/ejeE8UFwA1hMipkiq8c3wBh3w
IBW4B4UshQenYKintH2xnLAuMRw7s3yhMeofW19JN8NFAw6gKyJA3xvvoYoDxyy13q93RMbde3BB
eANlLuLyKo6k5Df4VcTsJsPj96gZ2eyI4ce3lJQlMHeXthOfyrMpsJGZA2xA488MtNekXdYsoWjT
efhw6N3LRmVgrEONgagCbUL/wV2kIgG3FLobXMYLKZQS/O7aMp+3WO8vDhN3alf6dUhL5kxAqV2G
VZlDOxsy5mbtcg+IG+8oJiDzuKLizQPNw71cluSxWw5s0v/dRk+Htbb+aDFGYSFsvbM//WfBD9HN
9Zt5f2WlW1hDvu0mFt0M5mZnatyjlLL+dteDKoV3ogX2RH+tzIPP65CgkoiF6b1+WLpyrvdPgcyV
P9lYAzJ5CfNFTRGTX7XTVpJaKuyMzmopXhkfo+cBKCctFCIw4q0eULnmOwYqDir8t6cvKa9Lj6rj
myoh2lqBXK0jdfPRj/WK0PKNAz5YccG3SLI8WYrS9KbqXbgIRE4c0PIr2uWujB5v4thJClLzxyS9
UtZDNuWh6m6e7u0Dg3+j35wQV1f/ynZJTbtyORFkhegNdT+RxUjIuuf3XKZP99r0ox04lu7RKxvh
FeSU1T9e4aTAgk7R8tgRU+lVgZbzD5yUWGw1ZqEyz4QgRiV6uxL9yE69tUslvjZt2O78J4fHTYnI
MV5kxvCYUYECu9LI9/XTpHq/niuZnoyPJw5sPEN7OMa2FYNM2Dx2tBFRfDLCpuVFAYQUaPIUbgWT
3Dc18zveN+yIDn+NjRLCFoyC5/GxEVPtp8+bvG5mK5ntg8H5TrUiVOUhZh5hkc6hPpobWAgnmsYz
QWnDpxJEdjHo4Amsmt2WaZDLYERHV6yhaIvVs/UHmR3mPCIl+mmxIk4bPPf9xZRLGOq9qEizWjBn
TFB8qByYNmeatjiYLGM9FOnFjWGU64ShmlmtGaSWmt4bd8sp9cjpMz7dlMxZfD+Pwa3y9Mx7Z6Xe
rru4Pm25ByoZUemYiD3FriDGfDjm6SGXnwMc1B2cVyIeFikKfHhn8w1iVglyBRZ0X8qLvYlek0Ys
xMwakJ3S6bEGAlRs1Gphk+5K+DP2mu+tGJMezwpghBieF2Krq7mHZBvJjPoj1P1JIRmRpJ/xzFxm
D5iq+SJEZoGzEtUM6HvSYvlp8f7i2ojCLwU6Ho6VAiTkGSiRhV6C5iyuukUfuhejcWsWnELMauv9
e637+uo2BhFEqg4wLeQApNDMwmLP8woYxoRVmqyn/9u51bwIYS7DTlf9LlR/lOtSDXml112yilgR
A5uu8tPCLqnYXndDL3KrC/2Q252nKExmrDeTimOPaaRb097gKB7F0XJp/ydK4zh7FsesJftU62u9
uRC53ww1u5zXtOgr2IzMznBzs4Rv/Mn+PCi7V6pWlolEagH40BtYifA+RZhcfx499EoL81M81XrY
z6TcGoyy/rbhA4APqoRZu9kARnTtmO7BzTT8ElvI9tro++/c2NiT3aVEav9S8eQWKJgOQvqZxkTy
KNapVmJ0Cg/aO5rNPwIMVnx2Umqvp3HMkk+A3ZaMHQSEk1zw/vo8L1ob6YMAJRecGzAcgnB/iDyB
wrcQD38yNu9d0ciHet/PiJMuW+qkTfhZw3pD4dM7szjiA0+V4oQ88ajkzrbdFFpKBy3p77TWbHaO
6QKr67TK3B0PbTsnq9vaK2Q8wJ1Nzg+zSdJBFTGGvaOmyDutA7KV12dmmrpeBad/OLmj1C4VVG/e
zfvvOYSdXQ9M8mtPtYL8kLq2xgiK2BB8HyitSG/uviUiG0DvAJL3U+TphJNdT80N7jNmTMdF3awc
PaUAUEjko5xSlV9wsFBwscEqHiZMR6YtIdRqA1NY20VAxviVMcidLZdn04XAhoaatgdxWldVfvDu
wjRc5WA6jBnKMR+YUPXEwtUsqdWAapEjsIXHw6O8XfZN8WVixZ1G1TMPxFh2FdEeYgL6h/g/ZcBr
3L4DcBUOmdGaH1x2EjFvHLQ/bt2vYbUD0FnOMGPKgujJljGgK0y/9GPTINN0EZIBw3a5ycr2F7rW
AzPcqEcHH/8k7J2Z4EPOdfqCn7YbceI9b/TWiaQX49QC3NNTTVwiCjEUdII/kUprctu7mPEvn6y9
69uNcp7uml721xXFS7Gq0TLoNu4JZ2vonsngGaCCrGGJiMzHQw068aQH9e9EWx1dOWQNvfSvv4+7
uAcophB2hMSDzRdCGP9bu48CRy26wTp3qLodYmW1Mhht7QzwPqCCCI6VMInZ5IL3LDIzPOrBxrpk
ACpfBe0vp08A4CKcY9k39+AdWjUgZctY0k6QVKceIQIy9d/1Zw7Cuh3sFvoR89V8JM+JJQsBPOVK
IbFUAwOraxjg8cfJO5LkEFbB7bIi2gZ82ijuyaWlYojD7V5lvuTnaIN2UFGD2BkLtQq+gkW7Y/he
F/vQ0OshoJZY7OdnZhuSQlljNb4AK4Bmb/74Xi1Ye31+/i6hcsKrYJ5ZBm81PqUbmfLlp776mn7L
Hd6Z72YVob42fLvgbXrX9yo7ctxihV1BmtZi/55z+hyCCJ8FhYWSLlTqlTk/uZfZPGR5pMxzUk+o
fXETYsrAZEspcPE+FtrO2OCzsIemHQ2f6SxV0VJZP7G7j4uWDpiJqyOxnRH7KCqdokVLrqXim1rD
NKc8wRk64nQnekx+7z2liFil4dGCc9lcqnzi+Y8pOYcOob0shJQfsYfAH1BQAL/6CrplXiBLaWm/
9bZKrtZllBMSv8OZlT1CwjQy3S0OcdE2cTwkEkebvK43o6orOSqOAA0JJ6+vjA6p5vKY9Xwz9mPX
Ub1ZtM0L4zlP3b7oDGWUY4RcutSIN8Ytwf92cibV10EVppnfMZlcBeVeFNe4i8W8qQ2yIgYIaPwy
D6FfK62GvuqR+nne5vaJS435zeZ+DdwFBIDsHZPZNvx5nXK6soAcCQrfbfmG1syCUVoMOWD+57y5
al3mf6G7MSqBbnzPI9CDAGHow9GlvrDVCXrn560sSjbYTB8NT3TE+cQ8aBPsbcLaYp08SjiWGAcy
dkb4OVaeRCYQT2AbGtX9cwVAeuvEo+Nq/JVSxNy6Cg6Iyc01lbgPwXhSfre0d062T4RnX3lfwFV1
jlwBNec677EIFX9m6EDxGkVA99/F7kN6c6IVYUmWKZnM07ajVAdGjgqawkrXkDVsfPtSBXqnE2B/
TjguIXT79tIUeHwvTdwOynmsuvsIly6sGX9hN/QGkbpqWcHDfAJng1HUSgnsYifO59C6gQUOvgqn
5FIp1PkCgMuKa4RUNolMJWd58p6fS7cq6dg0RvrvXAMBgUtmFK+Wy42Y18aHbZhzypD1mV0c/7oL
N1mp7DEk1eO5TuokQE+2iNhvHaUj310vbzH9ZEYY3XMMZfCZD3zp9mmKmpjiBlerh7SG/8rgoD7b
aABgR2nPoBKljCKIkRi7UDncNcrdtTzf02cZBYztbAOfJJAhjWWeV0TTOsG0G7Fv0AfWtQ/OMVhu
F8JJp92S1KnuYtDz9lTjwxyNrC4iIutyhHokgOfJlVjKOjC5+yYgD6SqqlmWLxV+3Yb6lzABw08Q
93r/DSwJKIRIggN+rJ6ja0ZLpK7CoQm0QcxYPK4v3gVl1JNxr14TNxRA8ogF9bGHnEam0sANXEqB
uB3nnFiANiZryQFSYwNLhts2Cj6QKcAYlZWi6WzgXY1dGxLwa6s3PpgG7J5YYudtzn3u55befpk/
RacR25gJqaDmtRmlwX1C155TjBUXC6TQPfA52oqTtvrdcvtsAwAuE3xbZziySlPsHIXGb7V+m44v
Y00oUpANyv4c82G1wlpatJAysl6uoE06MRee37MyrgXRSH2EI7H3JWDM78Q+QYBCPGRaet5DFNf8
19kJKCBnvJy3C4ucpaUmSyfxNoSC1gpYZVzyTSeoXaWXlLb8Y5Uez37lFbopLGZLLDg6vEIUeKHr
zehhF+ne0OQpvXqpPW3gqUPMVjBaf/TpYg4u5Bx3VXp43vmhl6HQvdKt62opodnvGzMjorcBAjuk
NqDrTSDnConRtVNIqvaSXJ6clqT5qMZBiZ4/W/i9jqUAiiBd0z6sLB5tqNSXaHJ3znDsQzJEEZTn
YwXhvrJzNxPOPyn3y2gpaJrPhi3senhbK8ThqxBDVDnPR9E4cKU7Tk+o8SQ8dfNMkgwf6P1CNgAL
GFRpDgG3rH36kEI+N9s4XJ9LnQmapqJufxR+GtCqoEUAfjFrH+ymOi7WK/mI7hUEZQwphfoaUYBW
zeguetSbMuh7+Teiv1Tsgh2aaKgsTK9NOfrC54LjUuTILErBkQCUwHP6Z5GFR25yJfdfA+z/dq1j
Hy6fQ61v6ui6+eCIq+GoCoxkV38T/YENIyHXpgFiotPRIZKzjhNj7adkKDBTy4o8/jLUYJ+4NpmW
GULZL2HwxL1ae1VQwZI01PfvvZQcOGEBr3OnWC9bNPExa3q/3m4497gAsYYQ/unmGBGr0Fxvi37u
xYz2CqehE2fM14c4m0AGkhf6YNaSqm4O7eY9uN91d+9CukByTLe+NGIcHA3TNd7Ytq0yfev64SZo
fXdcm2/Pgrv99ZABMnOKLX0xVpFEOunNV+e0w8/aUa3pdmZtmiG9YYwm88dgwYf2erTT33HZxbvC
knvYXWrBnqcUoSE4pyBgW58HFsEWyeMUne5XtRWtYKQZCSkxvyavMbrUa1yFjieibTMk5vyJRri8
XyIjoAi3YvpZEHomtbyGgiUJpFA+W86jfoSLX18su2C33GYY0/NP+X41vK3wgUWfAxk4M4Qtpr3q
DtNwdY4xSGjPS/jX3M376BgrzdDlv26JESULCG0ARH3GzJKjTj7oPz2GRYADP8D6UIyO1jN9smto
NBSzIj8TF5CFWQnqFmyfc5nGJoLLdf+c35DZXm8QqsXc39YSKcNFf5p660S2hZXIgyibZ6BAMl9p
4RJisth3A0OYXU/jJQstjOisPt01dECBmmYqDUzL12wYjzQzQpXcZ6MW4NOuPhO9sepiuyLfFHsC
Q6ohfcNIIUnaFzIaPUmgYvE1V+o6gyN56Cm7C/YdwzzmOgqR/bmqozNrM+RUz2YekVu2HDJFPZ6K
+AhrwsyAE93+QHpRWEpyVJnTqBqNtA4JsKGhZ2KrWUw8TMcUepvWpe2uHtF4vOux8f7Fqufd40IP
5I3GWrpwj97mrVKrIBs1YCLBQ5vd9i2rnYznVSrxwZvQoyqIWmA20jqJMOicpq+d82lbpopUQLWM
jjilG8gCqLK2hHQuUt1GRV3a96ZI30YPkqoh4f468NteEagZBmcYnYSoKMUsuCwtpx4vWgz36XDN
JoK9F9FwBX4XdiOhMXNHybwXGduywU/JhQK4cKQRBWQkfk9CfQgByoJzU4iWoJAi4UR/mEzI5w7X
4W/kb8dTO2wQDDXCMb2w2uslibmNf121Ik2US2Nbp3mfpqhEnmSzZl41xYaWytfV7iyj+gzMaM38
8ETcaFp/Yp4FnTS+iEJCd768c2w6N+bfJL8ON6GaYZYBePN/AJxRn7ZfzT7BXuM8lg8tL/LFDyuz
D8sstosyB/v5UrNaN4uHG2Pp4ViUp72N6nRvY0lFYHzeH8zHnQ/9cVpeXFUWSdZMbsyeXmZ8cnPI
nqTQya1tpwkZsQfUSVbPPjrzob5kdFgyROizjvaQOHJQiS1db7hW8ylw/fgfig9G/vhf/g9FzXIs
dNG4ht1BxsY+kvmq7Mnn5YBdd4k3eUWYC03eb5AMuBd1kOb3M2i84wTuuhWKaY4xgI2gZp2XpMlF
D73fqp1Vd7+NR2WQoyzkA8RfCXfoMiuCN9NtyLKcu8l+oIyr4hk85ma659fAtWQvk6VqsEyMBRzS
Guv4VLNKmnvICDfyyQDuWJfF7geaFpECoj2C47AeRNV82e7+DuqW7KUvGcf0hgopd70IsIV0jJkd
oLPGCK4EdiYJTzI2OyJnJSFtvPK28amu3FgN9JlllSyVT102CYFh73grXVnitMdRHDptvDxcnBHZ
tegOGCRetADbDBM6lCW2HPrNSeUr2mFOmmWpkJBhnDCIqpihQP68H1tMLLNOE5IW+oYveMC7icCy
H5Ok0/lMgqWh4cEkEtorTyp9gkRLWL+WafrxhtgkCCMfG0FLmBxc8ZBgB5agvY7ZDxq3s0K8NRlR
kQoAx0Hm1I2eMyJM7eOkdcd/fmsIMrhlS5X+T5guBd6ACwdzRIXNRwIgxkvb8gYUFHdAUhossxIl
GaIWvXkz2PPs5MHEXexZm30huqU7DMunR6esgAjjr8wC8e0ybuTeey1hbqW1awjPSjA0Y6zXthEu
bHd3dvHQzQhzLkHVHlEoXF+M+YSSGpRvdywRlENrdQ3x30rJJzX2e4QNrLmFNBfOd+Ujg7KkMkFp
25j0iibAc3Ccl+GNOFv3kRGP6/7faq0H2DVF0BXQRfzNIeltBr1dofhpsZOcSQuVV5cVqjb/QVhx
9emhWIBhwisJh5LL0TOHixO32zyLkjrS/a7ndz6RaUy0vDuaaVcSv+n3CM2X+whOxHQozzKYi7u6
RCl/moRAg2wEHANtIpc+OO5Ts+H9GeXY9/C79PW6CltUJZGfbb+Kiqz1eUmliq0xyrbZu8DLTcoY
WajJ9qqZn82FnEnU8vc5kZEidd/uwGGXzSOtXRImYGL4ytWhXSiGO7eCH8m6++FLMLjbFlgNL9KC
vjHMlDQ+IxCcdkAX3dEwhKJro+kBl+/gj9tRfxM3pen4c1RsEfIhXo6Tm2nCXF1SwjSzR20Lgptx
81ZOPRgZiVk/ZnQOyNst1cdxdpnlC72VVTq86cezLgUmw2KOaXeL6jAwGuycZVRZ5VOE+g8kWvUX
RiZa/uQi+BGa2QKG64SNovmAjWFGE80nGLsJ/7+drWRpsG8V2WIMkehKkFJZxdiDyy84LzvmLhmT
8zPdAj84Wwss8gyZnl8uwEL1hZ8BVrOcyBwezLkT8/kRRO42PBr64yGiYPJgJ0Et5bmXsXKvHK5t
FU6ULk7m3pv7CmE+rbE6I0CN2JTPGEQNUnbGV5cNhxrOY5xtrGT46OQ8XXTve/DCYxvW9gk67rL9
PzZ7p/xUZmFenSOU0nGY6XuNgd/AQsOZU4iuJRr4E2tDIu+CETglTy4Uus7tdK1K+0J5LHx4VIuI
dpCyUrktqZCKK1smgJxopPwcJjRR8QAWmTLhOQZDLVivUvhMrUCzJtP4IVuM5lYDNjz0EoCFTmPX
3s8wIFkZ2jPmRABYbtFbUZKd8aD9r/kYPzrtjNlV6DDmJzJZXjhCglxi38rN7KsVI7U1g7d8piyv
5QITqlN+ZZxx304gpYKsI5+5aQf3dm4+WgARNeZr/97xhnzNS75EbrC1u3kMST9lTUqc9gul38l9
F62FJN1inB/EkS8YKdJ+BVXF7G3xGTu4K4/ozHLYIzLrAerxYnunGsN69yNJAWCmRu++NA1bzsvs
c03ho1Y8kEDjpxgGcL68h+BfqOF+ipKk4SNe6QWAdo5U/+QbbLx6L+1EGP7enYwBBz3KJlF6ac+j
gzE0Q7KkQQVaha04f6wkp3PcsBV05l5e1ZWCo8ecrcn0NGI2H5LqHsR8pjo+nD2kFRj6uyd1h/RC
VHmiHaCf99PMGyquhg1ovWhPEX4LaX9kNA/Wd+5WaHcFxx4/vNb4OZmE8arFqeCtP9olAkEitz9V
w75gSoXGWCWp19pvtAlafqw1xQlA42pISxRxJcc6Oj8tNTRT/a8tVLvYHNZb8tYRPMWi3A1vp4zc
OrbJvMWO/J8CuTUJJ1dEHZpglk3Lf2mjhdYjpSFUrV7Fpwh7aJkCy1a1AN94w4Ow9gz22DnJzRN9
dF0v/Ebnw5q8dJf1sl8/nhABuiOTOCVsptl9ifbbFZYXsHmIoEiFK2djh3MeZwOvd9/TsEdI/cWK
6PjLcsjie9q22kKlR0S7uO6L4Dm7GmE3wTVI9dWw1tBNHpqJyNC8GdAedwf+ktucTM0pdivTItQM
CCZVf2DkW0GcTN/h9hprsuzVMgUqQCU1aWhZDc4bZvkaVQA/CfMmy/dXXHgdvMrCP1fwXGuVX1kj
bHsdLv5gPKOU6i2i0Rr4kVqjF0Utr3zqMuBGp7QghKbD6H8dSkHXHYkilwAACulWI2y6nnPwNN9O
xtyggI9J6WZl5W5WBhwPdb08YzguKi6Fc0gD1zaC6p5hUxzMpeUEFtUrYLUdlGkmXfwmrEp4ug2J
x6W32dMRTWcJ1ik5IBm2aVj66WLdLzW7wTrJUNNn+q+IQ+Q1niiDez+8jjpP+vsqd94Hm25ToE+v
allxYVq/LpCQJEbqID73NqDYQVCCSE9pAloU4zSrHX+ASNTUKwQxSVH7e/oxSQ4s48+eDtp1fo7l
xBMxz0iLqR+m5fCV/UteBUVqSQBMZRspeuN9lDdhP4LLr2tEMcaFFXdGnvH1iCj4V4TBH83VrHoI
jgmY3jh7614OUfNVIpTZcFz4jGA/3NV+aXQAR55elvCjIc9YbZ1BGePcHIdxlLoL5BiXwHh8hhd4
06Y3C1Arwv49lxHsGQGQFUNo0gofjuE4HWrl69EU18i6YqaHS8fmHrV0iZDsxogDO+AVcDorPByy
9mgIoqBXQTeXZRAMjQFcuMqTyP5b+koAQOZjpJdxLl0pbIYEEAQZuRsfa16mlGze0xZErUok+L0U
ndf9CWsztBd41o9f2t7e+75aUdApGr+wqHe3yvvNsCw0ans4aWhc1esPErBaiIpix19DX+cGrr53
U1W0xo88V49Ry8ldT4uxnyzNd54M/jQ33E/UDQ00OpYmbV8g82HfoPc1coz5qMmFS+XtFHh++DXa
5n8Bud/nv3nSzHjsgLasizcJlHpgW2iCumUlmBoEr5w2/dOt3CFK8CiHRWNyK/0nLnq9xzdhYtUP
Ru67mQ+z/dvcfPgN+LpuqficE3tpH9EmoUxuZ56izGVpJaEVijl5tnZnLKBYCP07Vd5Dmy3QmzBS
Q4BWeaHx0bVT1ok/DX7mtg1NQwO/CHLs8rBjl1k4Z3F0qR3suMGNCGHIrh5BGQs3DeoOlWb7cx89
RSdfern+OZDDKVOY9vXfoHWbD9111X4iDZIGXyO6pYh1BiKMyZzx9/alosyMJj1/cXTAJFbUmOZN
34HsdEzM/GLRRn/kWY/9iJ2tIoWPG7osM2TapvMGWFXHbJR+hmlWTWeptkJAySFJp22qTR1oOJ/K
kUOTJscHqYDialhs62liavnf4PphPDQ3PvXMigQASJo8J+kbShq1UV2ix7p5JraP6s6qc9Id7DMa
vuPxuRsB9eGdtpSAW2oi/lk4U5rv631eH37LVBiPSNyEC2HtzFMJIqh9ckEoJXBdYz44NW4uz4PH
w3p84uJfPD51Dz9jlGGZfd0P7npW42RaaGxRl+Hy9s4t/S5OXxCAmvRyf+626jkFyGwXYbmSl9Gi
3656MlS2/3NJ8AiTY04e8V4lI5iViCBRLq0k4hmd2V/iHFS/BnVSu0mBUgykQHYxiQOH2dQCLIoZ
doOnR5k8BJwcNrV2nVRabxSPSSjs4XzKQ/+KSEYkKxI3WHBXqgzLdCybC5H3k4vsJDykZuiWJ80S
9+LB15p9SQe6zQ2NQSdF9YWatTwsbXdiOQ/dyZmPSVfx84CQiEsfcr94SYhkW6kt6TOkmexopH30
z8L16ooqeFr7i4lUGP9dyz5heibt8W/2RojLX1CVxbpnbneZ+g01YszXldlEhQBFgOZt5icvvOQn
zfalZRtVyX9YcDeZ04fVfsmV5VKKkAzpuOyTAxvtCh9pORb/AGw6w6kH8j5CjweVM4KUtyyNiCgB
0ayfMZQQ95UBSvDzLb5OgzmHLvzu1x8pt5gRNsoPZnALU+rorsK9GJ7iscC3+HV78BwL2QhenAje
ecWISF1MhND8kbVepwmv7j+LnX41KoFAN7P99cYwye6MLyyaS3HF+fHa0k+6yjmOmoC2h21oR6tz
W3Aov3cV1ypBmms6lWCLCi8G0nu0EeXPxIJUpF5CsImTHyv7GMYhKNiEhoV06jgCTDRc+V40UZ7j
2nHcjfRBguWvGkafNFgemwFHfVrKC+GPaULRpwaUcdOoNKz4TewhoxXqWboL2726Er4voId3KKJ/
jN95ron1QBUaWXqf/bloJSwrVRYrO6ufk/ASFoG4EX09JGlFYgJWIr4jR6PaLCqqYPnzl30XLcJC
+B0m+RRMUxE/x43LWNd0zPePt2gVWpUfUBlH+BNAFtxLCzVV+D0VCkEK1NvRjwibwPLQGd3KYkTN
Q9rTGmSYXhyjf5/6s2v+KawR1D456V5k57aRif20xrPVtzfq7hKFBSJuO0m9mw/s88iuFTXrfa4C
LdjngaeQSYTzVqn9lREJY+fvHXCLXjmVhjO2O6cKmxtivUnWVubm/+5hd1hwr6OfFvHxmSKvRFGT
IBi+h8rz/cS+GgKy2jI036S12VXgSI12uJFB6q/SU8J/9Xb6ZTg8lZD6cWVQUNrbp/ZMkjV6wbr2
hOKXLgxN6kSj+RPrQPXQHQvTxOW8O98OstKxVSGwGf6dWiw9sOYtkQMjhMFKcc86B6db6hfHHJqk
05CQdbcEttKqiT6NnzugOFZq9QOI7QzEktzJMtvBggK3Co8DoSELs4XaEtMbB1yjFoGj625OpYkU
skqUO+5B97vAGmvYSYtV8Pllmw9TfYYIxuLAdd9mshl9/knTz7ixncOKb9IGQeYLR+W79i5Zhrfb
fYtzZsXQWnvwPoZ9SrF/I9XUQqmpX7FsRs088kAC2cV31VoFm99zmBvi97u8v2+IVoc0gbG8DvE4
ypkbYRgK5CQdFHRRpHYmT4piboLB1bEeY8jS9gikqlO33XNsaLrHM1GROvgAgoRHayrqjlIBksJE
rGpJMQX4sakldHSGJwtektcEZFQrCcu6wY8S2D3ZxGEsyQAcLJV93pmWOxI3fHLohmETq1eIAnhl
bNe6krUJSkF2u5kqcDIMtSsOiJ17yb2V5AM6AnW2pDgMFiRjHpQ+tCw8ra6Tl7dyjzCBFujZp7Pp
7wEga/d9ciHRdwDfaRKOcee5YRdtfT6/h7X7Okt/0wTSL7bLzuPWX39OzHzBMJ6DkAeYdKjsuLeL
rwsfH/2fIRp441J2g6FXczEqysfnbLBsjxoGE1zsXV+Rmo7/YzsaLhJfqq/cCsD1PmloFKyawQzQ
oA2Bahdh2+VB92TvrgaZcuO3smh89XnYUHVf2acliqPssiBEWLIlGdy6ydQnsiFA9hIXmyTYID7G
7uOGNfhINmhhtMmS1Y20Azq/wxjqZBnR6FjDP6WCqLJuOwFEx2uRWJQqe7tsWHafU8tKPNwN283o
xtbcvwdlVA6/ohJnx53PVbSppDzpY8n9QIx4GwCaVMI0La4ZSZfPLbxLBVzPRCQ9bpMJKfsOzZhm
BOrvDOgVBZQw2GfUkeDj3WxvoWd1PIVARGV19IN0cVWQvpJoWZhbsSQ9yqmodAIv+oQjENIzFcrw
ZYpY6zogwuoZGhDMkV/73RXa+VUh+QEnG4S2CruI8G8ngYUmm6pRblvX/10EtGGU1EuxtbV8EoEH
5pjFwYIc1M0pD2MLW3jh638KmzKa2zjFf0JMsL5FDAjobuXrW9vr7/zx7pLTEtbV7iP8YIguuhDJ
QPjP5iukapLP5rhOsdudCDFYmzAe4fm84fKvel2FbebL4VndA74LRtkzipnbKIOuZXsVJO934fBA
GSwCBzFw0PekGPRMDFV9wKnCHnciF2UEVNwl1cLT9XWD92IbU89zgUIKHiKZeJd8XeWlS9Pw1HPP
CPERVdWi+ShYdurQ8CB+fUaPusiVjEMrrfW6QrTBwt7ZW/4UfFVdl/jrvnpBd9OS+Rgyt5gcHyoC
bw9hfo5lVqME66K35W/hu8Zic39Y2FMuB0opO2GceOw4gsJGUEBdRFpVbg5ydo+gMFp+enb9LyCD
y2lYt5Railaj4KG84Bk2qZH16Gf0mF3NI56CZdJBXgiRcR9vJhhJAHHXOTB3ftPBeBRuJ8EGL1az
OwJp2J9IasASpUCzelZSr5mhsHiWwQZbFLbqUNtKnuuJQh1NmhTyYmvB05m1ltOhqPdRHmW5rXtW
TV5RZqpNH2lK6iDAad9Dus6RftJ3XiNrGiPtHj5ld547NZ4oLVKt8wZR+al0IfxqDNUSjbEvDscj
BrNE7HFUxsKykPb1qIFDrh8AME7mTrlhHI0XeTjmwVK3qWWiDqyKTpzvCG5t5ZSfUZdNGw5MTgSk
ZtXQutmfZSkY496aZ9buSuwODw1Vtml5OQ7vjeDVJpK/rOuA0ybDLvSqOZ/kkGK2uJvrG+ikPuO5
gvwur/RsKO2pSYo9mu44A+78Ba4mHW1DBrNpH9Ln0UNoBEMYcyPyX/T4RaLZQnDbikNigKOlZdVj
OvwNwXfornF3dsd4wFr6sIzLpPlapQeCmevlG+2dCzxzXDuFkYU2USx3yOmtJGrrP1qY4PxYFWKk
gW3EidMig6WVIE4Q0wVliLCo56GA58mzHuWKpcFDKHqAixQpX/jtyJiOHyRaB+nUy3TpIOD7+0z0
wTYLgEs2TdSNH34VmmybsbUtFhYOpL0pnYeODV4nk8DfC+iyHBI9CbthDv2Ixab5DtBlvq02LGjj
8ptR7Poh/I2QYjaooRjmGFamX4PoWvrQRDSO629jBdvHyOebeApjzUGgxxbzRZJwSx6wGI0szt3n
lIT2TKvSveevQ3ya/UlzMs+zNBCFKT+1LMXroQM18JqK8ApQb5JMDsLbW8zxV+OfV1aMd+vyQi4v
Uby5J4zhCWYgiHg8Zeh2zK2H1+bPy2dxIkWtcbBOcoypRxFQAMpb1nfaidZ+yJrovmEAgmd7cWT4
eLvu11xEoDIaEDNBTJRsAyKXttR0UY4wwlHCoKU3RuT0HvL8c0r2Qmm5PjMdgQSjsGt/qAyDNdva
JNgQ2FFF6Kkth0o2LTX4i8o9ergEyoxwryZNpbjlZahUL4XquCzvPokQujTSiRpiRbmPL/2uik+Y
jUasPgnDMq9dXTXb+y2nR21n+/T6viRqERrGC+pwIOxK2TS8kXys9jReNaYd8cDT5ZEJ20+v9DUf
sz0QXueAGfWdlAVcpb/7ZLyDHvZaIPb6mch9LD+VQ8t6ZPI3DbKHqqb46tTk2H/fViwa6GacYTI+
+hvEbEH5Mkql8TMAhFMHGMI2DfgO0VFVEMu0dity9hJGCETrZXvl80JGbENtdWsYm/kfABkujCB0
sbCk/0CKBuO0/7ajRbkAV5idJojIZdfq1cg6F6kSMjlXleASYgW7QobQ2hf49N25AhWqA/joYYeM
3zl3/YCQv6V86GsSC3VD4WK3yXkAdl0ZH/dL9K4v+2MilLwVdz8agaRlvVz7/k8ZQRtT6sOe/40g
8VZqujLtvgY0t3KmmIIEG+DKc+dzW9WbF44lFK+0oxk0lk+mC/O/LS5YeBiHe2eGLzdLOegKm0IX
Np+m2nGnLhpqVU4K3mCEkxjOA37BKEw/ytzxb6eAioAkuCqz1oqkeOBGSka1YaoDU6BS8XAfI6U1
YvvVgcSKnY6+TiS2ua/d41EUj8FRTTiVlz/DqkBQDFPVJAfvV0EkO2FW/Vhv877XlKqNnRiIpx7U
l9s7mRBkkO5loEow1BrgARWFzXLzncdYnY6++Ey42i5XFLi2ltarS4NHekwKAD5ttmcziLoImiII
MQRLwsXZrs5dcFJkqiPnNTpDlynbsCi9VODV7uzUYi2PS5qv1k9XmhEm/qalIdvB0t+u8lyotbkx
Sw5iGGMrm8ctJqbzP6sIUjdVUJGIHymCjmMFDHjTbNl2aUdr+1E+o0DZvSTWG93dDi4So4No89md
Ty83aN9kzBjT4cxQDH7fSvmygKYPoVCdD88QQPNhU40GLzAX6bIY83skB679GIxp1eGgC0q8PmPO
8hcpdqWcBYbFZHlqD6SGVT9CZhpO7TUETbLDXcvRiwCYg6HJsY5VJV4HRIG/6ahMJFUoWJZLXsYs
1DZBiuzH3fVBzlZ0h5OpGZX/mGkJGjd9hXymufJ6OlQlBmRn2bBx1A33gZEK59eSR3VIyDQAztuc
CrK0wE1Wag8yhElvYUxzV9ZCGlkMaOhafApmmcw/LSCzvERKRUyGgJOCktRtOno1r/fICHFlprNL
qpVCwf4D08Rji0+BHoQ2WxURX20E+JqIaFiQX3fOOm5ltZj7PnKu7zqz3V9VR72vwNpNgGGwAqbK
YJCZ1n9PBsuycLsCO++Hp2i4Qp888sMGizbIPXbs3eKvJJ9nnV65Aq3u2GIi8DlCcC3scxH/jW0X
R4hokk0QFrAjs4OyhzTqoAeyCKerGRYqD5x7lznCf8MsxRBEMKHEqFLozbXVVinn9OitcsDIG6p7
RHkR81v8VM4jTW66Y15gYJJlI+yuGMKn1JuThd9iMq/+TcN7SUU59T1bRppB7hed6BZR0zgt9SxD
aTZLcE9UzG3KP7ifRVsZ+VYsvfEUtgfEXyo/Ulvn7zC9Ss4Eemwp2wlHlZzqVGaMmbHzYCFKXXP9
wmNjRR8fONrYLoZWbrUWN4rCU6KRpJUUM321A63TYgjcK4USKa+tFGtQN5FbP0RIJbWK6tBmBLAH
k8X0ROKTo93AanKQ1LJUfJDKPP5bifdUBsNlMszv4pMDQKKpfgXkhlkDa8KKvboMSiwP8Sb8ijZa
svXG2532NYOzlnb6cQA+cu1pFe3wf7yCVmzPcMj4KfvBWvyZFivcu8Il5XdaKDmzmrs34zMxyx64
V39CIYLAbqyF+CK/hAi6/qqEcaS98F88osg0kkn4ow3gMiA+QLCdtkpFC13Vw40/QFRN3Isc/8e5
tYTZ6rltPs/f+UbIm38HCLWwd+udfUUeHfLZY+Yxkp8JWJQFHooCgNOpaHIXhnC7wnCcImrxPcP4
1daTAhcP2sqRtG0p2i7EBLPr2v20KAqi3iQWgboX3drNqQPwDktMY5cUPnsnNDs9uxmSy3wsX/G4
cPKZjb7j7/IYY1XQa8+TK+yMcdSaWnPQkRZZ+e4Uw6hqXMCWv1V2QKXi/XjRj6hD59bN57dJA5VG
3CiKuUy+Lc9ptmjiuvn/upRbVrgfoc6oSUc8DREuv3auTMOHqAzApam7WgMYXhick+SgL0OSSbh1
6UeL9WPNLDMJ7d3dnmU/39S734rR0Krrke4YsVoiMwha5Qdzzo20rU1T9gXc+2n4Ip0rtV/e+G9b
qH9nxv63Yn27W0iXETd9LOn0DhaDToF6M3lzUxKVe8Uc3J3L0E4WYvIUqTm7q84FJ0IUnv1zUzp9
sJsUAiMsRvqfARHxg+w09Lk8j5CNY/DAzad+MiQCA1Txxxx3AppUldqjIi/X3vStxrHmvksMh60a
aRMCu+06jM9QZ/P3WC9aIRIeE6UELoU6om1FtAFx1g9UhX5OHBsKoLAl3f0cc8/PX0+wJB2cqTuN
Bfe8zaDAEFW7Z7JPh4j/0IerQ1fUZL5jZc3kYa78dwr2uy5G/ZUYQP8ftuVI9kOy+IVnil5m5MTA
gUeEzEXaRMXdJrWbar5cLrQ0npuoE6VoVhAfK1CLSGAtcfb5HzJVOzJNMH+WFoCsYAeOTlndc7ds
jHUg7gInjDKzkqDG4kd3R8p68BWu4BA0pB4aRXPKgk1eRQHEOkui7HudTHOIcAUVr1TAVHpwqfce
R/VHn6XImNshf2VILEb9oJNhaWXCkiip0wEUHlURY3y13I86OM2DBhuIn4Zpl9d6IcA5Hpa05AeY
UzcNkfvbAVV5hijQgHDRIviF3RAIRW0l8/55lLlXuoNWyosPjC/rh7acPTUO0wy5Pl2kEtpPC0i1
tymw7YGYMWZMGAH3vlpcea98RuFIFnensc5wrYXb/bA1aBjELeDLWjc4VS7ynOYHGHsTdXvhju7w
uoNHXCWIXEtpp4hF+MMC5hc5/rIKSQr28khrOY2PMw6bpfF2ZRltTtM09boKJVZmczjdQZfAFUm/
DC+cgcVygaPyIq0wVSO37wwINrHMITAH6lUmu6gU2JSTRr9QumcO93BabVL51Y+bkkACK45WQTNu
1YnexJZs6OiXMd1Ftmu2agRKEfknzJAlpames9/5FF8dhAae4FgLtCixlLQF9O+zqObifwOyE6s7
O/X90LvnU7YwsFy2hqLyStPeygx6zb3P6mCsF4dH4UjGjJc2t1WNObJ8Ka7PL+asILeGC36bOXDs
SJC3e9kumSYTiu2UA/gnHlFNA3GP4KrHUEZ17BiYTIbuprG+PR4XgrC0/0NOxoiGYjuXVGts7uch
+5b6/+5EhpdUbwQ4Yzx8Sv0xs9rPpVwMZs3m5RegectTekEk3MvjeDegMeD17HlHEtf+ZAsmIK0g
cVW7PpGzf8Tp0qTQ7RnLQ761zwSbFm6fCjO6q01kSdzdxh/BE3vn3xAXBCWAaTCgIl3sLa2nMZSG
WVGFwGeUegAOcuVR+lCDKtQG6/cy4OuA1LPaKGIyHetw+glAc2TIDM60guASiGpd1+yFqJlGSTIt
nsFo8b5msSkr34JzIrrSzqWAiH6FvbcpiTlXmylQ8LlkFbMIe9tsdIPWB3gr6me977W2do2CL1K6
wd5gz5GXJEGJDPOSUjd2VQuieRLzA0Qo/+UdoYQpQ+2tFcBRiwH5GI9U5zgz2g4fUdS9hiXStwbz
58KpiTtUzFF9NM/daEy+3WceUGbDHRTpwF7ATyqt3nfo3HY+vbnp6jQC3GSxGC4pNS/VR6wQlpp8
v+ui6GyIpY+20uKg5FKCARi/vXb40TuXCZC6zG7QaQvm86TbGfRK4LHhHq+pBwA0ip4ppTICkX6c
hnDoQUxENpwd3T+cu17IsqYISi1FWcE/aKL2Gb8twPErjC5Zqi7xaE3xrOgnUE5IuPa+D8G4oowb
6n43GmGlu/yu0qsIgBXSGCmvzGYsKMF9JAjMx4OYP3QBuQL1YF4fUmPMsCTzMtZpf4xv5oy2Qr/7
UBhqhox841H3nRjGQKUPFdOB1vkKWEZId+fRxUAaT+3CnrWDGAWZaQFuwEdfump6vj9EF3VFBNSK
SEuM+pm/zwpAl9e+2LlCdiogn23TbrSF+k12UHUOwcw11mN1MDoMJs9jMuwismvqGbRC0kYXmBl3
IyzV6lBbIFvAwVbiOHTZiwZ1U19zydS1gpj+uyCysRPW5qIgdX9w1AMvX5rsqxHwCOV/NgnuglUJ
5KtuLE7IYjox0pzRAQpXO9PG8JlBD0WZtADvQrRYNwXaf1T3lh07eQLIYMr7sCexZJWbPjG33uoA
/63qcsvB2Y0XJXBpxTPMU1PyKZy8Ix1Ur8m+WAEPBp36Jn3Eweqn4om+m7FhPO7tmk6OCnhtsGjQ
ElzpV8Ii+wrOC8NsHfM4fsyUycfQgNP4gSA6UaupsEkHPdTbSULs85/L9WWYVCqqwzWk8KWeVKHr
2p1nLNilk2AoJqMym9yrBSBBiU30ecTczg3/83SnMZZZjMJWsED2mHfQyYx8dXBTcfcaZ3Aoaxbf
XbZ6t8tIbqRF1t78hU+5YDiV1lCYbkIXPPM6YRjvJ6bHNC2kI9E8pmvoXVogMAM8YKhMHCnF0BMW
Nr02Lr16//Otl9aFGNqDkY8CVj8rIcvbWduVjcAJcKgyeghfZhluaKsNrmV0tccREJoilOO6cihN
G9rZNzJjQ+apL05qXxVs8jsr00arGMbv3JXMkOd4+ChEJAmURXIsvEzoPHtJxEre0e/wezgCQ1XF
3rPxm9j3TGWSyCJpkwptYGh4UH+i9p3Y1XWi2Qsccsp9hWsn30ywqJAv0b7FkjYyWvcceRiZWTF7
ZHonOloHFLvfkwxddBaLsc7X4R5Knnejo2ygxQt9RLhcvu0cDsc0PHlO2IHcsEV41fYKre8uAafM
Zntk0NX+cx6ST/7PZQYwjaeOmZlRrblFRAEESx09FJ7nUlOEEDEqRDrjKLjvBPr0a65nmQ5zyB+A
V/dmDmHmDP1efDt64BcSo+OtreDioX++w2vhRHt1es05Vy6mWhBm8Ra2/j//VjdA4SZr7t/9PSQ+
5QNPo5aAF0lp5gPC3OhUojk4bwunnOsjGsXWU1feP8B9mPXaiJHWTyLf0LyCFnQJJKhL0ZZeugwE
Bjj8laM6UG0VfkIkcYIQQZ38Uha1kfeypIo9uZCQJuZEaqaGFYUr43eo94BwDsO65Aoo/pA5ivrA
qitNqKHHhvU9/Qp+q87MsG+iuJvdkan3G98Qha53v8VrA/UTvmFHyEHUtsCRfwVJ4FUSXO6J9cDH
xfGzbIlxFr165PNf3MtTCbuYjtQhV2kuOqwx7WvO166uWyzbMy12+o7Z3PjRUIabVKfzA5Pbveh0
wlqSqoS2/tO4KnQfs/BAJ51WhxrAUT2sFFEYVUmcY7jEfrKfewXc2p+T3feeaimwCr54CnvcPnXv
TN9wgw/4h7qo3v8BROrGVX/uk2cNcb500dCH2TzwQ3qf6WiA/xm6UtizirYE9hZ33oxaZmdRzzfF
vAABG7k4gVk/Y+vmsBUT1pZd2gAasZRGoIntMcc3FiIFFQR9Rimsk4P95VX1l27GI0LJZ14vD9gK
z/TZoYPeWOoaIqL9aYv8hGw+Sdi7EcCFGl00tilYxHKStOLozaRp5g2+fBZ17mmjn+AdZzqIFk79
7hlBVtGOLtn9IT4GPkL2whd76OuQgITN3QauFSRgDb45kp1Z9b6TW5jocOVehSftUqPKVRSFjhEU
yQw/RdJtE+CNmpKFaYghMn+kxdktJULDuyxTEpcNLsqZm4OZcxaL3O5mokeEjXiE4X+MvH4dRjTZ
4vX1BMfZYOSE5BqwqjOuTi4Q59gjs0XxKc6JSWLTD8Q0FsoRgfavfKTmxOWAn85ouSp8xScvL6MX
COdeRvx1rM7b7UClrnWQJzDE7RL5jdsJIVofsUutscMXmcZcMCzaY6dMPpt7kZKZv5MDBY7gvP5+
WT3QgLBqclrFpZkPMzmslS/2jP/V/mh7ZIBXM/7oSicVfq+7WIxWQjBZpAyNTsJoNB//IZv2p5f7
+bWJgdEy1B8kjtOU7XOZuQlz5NL+Ldkc3EOwyUhPs2qatKp+KMKZ6pHIlcSLpZMl7cCPQ1YPvffK
xvxwqYlep2uo+G1ot10VLpA4HVapP7bxUCK8HfO+jZu4ADIUJC5oW8f2YSPtKfmi70oJRIGK3j9v
koZKr9sLffjKNy1g8mp8XcqgBY/NRua1T9qfRI+UJ29Q4WouI/VUxzlNb46YRvsf1ztm6a8cIdTZ
fJNr3PPJurniZNCvTQlvJzCJZuXw0Jqtf7LGJUO7Jjv3YiYJgfqCQ4c9FguT+yew92Mo2SbV+Np+
0j5J2hqoxhM9YMIcqPVm9j7l9zGEy2j9kqyCNJfHhYnWkG019QN01fSz1dfTghx4HtzEywzPxw3W
l/K1+ffKxo92AM+5KdGvh1CRd4KUYtIPGaGPPde9turjTeBc2161ltXE57ukx1Ri8U2Viq2D7YGv
uGsU0OykLiIb1wnpRTUtoeWeNt90Rdo7CdwnzDiYt43AgjjlFZO3jS7rEM+0rcxHEtjAwInUiiub
xkigHux281cq6UoB+Hpl0bU70qc4HemQxFV6cIh13MosaJkjrK8CugIG8wSWMr++8Y7bvuadJH7m
/odMYUft7BWu5HI2WXwDG44E10IcuvCaGNtqFJHNNYWkifAZkBgJNTGtIM7Gk/1NNr4qz8o0wSTh
3JPNxpxQwnOkNNgBjS8kxUQtJTc/LZOu+UO824CQs5yNBEVUiR6qH8wRT1JYAr5XQCF/PxSx0vzp
yXs+b4myQUbLr8BDBjekbbfMrchrijmWhEs4mU4l7dJE5l1cBeYt/Fu7VW9cJ+udSoXQW0y8WFsL
H1zrcEDgT+21fbw/QM7fNfShw/3LEJeQBkbLA8+gX5DSHRD86/CXf1vjv7QOPPIIKgaEu/1FPYUv
Q5MJv96RlEp6+fiTH9iSUl89wXFxNVG/5bY7H9KCApHP8SjQ8WgTj2ReH6fR9BVJCZzogVrgKt2O
lQDeSbt29ZaZY2DwHg+P8VrQ27Xwp9ygeVZVUQdMWQy4x0QurNVOzDY2I0dy1bpnpV81iaXK4oo7
WUmta6SKCYQSYUFK0kjnoNWxIugdMUZ8AGXPC9xR2SA3k3+jQ8qPGK6e2AEpN2FiJ01QzqUU6QOC
mTWTOOjtSPbux96OaCbFNL7x4YTVxtfiD2l9nY6HBik2QvM8IyLf71rIbxd1JbIMbhjktlaKR8ea
bYKN+XP1AdadL+H0Kxj0gJXnqX4V78xZHrcQKIGD30FISqHbFXZFUqKu1WC2jqkc8xQRS9hTkVoC
lDGiX89kvfqkvLBkVI5e6ocgmzmyKEti5mROf09EGm4GJqBUM1uBaVehiyNc9yoYCFloOCy+AfY1
GcI17PeFqE6lRE2Swq0XhXA6rR4O189VAX4WkitgdkhRXNgGNPYVGzd8n4PFMDggZSK3uOA95LN+
1S9J3nhA9SnBhimiXXVeJnLSEOVZEUXNw/TRZmEmw7NC5i38Pwofs1UO7GnTeKJDIh34os1G08uB
uo0JZMCdzPgO8mgrf3oDQToB5+ErKIOCX4jUSBkndj6k0NnCU6HIBoY5i8xW9+iMZFpiiDZNHayo
B/u2SmGe9O4Dnjjf6JyXzznQz4wUL7zbor9eBvgTnTp9wD1a8kns1rPjNBtu4HiqCfwZC+OJCnBv
jwTsEz47KlQkAuqwY9f88kHYp+o8QX+wS0Qw0vuk6B+GzuImmyfBidIyyE5yBfRhIq8SAyR1gRSu
N7fpsEZ1OqHKmO/C6utlMhfWz5gVyIz+/NXhGE8a5eJDYZWqLcXfnW4zVNFJzaVADT68FAV1NbvP
6Cp9IcoBk/TE48n6VJhUXWuIyRVvGPojxznAAkFKSAFT/LVEb3dTC4Bu+T/LMGrAhIJLQPhKo3yI
yGZjbVBtZpiQB6s1LlDxQsycPP+YJ+cjWc19YXH5EPIDQg8+btlcfU8/yc0ivhCFd3l/7C6YK5BT
su610kASRdbGuyDnoSpfO+YPq8FYY7ZbB1N/4uMLgY2QZh73LhYmRfsfDwcVm9SnjmWTYowUdV5O
JPnmcIabbW0rVbxuf49sR/v2sSrioNM6WwOqPzPqMT8hk1ngTILFlqmlYZStuYxmKbhRmsoN30T9
wmv6Guxcl645KmBJwPFsHPXR7X5tXYZKtlL8JqUn+eNJG63dWo08G2426avQYn/Kj8Tw0mdIZqu4
pGSs66VnkUOOgvGFrxIThB6LLH704Qj52odFzXFioT3xrmBHwci3Vf2kvgBYKoV7/FI6G2lxqdux
alC88Ur5m28nkrDeEnOp85XWNUa1OruwwE08dfNNa/MRoFOFVWbG+9z5L5p7XYzlALgHW0ezHWH8
oX/lTfDGeHeIz6dxdzh5s4MP4bws8EftXN+z3v5srFRb4tPIB8x7GLOqWE/YdeVdm7rGY0tYis7D
9MbADPlVBQx7JOZTrbmYdBVlQhscsgezTZD5g4Q2R2w4oa/SdzUU0Ad/wa77egi61Z4puOowVywX
GEsteL8i3eBdkEI+gjTCEXHZHmQlhzNWPIY0sH7FsYb/kY9hTlz5Rp0YPwzjUbdNnf14apel7EzM
GvqXnK2z7RVgLv6SmgneAlXH/vWTaGukh7vqNEvX7yT1pzgFGtrCoHOocVLsO8c2HNkVf5eoviZd
sWxOv++03kqgseYM1PPD44t+3JqW9wnavB/z9lnqfr9OaXTZ7byOHqok59rvFtmETOEXgMITn24N
87NG3zDuAvr46BY0CClrGw6HfsqSlVS8tVVnSRgGg/ixlloAi8OCFxCnUDFW8XkxVr8Z97avlBih
6J7fJ24O8gL4rgcik3jr92wl4EubpH7d7B88bNuP6CSYVWzOOCk51rilvElo+aRzmgEr9kZWAYqO
Eo8iBZhRspvlk4VpV9BOk2SHf+hPg7wwbIj/rYdqMyF+j2+1a98o/zN2FJ2/q9jIIp9WAKsbypCO
WoASHaRxqGLJHS85jOq0xlfBECrU0yCG8L6FPZjF6YABtnFNCAzZ33Wvpb9I/0le2Dh9xjoQ9xS2
6aGXv74YjLtAQqMQrFLFQ64hoD9USgpCle8jLxMDPtdj+WredvlhlH9auefR3ttqazHVpmqcISjd
qfi1m7SFdKhbaEkfcNS9JHVxbtzPVBtWSEXGOFXb/Z9onmWlswfX1DH5SiZxdIWZ8Vy/0pvVPpI2
/TRu3fFN1g3oFH5p++8NQCScoxUFQOcg4ghzGUp6ywXvUV6VcSHkc5YX5TwKiLzGk/wJwr1rcLKG
g16FybN4Y7Hn6OMXKNs5zIufd4hgjovIuEqucTw1aln1klxBbXpRojjsms0wpcxWAvBLbC38IXJ6
uQ/cyyWCb/IGpSE8KaKLMA6m1/Lh0rkJ3aj6uDNf4oYUGvMYWQSM4YoGB/N7+fpgMM1vxSU1zB3L
cg/B4KyQtXk2tvC6gRVTYjsRQ+vDZQr3iwhubWY6yVsxZymKODtqM3awLQ5OEC1SNGynRr6CKWza
2OmmEHGq2i6HdNCCqVpGEdpKeVhzlWu5Y+Xf5n8iWaKPk8ceqVgIbDhIhRAOHgdtW5IGc++n+lbT
N1sHA8NgmEc9YeSKgPo4HDJneQjzXBDcza9jGLR80+Y2wdGV5Q4VBdOlUMpxxQBUovIyRM7LHzGa
mgBJEppwNEi93OaiynnmBs5uvFhsk6+PiMXDCk5eQWls55hRDkWHkRyMG4fwotHdfM2qzTOTz3ju
+kn+rJ+RGVGF2WecPp4/E0nyk2BUxQwMl58nyyb08VdpnTNtbV/5TqPwMOq90qGXOqJrv+Cd5dAk
xCIrPR9C9j8cpacUi22/gR4ebw9aTwbjw+YBoGPJRGAKuly25L4UX076NNNew3pzdUtGLYYSF18C
faQHejND/YOWjapZsPlJ2L9LBxHkRmtcDtad99RYHYghCClAmEGpTCYJ9oAdpfZPrZYR7doyeh1N
vKVJBUDJeqbKpsOPoASqkuRpyY0NVFR+vwu3rsbsedBQ5X0wGpySXFEhuXdeEFhqSVBhboU7lDRs
ba1R0u5Yo2Jc4FMjBz41Fj7SntN42X8T5uslIckP1qwIi/d8E5ORZXDJbBBLselVDYhH6aE52ZxG
d08WJSgY6BbtOeocBr0h7rfQ26DT4TlrNaNdp4LE4TNMb3BRTTzXgIMFKK7o5WeT8sCxP9ErJ5Nf
sXBjxRMqOwmcxaSxofpoaeLpV71Zsnc0Cj188EacGfD7uU7oIdsB/1mHea/NRC5kFUFKsF6DjZ3+
qwy2ycmO/pjv1+3aqXp2MjUNiqEHRzA8UuRsns5dVRcajsySpnxCRLDrhbhQ2naHFSIpcnF7cwjv
5ziLo2QAGTZroOdiqCu2jD521s5hV5slfCTv1QybEtw4ebYxaiiOnkJabtLsjqOkyQg2s/GVqYKc
rOyeRw3f4ILzDeGXy9NpVCwfBdEj+IPweSWWt3V5bGWfo7lkjmVnE8LZVysznP7PRbRs393jTw0/
JHXMbvEvjIIKhJU2NAtuUc2+EmRdWH+UCTZM9lA/cORycIfWLzL6xzrds1etCKOMTkoX8yoxyl4v
IIz+dR4uiKNqOLPMrmJMU1ybb7+H3XiA/94LLa6VBjbJqcE/a4FQcIUbR3cAOqZq2ii+AuKlbb/1
aD/tYL8ArPDNr+Z0p+iU0aNNbV6XBCU/3E3KyxGRpJA/wmqzn73Po2OfKRkR1HTdw7ItlDOLu9Xh
O1xDBIK2vi+Ta1yrkRDyVAz5Lu3INHRY67vHq6WK15B8oGE603Lo3CuHjlaC6RTxd+FbO0Tb/hFA
+TtOZhRFXK9JITArEAD/2ckGd7PPdkumcy8UGhr/OvmXKHmtTzAFSG44OfVJGi23g90NwND7tgi2
+YXNABkG4kZuB+EFKMVQ0afr86lSV3CPEhFjbPQIunhpUZ5SBaYz/dFSbSOOj7cVajakAoXlnQcw
JpngfTBB/aWNDP9OEAZiJ0b0+JjGXUx4RsGnD5r3uGbqEHcwyjtP0kjXU+GVZmQj6WJP4EWXud7h
FtSHENvLfmFRmRGsp0lEySwQe+CnCpf/OMp4/P1oSZV5BSkmUkcRYdk6uJgREFV8llFbAMS4gjhx
aFbTD1qNKIXyvYnAwnoHkUQDB63JGQSIy/bpj3ZhDt/xMznHZst0osE0gl660DlHNKqey5wREatG
Xc5WaQ8XmAqDlZCbKsC3VD+lTghWU29i+p01Hwfb/gypvpPddPh8y015JYzWXgocvoU9XPYNW41J
3dSoT8J/wwveYbxSx62jzxlBnGHFtyE2uWhf08Dhhfkqd0OmCAig4/0906hGvPl2/ktiNRyYe+aN
s/HMU3PlanG0CumlAflr1M9/u8EU4uNTCqQB5/cuLZGPdm47W2D1PN8DSuJXPQ9vnFNbIYkc+Xmj
bxQMkkhrwcwKufT5HIR9M+pzMLycmfygAX17zp1WLKdaPaYWDp0WdIIkk7OqMalXSCscB7WjLDBK
NkwPhnwJmJwHaKRqHP9RR4AVwy3OyRfdkmrThNAEQkx9DchXiHqahEmr8VEMLcwNYOpeBIWTeXWv
CSajJxUuDydAK3x9pl7ITO4EHOQrxjvsBR8wpf9fikF4EiyawO81JjR6fdBKac5Z8TI8Bs0MrLoJ
esE/kn06djQDinVezZL7kwrrcIWHQk2WYJxl73YcaARhjW+DCSg+wI4RSvz4TZ3FR0MFTArvfvJ9
kCc29lDecMFyy/MmFcLSLr6Bd3nHqZNODEFJ8qYHae6jupJHeTAreXBAVi73kmksHR9tsIQzZqD9
qBFL7TrfVyGtWuIYHwImbGW/StN0LGzoalp0C9Meb34iO4rLgUkJf0Q2PgnMcEQ/YZ6UBsrkNh06
NsnGPAYSGAZpWTMPICthHarw34vvyUVwejAICPEWkaZJ8ziUomhENQy9exzT3jVHa/aQu3VnA1bl
mz935bo/Ug8dzv0je4V2Dn7M7M9TRjEG6N0OZRvYoVVDceepvKDqIM7hFol3UMKxCIzt423QAcxU
Z+VMQXDzGP8iO3H18W84eTcYUHED/Jt4sOzA1kNVuO8MwGHxEhIvNnuqpueEg1EitlcfdWTCiyqp
E8sPhNe/ZoApiG7LSVebH9XpMb87UNrnekTIlBndXZ43hB+HDQlf7ETEBO5e7OPXesBjq/Ctb1vL
Z9Qu3L/CY+SaTvHVaSNX8Ai2l5kV/0pwe3U07NvHawGIkLfqAXGLgxDkcqBzsrZnFkSsDMP8BIwH
DOkNXy1fjPw0mDl+VvJW7hPLJRiHspoiGccBMmkaGEQWCB3A49LNmTdF8NH7buHgvRpau+efSkU3
mqkpyAzaDvbHsQZPZp64lmUhJRljsmfjxR1ysKOOQPS0dr6Y1a2ErrVh7s7mypMMPZXgNP7h4YRn
p9XJ87Ds+uAWb86Jnk81bDbLH9N2CG/8HRbzwPUX7lkIYQgtADX9EvDn9kH3cWOLpQ+G1Q0/K3vF
hHHuzjtP9KxV7TFyBnO+3hx39l6C2GU5wcA8O6p09veG7HsO/YDrY9vzTsw8AiZMDul6zCfB6XaJ
deZ5iOoKlGnuacUjXP69sBQ+OCNCrEfFN3bP5F8ena33hmsXJBzhta2Ind7TN19H/PCOq81/GXJV
MjhjZJMweLdOMvH0O0LPVnwtfJVJ7hmjePUsHymq7dkUdo0gZZUagXaKpB6thdRZZJKi3EECsCjP
CWA1Zyck1o0bQ1QxQ6nJ/rl2crYQOUG6jWngaqBPMfQGN5a9wjOnBDyciRav64oPYXza5s5TznR6
fnas5u320Y/hDFJB+vpDJDBn01YJjTcAMoZ6Ho5TFQ9pxhZI8eg9HjLxM0UFPc3fPNP8PfZlwZ1o
ucUQtBu/i+YfC2KCQu/xCGvflmBmS1wIZYrM7CEBois6rgjK5jRnPxVI0EbmfZ+bziouaLCKz2iL
4knHT+Oc40+yyvVUCeEOno04XVr1vIfMhJN6jLzxJn34RaSf6U9ntQbnmcz5jU4yKyY1gC5JX9Sb
p1njzO513/iXnBlhgDfRP8Uu+NAPRWiqrcYffohexqufD4d7+a/VoEJuChtDSjQW2w+UYwQ2SWWD
81UjwPLNslf9EtUb3hSr9YAlVEZOMF81CbFyI/ze6faxjz81JcnN800UhLeFt61PYLHvwpDB1We3
ZD/3AXhwXFw3PAHol96paZ38eUS3g5w6zwIoyZj1HgEHCoPqAEVptYPcu24OPYbrIBPWD28Kf0h/
cUb+j0L/hBRdsyJNTsagTF+BxiYmIha+Pe+0QSfl5tUfuQfgAmT4tzYRbdBvf5RAl3HPMSZgAd+7
5eN+YCRIuYSYpQtSggMbgF4jPn8aJoi5T0UgieP3qSkSTI5Y+VnivGV0+6Nb5UbfYE8R38bebdi3
P2T5mNt0RWv+D2LPpmACwzOQyeGToKjD1hP5hW1owtiU3Kh9BaXG9LjIme/kcMyULZkmUvcfvM9P
/Olmz+Pk0hzrtyViyEySxZW2MdmmJ2c9FRiuvFP7btzEBXWCzp7kVO1+5zw+OlD0K8rLvWqwUBRQ
z9KBySb4HyMhUsDkimEHAoPAQ/AonQwJgicQVyQf+YXbmXE5V8lOLdWHqXn6kBYeCjOTc25Ie6kR
FTK+iHfYjvYpo79jy+bQXNnEqGENPcKR7pi4prU0gXJlJzSKWoWhSeLDq5xePhZpHYA4XaADb+GS
yt9NuSOKzq+YAHgzq0M0YDFBLXfLTV7jfWRNDHyynEmeh+EnUx25waIJL2+YgHGLCSJg0sX1gEdV
3+nNYvydAXp0pDy0dQRq79nXcI0ItgOLJY5PPcZ3RGWNxcnj9A66BZlP/8v5WZQPvVZ08lQJCrM5
JvW/S9arG4gvInKT5O92eEFvBP5HdTeKDhvE6Ge/KEBJbgT0kaO03Z+aYkgx0iA9/hum/gohN3uI
Dz8qEukpC3wn0NtkSQMCE8LXAwUjgx3wq9DnDy9iTgZQnuXOstGbp1ukl0fZJNC0XnHhs0zge3sI
46V3wQnr78MlpJEZd2E9XWCRBvpd5O5H7y7Sua0AFqSY/za1CPkEfy5vxL+iCr1RtGXxdgml6vku
pbsHlurx9EchsfT3WJgHPPm8GQXVZPSDb8UPHHViMsvfeIJBlu/f3k/dZlEb6HWlUpudFiTbVNgB
hlHVt3+FefpDrqPiPJtINq0hBz0iEwG2YnrcpXVcoFmjfNC9hz2PINg3LI9Mg1mMVyYQBc0WJAjd
5/Pn27v+SQpsG9eBeiuxjbnrqxE41mTMz4XQU3VmUbm4sdtZCZSX6Ihq8QKvHSUcrkxJo2CMb/ii
7UuOZzQKLSJAFVs4WcTYQJpvAWjxsWz5xDyOs+dWwtxLYNjgHND/Wz7ytLf2ZIk1igR0KidkjWsv
sovWlnZyEj+vnEEooymdRtObm7pnSWhJcuxB50G+1kOeawDvC0y8dXHvniAvla03blqf9rmFWQf8
ZxuvqUbYwAg4hheeOjdJKgT+hW3Z8gOqNpKuqyaZcvIzMS8M3cS3Z5pdfO+0rJoyuwKmpnWOfCHJ
ysb7664q8nNnox6Z6WnEoF9JHAvKD5Qy5Kg2g142oLSoQEpB+AAsiEVj+hgEQtZj1el9yhnu1DNB
u4bNuAWvrTa0MdAVVTiU5RQKK0ujpNrlaWsViLHe0LNIUf/XK9DCbz1ngLizGiqVoWWUwHrtWA0J
XXfzj/9d4paAgKrU8chxKIM46z4g3PF+QUDvAOkZGcz8bKRj7/5Z4CE0v+Q+lMc545wntWRJcmh3
X19Rlu+B+/UFvj3UFmzP51KJrCw0tYYZt+F75CuwxcfFAgWT9ZGmRHVmhGw6QGFtR3YqTtEx+xfX
WE3QAHPRf1aGLzRpffnzcU/VtkXrQr3SHPAlYmz2zKAe032fhq/BZEEwywdmghYsWajnJX8AtzJ5
oSL/nMMhoS3+LCTQ5fI1uUpdkL0Yc87ZRJvq66NezWI3HDybDakG44tmDy+m0k/36pVudm60czOq
zWphZSCUmmVMJr+umRIzQ73rLkQEh4fv1q/IVC4vUkMYg0L0fpuXUigrcfjzflEr8ZVpcQSBHcZT
RdncXEhccN3mzrWWHE30KrkaJIGmd8ntqBEGa1WtC8mF+sPZcgXMHLB25miWPdkl4wnuLIS1Nusw
kQVlVZ/aSxB22+DXAICTmTggjIqaAgg0hrsyyvq91k5WQQYDokMH1AT1gdz4W9oh3RS8cogoT17Q
mm7V9td6u092rIRTEIORcVlvyOt0STsEH04LxZ29IYSzNClh9eXDqUS7C0GJ4GoeKTgBeUAYv5bY
ncZK0OAtuvMMnQUtO4KHS8ds9dKLv6A5kb+Cj9m+kPylLvIch44zI6N3vw09Lppibj2zQZsN312L
/baWW6aGGwp30HdnojiDg5uuu/U4yNO4cvvd7hcstnF6QMuToFhM+vBrrc9g2xj6GKT9L1WJtTcI
Quk93ZMlf82wCH/iLnq6B+fWqz81Rb6nISljo3M2U/xh6ve3RNNy4xHlt3X1kWbLTF8zbPzMfNPr
j4GKdaQCAZf/rb/yubBJJ8JAfLSB2MXabOdcA2/VWGbHK0z2adfelj0SRMk2nHWTzXBQNWz785v1
kqbZKjQmIuBxB3xO3EQFOJ56jgVGyJnLMogMt2Q4IlsQ1n1oNb8H1zucnKM3Y/DIAi6GaQjYoUnd
6YjJnH9iU99VsHzqp9BsuA9zErIHEpNJ8P0iFLNHFmlEAp0jg987af7OOsSFxHLnkRkSpdAGHFVO
1RJmjqP76iGNI2FZKZjJZaDwvRwnfRs54RHIc9lc1bvCAP5lVb9LgMKUMFpe0zGyHzU/F/tRJuFH
/UD+SRDtQD4xJSUthxRW/HcVP1F5tL09a6C60G9C6PTBPd7O9nysu21Am92V0vDnNAu8X+KjfMU7
TxjKcQIV8mQMZmpmoU4Xa+glNR6qIlD3f0WlbrqhRErNZNw2pomZORyAPCe3qTMKnGheXBaE2uI4
jjd1KrIe+5R4EcM4jVyxUjhke3N3u5JUbRgZMX8ErsnRPHp543cv9rwUirhVMtLttZZA0FkYaIBW
UhpCaOOMAZ2io7VmHzggTCpO8Wh7cRp++/4gGkxyNgjuq5vmlcgOpRz/156vjGPN+Qfoiw/kOGdm
XRLqePpWEgGzYhNaf2o3ZF05yJxctpj2+2jPpoCXDKo+pPV80Y/u6fBT5awlt3WwT8SAauGRSZMv
YuknnHPjeLvVM3BNadb0JEdfd+3NEfMjXqekLTfWtHGWpX+kksB9P2e/0j6UEtS3zJeh6ylvM7CP
lwayEqaF0v/h1BxkKzJJ989+bftO0vlYfX9m8ejvF3EYvzH+FgWFuV7mEXJBY4XvWf5ip4pqTZ4y
UEOXtq8iA5w0ai7/U/Z9Uhfz3usD5lTI/ROgVAJZE4Yq5T1q6rx7sfNHXXt0iyVkEEPJq+35x2/f
Yi2OvynPZgPnEK20KN2zY2NT/tNR5GeI+I8Th8S1ndx/wThW9slyO5oYpJH29mUeWd5ypEA+OK+9
SrtoG9+uRcbiA+HwqEko7uykiuVwkp7FYsuwnPTurNZehliiwJl1eQQldWayPDgVgUcf2JjtpIkz
XUdFVrnK441oqcRlG1vKrqU7pQAO3FlSLyTxBEiP/To8ZdISLueLnQEBEe678bbxpx5nwfxVF7XN
G35WHoZM9cF/ZVPlDyk4xSOxfmMTe1oFJ1jJfEi3FWEzM6Fe21+tmsX4xuecioIVeTebA4X0D1PW
a9Zj9RJT+Jv1aeM383bxiOp3J+AO7sM6r1+xrhV7vz8agIvPK/KD/Nedi3salu411Ow7qM0NP/wY
dmicFt+S/lM/LPZejB3epuhJnMxGeLXRlko+WpZcigucuV4gnn8nx2yVZF6j5kRG9an7H9SMLBJ+
5hSP2GjaUkAXp8n9+Via+XLozK1bXV51Ph8J4b5OR9lmQrMVaD37MF8/Luj+9uJCkLe8jzep+DLh
mG735+Yv/ffp2dag8OARVokv0N1ng+LwUXmyUeO8jw8Fb0aSRHsOaRE7tBy3ZZeFV+N8NfMMEaJY
pQQXgYpTr07kntucmN3JgyJXlInHqrCvTxQmXSG2GoYU2CI+NnWH86ljTrKxhFI6fVhoJ/FcyZsg
W6kBllSzkVxLBrQdfSdSAlRpx9ktLLcxJZHqlyVf9fbS9J/GTAtEX7qybh2aaRY7++lc9wDUb4bQ
IbNORo0X7ScUHOC1ktk4S/7M/4pPLzukyfPeukSshZozm3veUmwH7hvDxIaMhIi0eRJIJ0Ydx/A8
N+Y+2+ofBDNXFhW0iuIVFFJpvkjsRUfoxk0nopGjeRIsvac8bM4QgmIq2MLXEd8eGYgtpHTcUP1B
YUOhJ+ZgBB5h7PohB9rzJC5dedyQ+tPUNJIaHyTcKd7RuhUxTZxhaSIGpoCocUgL4ffngK7A04XN
xrAatJbOiePnF7+rxjg63rXnThCxhpvtc1oh0quBRCp9zzkmakiAWP83/ja90/z5oxRkk7yQwaKW
PWhznwsMocxUVtdqR2yCXtD7gqSw7WK5hT6bkvSxOIszvnjuxfLg+HXwFuMbMLTt7xw0oXhQbuOC
SV9a5hzUBbw6UgcoMX2XpFVXgtVwOArxNVY6YgEyleE1uO6eALZ5jhvSR1AJ+2kyouJ119hbS7uT
gFe2V8xhyJR3Mp+4d46dH0M1Hrps9zdP2Hf6OKQ5B/Pko61WTruGIgnmoFG7PFXmxXaqCl62wW9r
iTwsxB1WBiQjLsCH/DbgNds/4M+jALgl2z5voqOC9F67xpewOJ/oZkLGEojoRtSe02w8i1e82q7e
qzGXsLWfFuJKJO2TBB2CzIsMbGfS5YnC4vgsXnec+I3bwzH39RiD2eHbzw3gJH9mq/EFhnAthb5V
LxgR08D+wIttP9PCor3oQha5X6X8jglnOs5JHsi/5FWhH1P31pQIEg1OvKpFX9uqZm1NIbmOOsYK
mSf1/GFRzUmOO9o2I9ZJHZEj8bnIkxbSxSX7+Wk3I5mBDo4bFl7S8tA9akAVNR1Em1cxgWicvi1q
HSbfyLgv1GLf7vVhB9IfZmHMCml7qlwSpHnrwvWgIda7ghApnNPZ4NrmZazDEpZKcPias9aBQXrP
Ry0lIeeUjfiaIiGdJuAYDCbzCLT6Tq43EMxiMCGLkjAsfJI8zOG5URTA6EbP7/7rU5NJS66DGQMX
wB+PFDd/5BSu9cu7Jt5pAvEOyHbsQ+638B1g3nEc6A3QvPn5wYK63xIlc42mzoR64sMCtIPtUcYV
oROPCd9vtO5lOlMt9tETVzYBmV68oVGqsZtqkhwJ2/7cV+FHFQysYwyFZdBdmjm5FGxGfOH9NwwM
rIVLGUr49sz+bfuyK97BStf9rJz5IpvPTMNcvW+m60Pxo9ovZ/xCbgOqaEaVKDL/0uC6qybkZkLk
K9NTushWDixoHxtw2yZd33NrejB36ck7I8O9xH+3QkEVhyfjG1XtF7iMMocbI4vimzTCAj85n2Hz
4fengHEai5M/siD3A0VWBWhuycu3fat6hAZx2IMdVgnen7GV7eSdo1XZvEg4rNIZzwhYGMtHIm0d
J8DxBTcaws0hUOR41wDsG+jwV/rlNwAN0x0Y4IUSKnzA/d65h05CwAG/UF+ZtffPfM7CqAjbO1uK
Oj2Donht/BJamYKTo0xyToYWPJecvwNSbjd2YBqirmSwD7xJpS2HXhkkwqEE+LbKG66TQ2xfIq1g
a8JPSviZ2PFxFMMCQX6+iZxnepdAUX0vVoElikQ1WiiKtteCmFdKP3LfCPBOmoVt8bi88s9vH7yJ
uDLJOMauvSYvlXVL8WOFXBjW3CG5RBRsxWQJ+eMf0AlE0S/xS0M8V36KHURwK5+27vdZce2uQbAo
+//IcQExpHoPhHx0VbofKjriKyg7WI7qj15lRjSqvkwCqFfj6cGS0kOVqCC3Q2dV5v483OcMvCiQ
JMkxKfH2HtqhZmb8Eiq553gwIJWMybvPQbQLYub2rdwDpOmszBtq7JKCpXRt3MY8muou+wf9l93G
5hYuLBnk4CggL2c3SgxHiZt+FA3N0uK0LkVScpAHaI1GWmPWIsT3oh89Ta+s2nYV5XgJNRGnJnS+
/XpcvBEcHx0L4kTxvbnq1Oze2sfkqRu0Y3Rp3F51/kIO7YT2oiAKRo8e1UBNTNvEob6ppsg1+hTZ
Hvhl/n7Y/NE=

`protect end_protected
