`protect begin_protected
`protect version=1
`protect encrypt_agent="FMSH Encrypt Tool"
`protect encrypt_agent_info="FMSH Encrypt Version 1.0"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2017_05", key_method="rsa"
`protect key_block
nSz/MG4XYeL3rO0ZHnUDno/pRGhSnqJ+0T80MXbOOjNgHQyHZLLyO41BjofGWLQ0jlPux/yMg9b7
hvFvuUZMH/Pix5UusR3QE1kvPG0Byea8f/8QpIFdFnqgtIDsrLdtOdCNxcfhmJX4hAyt1p/D8yDB
wJKrepso24pbw/I6TmH26m/F+MfncIYYIcU3/ODv1/jWctGnadOnxtCGIZuQuv/qILWzn09tveaG
GVClDrxbNhCIinGivnrbx8V9vhsLreMdoEzRyUsLKym9DICsSTTKy+ghlcz3HkAQCyUEqg2FAbR+
a1qwIZtdsHedU1TcP/+3zeyr0IGIKLsF9mMnQQ==

`protect data_method="aes256-cbc"
`protect encoding=(enctype="base64", line_length=76, bytes=680624)
`protect data_block
wmLIrQq7aEFVI+347VdEVS17ib9QCA6ASVx0YvbEMhp0fsCd4KppT/SMz5rehCF2DVNXkulk+bxS
1XgpJXoMKhcS+8bwcaxr44Vuu0KEb25VUEAK8tbR9j0RbO8zctZbrGEpUnpvsnulc5FZzp2EzolN
1R/Gsht+NmrOyYbiBgIWwSWmxLIZGRfhhzPK6TRPX8RxjNJ7OC0jNR+PCDQKIhFD+VI9+3F0nQsB
yNorPSb8JheIYVUC3yhUQqrKcQx/h7VyVtoRAOY0wtLw5D9v1+J5k/gRAFApP+oQivaE1I0vpsHW
7jAlzEjlwIdHQyGsC+NStisxPiWepds4SuEtSPqmREClmPx5kOe5+ofvaKWoAOb+/n66ja95QA3L
aDOFF/8GnQOrINmb5fb5aShsO0dytDT9JOj2nXxQl0Yini3+hAeGv+MEoOWZue6XY/ws1mvvWq9U
BjWTRNxkxdTnAgOHJShFpsrhtJ0163j8J4N6KfxImMgZCoSnGZ4KXFgWbb4C3w7eczZf8LzmZGti
riTUABEbnOlCOPji9SgB6bQaXGabs39m12AudkJn+E10bVxoiLhn7YBTTYHlp1ly3QRHTf9zKt+/
CT7kEbAdzxWYNpCptUkJEpGHjhf9zjLtoFnLRgbL95M1UvVA6lZg95hdaC/tRamAJpMvsbyt+jBq
wU3BHGNC83Di95vCUctcPD1Tq1EijOIZ3tmsa8Sr+otHd40TeYXHHHFjv8cdwBruncZM4UzmuflO
VkAwawdZbZR6mZleb9s8gGqkE9slUOeI0j9TyjnDokseesfS4cCyvzWDcVWV1AzuKmyU+AdkaNle
NaPtg9mL2FVgb46z+GDdL1/CNDGawQMHrDRcwMZkIGinQ2wct8Qx0TghD0IZUGaSdJiGwWCUhLWm
E8uMAAiSg3ZAFYRUEj33my6gUNsjb9yBqwNgNMjYOqdEnexxUeiJ3rbVkARwkJajS09VQiARUz3I
xUQ4tkM+B6P/VzrjkEcz7/z42AneU1jJtryslNze7vLe/utIThSKQKCnvCbSEK0tliValjFtC5GN
lXjdD3xXNsXrKf/eiAh0Dve5rYSRYdZ13mZ/rPlYYvaTlLZ81Zxhq6l79Prk6xc6mUJrm/zY+64X
7Gl16njSUexJqhCtkPV/EwpJutTZDsX4AQBoBYVXo28JNb10u86jaJyVVYhKB7IlVAoP94fT6Rdw
eKK7KzR194kQ1Ei9di13OLxSlACdoaWJ9AvirEQCjQy57d2a9VCZbYIaCS2n9JVgJLdlW0ulfJ6/
rMmtv79QRDi2Kg1iFuM/dkvFaS3Lb0DQIoft8DcAJniyKCIi9+2Yg6MVnT7ykiT0d4bi5XNFLo3v
/bwpDQw+OhUMANsBpYXeA+Ynf4LXlJz/N/wW1qsvEwTyStdXM/e8uGlyteCKvOMc6u4DZBBUY832
nxMROaLTA/+ts5htbtznbHJZeS/86KbKMxXsABCtNnEFlHsuIv8BdUv5j3PsIDUAOqaPIFFE7jpu
9YzW4Lq9g3AdPYV9yZw795dQyyfOkoBwTO/g2nHrDOT8lMHCQxRfY1vpbyL+IHVqN0nW9VV5uYGr
U8HYLgGHfGvoNS/r8RnNticdZZO2r7nxDfM6eZbIa1QIUoN8v/S//LN5YcFOBA3H1fBhGAIylxQy
ZKwv654VVtQb5W1xfr11FzUWC9b8rU9bUkwhBwmuluCcXCKeyzqG4yPAw0RaUZfGdcIhSsRx11Yv
3OkfBh2B6OezfPNrrlSNeCZPbGcLibL1QhJi2Im/HjzOU0epb6M7nJMpO5QauILpGwCP4K1aknhB
cnsjOcWQ48DLSJ4LYbxe8xTjjXtNlylqxWwNYqheQPKIua7AHzJVhKA3fZpp0c4y8BFe/QZ6NaCO
44bbNGwNix9MVxZwGIWc/MNqwqG/4OsyI4XOJx9bLpW8OkGEJebJF9QFwwIVqjgRk2LT76ZxK3jH
Q0xM5CwAobfrpU1ArDBFfjDfUta46vbYgZTENKT6KTItVYf+kNTWVK9M6S8bYbeuGTTR7nc9a9QJ
rAdYonRhsGc9UWor5ZlEWXIHF30NpXNdMKfYOOevFdG4rpiyZhoK8j4QHVV0NarQxvrke4hgUryx
nnbxPHuGJwjgLi6JCG6BhPallqW02fG47rMlbO5CImKRT2Inn16sAVuY+OIE794nddJIkKJeuseM
OzRMK2ZqugsJ4cIVLhfxGU/U/a8Dj/DI0Clqzkfv/zUaW8vx8WO0bnM2sKzSBlsHc/IV4nrfJrmY
lL4R6teJqJoHJB9JaqmGtUmGxgtiQTm87WkyG+eQAC00s9a8qyDG5tzwK7+wF/DfyekTOeGymXOq
4/wE2pVWjdZ/JqtR0mhHvJRwMY7tXYTc2iJbt7zNrQlx5n4RL64LSJnDDXxVk2Voqg72LRMOkxsw
o/xNOfW6/5CL+NZDufEUm+CmQcIw4CWKEk/nvpG85zDDZCB7p8yhICwmjWj5yYFY8mFOFNLpqIX7
Dvn4AbfS7aumYU2DZL/WVNE4o+C9O02QOHSEVVg1yzRRbqq9ShBLo/e5WXq3POksDymurzPAzoey
LGtlJZ/L1tQsrX7tIhsPsv2Q49XqN0KXMOVlIxC3mXzTWnCvpwDzWchVS9GrwuLjjE5tO4Tsvj9I
jHQXfp0jrOK3EI3OkGcf+iDuIBl3zRPtpwq9jqUaA/N8Ti6gaw9/vZwUqIfVV9pTsb7Ltr+UfSsb
ZNnAWYHr/eFo5Q2u54oG4O9YneLrN7hsrFVDIShI3F+QFt6AI3E5Wa/vbx3kuG3NjtYo5Lvdygsz
+ECiH34vOuetx4znXTtWOkQOHwjKdB7vldfHlBlIJ8r7TKxyWkrfvT1onaD6J0xeemMpQW9cmW+T
/8vELPCjdcsVjGQ9vohTfa2If8H1A1Xaj712io9A02z6BhXykj2azKW8RcbCXNt50XGu8pr2EiBc
WFHuP7HsbXerMQ/pGsTnD3sGxOc2ttfUtWGywwhFRiG6c9lN9L80XPuOwYYY7XCXSgRVJuiw41wM
crrAFzXcHWWJvpv0e24i3TU0xsH7hc+ExQ1sevi9URukk0aDF0N3MltWF4ahTFZlH1e8qrmeExZj
DE4cVeiCQOf5t2BqE4CkA1h2bNN07FBvJTaAnnAf2XUGILTuiHip562kyQOTVhxQ9xnx9lmnWT32
SrwDSf/xXuvEqbAAm+w/Ek7wq594vAfgK9xm913F38VmmZOw9uDvWFl6P7s/D+/bcWviDQ3OWC7t
24oWxKagtUmLHV0qETjwI/4gnSDOlaWwRKHCGqzlVEO0/jx6cf7yNmoRepvuGieYowJcA0SCX97T
jpfQ3pclHXz++uSGTD+1n19xxY1yBNWjVnaHaFMtB4VGqTUxU9uk5mDgev1qTe06cXAeu9bnaoCe
VNqfiEPnpNO5LjHTsGF0H/T9DYcUda3CFCmrZfC1WFVVqqXWrjm4BmgQK1n39MU2oalX78ESs5xD
Iu87Cn1KaM3adJTrX9DR17fwlJaotd+X6g4hXZONPOxKZb8oR4c7Qc/f9R65INLq7SIIBb5lrz2n
IuTCGO+oS8TA7zjRegxGWpN/AIoRZGg8q/ymY+eYYyM6+BAIl3yiYXAo2AinLWjy9cc557ex/Wco
9kEizJCZi02JxVTIRoAtgvavP8q+aXU3cNMbcnJ8Akr2M3LVDN9aPcYOxOijG0IOonOZ8jI07kW5
k76yTBB2CjonsDb1kl/LMvdyIyIL4q04yCFYfyVMkNEIqyeEALIk8VKVC/iblIbcQc26/WqzzsJY
01Z/c40dpkGJwIdAX4K5gYzotnPkC2/ZOrzCreZzMvssNkZ7k+beEVljYi932GfxVrKb4/LoE3qz
aozBZtAhXvF6qL0nEI6uovkd7+K5Log8qpEicmqnDwllUZDCe3f1VZRXLSjt2it3fsS37NNq+bmW
sIDoyLytCuZXK57UXV8x0gjh/a3H/EgA4019/5SqmLHEKw5Wk9e+ojPmHSe2pQVQiV82tqIcizh0
k+E9ew3PSr/II6ClMiGUvc9HIH6R920mM7mCL7J93azNEBkTPAqxBk+VDIBgcLgwnF6kGN0iJM/0
NFin1lN2ec2/hKsKTmTuxELWin8cEKWpUjuZrVH0bBooCFhF+5588wy3JLAGh1n5kTm+h7Gn1jIa
4t7XhC8rhX96Ga6XpD+vh/zCZwrsEGbqD87t8n1unTlde1ShIh+ELcMB9tBGoO78IukDbSlVFgJM
/OWPfSal7RPR90ytfB94JbRMcWHWVcLJZUVYsw1eZjYNXnVw8O471G4ODlHwZun3HItzwpUy5Air
leZQ/xqJUyqYVl5UkL314AIQPrvTZit0zs3i6/DC8APcThA/P+lfiobF7zQYjem5vn14fhf9O0I+
o1xR4C/vGUzq335eGqUnLt1VwfmmAosF5qwqv1vGNGKLsTjec7s9P2VuhYVm3OEri4r+brfS/I32
BUyXeOU1IOKcyGF0SxBvUiHMmGJOOYLW7EDbj4JNc8SOlQdpp8bFKqPzr538ZfRPN0POBDrVfshy
JXg8iVzu6DYqavnaW7YLNMzyXy/v5l4uxc1zA7gLCed2m/2JdAe0vShpjzOftM27OVsJDCmKWIwf
nyarfm2alGVzUftrZ/fQdjHS1DXkow3QYeBbAOudhV6BfU6g6zz5lCREkv0hwJi7rn7WBdWYEvSI
BMh7EDbdBITXInTuHOxrzA+XTQLegwHxtJcuXsXKzFGj0MhYOnP3j055stXgm0Vsh7E+E7ZYCog1
qFafgbHkOvG75mu8khiA8V70Rtxh/xYSQLV61ejl5vM+Iqc2IW1Upmikh3DRkKDzwsmMBUhIBErR
znPr7RhR6KvalQNkQcN/GM6WPkSs+VIRZcY2SlwZR5q9jS7QF9d/+7YFns8nM9Te5SD5TiftjBEE
xoCcT4kgif5/hpV+ksYtx8z1vW36iajdwCgMzL/7Vca4M2WimA75FifCXsspXzt5VIgdI4FNQ2lD
QyjSQs1Po0FAfh0WkbkqficAH4jnvltbzf0gBxDkhM3tbYvx2TKWsvMgii3ZXwO/djYeLiA53gCA
H8mAp3+xx1L1szNKqsQy7nnHuTez1g3VQdACifJwR7apCY9WhlspzN5P+xFjjDHava7GxVsucjk1
z4zDGole25Bkl3h5lD13SI+ETOGVexG9yO06JAfiJy09uoXAKXHDNeEY6+W8r2e+DUVScZy9JF4m
+Dj4uyX37ACeUwgwgX2njZ6b53dZEFsI3CSj1EZpDS9MeUZxTKc/OjljPsgZrwThXPDHZLqUuDm6
yk6ZDpPEo8WIwIcjkH0KM5QsEyF7R+YHWEOrJmJoNZZFb+djY54MXBqrs30DkuJAMXc7z5VCPSGQ
M71/D9rHjAcPnIzvenN7q2LseFERcTKAzDP3Pg9zYTvJPcKArObzSYHNEvSZmF7TYnHWjiVZfqJM
c+5hu0fRRdfK9iDCiZLZHcfnYZPxNoM+BHRwU6MIV3a5/7I2B+Bou/h2P2RJAuWeTcIyuBV2HYVD
N2RR4f/wTVi5CLW2hqyRnoWfTxl2wCEC1bG5Zkv0Q+WI6IiY/kMlhCLB4saz9/J8OkAnuJq7dAhH
CPes/JmajeaboyX5Ylf5o4tTUonH3rjnznQtqTQi9TilfxsTqIdwZ6XEfZ1TUAO8tUMM923XBL33
wsnxWrWYwIlSzSwHWd/0gBYOZ36weQEXW0SzesODVW8rAM53ei9gtx2lzOgVTMBi4FBEp/kyGObA
eK6z/BbkeqGLwJJSBnC5IVCDMLcJEifkQ5Xg+SbDmXaOA86bnrZPVqQm3s24FzwWs3lKN41b4RiJ
tTYLEuYXMKYUF0Ho22agYvDgEB5bKWCRYDaf+tVuzgjEpf6vsILtlEdPvGHGvYNC7MTE1MUU9BLm
DeIJv2Ok3Wy09SKUdv1EnL7zoc6w5zD8tV377TCrDw5JEDMaQ5A3i4lmw8vViZPYhEC+difHydC9
weSL+6tN2Wk4W+hRVymMY514/eGv5Gb1NHqeWaejl/CqRiW3fqcL8qYMgqsF4RqBWvV4ON7UtMMC
+owSTbn2ZIX95ubhhPmYdraCR6Dhc9ZNe3ZYJjdtDD/CT4oA7/53sLf82lPr6giaUniVBvSj/N7S
ECc9se1aA5b/xhjImpk0AGo6W360XguFlboLcSsrYrRoIqFpmo4OdQ01wgCheUnegjtKRc6nJnUT
SPp5LwRlJwxdXqPma1xPbku0t+MuesnlLvpgvwD56dG99UqikzPFTVlyhCZM9k55SlNEPEi7qr2m
1C+uYvhRFs05S/Wl2t55DtsdASffKmE6YFzFNd4z9kHdrzr0gKUNHhmkq3IhEu91j4ZliZOGzVYH
TgJcvcnzNlh3zuuZTOSr/CmAMv06CFwraTAhA2C0TbwfvO5KOrPfJl8az1Wi8LbVEezuGRztVVmv
hRquDIm8PygPBPidoWb2HeT9FNVuo2Lita9RSczbGQ3aSS/8tVpQKtmRT3FIpWKx28lST+o/qLzn
ICv2/rUPlpAm17FP1OqXSdUGXT+auAyHQRAKTJsgVA0JLcFsx8WMlTTC2MnWW3VSslaNIj5WxIJQ
8wlQJGDXP7eBeESFJa8Sb4AHXQfoN9ivoh+16I6dnbVlV0uRRevkOZPzfuXMiopwa+kUFa3vaaql
8Nkj7UBiyeXFsog/iOay2Wb8zqM0AnmOmcXmIfOTkcR9/8ZWaslXIQiydQfaXuGL2XOfsGo1lbT3
slUSClgcRheTTmtCc6+XxOdK2fHFebRpfLsZmZ3wkn5xRCbB9PB9PBkVeYN8H8ncl4hIXUCFTkJ5
+mALgs0ucbBN/eKm9dE6B80KUj9zBzuSbeH6wSpCkD842PreBhQ9lxhPafmD+ButsbCC6SHnkcEy
d2Sd24ixrM4+C4VZqbduWP2KV0nGCmSr3ojvUTWRndTn9LHuEbN/oEZsx4PLnt5iEF2R2O0Y+aea
qQOUkNEVFNlVsSsvlgTLBAo6oG9jWKh5wggpcCB5Fe3PqLmxrZypWYMYNneEnRbhDoQuNNQD90tt
JOachNTV6Wi385Apb7oindYPVYUfGqAi0RUXlQ4kHBRUPC7uevGru7TqQ4iBlobXrbDlOEKnUvqx
Vp0OueToc/V8ojJB+8rIufHLiP7jN/krbjZqIDqwECpGdI03wZ/ADhAJWcrq2yds/GdR+iKVjP65
U9zhqF5A5KCHF9uDuN1bqTxXdegFfZXnvlDoS3onvOWCH9tbcGo8q28e3P8FCCOTV9RqukMeifdO
Aqp7/WtbQyBjRInz93SIrGBhb9S0qqVnYdmaJYI840yus77IIc0WL44cNZqfILGcF6FWSzSoGg1m
Q2RDqNgxmezaxTjVJ8kcZSpUYFmx3GlX5jhnyDAWNxToRLfZsQRSE/uYaqF19Z+yYIOG8f5+DCdM
/9blO4ZSKJ9oNZm1fohCgINC5ke7t2bsmVDRbOnAQ999hE/VBCsxCrhlWXKmSXgrJfM26M7Cnl1A
tHtNli13VdSraKhnAyP1zlRjDFSt6g4LhzTo7luDUUktMyUq+XE4ZFuO8pQzriU4bLLwI0SttfYF
HB0dKEq3E4FJlpIfUS6aAb0670iXx+bd2+PZ85ux3ghar7cPIusQReSzhoE4A7pI5q3RYrfzDclK
4bg8Jj82eZRW5OhSOU3QjVovUi6rgVFmlH7SnnnhZ8R9tNg6sN0htz6rkyi/JT8//p5poMetZRx2
KIpG/DJytQDG87U5iHCJF55hczVvj0O8F2NrpuHOzArvdKiFE8rL4sLzQIP3xOJiQ3nEY/nM+SXh
DhfsOXaGz7NiuObc4efFi3UJwYBMuqZ1BerqL7YbktSuXgRH3NSmlv36LJ5Ci43/u3zVlSKKgbxy
MgQUUaIfiYG723W2RuwDoVqKEG8rj/UcXWh4+8WuMWzO3BQvUBjS9ebGhAE08Zyv/zdf8hEm05+x
PpTenl//sMXLMveppX19WjbTtEoNSvXfgajwBQgYizZ4YTaJuJHEqZkIS9Rvdy4V9aY2uM/RvIR0
GJiqN6yn6Gji1LH+2cq5x1Tu9Ns+FDI4Bnp1PBEFMUcbzh2wyWjTGN/HCWKYMxhKmzpJi38W6y2e
B5mC2Lqw1+2mjkq9Kx87mq1SNOJmp6gmIzKyRMgN1edIRUGk5LwrCv6VZrer/57b2z1EgQDgUHq2
THhfb/mmsOd0AOEtRgwWQlzNnezk06fOQrQf2rlqMKkoO32+CQ3QoJcIUGvC7zp7NBeBOeLtoxIu
gr/T3P2bljfevBM4szKdcfeKNH+UYKYfIU6bJWea2sjw8qEjmC/wK5dcRhPq2KOcwYxf1Iznb9r1
KtBJYicC3YQmARUM0zA4U9JVMUNq1FIRwbBdbBxIlxCxKdrYcxDo1+fc9s8OVWUwhbsL4EZA2q2s
ffe0n/XUS2F/pZH5ygD438IPQPhgyEk7l/bmqicZRkzdjpr3QGrc7Y6AMwICapyvUlRRu/ub36i9
wm031uEUYOWq1JbuJqtU24/Rb3NT13ztUdxMPcTZcJad87hphVB/cBLdgmpSsXg3Oh/fyPY46KKX
FYi3sjeNIoa4xB3jxF5nUU99SnWqdJ20kLrJaMjXGtSJ+K51OZNrvxxiBdKUXvP371ekcmhl6Fk4
wWhUEnNa59CvwmjaST92I1iVsKJ8t1oq099sDezUXyisYG30q23PEsTlGa1apEbG0nBU5+JTXHNr
H4MOloe9dXLPREZjJ14SKZbBWUupFuznNTY/fkL0CqLGoSdN+Jl3JCqcFqV1QGr7W3ORxEg8K9FP
YwTwd1G2FtRxQItx9IC3vvXk8CG9vLj/v+8s5JswrpifZ9SEDJYA2Ix14MQ/Ky9qyY+qRl0RyUdw
1MBDBo5yohCgGtQzHmBOhAlnnce5JEMqiFRcmYMKCL2nXvz3ny8T3heccx5nHocx/Bak6Yo2g5Bb
QoYWFaz6FU1zLdOOjo73oATPUR7twW68OJdcxpnSa8HkKSUeM6F+oBtN8KRzQEZxnggZY+cLQwUW
CyVqasZAKehFM/y4YYuxMki2Wzlw+nv48efit++GY+1l3yyiZv6CDVs3Onv2O+7irheX2QPvfqR7
y/jzlDUEa2lE1Dqi0WrM++0DCVPg3fSHpZyuw5eBs5Z4BkWjTVqGa4ZKUh/HphslxRQ8S4HgiEg2
mwaLRbe7t13KZF2pVNYbRdT6QAxw90UY7/rejCpXL4vlg8rT7T1tAiKAcf2JuU5mxb8AwHWcrbKT
n3zsCF8O+/arPQ8ta36NNJ08ElSlfJ0vj0rd7O7F3GkE5PUXRPCot+xT2awET4gzzYG8SrvV8+2L
LtiaJhprkhaJfXplw/PLAq3H90nRgZTFXzWUJinGHALA1pCgZb3U81fzhxxOyblNK5TABswHpu68
Fi53/m4C2zG/9C0xRVnwa3FWCKiL6K+gRxkbhLH6i9PWO2eCmD36eKgz0npgQRr+w46OmFlPKNM1
t5RYYvag2QGjh+5+MMUUxfg9cLrWCyEHax8fcQ+J9FgfkmJTOyIz6dTHySjlyV4ZGbouZUSQqIeM
ae05Y3tJpPbTO8DQs3Re5CwYt4iE3+UnfVxWxZWJg+l2PMQYAm81gH8Cfz/ncoZij+9EUXsvP3sf
kx4pBQWBbYvmfIBGv7HwC+8d32HVScANabd7HV28bPg94+brKolr80jJmSGdUg4LoS+Yt3WrFpev
bqZOJZhza9ZOIWr8nTdgp9rPmXbjzpk13fxGXkn+3Y802vQzIUepwamlEDh7TsjzN3rleIHRTKOG
aenUTXhx0Cg3swc6F3W+ZvTFGIPsa4JrQgPFv8USzz+BrJ5RyuRhGpeThCPTalrbvRF0WU0aF0wj
+aN4qiAf1QVDJkEUh+Vss+Lzcs1aJu9JvQzBmAD88voEYlExzZBKlNibPo4jpeUhw0J6MZGg+kv7
TiGcE4avDhzlD5sa8d5/v98/h5DQcnfj/I5bhWlqyznIgCl435ywvntbqLxI1DvR53r3u8SEDfJa
SJYhjezz8g0we/3ue+kYQIvexH67r4S4Sq026fKiOwWBdC2ZiMtfR632nyQJh9f+OJcLzza705Es
c+kfpKIGesrGInCOJs3opygaWp9GJs8XlsRB3K+d4IZtvEgsuDgyuThTEvkIhQqLQNkDl3unTd2k
X8v6lCYQh1n62wMJk6i3aUQv+KHk/7BzrE/nU26NmFutL4J6U7ayQhDCxXBYYb8dQoE7BmI0iQJI
EBbgqqpAmcPSPBiQ6ubAIcijep6SJ4KMEUs4Eap5DxH8+vk+7i2yEYtF5xFENBdXHiGRdxBhIuJv
DCzXI+pRKcmWL3wBdcSgVzw3EnmB6vdUAgYXBb+Gx2kVpVrAT1akNF9epYNgKZ41UJL5D7Boqg27
ZZeMQlCsOL5gDYIDsFXDPpIzjhqdpT4Ud/qFjdUMNx8MdM0xR4UomhhhIzw8jueIX6rkbbjrqPb2
Wo036PQ6waRSe71jsBauF7+PAvP7BMiluBg3Nb3Z20WXHojnPggqoi5bSJ3Nq1FkjB5m/MCGeL+b
L/aMyDmJCXg4CjCSCd9FtuYyKCjXLGSCnRsXTwAknrAnl7qubXgmMHm9O2yWfEt75PEnaug1YCib
igk3/nh1b4vfqomo4yIpsHQyTr29sdtgTUcFrmjNQY9FF0WG/U8cEcGGX2soU9mtDM4I3ae3Apwl
hN4FuaVQEzlgjQ4c9FGrYwwIaUa9h7uOtRRoTa+MDG+F9GCw4mAur++z9yTpmviJtcBBENL5B3M0
A5UaQksJsxNA5ZCyfqa6h6rBZvFc7GLn1cbcWXsRhuZZVf6uuulYfaB3lZq4exHBRoVTxzIyJ/s6
e5rKctfDK1LPZL62jyPSJfR44LYtXwCf9YiD0GPtBP2WGtV/8xHNFANjmvnzYj75pfSjo900xodr
fcB7EqQQ1q7Fca9uFADqaSHJaulDD0rGGN7e7U8UIutqRv2+2Y5xe84EoYnVGElXpiQjmBO4ZIcO
KC4PygDt7cPn8d6H/nak9PWG9BhFkZt911PUdR1QdNsjoxjX3D+ztBOyh8UY5QxMTme0v7EmRExw
cEec/rTucQQVdRQ5EHtnep9NG3oLbxN/MXfz70F+SriDshw7KOvoRk6BVZVG+TemopOjKVUolT6r
13/oIet8AurGm3GeVXrPL8Evkw5pp3zZnticLU1bu6MBszu7ClTYvy5T6rvJjl2ydmCzZbiO7Gyv
wWgKjl+9WXwdQHefreWsL7e+uHOqN58aDbaHmmdul+aGOhpFyhuzw+jhsnKIVvof8PaxQIT0XM7M
sSbdnI7r7JKFsf0pCEKZzLQzQcvaTDvfkK9Kre42GFrcod0Xan+oBYwMIQHluX8ED92IXDCWQN6k
LMM43irc2mQkaPy89UiLzFLxGCPbMWWwyHojWMzGf9qq5/pdnAS1/gcmVDRI+MAuP1xOSQW4Zvf3
BXuvj0Fwa8ZMVzAbSYCwre5wkYRJiNJGVojK1WjwwQPYiMilD1XSBJNQM6v3O4ozcAD4caCEGjtl
VNXwIRxvWIbRJihr0ySCpnO4RWeEFhjiF/hQoc/Hk/u5UJwpfUjgc3IPM0pfA5KtVjk+jVEQbcgm
uMq92rsXFpgBFkPj/Tre51YHDX2QvWPMsQXfJT7SooUQJ7/3rYxDKGrYdhKyt4VB9TkTKqqjPjSu
/ymXKAetWPeks3e3cRFZJLDHCaXGX2ve23rYmBRxLHkSaU4vXbOTRMSWM/lh5Njp90WHOFFV3ZDZ
Rc4Izo3qok1GQ44C5YVfrHYuZENtD7B6G+eO4HdabiuCdhv8YJtAnZxWHp+2dXMEkiHXncNQxMLi
1YqvAzrEv1FQINAU5VnnI1qKYOghcRSS5Lrxon/LgIAoyBiES6RvcT0RK/vuRJXA5F2Z8ZdCU/NF
0g0tqB7Z8UISot/1dzb1KPwZ96RT8gOKJ9sbCvZMo9XDyKFE2rtS2sn4z6UpiuC8qJe005MEdEk6
Zbrdxrcfvu9MyIsF5Ect22TyieabpK19AkN2yG7R7oDFeqBQiP6iWxnVtHLNLFv3NvLujgtjl1ll
NzBokc2yCcvScxmyHPP4oHF+c6TKvlU635xggsyr4gXz+vIRBok2H4Xx66FJZRLa4R5IvpsYgDxw
rdAgw1idVHXOYL6RAmZFuJYp6O6sx9k8wnyBgd3yx8i2Vq2Zc9SWCvxIZ4xMWkMBniZhr2V7LXaI
avJEgrnod4P3t+EUcLajj1ZtOneicFEZWYgcYy5IgGnABy03Djnx9mFtH50u5xTCMuAYI/tmOH1O
Pwb1v7pwKheTpmeTfb2Mc+GsOqAKchbZPMfrL7PqUuIpusnwCJdWi6ScOOV73JYqXA/PhqEWDPOb
1mFk+nboEOPHg+bYJe9Nx6H9CdSjtQt2RufzDVl6+Eij8adSHjr/DjBYzJmfHvzobpunZQ7lljPV
MpmMwS+zCfEnCqiXciRxSSo6AJpXj7EM0qNQe51DzkZsMUlFTiz3HWPG6+aSWPFnDWrlnx5+mzv4
p1tJwLFazDLTmnTeHnG5uz7neLqyP9/VW27qg6uTTLvbd8O1Jraybq3vDHLQYVf1ydXYJ/ATwSaQ
QF7M/XwiFPPzi5jSuFSKrVH3IWxfJoXwdCtQQKgSt9ULLE9nWe+JHysvMgEPcrGMpekxwJ8vbSaX
2ZuezFRPbnh0ReoDW7vYHcnKWbD+lrn3hDXdZeDEanf5Z1yXcXP93S77ZdBUlRI7JaHFHTLGJCHt
MtXD0JUtD4hEN7k307aw/EL45Y2+g4hPFpjZjr8ld7K3JdG9RkoXW0dZGQ0W1SkGAX7VoX9/aKKM
P3s8I1SlZ40Qs/TXvtBESdLi4NZQxcmVIh4ptcX+CZRQeO0Ch71QgueTCCqvebym6r4IyWQwd9VZ
pAGrLsZN3AACL281Oggfkud6aQQ31XWOw6OQ7ukCo8Hk5a91NZhV6dyoXuHkIYwKFUVe5nxaJonS
BMgF+zvAAWB6QDvEIHTIOQuLBONMuKfLPM01m1EftgP4LQDhtB3HFimfLWQhZo2cPq9rzIuxJORA
UNFEnHkHW5yW9OvFvJk82lO/L4HYsYlOZAZzM9NwAauT73hHg8n8JaxrcmU1bm9+1UM85lUmdwhS
4uRRdbEybKWZnh9MUZKgYYsKbE9SZjgIAoPvV+RjGnRHVor4kypcWLUH1J+OvkaktcQb5o1Mr+7c
IX4x9XoQbB9hCLkfBceuiLIxS0Q9EXtXLxn6uQLOw+b4Jp1w3Q6+Q5K/csaRuApIDsAt8SsuOx1y
NUl5ejOsiaMT2yKPIvKqQd2XbtPSTPUV8XN4AaEgLwd2h9i7ZniKVSRtZPzg9xYOM/6H0wVV/Yzn
yMutk6DUAwizw4904/3hDJKvbk/Fg9KGGKrrAxgk5ozDFng+yB7zr6PU0bAGefXeHvArhWCY/Mcy
irTN2LD6E3WU/jb91rwyLvTXNc5Qt31sCIq1BOD5cxAK+4VX9p4021GBQs+f4Dv1U7zaWLOBRb2C
VARslJvH2QAD3lmHXxONxIejEZQFtr1DMu0e2faWMF0VUQdA/AnKtBahGknPhLEm+41VfwcwFUv7
AM8earmjIgzaUnOLJxEeccnJ7EEmcyvhpZMeOmZJ+ykzXztR0TBeami/+/NA/8tBTQw6e+hy/VPS
Z3nWGQz+bgV7eWt26ZlSHxqySnRp3jjrEPdayJ21WuV0WELO/heBcq4h7ComdiYrH8DVQz868j90
sBRfu70xKqrH13q5yMu4H4b5Nf2c0PpLy0lDn6fETtrZ+rITPS/9IaBf6crG0Ta7PTwiBJPyYkR3
Jmd/SQXj7P6cEqmd3xIei2aXi0LoFuP3cMbk96+SrgRQBI4QLlltRzpyZHxQBY3iuXGcap5M4/6U
cHeVH8oFOmA5hRzn64d+IlsbjBDkcm99wI2tUqvb1eBJXGungyDl+v4K2NrG1nbduEfcvgJhzclT
NixmrvpklCsxpsQoJ2IO7xioS4AyXkrYPmAq83C3UNq7xctM8wzomaHVyUR33PmHahyApLOcnQQy
o3Y49C5556ke0fPyKm+f6D+zfS53G8kpQf46cePT8EjHR5kNFHV8zNuY1sdsu2u/NSyi6WAOgEjO
dt5n123szB9UDU097+vaoPyfDAwgUH0+eusZJsA1zlG+kKvCNW4DfHni38gc+K2KcT+ozP+EnK07
RYzKofFapwd0hwJUIt/9yk9UHsM72juxyaZA4YBCFBFkInIKOnd4YeKq3Q1f+aWBCqa9QTN46pAP
qyIIZs5gKqrErBzYBouHAGohHpK6OkUUGIJzAR3mJyfNky5LDvanTQJHtwaV1IYv5zp0CpY51+uu
NRkIbgoHpmbfAevqPhdw8noH/zg0snDpougrKk5NHn2v2PgWsAuAhSsXOG3w3RmaZFj6kXMywhhk
SK4UGLYc0xh+vQCtl/IDTQ20fjFU3limKdpfj2fde+HVL6AYwNsHMYNSXUSJGfX7EcGb7qpqmvu+
k+fY4BsAc+4rDgw1YVATQY3Exzm4p5uT8dfRPCxz0fd62Ad4H4JLX0MwQmG+GAJVYZ1pPsXZN3mH
wddArVtERnrLbm/Tl/+wJA6T58+Nf4WcP4tE0gM3h6QIcvavclE3ldHGaYbR7Pva5X9e9uars8BH
C+4ZJGtNqKP4POgrDYgRZ1lNmqp++D5ECtug/pc8Ugax5r1JL0jzBRSuhYkWGG6wtZU0lON1V8p2
g5vaJ9ogpJDkZRwK7sxii/z2xBUbg+rhKl3DyB5E0qs/ujQlIU8nQ4d4cr/l1r/X7lQAX/R7l+t4
btIUFRw69/u3kAPPFUYTiiK2v56MNERojJcU0Py9WkJ6z72CKlXo/upt0wYdXc4r8SGujsnN0GkW
KxzXMVa3SWripQP2ps8JZwyVlRyIuDQ8/PYELt+bKcKzkAdyj0dv8Xw/Tep/pq/yg5udVgBdS9ac
4jGnfBPT6xVnj64NCYadbdlNX2gNXD57lubnjWBLmZxeKuj0ATkwADV82PcWJxV2rYb6YK2KMQyp
xvvxcG+d5iWZMiDFY3FVmgikXkwBhRF0RTs7DRIZdWrSv/VYl7st6QyW1FDYZ5PcWBRzES5lQtNr
ESjwEWwOawOLEciLcyUF2GxZB7SbaNcRJ4auwHD8RbUbOmJVYc0r6Hna6E8P9mNhFzQsd39Z0bfN
i+OSv8OtcHHDkqXEzxU8iYz3zDwASyv4mJuiiVAgFVnLJC+RCQGPlguXA7as3Km2kyn4pJXrogWA
80CdXD27LkgffGC2Rjz3Rh1fjA9kKpaNuB45IiUPJeKv8T4R0hCLgxyfP57Mv4QxXKl/bbyzYWv6
5Yq8+E+ogd+0l52/0cPO1IM9N+2ggsKHvWdnWrRh8dqd2mAQJkFFY5BSjxpJfQJHHfYaJIuvewcw
burI98EyBHFCRxCNwga3Yov6YjIKUCChmb/g+WQXsQx+K2wKLkFU8IPXL+e+mERqzeHokEFEqWQ+
9H21xB04zACYahF+eFSZNoAJJEtwcg5hvIxVytORju0fjmwIi7VkHO4RTQA7HmlTUZGg0iGlzVIM
QYJQBTy7dJBE1r9gYB8cRyVm0vbPqAjIJ9SyTmACAlUJ0/O3B94Dk1k27+Es9scn51WQu3xW8gwQ
XYnaAhJZ7acyC7aYbD2tfXXIQpwPiJaG+GBN8ekpyIyWGPuQf2V0sTFRAjFaN/MPxjWs9rc8XsIT
lvh0opUKsoRyw+69+MdQouSVcTfxJvAME7OKoZZVpW42zifEURhWEeYp1LFVdPBYTZ8hv33Ph/jG
NaDMbkc1W+f8nX/HQHD8nlKy7YA5Hr6q5OCLbJs4SkI8PX9mHj9bAcy2pCxcRURcwHZ5wV6ms9h5
hbC9XpT+tv+YLr9x2evJWZkaRpuDZUp6FeUelXvB/GhKxNHsozIgV3uEST7vc0Ith7qRwXkNEfUF
n7TJGyIjGEIztC5KlAe6oEskLaqyQ7Oy5knDvFlsVevy+sqE/s9F5iNMA3LVJRfOSD7c6znOZ6TI
4e6Zpqte9EoxP1lmPCEQjGT7BgjKmM/junflyqgWATGYnUdyvwxBZFf7m9mUW+9qqlj9uDwwX/0Z
nzzfhJvuWfLo9GCdO7Q6mtk5w2Hio1SF9wuJ6A3cNm98G+ravP9yFyqTRKj9kWWkCKMgKbrRjZHf
e2fG+27cRmenDMLgz7V9h/UZuhO4T5BMfwzU5D+kvfV9NRsEsE3N/zVgYtsQ0hZ/cNB4Z/kMvSDo
0Bnv2IZ/8yCJpCnjHjoYhYZ8Px6Ejuqm1rDkwB/1lv4Xg197T71Sa07fTgn4gZ3zzk6T47f67FxG
N/bfXiCKCLDpz68O720Rl4IpNsifagB7qWT0+FGgaoH76D5w4J7DNEa2JhKj4gGt5mxrYpPsRigC
DLL1I0ybHAPW4J2HybalYzoI+GW+vPsN1rauM0D3uMtZ+cMjpfDXfVVKBf4CTy5mVkc1iOyD3Dib
s3FuvW10+WiKDZuZ4+Y4237c6sdToiJMCP2gdPNbZ4ej+Mp28pRZ8K9M53bxG6DUkOjcCniLAzQ0
Mf9IS8a3Mv2euSA28mvG7sGjssr4j0rNF+wsV9IAV4DHJf+6gOg1DTAgz7qqGGufX+PmTa41G1PR
3CUcDJiLVaxyGxo6PDJtuFWEA4MaZUILor7AMs52xZuWWKuWEnsgch25ulTzNCex+ew5YDKSmyx4
QcvJrl/JLbayanDm3wrfceejwKy1qmHq61UgW2P7z8mBRo+K/mW9w8cdw6cl7s7ad2cZtRfWaAPU
HXH8goGYZiiZz2Wjn/WYdGS2U9Ol1aH6E7tQDy0DKbsmdCqjTp0Blhsk+A+rGl2qRPqneNHUwm0a
awaP9XM/PvMkN+VhW60CfA22R7nkBIdIHgOp1nUpL21+9P6P2FMe0irIepR+TGW+Fv5YnHjIdFXk
xnGjH8jdeUYiX1WusaTxsd2IPwPpCB7eGyu2+IOwXdxSp3TuiTEz3BxsbyEpF3ozQbZLI/cCOksN
VT3Gb3L7V5U/sCS+mp/MTNff+NcStwQ8T5fJ7lZNaPpAr2ZBjyrtfWczBQpKxatibnNdTNqP1vPm
JK137WdUhbC3yVheODck5rfKHQZ+H4OoZ0WylQShLcJeLj+86r72LbZsA/U1IyzWmFmZTF32dFY5
BdBanT6l2ZFh24KakvDAfPHxLuGQdWVmmRU6soAqAGfwUXBTWSiN9TLzN9D2pXwfGJ0JCAoIlb+4
sx6+dGxPhondSxFqvCe1jg0X5R2xMXZMVTrkxzo+JYnj6nz97e6oMvh/OYhNeaQYAq9RfdmVm4zi
LDRe/f0T54lrhZlNui77vvc+0pMAhAgIp2ufE0ZSEnoKuspor5FOVoR73vwEqW+tzDlDlWMXZXSw
cUlnfZJ3Iar16SamlxBWwdV/3c23766sAgj1nhd5kkW9pBM2HcGvgCJGn0AlhU5QXwiXz24D/B8t
EJfvLqWN/3axr+CtLm2T95FT7Y0uc0reMuAAblBUpolW2IaJ+uWnyBrKo5eSOHwLtModN8IXJk4O
U7LI1Z4Z40XdQdFIRzk8U+S942M9KNkwMSBJikHE3vU+6WmZ2Q4Ze2/o1ecGwj5z3+qFXkDfHYX3
5kzMafVu9szd/IN+K7njpERjBWPc7W+MI4TAKkVj8lSo0JPHOky1HnCDBt26ZarPBOpN0bn7m3eY
SkATyHv8666kDqJFMcx3Lyv95aIvHb/pPzeLMK/0rPMiqVmGtQ/ij0sdKnxBJcgGVjasuVyuqeW0
jitGNztkxPOSYlY6scSS9F53qU5LNxj4EysUEM1K5k6jIsK5heI6tERpwSBIbfaQZRh898IAUdJb
sECSnsCgiiBmOLK4HuX5pLdJ3Dlqe+BC7QxtyJpJyNsLrJEyT0os8OiJ1Hf/GHsLAn5vnVGfaOOp
O6l9P2BCc6zfmLv6YDhgMl7H3pm3yVawiQ5LoFKRAS2jLtFD0h5jrdTIc1g7VtvK6umn+4xP885p
CH5T2c9/vJje2iR4RoL8HFW+LsyRgLmtKFK3gEA58mwp/qMCmkVZKk3RoWv9W8FrUKyr3u3jdqOk
gdFNcfOdAEer/zC2/P0X8LHlegMfYH2fbZ3u1QxbCAQ/Sdm9eOxg77C08VFTBXZYqk5FCRFA3R1E
rfF3cI05oJAzZF5rf8hUa/fC1Ei6T0czlRr1N3dxL8ijkjJVGgzw5cKC5Tbk/9V8YazaU/PKQr9y
5vo7U/s9+G4RF2dck9pyYzj1CO/eLc4+6Ct/ON8OcVbyqqEjZInfbVIgH1h1MPmb+nhYy28SOP7j
VlPU+AZw9tZ8XTXj7HZKBZfv/FtMlPc9A8BzOxd39qi7sam8kmYvpSqdgX8w+puES3PFf+CXX6Md
wuQcylKnzwf/iEZT4IeTGyjUuYTLoFNGUsaRZJZvlWvKsfral1o4banzeFqoVkyPMqrO6fBzA8q9
+8Cvb0YceTMJcwT7nWiEaaXvORztsX/9U/uyTzr8e/XVXi+ItDAHxpOqFsoQ1ld5frYMgwnlrUco
I8jOllh3iqHfFuJRS6Z5xuIp8hlB3auObs/vrjIqYVwbSkQZ64uM7RAmf1iUoM9RNSgDQTp0soyF
CnMQOot5bh+HjvL+l3mavMQsv6PrH/NnIsXCn3td/b8j/PUlpoY8XqAWhStPJT101LNLzoxgUu4t
XzHPJani+a8lsTpBqi2ftT/KXNxrDOQj8RmjdQDrINw0D8KfWPR1X9GWP3qmjB6R1+6TpQBaR6PC
voAzZpkahwlJfKrMkNTIBsiAemd3A1+eXWP8MIzxHPdm15KA+fdgl7YNiLXsheuz6OEGRJpR0Q3S
F6AitcewxDSIpJWlJOnIOQwR4u53Fb/rGKod1wCsg/KvGnyULtdodj7AGxPOBUAOPo30XezEkq21
2DB9uj4ZHyVGKSWNzhyOTA2UGLWnu5M7bu8ZJgd3GAqNRhYDoKpFQ/MqqsxXx4dMD6dGkfK6xQ3K
GutMSlDKoDtBtBnd2KxaG05OFWgSKiVsOFgnxPjt5xbDjhPP095Im6InFWagGgVNyWMgmw3a2+Ai
EjvVqoAqA5SToBPhqQrtV4oZcjJAB382yZHdpAotxz//9H2cfs3PwJrJDDxF80U0gUlpA4pVEdOc
0MoW8FddMkJltrJOabIjbGTBW1Fk+lJwYMx1UW8c7wcmvgjBCnTzA6D9RE+nuhFjgam3dtZ3pFHc
rD043VdMutu3EPM185oQakPVSHjIJJEjOBrTErYweYCiy+T1G1Sj6h9qdGHiBYFE9zEcZg7v39fa
xoUZVPOV31fARq2MCAilFocqFCC+OBcg6NAZ5RidADvYrnIWCwkefit5w08NccgZ0racoWCbI24D
Za50wkWCe4HtIgyYwlcTYOa9C0V1IODHUDMfr7k+PT8Iq9zaiFmwiwPMpa14jBkkffYOZRxCN9Gp
IElTLIamv0W4OHekMq+jgwTiC2TYBR8hvPOef2a3EO9b/WotKz+1D0iJC3Ilkq5s2BeWAskpt967
lVRzyUY94LbAUVQ2ekWyxErVrgggdZghRO33w8apLgCJSrF++v15dyHPyj9nLPqjiGd3VtFMdr0P
EJ/XhJ8EI8H08Pwygcc7vbUgHV9v6p/b3Kyh3nmNUdyYYOgpeGCDJu++w59amKAhbbVM9+aADQUU
c1ddus1HooMpcEMTKK3qTIo3wVEHp132Jt4IQtAPC6tVC3IdRdy5jF04e1YglUGd8gpAJtiyjggM
ajWEZyh4CAvhXK3Uvr5b2n2iKy8uYyIBDGc6WlEhW9nDqI1wTmTihXqlNna44ictHbgOWQxxfEWn
9kotU/G3u3AUi6gRKIbNxQn6X+l5E74H8dWSx7WDDMILWJwSFgigrRl+CmxjWsccLIDb28rHNEES
Feob9tAOTYonNXHJFPmvQsEhv1bj/+YY3dMNm4EiGjr4eN6hgqejxPZsN2sNC21zIhKSPsmh8bEE
vVWA9DaT94IFfzqgREmlWAVPRz8KDSl5nZEHhZLhDt5mb50qOfmt+TNWdZAup2WxgDwQpkNORUkw
6/SNPSZxF5Mjh8CEiBfQDM7OQ0b5yJ1X4h2w5KK2vg6jmgNtqd6trb/7831R3msyP1hCpZLf54FV
iKVig0UvHaXSr59s+EIRzJibhg8zgUtkJvNp2idEEztW0urMYA4RASHPQ1x3rK/yz6MpZe7jHec3
lvKYW0n0nS/oZTOFmq5lMhXysz164SzW1GOfBzuvcLdCr36Z7zGZ8SMlkYSykCo8vGS0xWd7xkpH
UKN002Lkp0Bj5cg+QaDrMqxTmli3zUKbnkKe0Vsnlt701gTc+yzFeLwCvZt4v2Vy4V+BCGNjhGLu
rb7K2oRTn2dqwTJjh0kNO6xQAIm18LkklHAq1i8TdcXMsFXUcXB5o8BiGqbh+KIxsjq3NFnx7Us3
shn5Kk8YGaeFwTEXyN8iAQsTW7wr3tKE5NfXxC6UWExplKkJWd48AYXAqFrW40UbM0Bq8Wp3r9el
kFFR1RmqFmOX7xylbAgJmsRZx23LrZLslqZUiNXduzLzmPeH+WsgHpqIITlzJ9HSNjh1oQ1I6ykL
hcdp5kibX9owqvIWom8n0jyqyQz7jw0qS8TCZ0mOwCg6wumrxa46JleIiT4UysqWInAPJERH1XfV
3SFMvGs7rII1DPREFg9ri4eRlDCI+OX4KiJgCVDmBi45vZJOHTscvSwQqbG/pYhbdhRuvV1QftiN
v8jv3yHRdtxs8bPP6djothuTxZkUxE/gcmwJerXWsdoJQFpptjWhqDzZSONmEIm/NjrO6WDJlsBe
AaB4cHZRlTpRotFzDS4AOevenU4H/ZaMTp8XXu4kShtyNtZjDBrmzqJ+C4mWsI2t9k+tJCUIMMSA
ypkDuAtmL4EOyjPzKLIH2rN0jahIvzJuxfW4b+hjxcFRWXz9lEYeiSUDACDvt68lup+chZxF8OK5
fnsNLjAJ+6mnSFCjx3KoXSU2D8bN/uayKCH4RgDHUEREZdwDP/4kn7XVhyT5QHrhs4FmuHq2DMj6
AmUsg2QBIHK8q1nVOrRpEut/RJU28+Yd2ndNP0+X0uAKOBEEmKwjPymMqTqxBGoAdFzOS9Dv8Vp4
ic15maW9BTobQRujMcoCcSXOe3clDwTz0WFhIIVYdgsb2ZM+LNQrinpCR7wMpBfuRTysoG3YEclD
/aGDTGwWJT87umJQ6eJewAVSj6JxqI5eTERZ+0Jtbn3L3V2kC507ihqEp2ybrj+SSjsJ/G6TVASw
1e4iuotWXGKQriNCGC7DlWozyEJjpfjyBAF8y2Jq46pUOsi9fefwAPr/W8TweprqQK02uRGwqOw6
JTMh6ul+8ymkUzs5mHOd2kifs3E8TuHgk5NnY1XV9VZElrX3mc5U0DqYHm4PuyqHrhDY1vbtPynr
SLjT/8Q3U4sqFeSDn0lwa+PpsDQ6WGBdpkRFsPtiSLcQfkruDVUOgwRJ+dm4twc14I/9BEPOG7IL
tbEYYw9EsaFdrqQ/WElfrZX1oRJ41AKvsuibC8MMdIuPsl0MEgTxrOdJJ1DipPwuirFrAQQR3asK
a9L4G1qfJu29xCB1CfMnhNYg2+b/N7bYc0YsIbccS7s2YK7G8l899p3vEKuA4GeaGovLlXXJTXXq
luI+vBCdpL3MgsmuqwQH029AJrR2TQ+JMRHjtHcfTdqzek2GrnzqlS6+OJyfpZ+Wj9WSSj+EzpTT
qUp+5uVqZg5eP065+gyiOLZvdThh342WltYkM7RqRhAzuAek20479IlIhR0RVfHbPwl50hl3cS4T
bTbsevYMa0drw9ABX4LoIxzYsYshr9k2Gm8GQYA5bJHGoRBzTq8lXOtjOXp5RsRtLWW4QtoJnJl3
KR3NSn0alYB3rLSh23mpDcXdL5Pahk05TiAq5fSzZ2aVNd0BKny/YzEJGv7dHap4rrqj3WaqURIx
oKB7DQJ5nY3SK/nZkx0/p2odpD+7MCloEqPtJSc2Ad3D26YWKTzFI8TbzDsqBVF7RufZTC3TaulH
dZs3Do0xvubuljL9E9XIpe/qdNrrBtTLvWi4h5PXaA4asQexHdZxxhjJcxb9ohAZpW7eY2CGEHYl
Zc9XdUaO39DidYf4ujRvpF1Z52IZ7zWSmL2hvGOln6fbySYhGbiWD61dY/q1d5JlYK+ciAZQMz98
OUDMLFSEs5c52TQoHAmKFPg22z0B0saBFSvoWgVIzQeZftnUXkC47pVMRNAjPKV26w3GpwdyFTrj
DIEWrBHE+3X9MHOFxb1lV6jdtG7G6AnB4+8yE+DasG0TKLLMhNgfJqjyCf1iD3xOuLIxHnaLEO25
+HloMGTHHa9Qdlc5TefhWdk6ywR/OeSFqdk8PB1wjjE/+35PSy6dluSQt5owGd7fKP017j5XZoGA
/kbieAdV3AKxP3EW/E/yD5ccJvHGvK221Y9c3gokO3OWE9OH2YDRy9HTHp+gXMbC5fF3LxUej6Nm
DDlkVkrkc+snxJl86N26/xCQK5UzSircPsjaCsxvm6HEoabLykoomDwMJXvm0cMVTYJhUCDaPMvy
5HmgZ+MB3xiT33OLQSuLGMQdDDScgYEpLczcgBsrUf6JlRGH1QIeuxxgzDzQsIwAPLCYPJemU5vf
KLZ/MuxrfpgIADQ1l3n/Av/Siydd9X7CVWrdcowA7/KLLQOVPY0K+jLfSek+nr/RxjuU4Gnp0DFW
0GxEXigX5JV/9WvYEurzC87e8XCnmSTq7bB5eCh9ysTT4daml8n8wXElwZXfF4bv3cRX5dWw+GTM
O2/IKhSKQMvDR8czIMKy6b9KNkuNKF883f1M76AUxK05Of50rUoVEup8gbE0Bcxv+GsFyEl0/0t2
iZblgsP0psvRWk3F/VrkiqqmiOqFlQYaylePDHJv/7OdX+tooU1AB7yM6Q2ickcTcOrAZNugRDii
v4DHbOT9pJ6bWCjG4kLlGIYtJ1BueUZxrXnrw+3QJBlS5580S3xgFQS+9TerP9UfvpCcQxOU2YJQ
/9D3Yj2XlLzjw2chRTcNcjD3fCio954/WqrwZEYuSE2jlXHvGHyWSndslFx7Kwt16/R/fe76duQ0
xZwOM+Rn5mlek+B1S9irvu1NTCWmytGUI82JGqJZAF7rueukqXntnhRfu9dmDHJ37/SzRU9vOIR8
qDNbNYlhIn+1RlIoLgzuW899dtng1dILJ82cpvL4n4IfS9dwkWXDcExoSVy8iFRwW+NYN6lvcHoE
BVXKWSgQWYEZ+7gbV6GuTltpQTeENbeqxCC5GRxaYc6GtiiPFkxSfbZABTJwFx0o2lcvu/oGlznp
n3r4wuxySf5cOK/pzsEz0y018EVAE6pmucGZQMJ3ND69LK5vJKGo7m1btYORJK6qX+frm7qrK+nf
c6/b8HJUQq8cjlHumblFDrB8SG6IjVp/gAFD8OFpKOr0Agqzycl4Q13j2vfSE2NlNUS2FC8k8F99
qun24gEgVuEOdwc0OXoDFwJq6PdROQUbZbZoEy1NjPAZDu/7omEQDFxYJnpXWZDD56mwUGH9fjZr
OtPj4IuyJSHOKTjeBhAVqxmIdRJx52lU2aVBF9CWT0CxBYiOJxkCYVgaIk1Ot4H4pSLUUCVtaf1C
0aDopNR8BD9/Ndr9ey1naZlJ2jsWe/xTOFnxGzLDx5ofuCj4LV3EnUoFWyu5Wg2R6e/iJAjCgGOP
g4tSJ7TUSiruf8j0yy3Q5ckesaGQPCXeRaZsbZGqOGLYCOD9tPOcpBPao3vbCGX5KM0tCV7kHbQi
wTv8u80iCfQp9UTbj/mejxf44BAHhLCjycTCxO3rgXvlo086mIsHmu/p2G+jWm/+jlzJ2swQSsxJ
45lWOkWc2VU20kwTOpE+KlNiYfoOzxGPmnSK8mR4tOYcUyWKi4TJL2NcYni/uQh3DWb3L+GNMCh4
uEHeCZBXhoqlSpEUiXhlFMpkwZKMZUo8t2BkVy/oZsXHnILV9Hbkpw5T1IAkkdBUyIhqJiJ+gej5
JXgjO+5tra5bKPVG7gZ7nEMb0HnhoGcKvH+MNbhM/seRL/SndMnakLKXgszXPSeo/8Q1yzdZ4pe2
ir+lwhAY6fGvHvXfVtQ7+cUksTYES6LfIpcnt3abjg00RI6TWTTJajtQjE+WtBXzWfY2uLOcce1v
kr55UbVmEHDMXDH4Rw/AECk1GEjnmkmH/ig6c5WVy4ROhU0hYR31xKhEKWBDzXMK3rMzmNxoLrZ4
oUV5D8UI5qLwfyLdGidZknXaz7SmJwpDqG4rvoklWJPkX9+guXEHj9REKKmykskhBPijmH7Jd9jN
U2/IgWnA6HlAd2QFTzmWAZCFR/niOxndNQP+7rNZmecDEeiN32wuh1W5nGIhj0LnfQpPSCz0s0HH
oCeLOCoaxG1juSyDu7Gpj8YHhagZI7fqBwjqc9/FmovPfmMdq6HUMKb7T60go9PIH3ASaSbO+ZjV
X0X4VIW1Edg2kw723BX52+oqz3P2xhO54kwMnFkdiKTQqk79AYPIEnbb7d2TVo4/d9Pi21UHFNSA
CqcZqjDGChnf21E0KE7awxoUDVjMMLnixX75HSmBz7JpDVreBiuu/+T9hWmJlim6PanO1wfc1KWr
InKPw9rVquR9Y5QaIEtbLkJe/f6b1Vsk16qgHSFz4lbXhXyA9YFzqS4EBHw2J7IZw0zuOhduyTkH
0KgN5TVChzA7lJmrsafYTyMq7HeBlR8OXMw8kXTT3C6h4lIBnZkFtoSj18ik62FnBpMLmcNBOosf
VaGD0AsWh4GQ47FF8YKHsQWBimtm7XHgfU2erKd7AsoCuJ+rdTufHopAWFTaj6KLoCKtHNttPnX0
KsGLo7Wq2EvWE61vQgW2xJNWqi2G3eHW4N8yhOgOPBOjvD4BPHYgiUACBXfsWd6B/LY/mk8rbQGz
up1MZ+d55RRbO7cPFeccYVwaIgrd9POhhcAwAycXGuWEeiLrbNACXTuNSSpkYjaVcwsmw0HBju6w
F1aRF6D/fkDGfZaAMm9XIlxSHNr2yXyy9TJTyStp7pLNUveJGKPQXjn6gDLsgjbqBrgp9qcyrmHJ
3k516vd6S3okhlQx25nMnT27ZUaGy+mDP6OSSU25UlkOe4YhWdeMHrBTEWQEW/M8vnelGdPBNAlf
0H4laTViDU1JxaNMXjgJW3CR6BNDfHRC5n/KzAiRmNYVQikG0rPoYIQ3kWiJK2U3tPZzm7c09gZG
hmEtOE9zpx7O5SgmNmGRNxyIkYPR2EiByagUa8awkm10JQH2zixTd/KuIDxPDsfjSw52U+iy0lEf
ak8NIaZ1zPmQCLoZT0j6MRprIl3OiNtRzv6Hyxo5XgA7PKtw3+nPBg99PGAP2HR+HetdZUTgco/n
xQZxxhmo1mOGvIuZKtPBAPbpRCniHwoVUVmeO2vFJAnbuM3RANQcP4yThBCKVHoKk9DRlKRz11L0
GQi2DUhWp8CBi1P3aa+us6K2SBmadpte2oDwT2W9ebpbrVPp0xIaON4we2iB/xOYslTwD/dS55WK
HP9SMrNvCQ6Umtkl+lsYVNegJLrNB1aNUMRXygYdWST6++EeLOYavI+cX+bKMgqCjJP2PP7EE/ga
OG7COWkvUByGDGgTMVYyWPvyRH3GJslUNiLsMKemhi9tAKjtsqBsKFlrW+aP5jsWC1UaYEQM2JIp
mdn2B6w/lHxNRJR4bjH01NKe6Ys9YbtNb8Jbj1PthAP7oVYfYtIwxHIBkYHgAsloekkO1NdO8j5e
m7A2R/xWQ61bQyMWFVYAVcCP7nvIWmueoP3rYt0aYlY+dtYE7juzkQIiCNxN2Wu1uqFjc4PvV+6o
kEGd1pm24U2ORPrMJXrSNODgJ4NKUz7nEB5p6pKE1fQFyqf4F3CgfGRvFTZJqdsxvLDV4+mUDNNo
PLoRJCyO19z+7DMd/8OR9asm1O+5+yy52OrnOky7Z8zDpTJf36WYA/XNmS13kOhKmAKVIOq79plJ
05tAXZ3SUxgdrVDPc4/rzhVDYNDEVm1urCvd83dweqQw3SgmAHaHnlyr+Xki1WvY7Kb6atpZkfEf
1DH8wLHmEl3Rpvzny8TH27XQkHvsLMyo6eFO53CFidWui71CMK110ZFFLVt/Ty9JP/vdK9SLNggq
iVORkNZYdb+asLjV8hIy9ZxBbCN6SvOdQx5FnXsel2wiD5EENKHCEDOe3fpxgY6yMZSrO/QOFraI
/eVLSn3viz4q8SX/mWplKoub7IPRw5R6g47t+7jnGknV2iZya81fuz66Ne7WXvL9XLFvZcVxHxrg
iMukMOqk64z5jXMhjg95nRnTHBVyU5awunniC8oyrqXJYiBN1vJ1/vtc0dSMCXlicKBqL1PqTMsU
Mjed+pkyVX+4cpWCO+KWNhIv2/m5ir2mN74427OTtjGJXPODagkcj6IntPq25HRNOX6fwPHfxiUW
ZRilSy0wFxZF++b8Avz4gj9beTJVIDUsoNMN0Pmy8OEini8aBMulMP1MWkJDth7LM/FrJWIGBbUD
xPv+cJ3WqTwnmfgFjf3Vu7vRCNlMfT+Qf6Q+DW+pt8fVGJ04VTunC8OhTA4OvZkMbhUj4zWj8y17
BCZl64UnNtOgfrSKKZGkt23LFqNDKDnlam7IOOhAj7fRSUOc1V0x6ph8SJwO4ipuYgfQk22Ymn1I
UWY6AVxR/9JZ7zlL96fgBEl73hSbqIuI7ObPYC8fLYjsGq1oA6HRN+JorkaR40N+/wUzXysiGBXM
O1vXd0jvPq0nSDaPnyXjWLBemCPw2rzmJD9qjw5+SVRSuiNevfetFOLQPo/pfLNNVT7eYRstKfKE
6UeF82UlGbbljo7BkDofAlXCSwaUIqzpoAHdO/Yeoy46M6x/hm0c6e4thA0r6kyq0F9YbVckB5lC
/u4d+kYTZkuIjF1pAbZPrdKJ9clMkwrTsRVgvTLwdCw0uoZ2/q0pYbyX1zGGLgCfM4IL7vIMApEG
qlUxtVp49nK34dbS4XHCfPSeRz7YdLKY78FHAS5BWoWWGppsvzP/ph5BSZ5bf4l3siu6RVtitf4N
p9jjOzvfNM23urFfJuR/72IiVU9ZYkYDYNQer47koX5K2hAWUvKbxi2OrOjNImgfF+dmeQCZgdUb
+4poZAzSKyPijwBfZjq+wwpXUwY2RXfwDudBQx6WqYFKxlXvfTLieXPDoSgoSNhU9emKfwCUUu36
m4CRlXMK7E6OvdI2HIh56Z3JJoXcLwWxlC9Yiu6RcctTVSwumAhpvuNt3h5Lsb8ZCbgDv7d513u/
gcmz5hKvNAsDgcL+0Pto5/DjEUHgqnUuUvkcloqYiiEWimYae/9NMHcicF/4fAK4O+UZQsvlzETj
T0JXDZ0ltQN7t3QLwVHHJ0zsTAuPecfV1VuNs63mKqXqCIYY9YBCAxmY1Sd26dA6usdLV7YIPt+B
nFtX1F5Qzoq/EzD1U25IXh7AcbJG2paQBh5VlnFWmv1yxmbPrM/aF59x+wflE3IfUk7msYETkzey
uj18iH+w2GTkF9gwKGtX5xQnfRSA5Xsgk+HLuNTy5ZNmOzd0OsZQ3AmluCQiB09a2VwZjlyNqFMF
uNKjZXEF/uR+QO9ARkGysSOQX4Jb+i/neEpKwprIzryfFoCAeU9FKIW3ub5F8lli1CUg/5gSrm/R
rRa/DcsyuMGs46+8HztcDKjSCOkEG9T134Nt80zDdt8zZlIFUsUDdo0V4PTvsgdlp4SUvlSiE03Q
BEeDAK04maTlIsmjbIOVrThrXz1CoIsyIz8gQ13y1nti4iLiNXLtFi/jZ24yG/6Ba+7pFo2MzkMH
J45U6on2jgQKfYHSu09XhrKkNwmvH6Kq2zDuXypVpi5VD/ggBJN8YX5NzZkAgQiMgEkdgNWgBl69
S9MnYi5FtU+FwIX9uzRKehHkFVqk4YUpjWsR5ninrKHIdNCOAhkTOgruvHgP/C3jpaWp9rNdbw1B
RNz/5yHKxycGeYHI2H8PLwILjDw7NFx5fx1RyBaCtcHAMZGotsldswkOR5miNSUj2DAr9anTchhU
v/LRtIDmyQJhJfSi8UuJSPUgWCr0QHZvwJbf6EPIcO2m++lmPNYRGsSBeqcSIaijGu7Nxu2Ji5Aa
5jkMLCJWXDBjDBMyKPc4TXR36u7o/4MpSO2uet70Wl068YA1doTZbic8xMxJLviqMwL2/XCef7MX
d3WHta+mwvmf19eL3jD1gU75NlxBGkUO5SzGh59kwUL8kkNT3rO5Mivqy3eHxUg17vYYn2JkR2GD
IgONkgczWopIOWswbnc22tgIMvaKHHK81/Gk16oAf5slOMknxs5yXMKT5aYP1z5aVgBmMHiscE0Y
Y0u2IK+2fatjTa2L4vWn7ERQzxnpZdEyRJoH7GMeJhyEJCM9ZnCp3Mts8jFwuoyxwfVn6Y7AvuAD
PY0OtM8s2JIPwkoalbFE5IFPnGSpaCeO7AKD+HbzQxyq24qGrtYzkpYvkRGWnYxQwWT4abSa0zTw
9lAzO/+TeMzJkVrHzg/emSkeItCTdQYqIK4XP0mos9eeID9D3QPEsiBzys0y20RwR89VxWZFw1ez
wSw7b7jU0R4McePD/5/nxaOP9bGRofjlDemyW5J0WigKaU776slePR10bicvBOCeONZYjAm/pFdw
KpHBv7iUuJDLDkcCudlNmAT+3R/VMGFFehJL2GziBroK9uE6cCUX9YBJdUiVurT/P//ZkrAcuIjm
/vgdMLqipmPsHm/t+O+jjeXijO1p5oN7xFm3jT3pmf5mUVNkb880mtQOmSwerHOEACxb4U7ikFP4
EvEKfaXBXLyppc3gU8rkm7q1kdFOi7Ewf1q7MgNOLxIsPZlUfbZ0PFkgH+J6+tUZurIrBgJx+tQf
wCsLovyZ27T2YVPOcQ89pe5bVdbxBtdS3Hc5nleISq6PY7KR9wUagFnPewQmTx7s+KmiYrK7z38d
39NP5UOB7jkY9kx202XrkfERIlGs1Qb0pKKL06u/9NgPPXGij/reCQ0N/M10/qhlzvd0YlYtNsyo
UOIJ2UOqd5oHpa7szdLR/G7/vX/xkz7t+CaUq5cBAs+tVnFZO6oGGlbpOYAUkIIKf2jKzLttX0lo
IqQUiCu3Y2+uYm8vzqhadwgR2hdN2+LjgYv0cMyqTdifUALMj0S4hikClUc78V5ANynCrHVCJN1L
qxvnS9i8y0FSCiBIg+TRojBQhxPW08ttEZdgN4qq9kY2FKE7hYP3oCE0ulkfidhZ6Z8PMsCZhBIs
tCZjMEu8dQ0zaWbxB0TVFpRt6HiXWRlk2Jq5+pr/9CaQ47xMY5KZu0y45f1P+p71oKLEBhWunXIq
VqQ9oN4QteAMlGkSkgDtYLoqs6KREOWdx7UD90uDtvTrjAwEUsNRFG2jYIax/XjA5ZLDt7SEWFRC
nLweaZJqud9jVWXd1cuVrJFcIwYg3ThdQty5Vxt8ULzAv1ojulbrbvLLS53BvGyWD6t0ouJVtMl7
PrQEZFttO9W5aOVoET6UTdJtPmjzcLnFOPGKzDJ69xK7FH2UbMKl+ZuXfEsaSfzQBLqpWCsgCxs/
TQII7Cevpm4BPMXJQoWFZwGDw1HUIHo3vY/zgGJUXPUPV0zmxbstP5us4DEf7/66lhPnPEf+Crw0
SXpjCggHR2V5AxhYD3GWtqt8ViKwK3Rs6+7pJdDoEslpccYGsOP8q4LWDMFy9cp1DhVgcEg9xxj6
ElvXvoLNYUhfihnKmhkly9XgKVoGzaiZ6ShYBWCe8WVOZIMHpisQh5yE4UVypLwdu0t43a5O/D/B
eobKyXhXxBxw4E9mUhLgk1B3MTHjgC8xSs2G53s5U19ZeuuTGu6yH52ksqCRqx4JbicyNvwEZSFY
L91bABTA9DV44du+LO/edqE1E4HWAUE3HcqbGZYWmc1S7wzBtIzkJmExj/WPt4ItNBaxgrrdFZVO
K7rHD4HSZh9GQ1Irj2E1u2oGptbw4KROTfS3nZeaWvtdZGTLxEe68US/x7tmTE2W9K7HMfMsgPyL
/rINbqFGmqn/G0z1/n52DOdFi1wvnf4mp676dqubWlvVw904yn4/aOQ7EAiZCe4QpHhOH3tU9PEN
39IGT3LIIlnKzERbrnZImRjNkmnYRvxdX/9cc/Z0SNSAtvie/rlXavof5DVO69wIWmCm7VJ9Ll6w
hItcyRT7O6f+R9tS2hj08xi9H3feDlYOWuwdPaV/ZqpPItn2YiI0mdkw4elOlqfxwfDJD0E/nKb9
O3y+TzrbdOlbzJN/c6PuWXZocHGx/P8WnPnMvAtzGn2zcQm9AwoE/CL8IsXN/ueNQ4cGolh9DlOR
p8kmQemqw2xMyV8Y6aZrWgn4WFWb+xM35dB5tSHde36iaJ4bkaC7gdmKyguy4eixKVHa+68ixGVi
2qZ/8pm3e4pg+b4Fa63i951KSC5Qlqmu0f3ajbK/kfWNqJKWt24iMo16Ugc/7Gxz0fhGDXKAbPuj
MLTSEYtz5dBTCEwPu3J4C7kkktoouvsLc0evypkm+c6OXGvP/BT8xDeMOEPBIK0rnmmRj3Mmx94O
mg6rAG2oqo44KjmR9AKIVkLrDWwh7Oo2XgtS1VKomNLpkk88S+i5E1Xc/yujNNIY2wkYieyss8CJ
Dwq0dykP5q6vhq2qbctPqUeQ1zWuFy0qlb+wqPvXKNMfx7D6GzPlod83OI0wUGngPisb4YIs5RaM
maw9360VNG2lVNuDnWDLmVjWluj4sWaUgT37/REL54WPrjQ5td+tkfreEn7BFc8yQ+wVaP7BdBok
M9Bqjwh/iKoNYLRUe8n1vDgHonB7+OrWyD1dsbz4TtHq5A47rU/3E8AcDU9a42LVvqbf54Y299r+
Ok9cwGjXJ8wBSRogpIg40VaWq8oF8P90AfrmrnxDNkflsQCYpqHrvxTDVGBIPDewoYPJo8TQRBaV
5JBSDYTIVLdJtqxn3pfZO/KWRTMIsxCqo6w0+aKe52vGgUKVwHpCrnMuct7vP2oscp5gR+hmCTJU
hs8zKXieOj69en56HhNWAaqZXdRdOuJ9TpUZbKTjijsaLtk5dPiSVUrHkuLARkv59RmfZKnPj/ql
L49g5029akXQAGY/d9k/FvLjSmCTYx5VkiNGHbIPeHU10qT7r7dFhDIiOvgirWXhIn/jLWn2oFW1
r7T1PMyvfL2hXpUJF6O3cxaut5XP1JuUoVwjA7WLXGleXFRmaJ4wuUlK90GDsH8ARzHRQhT1jai5
lOo1EkpWiBhOQb+snmPw3/crmVDD78GzSF8m0uuTBUw+4pRskjCNLkIjTPtyl+aRgjNy0mahhK6/
Cs3L55JrlqyoNnu1Q9X/kwZ3AF1fQnM4LfYPQpS6nNedFdarvd/b3yaQbyvN4fU8Rzplk9Tapc2V
nYa8CYj1wV8qbhK007E69AwREm+ncOAc6ov8vywpqL/bB24wyZTXezwBhQpq2rtPNV0N1s85e9K/
Ox24xnBv/ajygDTZjhdASn9N2gA/ZRfDofZroCcU3QjetQP/R09sWNm7Cv5CALEr34SxkxKD99q0
EyhN+hEkx2uGPU1vJPWomV8ThaTk7nWTHkwaXzZODbkIrpzxYJXQWe2+U8qNakXka5plvxwtIeTT
vWapfL12Pdws3WVr9vzchxq30LzvOukjz98YhPCIQvXjl//16twlbEIJeJTSX+g439SE5/N3hZie
9OmVpW4e1KQo64PvbWFVJdxbYw0/MSgHUVVCVoowNXIJdZCEPfb+41IFqM0FCgsab1eSVSa+JMkX
tI9OUTYuwbZ7R34TmOxaHgy4rzloazRzN5/Xg5OKGKpqNJq38ta8orRVgU63JKRKWFvqrRabcBGQ
k2pD47FNP5hOFKrotCx5aDF9SgiSnk1kl5vNwqGV5HbgLdFJR3XH4bIFsU5hgZBoD9m5l9ICl8OY
R/lyoUlNr+rt0gJN42U8r7F3BIDtq0HHSK+m107EvYH6h6Qpo8zBxftWs+DISYSYYsT7JO3jNsI4
N/YYbHMo9//f3IrnYBkhMs80pk5D6ssEXGOJOvmF5viCZbxvWfadfbDCCRT5vXJeSk3/LEGts9kp
AnAIKu532AyaqN2Dky2MD+ZVm1qgh1zy5twuRvVUpltwU19CRZvp7luJN4TwfdYPdC+cj6ZLoBwJ
iphPvEiYdKquJ16BPy8p+3wSkajmIJFiHBSu8iZFpfCP7qO/X99MtLwCOt3dMrO7taB5tLPNHJq5
OYz/lJXGNusmRo1wo+VmAASaOvczcRNHWqt7SvYdHZt1Lt297UN1m9Kr/LratGmUhvpSa9dQmvol
O3i2pGWFD2Co1fjxcoMytjdua0DacMYDD2ABkrN0ZYHBTdAZjWj3IZ4fJwfIEN16Bv4ThhcxiwkQ
a8nUVFgNhd13tcRkd4C9txdR1vewmNZzA5Cq0A+6AJ9TyKyzFZQO1/p6Y0RtJFVxmK9STNz5ZoqT
D+KMyGVgSFHisKNsexmV2pFcWhnFCpfMAoN4wdaGZPyp9Ir87rvTA1J7+oC0glVssX6vVNKG8HSa
2OqIYhFvNoR9huoc4lHaOXmluZ7p/MZs/bvSK+Xx8GGx+Znml37kop0PGVrAYEdkb1VFG8npa4cM
46gpsifRep7hcCK66+wXSJ5xil1dF+qVEg+FlCtQ+PtGyItILmx4o/OsT/ciDUs9KkrYUzqAZwJq
zU2CxvMkb+oItsYarmx2NVqwApmc/cRNeKgUawHwSDVsDDCngSSdvo9Xh5IH/vwW+w4JA2ooZAbA
DP+GxcPaCwL8T2U0hqRn/tEoeczug33bxVL++q+nFZuGM2YDLuv9u94CcK261JzxNdFQj8hcZCHd
px+b3k1IFpi7kl6iEXE5KCOXIRfGTlAMZgDdSfI0V4y0E2MRyyU8aQ0/PrWdMjEmM90BYeXiS5Un
caO+2Ul2ubiI1m7M0AwRnwkwYmWwIY2X8K7p5WmwWLiTJfi/3NfVmkcHFXkEa5rKEei7V1A7cPOc
xxHpGH7RhWV6Q8WObWD1jfzaM7EjO7w+E21tfFsDzOTNkpmOOyfnH4u0ZASQDALKM9zwbSvSo4/e
ymTR5Xm2AFZtb0+lcnRTxIDecMlP1moK9aUK5Ea1kBhhTedkIzo2d2dkKfu2+jaYY+C5LjIJX5vz
cG/FH0zRgTrtFaYQJIkr3JPe8XtSd7Zs4xkILlktiESekm4Ez5RNsCgPtsg3UO9qAyxZAJiaVt76
qp5zgHcXzcxOm//uwVuwCZe/Sw5hZcBCJeFoWOH1dOhLzma25iqAvbcuKIjRrHCdNcHsMp9DzvzD
vcjznRAaYer8o73LiKu4JgF9vl4ScsHnuQWmePPjBXnB822NkZz1vqMVZOUR6O7mNHfZ9RB8Qy2J
eUlYdB+S4j1fbIK4QEpBoIACrNN0/Mz5O6dDIlQCTcURqs9YRZdgC3pGoxU2sT+tasxBWnppUGfN
XktZPdzX/cz3GaAbZ+L+oN/LljwE9RlMM9pkx0QunhPZ0Xjx8O23K1Vj4GdY5v4EbAW4+1OvQKRW
YKcmVaRh2rSZEPVENo6v6fQSGBMSvT+0NZBwBdPVIRCww8MffEKHcI1EH2RhGpE7aD/NnmlkL64t
0PWBVeL2bNfvfEh6alH4TAoXXWSKPjMM9T+cjRO+tGVbi7TLI7TH/rkMOPvz6z2AnvYc/QKqP8Wq
e3czxwkryY/otBjU9pOYvfzCp+92fOkUEPvRJSZz1oZ0UHrGG41618S7uiiKjCDJ0pLmzaMSWlxs
4jegMR57fBpmVFr2zqVhG0njR9fb7j5fOWJs+pqIO+vL0JLtL00BYcCgtseqH6zFIAbU9IaaYida
vc8VFtNGQUN3D8a52SREE/O5qsDh61xhD+GlGJbALh8x4RKewVsJwS7HqX6fbYjkhYZT8TvezBb0
coCbiwlKpwVMeWBBa/Ajyc6FcOVFBsTq0Bqzz+fv1LO/Z5t2/cXuzaQR1Q03mDdKnfgufOok5NcY
/ohqQrgdS91B8DoVFRe8EtPDBUvf9VV0M6swLmHzmfFSvlNOCnXRwT3FwaBqWZWEvFm8mfa2OY1P
6WryzagGOsIG/H3Gij32xNLannHCKBqXN3EYVb5wP95/BiVWCMQVzYKDVpX8Sbde2/BUSLxqFJaa
gj8TVWKL1BleSqKd4tSYCY9rLL9IoOfOUk5wVApYZy0t2Y+QvzytZ/2+vl4uKey/m7VIFs0XY2/b
V+fvA3CE8ynGNxbgxYRhSs4Smhw7A534iTRvCqH/wKM9dL0vLsAOpmdGmzb56EOqis9cLXHn1RY1
Kn8U6OGLyqUJdFNLHMKgbpfucJ62xx3gzC8deApk9ImohIrKHAlyldr50FGE8mP+4fmeXwZ6Vavp
+snMi4nSIA16CioMVcvx3friNqfRPrQV9tivGjHm6g9gXhtsTqxaxJYXqXit7WvbMe2m4as4+Bvu
S/HsFHGguJ/TZJC6i3U+O0z3tJVSsa0H07m11Hi3/p8+BlBSgWrxQOHeMx77dfvcWL5MvCznQNZ0
NKNORvET7B4Ptfp3tRRNovwDUhuKvl0B3h8oUFz6jvva79ECQoVlyMH8phnKfeWhEfsCQ9uvBEby
CpySfyIsh7hkThCH+FVMp6BjpKCTb29P+TBGy64UYfUWm7rFyvKTnMuFWdxPIeejmKajqL6gxR9r
isqix/G5GHoCw5Z2WYrO2EyAOnC8FDd7zYUhcn8O00IhQ4gHo8Din+ZR5w0tr+jsWa6AsBRH4sv/
He50liAUXhdzjgjRBmmVlkhRz2B2DboC0cTd8do04SlnC7y3zDJVtdNY84qoOlAuTpcKQYYJvMco
zNVZAaenvtQTRZAFKFXxPo0g90GTgbuiAgXMYSFSeQPvszDM5+0bhNa+/7jiRp0YHkaVZOhTcStg
3AMBowMbQ3A2f2gaBAzROwJTR+1Y+1J/FEoAHUUdiMKrFcvbLmdUzys6G7yd+rVZgla8dzXa0FB3
fyiEVgsYv6LsoEXYFdV489hYqR2u4+KZ8nIpyaue/7HZ29aS4hK6OEMGjErlLfLF3uwjD4q6/uhS
52VI1+4u4r5YF+q9Jnj9S9dNSITTGNHVyTYJvs+DxogWwSgmUQCsWHKUlOUdcww1LATMgwwUzw/Y
AGyqYlLCzToBM09Yg8C6RxRotM/TZykVRqq0kaehPM8jw9B+iCxJeSQUN6vXNryWJnJMpP8ev+H9
ZvaESUI0pn8fXXjDY+BpO6IAt/N44Kk0si0Niis/b+K2/qm751aLoKwgkxB8QuFLWNkfqjn6FEba
18vzR5RI4zWDDLY6FPGXnZWZRb0fWmArUyr1uPE1wGwERttZsp1wEwYvTAYYK7py3wKSJTi2+NQW
w0VL6C+l1Ts3IaEGmvWsT+ezWj3O8XLwomtNAv0MxB+esxmp2JvA9LVb0kskvGnyciRqo8ybaP+X
bj7fSNAyvJ1e5BzHYJLGF8DLit4Pr7WzQSaf96XedeGLLd2L936pt+182GqgETlQ2mkzctsea4HY
cyPyDlWPxEoPpeUOhKU4lNABTYqO32kmznrMf2CVBk+JXyS8IRvuvJjbOtApFodncyaeUJpst5uO
4HX18CawYD38dVlrvyOQX/evYFZ170/AIk5p3T9DIvlRNlR0NqyPwn0IzKlMWFbKypCD8FLqVBN3
F0sIICqQ5YzXbeiCRsbjWaVftahfZ7w3R3aGFZDi0U/OTdjDoEo3KuzyFGG0PHYhFYWw9pgqV+sT
hlQSwcOM1TStSbo4RjU86EWqIVkVlAEB8Wn4Ou9nLSlf2KMI+JAXOhAubIIp4dnhLhCOxrjNt4dx
dgC2iv83CfE+HitxFml+wsMBm5gOOlafJp/oTSGGeiP6FO4JjTayNmIhNNhBXrCUIjSaEVgaLsb0
05FzFGWuJW4sojOYBy1QlM03mlkYB2emfO/0DBtu59egE+SIIXH+R4ITGj0yU04DN5uuKJz3IM3M
5tuXvSryQ9tD8kljBhuholeLRj11qngFvB92ojNFxSHkZqWevMr+M/JY8l/tGsYcaZfDSU3x/8Qh
vvHYoYer+7EwpUxqUeExuEylX5iCjzLx6rdIt1lpk8F1DJRwVCBMZrf6LBjwsRvfmEaz1+0g8v1H
pDJFD0RHxV7GVWVeKyEl7pxak3Jvw+mfj9+4OJU6ob5I9MPo9nlTXGLG2ku3lkTNKkRZy3YhzZSE
IVtV3saJElLDhyvBnndmgmHMO8P8hMAm3hgJrxRtOFv6jXUGgiY6OF3o9ZQhcIdzYwNg8JCo2CiH
2WPw9bMwV5xvKERZLH8sVpc6hYQjEV012AHC6BZJZ/RJCcRTU/+UE3r/DA0k7dpGb5auRXUVd97C
Bn8/Bgs7ZzaT9sAz9Fv0MQjbQeaWnoHVjeNgpsHed0o7+e8I3LsYcfDX3TUpmI7SYp0oYLYgNu1t
o/pa2gakmHNB/BJEUaf4Q2qKanL3SMQ9rgd8ZkSTGtggI++qIlJOo+WBHfS1mixrCMrV1Fz2l5/e
AxOiAU5zAkUN/Pe9tDIpdU+SMSGDkq0r1jWeCCm7ngdefu7PxnOHK5aOcoHVyBNjcISJT19PhqAE
aP45zriG3gpMItYEhGSTHBZT5ZNXhw2izCmPWUisWeQ+0rc2moZ4F024jmAVM1c4waZmVeH74Lsn
1Rmq7D1iuAVuYu9iMV+o71BhQ8XL0h8GDeAV/w0ZkMd0IrHXsbAFHvqEDRMqpJbtwsfRBs6u2ThF
+uqZBnABVU6A5tpIGElGNYtGuGncbgWG8h23HkLZYBNB+rV/+SDkGsfiv4V9d1oG3nhqtykgUse/
ifLbxnu58rTp/oNQOi8LoyeV0K8MrXVYxnWjSpUf2GOG2vXAbQ4EsVzJ9ij9+P+zntcaTmzVRGiX
4b7lLdWbBQE8ItwROV3h1tgqS0jnk0l3mxcwx2NGm2Em2zQ8KVQzBdOKcnLTJfOxVkk1UiCR5mMj
m8bclQ6Ve4fPZiBVghY1yfZzbJevV0IQxQ6ncp/cKOgOprPDAs7dCsP/7o8ZxsZDHwrk1fQjc/GT
oAYwlvO9DxnYNqQwS3Yw9EM5A9/mI5FP9VLBhscpnkHuBXpqwUc0Ib00Bq/+OqWOJSvXerUpSxNj
W8YrWH7xKEi1VYoCSYRe0HWA9l5I2rxwyAXB3iLnYii5vUgK2kB/0gS6Ktr42tdOeT5jVvSIrpKw
eqrWWFDRv3LlEhzMeylo47ezmrNvN1u02P84aTl0Vr6RP0Po0baRx8tzqPFqA+zvcK50CaB5IiXE
bGr5QZjP1dmsNNlZFGLFnIyhHcsfSXwaDWItOdbOzf9/frWAUa4JwxlGoeHkcMwFZjkZFaA/ZofX
NCONWkSL69PUms5eblXyIzrQkgikXpzXTLli33S9/HEYBMh8PFxIjAWHbeE4/nvpa1XVdqjsRfVj
l+NjjOHgFY15ZSDc/3DlxW2KktWFfE7+jVxvGrsB/CzFX5DziKXGXcIeFImfEz/EfMzFXHl3r78F
xcStS66uTsta8EbtkFvaasx188u7nee3ttJjszkThGgoZ1YY+UMwqLM2kCKa3oLhgugKJ59Zf0YF
D64Z0AlCR5Vp80YapxM07NV5sQOPzj3vCRmLdvJgxXDRLUU15f+cB1v5xZEavHgECf63n9lhRHiW
I7LNylL1A1581MaogE2qlh5cdjd+/UEQoUhVgJR1g9L6aQSCFMmWvaxWNLjGOHFA+Ti1dvAhRf2M
PJUyUvMo5fytZaXicrxAlTHHVHDk+otMwpWtBZGq3OPVd/oRKVntlO3jrpSzPY83XyRFawI/AwyX
1pq0mMyhdfPPQdVEZeH776SzrG4/vqVESTptkH/sbc18OYC7Ja3LbOQdJ+v17FdzPZSy3VAe79Hf
PJfKWOmg69haRxxZIUkn4xWXG71ybuFZIwtUJYusLiS05FFItiUovx/dxok7gypwzjJRbLBBWfci
+WWDFQariw8XODD0i/kBXLvWMDzYmBECWe7bsvN+hzSYI4pwtdYdi/cj4Ls0smgZfxnKD8AZPwU0
5IaJ6rt64OIICZTJS4+SYHcTLfx2uYpmajozna+AM4fMvmy4tSs5whPHiOx5xExBzsrGq1i87CJH
eXGrWGeONizYhxwxAYXoGU8ZkqE2bESb9lNRT4G6EvWFW2n1PNlH9/Syw6PIJI4h3uOwSRM3r6pS
ngisZmG8HWeqonri14XFbltE/lxt0pmIhKs98/CDadojDZ+Qgs9XwXIHU8CvzFQMu4TmAkT9LL3y
4z9nQdKZx/esnU5ysQbv5Do53NIJNo/1UEa1rLGTL4QlZ6HPOvZYZHgXBu7Mmg+pxC6cS6Xu+6Kq
h60ewisnXqQTsglY0IGjbZsnyd5azMbBhXOR7WzpLKNLAXA77+Brpbq9p5vJMf61ACkLL1yMPtfb
0q0A0k8gby/F8FrL0Eqgs12oJjtt3chcaAW35ZVIGFku0lcTRUUVHsNTEXo3qr1O0/DovY3eRR+z
tu4avS9PqH2vZuxnt2eAYw6P1cFNqfSnDXtKDlBSgQ99uoqiHnCnhOOK6s1z45ME3MpiK1UL4azn
cHqcrwX/HCMaWpQHXJ66B+VEz5ZO7YpnyqxckdQ1NJwMCBcjNw70sUrQpxawk52vzMCrwt1zpbCL
tnjzgOLdMn43xUUeztWN87TLuP/cQ9fIQRHh6iJOU2QOqQVlObh9GfFE0fAn4pa/6o4H6jZGfGZk
HC4lGv4qGFtcx1zLC2ElFunRqzg6inqm5Lu6/p+EOVhUUecSeOZF2Q7Dml1lxrIQYiKYrbl1+LIp
tVWEHopx8m3fy9KkO+HLCu7KSLSqHNriRW2RU9z5D6g3GlCrCR9jsVQUizsPVLmE6UHxSFLHdtmh
pEeU5lA8r/XGTNHHXYHtQAG3QDVZIm0KIsfwzYJMPlmd7ZA0k3vcYHOwOCmzMw6l5N3w+9iEWkA+
MKKm1OxF1ygLMtPD9pqPgjrT/OjpY/V/3apZI6z1nJJkeFzng1vK0tg+PXYrjxhZqi5q61UJUqZN
Oh3T4+iNbVmGDLm6xlYw561WMzSGZiNf7gwsXqHXiwfMTCvilQ/N9tq9x//ynsBTYqDe9/SWTbMq
iRyM/T+sHcm7/VsYLuc9rtV+iws+5Sy9h7rx7VE+tjZLPNL5974w6rUqiG6yMHkuT+r4G4cUdw54
sJBSU3fSp0VnqboUtDQ47XFdyiGpMl7vn208NwGtqRpNN/0pwvDQV/EHSZwdwWfYrrC5mnAM/KTM
LQQIWZU7ZDoQMoYLB8eEXDsTMxxRrHG+RC+hCZh24P8dKZVELWN3A8HIKYzB0he6M3gOR3Gv95cx
ie8BrxqPMb1PbRJqEXm0IZt7P8C/TfhY3lCQT+6qJiXQhk6+EQBNlgH4CGi0PHMZdClIbJRrTobP
LCx8BLI4Q+s5z/JjSp4vIujlCy8/ZquuOmV+nuB0hT2bjWAbEiut43mcePjqvc9XKRj9ljZSkHPW
hOEIVkaIdZRV3MukoEZWT76kXEXaC85TOOHX1tN/fRm5yycuPLNJtcOcrcto6qHQ3dHV1RW2RqzI
XWb8WZllWYfsGNyThcIH1g77sTtH57OonYXEDPepAPdesVLxBpXB0wco2mH3IX+Z0JTItJlJAI5q
wDapr3oRkFBhLUA/x/59PLnZqWD+gnuZQOS/vz8DHrUXVCMockRmZnKdyHiKSgl1ZfAB3mdDaFWn
jyj30aTrPUoJKjDCrjdIDI+Bfpx4WFZ0dpqt/1rz0BFmvG6+g0a+TjyYOqQJqyfv6KSFTPLFQ1P5
gl/W7w2vKHSUhVFdGq5WW2rBMEQ32MwQriJA3oSZ8EgmapMCi0lSft1Q6Cs9ctko2v1CK1Qlfnl2
lUAf90nkiQ772xuqcVIdMtddmGfGsIiZRBF9KiZLahNMzcYKMG05rLMfnkTqLcy7LXrgN+s3ZvL9
MkVL8zz1wwm9z4vPwvNAlihPhOB1YqtKYBqFO7s/uD/G/m96a2P+kOFOm1HgErziGqNsQ+K7DieL
m9fArDHuRn3lf6uDKXSTFqXPlVADKaQO6GlOu+Aucg8pkjh2sZG0WmWkMGEBmchn7t30KrMbN09V
aJWml0Di/fHHQPpHzOs9Xn691/WvHTSzVumP7CmxeULLosmrpwykLjXOtSZGgoxFv+AhhzXZv+L5
KoM1FGfgyrpavpwcjKMJRDQl1IglXyMcol1+diwYZo88wOsGqRHFy/FX11cR+fB2byN9Qx9NgdH/
WhP1XMkx7PAqQkaLpwOAcU5LS5AAzH44Ley2mZhdv+AOe9JLMuAZHnr442p4GBN8qTwCgQZfgVNb
pcUudBBfQ15zaOx9BzYaELHbc1+2Q2/DqZ+qlyEymVRs5rH1lsFR4sRGIwnzBQictXuNLL+Cj35R
y98dXEqlhLTQMOmVaCwhTJxP9ykA71pzF46J6QUXBakGs/Jo3rbCWPTlKMlOwkb/VWiITvZ0F2Ov
CthHF7/IQ7rq+NRhV5J4/xztPTaFt3+xbWU8gNimkA5kxLV7Ny/piyLdrnaIsUfFHRVS/oad/+s5
AyBU01wNnaxp0iY0CJPbZshO9/T/or7i6lJPlwCVlv3pC7l5sL4aDngu9gXADHIHVgcycKcReBNO
GzH+Y5rfyTsTZdYPpyUqefXsaZLMjFHcn+zITsIHMo2jx7j17C2838kK2u91DE3im8efcjFNn802
7S/zPl8tVM5PsKVhrTTOvxxlVF/WXwUeg2lpCx2pWRKP3Lvq9cJnUeewRAXs0HkA+4Qg0sq+mEiR
5d9kC7et7i4ofsaRSMfL1nNqmU+k1oOi4wALlC2hC4uP8eJEROdQMtiNpjbgfnPSytyl1fJx0fwS
FT/6VLEvRUi/77mz1uf+pIvpKb/8Zp3GjLQ79weeQMNWawEPsZwZJ+MSDcf04wrTRS+c7ENHohlH
B+2beegzNt3opqkbJ1DwTpqLTyi7JXeYIwfqvczqn/lJnBCiFZzJTHj/xDjMcL5q76TjutgMrej8
TaWNoMdFarOEaFuNKQN9ypH6sWmL0HVraQ8+wiABqL7i1FvKFlPkvlgFCJ1kV/7MMuklEQqQ6Fh4
Inr0conC7nhaiXt2zgLfrNbZUjdYI2jsFakLKIm6QdhgD/qvywsGgen9vtkiCo5r/OthSvNRN0Lf
gBGxqgzlIDwq/lGMLHYG2FnHby3dqBr/dMBfyTM4nl9/zYlawkA6NA2CMR4tOeZhJUsRR704getc
dGKoD0evtgH9N5/FVP/RjD3U6DPjMwZp24alP9J6rCFFjk4oYMXVYitmxn9PH9mLcQKld1AkjGjt
dLIp6NDugegS/j8vzdF7Swn+/WKltuWC6QZ+d2CX+a1SPpENO0hCNjxjvyY1f/fs+1j3Gj7ft3Zf
GwuqBvYmN6V+Y93XZen10Rsc7dV6Uv89kyh6pCK3PYxnOzRr3Xsdi7yjScClfAZGiiJF8lzwduUG
8ywJ0S5I/XiiDkS3EFYldwh4zUZ6vUFpC5Sm+GglY/V8NqSf4drq/kUBcDBNdwWNGkBnKRh1VESL
BZN/SW5YVBHAYfk9z+den1xW0yNn3D0bEy+D2rAov/jG8upWKaKIBtWsLNyF/XFu+2eqwrEm1Z3p
+LzXRVGYaItI/CpOxDw+Oe6n5nQOSBgfOX31JqD3cJthy4h5WB0TBIDFaVAsIK1kXyA5kR+Hbxce
Kpm6jC4u+hOx9i/MznORIgEQ9mU/mes/m6w1OrV9m7faPZ6tZs3PvWRLzwnrOlExz15yMm+3yRrF
5FAo9gWWQRwDFIn52TcVZAH45XExHFxJX85JjfmIfTBju0n8lm7WZ+9gb/HMm6gko33Cykz+ZcsY
eBZpt1Exbo/yi0Y3sUlZME3ST+6X2Jke4w26uuLtA39CWtZIe1lLcOoTU83v8ZbOInkpQv6jGF90
YmzZBEb0CzOcjANyqqxX3AbkAPI7kcsHPZf/HpvPl0xP/qPlZE+FRxJ6MM8r1WKg7+yx9UWtO3El
ld0pallF1zSn41Bd2Offpgtzb3b0mBauZerTdKiUecfepaZhCVALEs1W4rqeOsLiOgsFcWHqHhWn
Fuoukrh+zz6iFrv9doFnM8bKRmq4TSVc6gRz9TLdEDCscFrp9pug/fj5nZP19dVK67XmdSo+jSsQ
ZGqN39rDq6lyj5UGs/S8IFK4cBRkEjFuDs6B87UBWf9+qNLfiH9H2IRAzP5t1Eg3vf6p3pOcuRm1
np4enOonuU1Pp5KHlnLmyar0XM5nocEM6pQKW02s4lGKZPItqhJwoBGoUKA8zlfGzRVpTFGPcmJ+
ImjK56mYeR7BkSpQOnVXD45IkWfvTvNjno2zhEnR1d0Jc07X4iiBMfeMfO94CSf396c1kJ2MM+L+
3684YstwsCZug4PQRRGUJQDXC+2rZ3jm9sC9Jy4SHsislI7kJ+irrOxnCFaDg1UzF2Y3dB6i26Z0
gxJpLS7KC5IMyW+QBvzcT43lOS6ZcbWnrPTNn1ve56kSMuaz1YSJALqRWh0Qr2s7IH2CRma/w7fv
8ojjDcHKplLGDOipTQHjuO44TzpAQK74g6dn4W+0XQotkajLyuv1Chy/cmTFAGLg+wfv8gabiGDl
EigsRzxDpgHxWW9+0brsaqdQUW/Oefp1ZWfVo6D57Ba5/meLX3e287CXN4Wf0UjVoWYpdnbYlIgv
dGaLIIIq1sgmdyoNePfsvGYQgNRtmeE4r45tqfFnvOuE4U12ZefYkwX1JMfvmFzqpBiwBdiguPbw
Su/cKQdlicFMecd3ftVkt6R6rR9+RhUr9oDHLyxHvag6VjvFRn/MzlbVAMkpPnu6Fb9BhM1GQ4gI
L6QjnjdoG758pOgn3duHm0icuKOw8gjGyaM4Z030P7DBpS3PO+xGaiszeiBm9dPm+Uley8T7lDUe
xiBf6pa7tIoWr3wR1TehsyRsMV+qWbjctNUT6q/w7OSSHg5yylW+t+bO/UQ6zuMldr7cybekjnEy
qSK3iGqle+BowaLNWGFBoFuRr3nelbneyiCyWLQg6G5KJpxKHLmdkx70riTnql/cFfNkcDLIEvkE
u9H3mpDq0C+o8YZvcsK5kPSUYI+DBq8DLIAG5Q+8irQy2F8pCrib0zAFDyd91maGPeSLHgdscRTv
4BXYiuWVn7bodo1pFw4ByphPM4ZLCcs/LPT3w+EqyFACqTDbPvT+YSQbwpct8BX7+s0F27C5VHqh
P/aL4j/YCToejMKSxrZyQ4a2vM0NY1n7X/ZVSCoVmA4IzOxqrr1+MxJo/KL+oNTXe1hYE97inb3i
V8zhJgyEKu1z7umggylw41RQP7URVUDn5XScBffkIpEgBqOQqMskGTIFmk8lYfOD063EukrYLRga
jEUmAz0gYnXHKqBSHKowdqkFVdoME5Aa9+Ri6X5mTtwuQIFAemLEMJpeOQWZzZoh9MzSjSRbAWHA
DFqrqnwBn0D//3kdegtAGu2vjvUrgzH4jmC9mV0vBj2bTdqPyDQybIQqVH5umLx3ZXaYFE6w6Yfb
BtekSibRTIp6MoVeFXwoynBjlvpLwrl+D89GZ6gkWCYN3AvAivfkeDm+y/vPdiM4kLNdnvg7IBJ0
JYGKfATdkV5+ScidqwDdrqqj+JES9tanZ2d0iWlW8P1OXIg+aJ3yoDVBuOJflZKb243/TyrTrMGg
9jUsP7/D+lLWcDNroE5nHCyPt9D3A2Uzm878Kk14r6aoymuH/Tqpp/sFzBjbFqxLikCJPWRBrR2D
+ej5qMhn4kTiuWDjN6ovDBo4y1tezSifMRHDA8s3lTQV18hud6Me6EIwy5ZruPyFM8gfmgTSLKFU
xdC3IEIS+2UXN9azCYOnhMCbw2W3pCukGSWJk27LCleKuABAHajPZein4VAGTx4qnVtXeUqFrrr/
x20/6e1eRYf4+wiT8VLQu/YIEKI7z367Kuhp8IzqXFuHVTXPs/Jxrv6B7TYCQq+M/Mb2BaMYcJka
OvKC43D/lJjvTzCrpm8lfJsEZnLg1GTsgv4TrXU4DdXpvHtL5Qh9saKRsQrEl7fOTJYC7anu4iXj
ol4Sl72VGZX1ztFQT/EGuSs7HiZ3nd69RTrLr+uFkNqK9PSpPLBhsF59ZPLvxW922JoNyUculeoy
vK8mFsJFY23bpY14XaN2WGpqLyNlF7bmIa+TsmqZaN1w/uulT2EmEvURPlFnsR8v/836HaE1oRIX
W8KNF7uGUYlwPXSMSjUb6Ka5trP5iv+BmeBGyhXMKleNxdZThey1oKtGWrV2CpUt2lNM7lFqmYvg
riqbGhvQZMcdBT8uoancjrMH+Z9K80ONLf4TvAyn6A2R8Vai7D5FWgXPOG44y329X3cZGVKhJ3pw
uk2kaX/NRYPdFPbummyqMsPF7geYZPWjoFLOyml7kA6lY6C1m8HdrTTYz85YvSFhWCci+X7zMPxp
G9graD1dlMZ+HneKAzf4aVgOR8qFizCjapBJ3rfaqr5BsgIeWFofjS0CsPMCtGsfyphk0c4kTF6o
YTw9QLdEtfk4O1iU5ZS6STerOGkRbP2Cyccq4LlnpvEzca8rMfNwQJevmL/2qE/U1H4Cx/cfvaMs
uuQBpgLn0YcM7kdg1gnckUdfiar9SkhCXk0BsyH0etzSdp2B7vQHSeadbO6lR867lgcPLhD0qUKX
yptPGDYmc1nMxU6gKrqtt8X4NEr791KDplpeKbJlG+Fn0JTjAvMUexmSWusYfZhplXIYMm/BwXV9
Q7FM5JqmHEzkJ3UCkJs+A5OBDcHw5+gFBsowR2NaL34uFS4oC3qdv0Ojz+AVp/9Pd8Ar2TynYddV
MBXXCC6GS2u19BkNI7Lt7SXo0CATZGYX07/93bFpDlK2tEH09LWm+1efypJKJA7vdydKWVkQwLvq
6kYY2/qzMLpdRmdBsJ9It1WvJWo0pezx/aNETlHrHrzHl0LFs9vIvLAgjb605262RN51YpxGc1dO
t9oVp0MEY2uPR+2bzMIBEOwy038mI1neY0R2r22e9KvMKIjgmqTf5dz3QuTv9rTLlGKjEEiZrDWD
paAofosxcN3sBzzLxTFNOuCo83qh0FB0g19GoN0U2fsUqi+hH6WI7nUSrZgMRK3f3E7A52fbFB2/
fOryhtkHXkj45il5GofX7GJlwnJ3upCKueEtDEeiezdpWRzm98O2hnTY8gUzwDKAAi1r5/GG3/87
wr9TmKmV9sQA1YdHRQzO8TH4KtE/yh2wKmijz56rVCRV4ISyJUMjrdiVw5aC+6SBY7MhuKcNeTIo
WAgILRPfeyHlHPU+i/78sIVhHLEygrfIZ8SlBC2qAZygTTiiHSP6nzTExAczzXum/TcR6hs1nGOW
BJWjcgOmlZ+ZLSiCmel20InPWKaO1oV0FSAOqeGut+DtTC62xDBkOVd52PyTxUZmXSthDHxr9Kvo
58kE4i2sXklY2ohNqrlXQJCSvYwZvYnwqXr/BcWuqViTfdMye25HRMzXKfLkDCt14xweZiBUvz4R
PMbo/FMiCONIV0C6UU016sC3eZXrShjGNAVkrf4x4s7wXYdP1A6hO1L/QHbjq3qr/2ocVsYDyxhS
w2WK/1vts/uRBfIlj2NOq7ibEBPkzwwtPQhDSlKWrzlOlqGL/EzFO/11YrgHlAH+O3yE7ICDQEhF
+MZrmp4HPepd/FYGYzXTyGdK94eJkZN0UhZRspftdNqf1RoG9zLn5vL7scARaROcH10cHlm3+8He
oC4rg1VMOJ407A18Q3fob5MralQ62hpEoiVTEEkT77xG93j3hrSzLA9DxH664UEsDV3cP8g5hHYm
u1TcwK2VLsj8BzbQ27yh3Te4XB8s+G50OHqzheR0bIp2MMoGVNqJTczzJgybjQRp5kVMqypx2Fcj
WHNNhCi581JIZcwdwuRysGlieykwss4YgK/BumJOCwUgJ8tz1usOF6Q7OmK10YZYK19XZdWVUMGX
QJLJ5nnJdlvvDVxmBY+3ld2JMVDTHaOfPvJWz5r5uqjyBFde/gjivMRjYPKGBlhg1orTwFyDTvj0
Qe0wcgmz8kVJ3V8KMggjBegxWJhBbN2rgwdjw3CF4iijd2OSojz58kOC8NZBRIJyRN1mVm+d1mr+
ZMxeiysI+SvJ8IteUFKtPv1nCZ+bJvpIdR3YXIqmJ9BlePfoXd4idQMlaZm46elHwq2YAQrVn3Rz
VYkCmX/A5vjVASicbt3lwpgX7RfC6D3+NSKBPoORdoOP4LYee2APFOqerUTRzgOBEXmOZrV0GXnE
WAWSc2AZ8r2+cLIu3KmvYKzbVyx0HpLVYK4FXqWpg4135QU9FX0nFc2OPKntz+FnfX8DnZzMQ45K
fQc5mLTmR/5mlkj2og+0kIM2J6LIO7l8hWobkHHU/cAq0YJLdR+awusiHgCmCO3pNi7EMRNqpCeo
ePYps5ERErpTjOcrInQOpgdJiibnUB/aaI6EQ3ldtcRQg0q2xjPnJXlMm9wX0q1+DcxlfCYzQg3E
KjaC1iM4UuXct96mu5/s5ow8Pk89qjF9UMOonXK1oDVleiRqWYOhrUOb7TVYII3dlkr4+ZXm0ITu
ymMMzLb+dyi9nwBzYOwtUYI730c2KAtR3umzxzfIHjhyOzQxGTrhgiyF/Z3vavSqUkmOB6a+NUoF
cCHvkt11UEKYnTDqCy0m2CiL2G+KBGv/znhbFDFI9BBv+R0ZWHfCRNUOR/p/1npMIrW1tk4FsFVU
0D7muWYQjNZMi7vPYh7D/Pu6dp/Gn+Gv7gXR2LK7jAHaKpi9MLAVociqyOkw50HukNmPvZuXxnoO
nSv5dtt/Pq1g9F+QddeQRoolBkKnHy8PUxP78MkhXI4u/MfGDq9dztHXKcN+dudYRhc97OoXya+G
mUBXJdEJv+Ir+E7+T5u9iQszBlkna9jKscyi7HIumLH8Unjgyrgb1Rx06Ok6K+c33QgPrWK17H88
SC2wBcZPhu98j5PzQPA7ikvo+UiktPRZrv7PaO8p64SJsaQLrkXKwU/MNkHyYFRPoRDj+wyuCqy+
qp3B2M3dRx3RrIC8Z+3oeQdaDq6JZgNKQk2zu14LKcIMHc4MFxmDPkm1U4zRej/eJsARWcZcJaet
idIlO/xbeWuQPAW3VaMCqLYOeGBX1Owhl44aFiKOv1Z5qsCLO8rQzJS8HFmzvEse5437fwQIbQ8p
fpmtH/p5v0H3DmpZlcwSqejc01HVlJofPrq9ZwWXkbuLJ4+AClXRgTgyLxdpROR8UF3/NS3VaSAI
m4nOJdBGc+92cK8mvsBXDeCDJ31WMzxr5nl6mh1xLmN5p7nbsCt4yU148FWhCou9DOVq0XWFBK0Q
IIGvdWLNIXuO40DITDak7/tiuawC12eHJT7tRcM7anq7uWi6MF+BiD45MANPynxbDU7zGboGSzJf
xuyogoBCFhSpntIrijjkoP21F52QKxREz0bmgZpaT9QUIAGeD0XlF+XLb3sbWg3XBpiyjw+6n55R
+HD6QnuSsBjyrBQE49sr+DOGB+hmzxxVGm1kN9hbOsyDp5X3wghQ66DqS7xKF3qNo1qvJhcoZBwd
1HCMxw+92qpqXoOPm1zii/eSvFZzIDFQxVo8AULDOfW7IyS3p59im1joiYaECs+00ifBt9Dzq6Xg
j0fe3Zm6Sii1O6UmVe7n9sUjRL2zHcKnCg7wKSG1TrmuaZ60LcD1OrlvgrXOuDt+MbcHr6sS9kmJ
j1KvPrAZzKp0G/yvPkcaV9V4U8O7qTOGt8GMOeMWzOLaRl0GAzzRDYfF6iwMvG83MxwflS7lQbQU
F565yW2Pm1luD+MzGTsTXAYd3BNRhY/itK1WceGJiXS2ueiliVdu/DkVw6nMpwiVJRXgJcu7/9if
DvypYT0oKYS7EmshY/0/quKfavSPlPooWuKD9rv9dMMKpER2y3ND+V7QMnlGV/r951tAtrYhi5iR
ZFQBsfHtuOJyZDi6DyNWyB+0W70k6UzSGk/C8apKI19gYHYMtiREnbKnxfgEZ12hm0w3qkICpLxp
YJKz1MTzD2pcpqZq925Fp+5uA20yOhEAUtlsMn1kl0RUDEDp0P4FKNOn2Mo+ZkXNLBgLx2lI+b6P
dBWNeRqQIRSRIk5zcQxo35urMEzaw99n91bEm9cLdEM9LLXFJDYWeVx8fIfGP7mvWXEuRFBM3zVV
wrp8LSCYNMhhL+184U+In5HXFXAqroNu+jxzYq8OUWXBPCTf90ORQAg+YDAaYzS6fc3YEWLIi3vs
nqL4oQio5GJZBm6Tj5jYurQiFoUae1XcnrOy8KmPMQMX8yZYyG66nsfzQ0FfzQ4sq7x+qOYK4fEo
LezZ7qJKwh3vM7HYqZyUopS3JXMd6kdhdDzakn6TSPjbvQUa9BZWI9PkLw4wvTq/hAMPV/9zsYe0
ZQeoBxunPAM6yiKpPM1qUeq3Du5XVYXK8tX2QyDsLUCH8q+wNj+TFsSdSivL4k2PLVZASBPIWWpL
yIrTQsKic64xXYP+T+TBucVzbsSTgOufknqcsuGTqofo/Ns4xon8jZ6WVfROOP9gMCnkEanLuhY9
zxeN7X9Ft/5waT+cGhbqqAPcGeY4lslak7PR0LSBXnrmEmQjA7QwOBeliRqq+UOn5xOO+aYX9Gy1
uGBeaFgf/vv3LqQ5rCA69jzDVRqWGegVWyCDGs+4mPRW5S1X04aAvSeSMSK9gjitzbTDtHY4yzU/
PXlvMy+DdtfuE0pND1P2NxtoNjAPou7qhwvrlRx38YmO7zTQ6agEMrsn73pq1Nxr2MDmemBInSwT
kwQ0XuLkQw+6Y22+Mh7SrASsnbSYhO59+q4sBpwX3MJftkKs1a6en8fw6uQ7ZIlnlx3S0fC4AdMf
n+h5I+htP7az4IGG639GQVbdePMylIV4aZFeJq4U5fGZZRIxixleKZNUCINhKX6aQr3937zUJapu
MQnyV8NMd2rFQOBwwuRQ2BI/5XpRjHHA8sLjtoGx+5fIj4BeIElprUvznPUojn/7HbdNqzvbcQFo
hWuRCQBgTqtPn4tKBSVZISDjpLv+WXGjuEdSpkQIg/zB61Tbhq5+3EhiEeYMKtPevP5WGqCJfjwt
oVXw0dnyQDL9s5kgVC11toiYirYn+ml56La41Nc1CfGNI6teWQxaEUzfInCBtJSzyeySg1GWm2Ui
Admj/xpzYV8xnIPRxHoJqwovf+nQzh4EDiDcHydX1ATP7DAnZyd20b0bodEWre79pGymmZLmpX5i
h9O++7OioKoFpsQqfGxdd6Ti45Z6E6pRBv2M0ZsjnI1XVXBE2XzH+w7Px/UeVeYwws48y6/i9TMj
wMULPhXkjl+VM524h5M16DqOJt1MML3uIHeUqJldx96TQJ+n26TdK9BiknNrKgfWVLvO4i3nnkl5
dBdBTMWipkWTCYZBqlB0uiGYMXVnzSGygpbDI5FX9bcEV5793DDcUciG8DEDGqgrXxrk7hltD9ZH
z5NQs84UEVDlL2oOMClPkkhrGztF/eu9uKo+L/fPHq9kzf/nGJlUpSBiAI1l2gpy/mvlrDyfmZ3y
CDk9zt0jmv6ARA4KZ9UjaczldJoJUZ+CMzBvIiiSU4G7uc1Eu90Qvk/lbwdpJLJ85Hp9QWu2RdD9
A3NQvF8VCEw9EmQJ+V2j8H71X9/Ny1iXVzCvBxwaOKAvNzAJ4vlGy/f85zRfPyxuYT5P7ysmYuoA
ILHQJZUvWHWeP4PLJhQw5+YXwsfZ9IaHoN++k2Wxu/peKC5Qu7BcTem4UirWr5G7F4fV4/m9Wjsc
Hj8DJyKVcrc8P5FNy24hv94zGBJI0lYMjNXdMjHMjak9xZbHX8bia23wPaa8DdQ8EdqrxbLVW3qB
+SczfGoa2BcLE0fUUAN9SvWpVCfiZ4Q6mAbFKuucPxoI1NyIElJZMIE+HRwj1Ld7RxQKU7qKZNDI
tL0qBYsnTVj8CJDFfxqsmbOgnz1jPfu2o5IAt+InWJb5di5kcjJg34ReofVXvXT3H9wCGn4w9Ei1
CTBRxQAxQbqOkOfB+pplUNBQ/atyxluQIZHynGoPt0OYLXK8VXpuqNwqRsaIoetacn3m1stwkZ47
Zx//J1GXbckytk7ypN5B6y/RSl+I4v2+fqj66jaf3uqEYKP4MigdqKK2egDj7fncUpjSyDaKVEeq
HbecfwGK57ViRIyC7CqszJ/M2mQVTRzvpJKZHtBk9RiAqJfcB3/UwbnRY2fNrGgMpiFmrQd2/71V
qJ6Ug9zguAfuCPZ+vSthLMKV544+HyK+JRjoWynafHpq9i0aB9syZDREhezbABrHQC87qv+PnhgV
pGL/SLuqMhTFvPDd3wA9p/Alu8BXm9JySa38akQNtH9bbLALHOCWaO4K9X9Su3EU5aWxAKN+AgUW
hZ3L2iIMjndYYy2yhKafW7RT+0qgP3QBwTvqqnGB4jsn3C2VvMcf5Zg2vOfnYTb0zoIDgVaIrDRF
Q9EZJIWXCjdT5Tp/p2OI0+FzkV9PQjhmPO7i7+golG2bxEcxtILC+NNWxErG/twGIxI6Kf7kiIxj
NKWmMO/OvzjbdRcJcwUtldPaYKc3OOops2LBIPod9JCxEXezbjSoxdd8VUlYg2EoN++WXvIt6KOb
uL3Bc0teNXGDZ5dowJ26v7fcmrfF1ft0myTatd7XwqDIvC6UJ+sZrNRNUHWuwT54gmh/XrCeNNFh
RUzPy5tCwPFCQUAmLStppcly9G4WUsqM9xZV0kH2qToRkArN6Aiqrs23zOuiOht5NxP21wmguNIL
hQqL324AfXwVfaZU/lm6r1o7j9Z+ETui9FbOw02z7Wt9vIOUkqwXzOPpcX8/UmSj1WFGdApg+vPU
yh3x0/udFc0uFZM30ThGlcDEToerTVcQ33C0XkkDDFuAppZosOKJbKLGtFjUuAgN/y6uzTXj31Py
6YfyA2NPyNkBR6DUNQtrBHfqyKJ4BDyDnEOGCxMe6RYjo7sL3NVP24OcMCpEsp9TbPLpclhRdVHW
b46voEALHFS3GDGRzqirUzXCHe3WKk9Sa04jiyjznBXDrsfIOPr9VUzVN/kUdnjPdANZdQpYfJFO
B6PiE95gcSA+3utGnUBhzpOoGFzSB+D3htO7Z46pvNPPHc/5+Hn1urc6+hVi31tp9IDuUvS+wXbD
aszoKazIoFXcesyjc3rKs4sMW4XhOFxZRFco54OAF59AJltNO9RH9eyj1y/wOUzyIXCDfyHSFcVb
y4Re/D4Pd+6ikc8y2XVnN3mztDVtOYdRfvqiIPNY1xqqmb+zXArSr32q6gDg8/qs9QbpNW8wiMiA
EGs4wWRyYX8GH8ILIh5UVBMVw+8TIrI79gCpMDKixxCwP0bBWgnmVn/5GpSf0g1IDR0JXLnOX4kf
7yHt5pbwRwSMVHa/DQ9BZnTlLYtpfrFoXoZYMvmQ2Z3kC+AuonLsSjceK59HtUZytkxw16Cpn1EN
JxGwXmN5v/JVJdygVFPYUaTe4gc9vppRhxHLEJ73UsBGxbJlfiReE56zFop9BnPiXiU1QrAyVkg0
slC5FRrFd+NAcJaymu90YGrrt4J1sxfVp9CGmxg1y5Dp/WnMtlHFs0WjdHkDUPkmMrGtQzRmX11G
tr4hBmhXoLWtk7h052cponMo/Oof3QnAOqEx+VaWL5kzqo2BsR/I0M4weCfb+v8Hyg8bmWSNjPSZ
8vT4Vdmen9AvadstSqFceinyN8NGmRrER9wzBr4M9RC889L/7nNL5lyi3I3H/gqkKWVeS1YYkLwm
fMX/BBPm24r46dX7ObIukaLbUPQ24wPnd/oSSHAUEZL23XtlvlkA09Y69wGDW5zvPsNzveluamak
bSC8KXNa7M6lEAgmkn9p7UObCgy0Y4JagWIN11Vl38mV+6Y4w0z4CCHtK8l/c/XGBBnazKboGLLm
Ye2cXVwTPDVWxaliL9CrlQRlMqkJ80n9GbZzvckI+opVgaHLdzl0ebdM8dzlhWuTw+8LYIEZ4kLo
FMdyAq3L4chd3TtSNXvqd75v/Xm0VxiT92GP1fU/ywYir7w+pyXILb/nlSjN7KlDCd3ZZlx9BrRz
4U6xAqSValZvYXyc2zYItb5QxUEBPN2nPjdpzkeRl4fjiOit1qMyvP+XTesO0xch0BiT0gB8wY5x
05VSHDVbucX+3Hu5mbAbajp+v/tOnXhjFQQntrdpL1qJ4HQj4+TJRAiany7lDKYY2W6Gz2rg9I4J
cbqtS9JV0OI4IOQM0odbJdpJB07zW+qHckytIssEQxiRwW1bvvHW1EZ+rCuDAJwOLMtANk0d4gMY
ZhrbpuMHiHxjYOazTRvwXKx2B5SiawD0apPloE2ztTwtdmP/ys5ffswIwPooY2LKdQ2YCofFSxsF
VFbVHv6XnVtyI1QfjxvMVtk7eUvp8NUgKm3D4K7nUpTI6DIHG96DrbOqcvqNOUku3YTC97eur43p
G6XF1xg4IClgjapPnvXF/x5thxcCeCxasgCz4dxDDEsK6vn+AKfe1gW/HyGWXdNjwFH//0hNlE4W
cyWySjPzjsZSzaLplTw+jDWVu073aVY/Hj0h1hs8zdPU/VUTDbxQUpe4ZfaBq/ASJnNV7I6ypKa1
YjKLXnB2hFUGqVeX8bzxeYqLjgcOYILStNQUVej2dgoalbb2IPcBN34HGgh+buDEZE5nyTDNkSa4
PcU4LPT8IYmjbuKOc8YmG+GtEPzlCwZgogKPvUs61giXIrIiUTYNjEItyfBAjxhTT8SeIsKRqW97
01nbxQmii44uZeXpZF0txsCRZGKwJWY3URRTjGBkaIZhPIUFVKpRLMXNxyeKMceU2OwmNJn/OQHD
EjbNyRBCojRu09l9o/lJ/4ia46SF+s+qQ4NeIGI+feezAxmxMECER2nZuEM9IflBSl/w5LY5v5tD
k52qF+AGDShfz5ivHnBF61DeQ17kt47FvnPRDA6FmPvpGU+heo1urkcIN+G3VdbL6UUPobQPBVVS
Yq0q/QglAb0fAFPM+tyc8qnfoJXWOOzV42R8YVDQSc98XlluNjktME515Oix+DTI3g1mLIWtscS9
/OewSMc6DScUlsZlB4ECzHuZCq5ECATGGSR1sANxWIH5P07a7XhfhCLCuoQ8hKBFGYEsckSn/b5v
f+7nuinySe0OerwGrSybiDvgW0CfPsoHLsSAhreupSIQ01MXYlmAoFmkpBbG51Bo4nfeEdOV2VCb
gDez6vxio8hTi4lH6RvUxD1Bh8YHLeJ4kyqf+CMvScbwkoYiNq4w8tsjE9x9r9v4Nt/WA2TfhY+a
NnV2EBCqMGjxq0KmFQkvtez0I6NFQ5gVUltjA31Ttvt5iJvexB+8iiycITvusqonxlUTTxvd9nOg
mrjE7ngXsWm5fpzSUf7EKv7m5dfmFOeUr+XaVjBE3VvmEASK3IqTMksFanzX4XQON/sfOVEg5PoX
dbc+S0GKRhztHIR2YWkF0o3/+AeV2Jqi60VnytMZC4rM7+v7G7xNDt1x7eB3eY9Iw1SjG6qBstcO
jTNyVk/QohCB0Aeel5AxYIXfXK2k41BsfPQWRNOtzcUBf4l3n8iC4zGfebRc05XltPKAHuyrKTz3
+0T31Ku4bY4ePnmK3vFj8WHcGBBmReD5dSuuE8sZA4pc1h2/kM768smqZaws7/nsGDIJhVdJfV59
manMQeB86h+y72xedld/ii/mAI05TYz5JSnl4e05+6KHB2xmU6fhQPG58C9kgmMy1xLo24OTyMVO
p57zhu5QU6ERcS3QHc/rrVq/XJJmVXntC9pCEKtV0Ue1A3OI5b929v7r6TxwHtvoEPPVgDT3sSdH
rFS9HrM+BAjtntr7C0FTs5f4FBTO9rBLnYfGpH1wf+dJtuFAa9GvAJD//l8/PkXxhoqxWbtM3mR3
j7t86uv7IIsw9+MaxuZw9OF0h7gs3aXZgy/dXMc6rFRy0wQcZwN0krMUrHx/UFY3eiK01bXuDC7s
qoZIJ3GDfdZ/8a28L7K0VYIth5zZ/Vy+QONKnju/hDVvanyXHI6a3odpdAQ/ZmY5mbna8bLC8uPa
4kiPWWEAEN1tXoVJeYy0XpggqYxlbRamWXuJPBMxU6OaAIREtQKkAuQ3YUiT9vK5v3JGvLs8VSDv
cEgIGORvXg3v6+jPahpomV0Vgegyq0VsMvCdV54OPY+52FVQ2vJpr4oxON6phduWuZb++ISIsmXL
BS8OgJWuL61i0Dr2bAyglkF/tx6UorumQUzIJMBZ2xjlXg8ADA7RSucrzcZWJuE1Aam/jXcHAyfW
frypcQHSBcMCiqY6MqFlKpuliQ7oE3lIyCih+tRIRAp37JlH/mgz7k3ppem7qC2FNVpxq6WURReE
+wuiBrCeiyr7DzTTVEc2KhDiyD2TEBLoIH0jD4ZuvcMkT3jcRwFkhvCRwjtwbg1IIn54rFqG4z7R
d/+uKBLrvbTXEsLZDZ+gMfdAed/Y3cYjKwmgTAVkG629pB0PyzX37rNruBukkqq7F6VI+HijELl6
7e6HfkwdgEPXAC7Yv2YmRbSrlxQR/KjuaTAQyvi+3YL8vYiVuB3nv93tE8oscCgEFOQXvBkIP9QT
7mnDF0qaDixte+ASEiRul0S20e7K4WKdFugArQHZU+Y1hH6r48GcILi7mJDAnPDEwnKfLjEsGS2B
VKMcV1pvO+Hv7ltXUghnHgj1QR8tLE2/5RDPANXXJI6oeqndXmNrdd3RFxKibFOtKLbRK7YglOmO
K/zW4ol/31cQM1RwEY6RJ+wqlON4E0p7W2BGzgXbdcdAsQPTbTIOJe3WeHSFM1wHsmcE9KeC7YhA
g7jzWRT4cR0g28h7l6Oej2Ozi3arI2RMUFt8er7a8j/Un3f3nuMJv4J7lRDLPrqi48oEyQ2rHDku
5qnYTqCud2hvn/zRNHxIJsnLklQX8QqqDGC0BcZWqvzsnW15s8Ass6ypYNuuB/0sx/bIgWUUqtCz
7Qv5mOBgB3f8KaYb2A+5n8bEIo9gz/kS1vff3NlcrmBGXftRc0ycPnb/PIREULoVPHyneCNAo7G1
I1k7F6htUIRfQC8ZYYa8C0hS5N3PASqcTgAvz+tU71a5Hu3eRSagz3tqfRPG5kTLCuuDGwr1ISFW
3yodCOVAJRGYtksow1ottk9GIWknD3PntpminhSfyY3yQtwKrDr8YAQ6rYB46MvAlBbcd5X89cdI
xkpPjTvQxY4wSAs4p7rrvu4Sy3gWCpHLLiaFOUsqeJ9U2UpXqU7/+EjRdNlQTyjDIlCpLwNNVtBY
J0pgVeFHqMlaFk8ZYToLCj1PwMieIl+awqHm6BhIbM0q0Qw5/7Qp38Rhe84I4F8fvR6koxIoimG6
qKwcwauh4uCUN4g2+u83KHQf7E4TuaGAdju9mQ7gAC363bMv+iiGf0qriKPklqlhLmE/H14mwRwt
dfK9uMRaBVWjmuKkLcpZrr0vgoYy2jnLxe1yV4YPB0YusoEsUwPuLVL1kLKQfmDnxZGrZ1rySeqP
lo982V6WMLz90O95hPWFL4Ss4QCC8c6MtXxh1YIjbG1xcY0UybWGntbG0gv9XEIKv4O44jeASRnK
Pd74/yt9r4cYFX5RSO0vt0/6eZigqHSbJc9uJ/n4r5bD4I4VFgwBlTo/+w6gT1DVStQ2+/sBtN/g
m+0nrWPOz+jUGCdi4GwLQ7i6JqGD3L8Te77u2jQGMylKDh/hAt5B77LMZqWouKaclYuZl7ogBUyA
AQD2d9lhkpzo17cfpvq8zVD+VmptIyfTpytSGT1sTEcBG+qLyFnBFj1QTYj/X/RtSUfnEMZwuAw5
L4Eu0FzHdk/gdhOKmWLl5hMmCEuxKNo1z8joinnAqI66gTFz3q4SXr6r+kTxr3WU+/J92huw++Zr
ThkDT1ZBVdUtgLVT7LF5dfzCQbcCPVMrvXeKePonb914jqBUh52ev0xHN0B8hOKGv7MBnv4VJVqF
/T1rkkdcnbIYDryZaFqOyKC2jN78EdqJKosxooL15ilaGf7vUqhgtjs5XyfOChJEkzc9At8SJhSI
6sz3EM8tXMdlVesDbJrO7GdWT/6Gb2NYy1NerAWK50l1ouRWgn5tb1CYw1hfUi38uBKOSjSCAk3X
hvuT9lCCTfpcMm6OZ4xNbLzEAR8RomZ9dgbbmEUsQsAs7xjB5Kt1u8IkhXjpWmQrxoZZCCWVVph7
KgCP+KG9bUll9MH1L6oZ77euhlBnrENckqgLje9swM7EBs2qTtV2k++PpvpBC9TCcmRcwSN23VHl
2tJAiXSI/l2/3VytrmHQSc0R64QcaNTX0nIDioHfEfssO0J3tXjlfAsipdY6tS62BYSG8Hu3g+9C
xUPpKboGiCuHEQV4PpzlpIMo4yXIyzWxXxx3+Bfwzmr4rfplSxp9Sl0TXAP3LmGl8y7CadqR/OCq
NbCksx/Avumx8l0iheFayW+OLBwMFeQnrUBuksc5JWY3ABAD3TkkYKwifAyMUne06+aXT16BVFoP
jjRcOLT6GVR891dZalEdt5RZLz6T0dMo6aHSa5Ft8MHQLX0C8ZlxLLYKtnGSmjAGoj8pfYzirZzo
ulIwRLLGuTng3T2jjgpTAfcgrwYJumFYJY7hRUq3NRDMAKVoH7WYHSV9QK2uVrTwLanLwcBWextH
4Ycj/cjCmUnMwgnI1L2LJpHj+LA4wKA1LEAyHPsv5tTxt1TFfNk5AwQLjNf4iDSCG64Z8uuDuaS4
BO4CtqDJ8TOA73j9nLZCKw8vH3z8tAxqiw9YGDkSgP+qNASK+QVXDhYBfMhvAhItAqqMyGJKu23u
gfU4QgHiHWYv4d5qgNuPCcu8Op/uq6poYjEMsdnspItGwX9G31AaSL/PV4LX17BZdUYjI2rzima7
MzqnjWvAJe2ZyOZIeBjj3Ao+uRZ0owRCKno7kDAnrwU/4jfHmS6mBr4EBekPCquKGWnMifNT/ocT
U/XPtmBhJSsj46acS0GZp7lrTj1qsMO+1HL9AoAZInacyGbQ8AHGbFPpvbPdWDOste+1tOSU0+TD
JoUACTxk0uR/a6DqUMiRzG003Q30Ki5C6c1AAjlNSJ1AYPbAeupsWR8s0IPD34aZ6jsrS8Y/iAiy
+B0PJjzucQO+S48uO3dhxwqfdd5KNvJQsE5SwZSyZJd9XjTdgZzN/D3Nc57lKbPF9rr2m20/6QHx
MynKTghCSCJ9cO5YRfHfUTmF5n2/ibPNktGjmOuIPj0OBVLLEJ0grJt+QdeU/ral9jUl7xpJSrsf
odZSWDza/ibKss/+zA5Wshblw6rRCcb/JbOQZequl88T2sapx8B+iunUdLX0DeVbj3sIkmmdq4dL
OtTKwcXxzr4Xxj5OWgudzI1Yf9vkIhRMCKerRZStHEMKY6AxjeYgylXi2J/xAbS+2rGgEqwBpEzv
X1RVwGpLrlWXJf+We2H17tbiOX5v5zoKuT3IPSASdFuTCpnw5FHLZWHhoDMLt3R6yLFQ4HNBDD7+
7LWBGsN+Q2XTnED2oevTib7XRVu2SWj2cCd19oSHkNNIyyNe1LRAPxfeYdYZa5Fih9g2uLP0jAYX
s5Dyi4raXBAGzNFaVo9h8nscy+r0XOsBwJFGkNab6dWr/A7ubm6no9zy2IRH2YJnPa7jJrdlyuwp
qfZr9S/DIoYz0UCyF6vj3sdg3YjdDrisoTqRAISDWhWeleX7TgIeYv2shquxZ6FchsINVpu7o3PU
xQan7j5AdhGZPeg6pnO9wUxit2ziKAUGo67njVWRmLkSQoehWTEXpYHNpplW2B+QwlAd0muZA6Ff
vaUZNrO/mHn0u6kvP4dgxrFu3jATLP/G8kDbevMhj0jSvLdhZBNRhdCzROssx9f0AGPMRDMuyJNg
6LbXVrEU2dChO8lq9fCdmBMeBXq9KTkz2gWkbtmLLK6Mf+T1d4tIzVPv1xbYHTLjvT2ufaHDu7h9
nkDLxncAuCrst0paerUDL/mgiMcoW3hW2rbJnpMZUwtS3ikqJ/auWkfi8rvVLVrcizKBooRT4O97
QnV7FL/AZ9+im+4qWhGi4AQG7GR2M3Oyw/hrc6qQdfsrh0BueQTJffv0KA5vgSI+xwhSv5Qj+fFA
grggfEvezefZ34RSYprxpKCKa6YjtGTwaYu4e47B3m5sSyXhD8S8zJMPvILm2cOTSj/iGMGl2kqu
BHSCPBngUsrD533MI0dDPDH72VXsIPkf0G78YqcHe3wE6x/gxSO4pcJ++ZxKPO/wJeWH7Z4LXyI/
ux5P31oPhCLjm0a2Ss1/EWQu9eRIhebh53zc3cdE2fbTqfrrqis6NOGf+gRcjgxnNLeREBt1MHxl
SEs06JFJKQsbpSEEQjjQCud99VBXXVhrLwbGPe7cIfSKzF9F3wsrNxcT7kipnEyKGYF4Q2GXABwY
FHs1S5HKXvEWjdDEYjxfQn0px7ueFiM7+OlqNAC5DWQ049n4I2AYbwsi9PfABkDDlaXXYAQEXsx3
TmW//DwZtFgnNVIIhzj7rDb2l69veRPCPlVErrsYWVnVmkOSuE7b05pzLsNfwU7Kfro28zbS3UnL
nLMHnbDMwM9SovrrTZ3mW2pNKugqAySXkAsg/lT/i2ZrcqtvEROXUxtHxczQBBVxwFSxa5RK6B4L
pZZryV1kJzqVPIM74ChuVdoQC6iMnf2DHcS/OZQqPdCbBs9HHL0tGyUaUgqlaTjf7n1/TCvIpVEl
/VHnChNFbiM4uQEwyyNJsttf5P3sX4Y2eWXnPvrOVbw06ftrmn7pWZDLgf8iFn3VNYlVHaqpX8Oq
Igb1t092u/dHguUQMyxuuLLnyrtFoXiP3Ms0Ze8B6YEL/xPyFrBai5pyXKOHjFXS3lBwcPWeW6tK
gYGS58J/XIvrHXV3m5RD+T02/jKJInxykZ+rD8f+qwtvyNl6C4xrGvESr8+dcjvWPx8uEMia2QQl
BB66d6LdkeGZARXQoI5gbycXlpIizCIQ0xHdpBC4V3WV2PreIJXrOyuCT6TGK4K8RbHL5y354yMI
U/567Gbd/tJoUpQV5vETyPpF+yS9QvxEPtXZh3dtJfldUXXL5E2ae8n/qUTodAK9UQSWXCcdx0jI
fzQbnea9FxprNnXaOU/1lnCM0aXICLe8AxFeOvFMflZ4EkiJaxWtflEbGufp1qK5uYAhZIw1/OAZ
e7AcqsewQ1uJJW+PIcqqp3hliWcyernBfT3Gg8ijTFnU4W7tNVdPdp1ph0B75pUR+idB5Ts4hIWJ
FrSROHAocrDUG33t0149xoK3dX7yGutu28dK/I5KxfbyJ3rnMS0DHjhcLUV/HP9sAmQeVp5JMauo
Bphn2KRwbp6hLrKMwk4of6UWXeyZyiJUOU1WE5nNrXzOY0Ubl/nkXCoto2rLZYEchStjpRAEuX6t
VfReGouQbRFbjo5qO5j9g5bWvT37F1TVG6NtrxTGDuHAV55VRL92uUlvbjZ5Q1XSzOSgUQhHT+Bf
e9tVE+L8cr3Ph39jiASPW1GxNBesJDRShowb8UTGr7AuO5vQAaBEddzmaV0VwXen+f+QND1m33UM
2fB9y/GHqVxog7x0WcMUiBqn0KQuI8dJ9sYAivkmORPzERBO9iyLK31kajYc47OHmzk3SPXWWkXR
Sgr+5RhycK6P4fLVH98x7yKGJVkimXPfeSfEU0HdpFiV3LFo5PPMTZt7XjCiPu3yyVLCefwpPOO+
B7GUIY22UAstV76XhOpbnTSObatI/C3IT8M44rDs9IUtayWfHwjcaUgochuh3/xXqyUnhHRv2tO6
mGYAKpdvAfZXp8+ev1BHlx0O2SDZSx+DLOITBnUuqZNM6JoPA9dkknT5v2/u3oQABQY9aUQWrugr
UzGgrJZqI0NB5SlWb0suq1rS1DjuMIF9sAvfZi6yeK2KGgGvMgVKJQ68L68t7XG6KQ99frWmqWdw
6/9nWUkxlHOuHEmh682QSfHUUn63itBGUwNxFmYyNRkV0jsFK9HLkrkZjklWXchkMqy1WAvNsl0W
/9EPANXkphYoh3b6hAfttaE8AGjMDGqIGWhrjGGL+RDRAxV48tozRcq0sVO3c+mjDzO+T8E3r1VU
gtBXKGa/WwIdQ4yu4ja7/Kj/DDK7vNoIyAtKiU4HhwHKN3eDlsiCU//rAjn/bFXD9oiaxVqyHeXX
Z29EllIURC6f3+A3e9e1Kqp/eOMwDTRN7YQKviwT7+03GsCSs64LzG0mi5tXhH+Xn0tdlsOTit+e
T1iMg4ZEXUK40qTso4s+XrGQHM6ECS+RcGGapxO+NnkfCj7bn6vBXQhMEcXd0wvUq9HL2JLVh2tH
Hm7KknAs12XlxZ8h1FiVCsiM2iM53dKLc6tJdNfa7oPA2FyuEcgRTWeZw2qE/7hCIBKfMourL6l9
6phLeorUWft97RYmoN7vGDRlnlO2A0LYZ3hhxkXWOu8xWtY4d0ZJlyqPM4bRJshcozLZlM4Im1S3
C65zFA+TTxtc7NEH1uTjsx4WnmR/1+8WpXJkHfP+EMAM0NkDrZK1+E0ygAk6RJEfD72mry8zy7Oz
GXo+4Gu7i2QB0X1TdX8YdEfcSWYt429y5ewOYtuTc5u4kxs/unVsAZqtE+th5ScY3yXkH0OlR8T8
wkjO1YYblHbXox1rM3VJnT68oAiyxURJ3MOzEWjaGVh4Mjbrxw+0/cmL/oJGNn2xmq04puFDd6BN
B6vttA4pdzmVo64r79ohVUCuZUWzPeESnLDlzhoZdad0rrRRIxmOvaS1CgqqYune6HIpDLYzUvN2
cGYIgxcFP2+/OcfiOu+nwxcrJZHXomDRqH2X2Vp3xMR1iYXYKuaJhEYjuYQFMfzCM127Vd3QXJOu
/zcxDiZp+TIk1YxRJiAGMgalRaThfdWdpTxBe55j892bqi8B44mxQ0ISAwUZfpAsdhECiW5Ou3XU
BLeZz7FP/oh9G50dzAr5y8qLzCGFntQilq/WfyrNuKLo5ZLW3z+n/Cu1ljYhawPOtnDIvAAk4XIv
3DY+th52G87sJ+YJ3r+GrlcsP/56VPrVfOr0ARlBqEfUWTj9KLk8vA+31bd+JqqrLbdWGHJHAzhS
ItGL1rSM0y+UvT2Hzia3Ozy7RLcZfK7AgGoksFaA1Y+nxKldYHyfVXtB53FZBQbtTOCx81K4bC8h
5gXbszn1z7XTN4UWwYNM/2QruYAY5FEZJvuYjelHsUTn15D8S0b5Kk8s/klAU096wi9Aei07/nRW
+xPuU/c2ykZ46YKJOKzIT9pr+VXcESyx58pEi3uZ+odZDIpKFb5e9p38SbMt1DJQcGdRclAH4+0Z
rcyN19IwXz2xgKeoY0HC59hpPXFEdB+xcpQFMq4klfH6CF2y9oCDrF91LF9Q8NccfAjEhWT4AhWl
4/l72lhJwkkspz5lmTcImEYpvVo3rWiI7q88fyeYt00St5S+w0+2XWmk48avkHOpvOnJZSiMlrIU
5TMnFFnwUVSiAqjVMlh5LWTDPy0OFlgkLn7tdjJZtWDo/8PvIen/+PxdD+b/NKmNGPDUp5awrHlH
gMP7fceMu9NcESLkR5d57UCS0I5SRar6m6MDs9n+EJdsvDnz/lhQuUcTcZhgcrpR5N4UVbnc/UQR
qzbaFf9TxHXXDFr6PweuM657Bd3f/xBhcemEqd2wAdMAE0GJbYarSO0xM+arEtYJSQABIxK7Blen
5BWtDQGzneyTmfBnpWibXqU/qAlMsvPyBlGuzxcFSw2BOsdbu/V8MDUizKRo7lDACk/u0hIF1UbT
sMyDgWZyJJKZnuuORMyYsxd0n0MwW9x49+pJzZ9taKLK+vf10Fp+kiuzD0J9hopMuV7nx8DH1CSe
Ren0I/tQrY7lqsiIjE84ix8QO0cIKvqoNuRJnyVct3JZCYlVOe0e0nLaMCsToyqV0xhWMM9qwdn1
G7VmnKh+TTiIoF7IGRP5sq25mtkU0/3BMfjpQ1Zovlseo3mMt4bbnRQ91GFTWNDLgljiHqgofuLl
Vx+CqB/ngTi2ifiI5rjRRaOg+DgQ5x1j2+WYhQ7+uF2hQ5bJeu0aBMN5KSejRELH3gGdQf9yYLHe
Y3n1oxP2HroeYf97P0iYXS094aJyl9niu8Y2GST5tR4ZBSzQFvInxIKTmjBYCpYgZDnLbk9GIGuK
nEaMw8ofmuiPLfZP5UuwNUTnx8hiwuG9UfZYTTuFszujmrSgOozDc0vBSFgED6Xzi2Fk2wzW285g
G4zmCQa/KIoEtuEadXpaL3PUB/22s42mWeyVCGKzFyNzjbRk2OkRkbf0rUDcOztc8kqin48Ng3wz
PvN6AlS1WXZYZV5hmuIJUia2WUBSB8dw7RGNAF9G7dkk9f9mO+jjbO7GF8lYj111xMY1WhKNEM4k
d2umw2aEqKvCv6CKqkhVruJJFiksfhoKi7Yg5vSYBevYBJb1XCvaWHHZGAEGC3HHhC/p9gSpKJ30
yUqdestOCWT5AwCd4EiMIURWCrCW9o1ceE1HkBCSoL8ydRGdBCU2C6f2oQxEyrAn/DJs7qf0a4bn
3JY7OgDlTYWjf4o74bGvK/CnVH0tbwu/AQAROXrouTCE6omqlk6sq8xBJYg6NIxTQKvHgQB8pQLE
q6OWQ0kTAjxDRH0P97gLXhbc+kHxkmR7Ju2LuveR9Eqc/zo8hu0wOJ8VaYn7h2Sg8EQlFQ3GDZfg
5MbZaUJqlmpYX20uW1viTvICLwElw91vjoKuJ7sErqmQGrIdufNhFGnfSfMNR3XmAvOiqN2WDz5p
EyprAcsypmCFiDOZyQQC0Ix2yfKwGgnMEdIKQxcb0rAbJeIF68fUAZLy2zORXJt0hvhDoPjb0G6x
zyCE63ba//FpSxyx6x7nrc7yBp+OxQhm7N3+QMOzZvh2sVtvgtJ+0DyKUKvhrIrI3K1cD/NYMUCZ
ItdSp87fMAfO5GaxA6KRY5lkMAxMVNTZjNpOOfYXXIHfGUPE+u6WKIXCWDasq7xhP+9NPI+dSaFp
9TCIbCQJzQAROZeRrDu1B0/H/gxFiKfVD0itv6yTvrUW81HHO/06E96cRagwLurouimsnO14tuCd
ymNuKY/Cfy+3ov9nwG0lNU6BQsuWKVbnDyMjmMGZJHnQIOOukMlBnLellmaY12FOUpirZD1xQNsg
gCAo344G/G42GjtpZlG0NGuuY6x8F0Jz3n4bdDZy3KH6/Cjz/x9yCxWDDtZ+y14/b3gfuGiGSYzB
pBJw2X/WMt0qwAUeTowRz+wz5atrMD99E4sweKra2u1LJcNG2kchPhb9/HRb5YL569d5+on6iNDN
8NoVq93xX9usb+pWPjpcRv4xjdRyXvdfZ7dNlMGTz98ickvhhK70IDpuWYCxXiuYftgCkfWPxY5F
7apWcjK6sz/FRRHiDyJEMhDxrsNGV2MUsoC0aWKSPuZmwK0UctOR1C/t0dEKARV+UeJ9ml6RUpQL
nKYILheS3Uoi1yjN5xqMlRBUY7Ew3Nm9dXtq4/XKxv2p6o3rNV9KdEOqrolLc9C+y2wxxgn4U5X0
kc61exSTCcDZ0GaAB18IDRXvLHK6j6bl4Su/xDx/+SLNaAaORumaFNIn3DkObIK3ia0bh2E2YT6F
ZLQfE7Bc9m4C+LiWL/HHpFpPScXLe6eu4GCVX8NekCT7mUVI8zG6fTmH475g/w3fWxrskhV0o+oc
ZqWwFijNcqvgsxSKhnjd9KKjP45EetItEorJJFfsNsFMR6lKo4dQmUMwnVgpB8Et4GhD8Px1dm+D
orxuxeepPmioz1Jm27iwF0B8EU1VwLGgc0vbuceOWQblTo8QAczPmoNhqJvEuhyrBbYnjK+LvyJh
32K5qx4Q6o7VADN7wN2vMc+lVc803QXTnmNbyfD0+ebrpe33QrBNzO6qC6UU83ZqdefR6hVjYH2J
+7dqr7edwS/4qdH4sw3D9pGmloyoJlkrMumQGdGH7dLzHms2Aqqry3KyvK4xm13+hQdMabuU+nNy
uLuxUJXUoKWe5L1/idI/EttVhkE+9RpjbsCXjcUqME+hLTNz+0VGkS5c3eI8Y+2mgmLXSEcA6lpY
AgUqpmIOon7h9q4D/z491ziUKhkdjPtm6yQSOUrZvRPWKiWiarYPeiHmasHm+tG19GKji30Bctuq
VTHWjPeE+uGDHz8AtG5XghDwKhxIBcEFVc43Y1OkPvufmZxruaNEZIkV/iLmVZBXxrLN9GvG43Lw
sxi5vWRUS1bhfSF6r2nKtvjHgc9b8t7qLTCXBnPJ+ZWD8WPU5I9lGg7X1Y2T75Evv+6OnnoN4Fda
Gi1yR69+0E/5U/9lTLW0c/hQ4Wcd2C00fLdlYP8ugNHd/BDywwdQU1IYT1OTT0gz5aH2++uHEibc
3gnmgXngcuVJS/zcR8vfcmNsKu9bcaxjHSmmNsmEUy1TaC1/CoMii12U13sg1a0lPAfarXUMm8sn
AW6q4FCIJR2jnd1W6wOUycrhpn655nyExAvak6LE9eBcVgGsQxUGUIc9e2SLEi8fSh2cjAGtRtFd
1zurvKa/jR5M2SB1hmQtEkUKHztpF9RIuJC2yj5+e7JmHgtUXmQg+1qlAcnUZpWZw9YlaC+f4bIj
OgQXz9PmDSrYcKK+CG5swxsaAURHEHCee7oU5Ux+RXgtCBJhd9jNSLwyr7G7bak7PX6k/cRZ2l+U
nZ71yN502cwR8DR7tRqP+Kx5FXsxsJdZyF+geZQ7J/fWoNzOisDroQi4IGOofX2oYgmHeE4frFpi
t8+tC3a/6LosxUGxzOPHGmf/1vgFeOcYZHujh/B6G11NVRphhxRo8hdUoJRiKgtoXkQSbXQNfFHQ
CZ7QokUkmI90N/54kSO3sx++BWA59HkJwNnYY4yM3Grm3M351fRM8vHrwmdAU/mssxSL8r2SXVnh
ZBgI4Hjci1QvCZ3w1H40sUHVmjf00Sm8mZRbKmJRIzS4uDI/3jVWrJzq0iX6eI3ruCpaxMj7RjSY
umRyd6qjfjbgPZVgDAvoyZ+KWU662EUeUUTjKz4kwTq1fcnGIVurbk2h8OBATd8afIQLGAhX+JU0
1VG9vrGBv+9ftUxuv+/Rp6qP9ueB0LEilIGh/y3t3VAznOPafIDx36LrVwTy+k8ms4ONt0jK6zJu
sAoNwvC8HwHk0bma7ryTctGD0cZ8CoKE/lPZzkGhBmotUO4BrlK/wJDoJB73g7DwrN7AsSYz26Ce
kJNoJhBl2WNYsqfy2NYXawUYsrTidEHjKR+u+Hg/se8WjCtS3MqgIbfPHRgcZPPxAx0va5O24oBC
bsCemIkQlkHUwnO/nv3BNEGAsY5WX3/LCwaxs2mbpWN5z6IjxU07K2K/0TIjB7Xl6fd8s/fT6XiG
rGss4Y3N+vWSoirjX9x0yM0VFuv0nTi+mxZpYGFuikaaMH3CYKlDyEMLmmviKvhHCSS/5JtpOnyF
/Pka7RBIRn2Q96Kxw/HQG+dlq+vVN9P+oqV+3/wSaU43fxWSok0F0sZheUyxc/o1ccePkj1Bk6Kf
IfR1nt5plSn46GL28AfqXgBWfLVyjAmJCX4139E/VfxBLj0Nny+N8QtYajafEJEjzWBy6TV3mezY
OuNMeC635xNP/lRCYZAe2fAMQMKHM5oYQB7t8HTyuvkckGD9huVMcTEjd6/4g1TpuLjwBrSVYIHj
saUuDD5xPzDHAJa45njAM8BuGpSWdPi+DZ2ZVtCQtKHMPyrjBQMuTn0YxPPEQOca5mvVjcDQif85
P+AjdOPrzLgCA7XfIvEKbMMDol7btivdjMeQZwI6G0H33YYvLEYy0NtvKUQswOKG1yjQR3IdNEYj
+lIuIudOJuWE6cWcZu4AVkko6SDH+GW7uCphQ4DADcFFxPz4TManK3VOXZPqQjFhSK/u5qMtwkeG
SlYrxY+4i5fOdIcPCvmLXY46tKhoYYGZjQLguq0edNL1ncT/p9qwepwuK+4ybv+2lAZMW1ERk85a
1mvxUydSgaV/Od7Kv0vu6TmY5IFSrcRTpqIHxSxOznOekFgvkDNjLt+aOpvBCd8hIE6VIURwt8bX
H8ik9zoXUNAOEWquvc0VZCGk3Efr/YzOKT0jsHUloKZfuO4+Ed11o/obd3B1cIj8wyxDWc+IFFlG
Xb5dNVf/BbEZr++Ga5hNrRfqxF6lw2VF9SKjceklu0evde8ju+yEIdXtLZR1nFQ9WuIF6pUCYrUX
P3Av2SaA8Nv5dpqfG+umuxeY3Sss0+kqWonU76CERsmGdGZCHbcsGf3MrCLu6yljYY3y1Dh+bftZ
5Ot3yLnilvAbmcR6ebjNyO1mlwul89nftaWNcVoTyXAFILTgc9C7aeShYLbe+ThcL8OFQOao+UMD
ugzZWpraAAX1co5Cra1AmfPUfLXfvY1sytc7zPrNxWsP+w+znMoyswPHndLFh1O2VpDnjGscx4aD
VKkFDBdDaE8tPxf5BVcL3/Bvl0VzelwIew+wS8ryoedy4oTIHClU+uF81R5nFVXFMZy/NANxG+Vz
/3PqBid5HNnHG9pkpO9nnEXhzZhPPT2STLLS8a5ZY3ibgHyxJBcaCbOhY5DnsPH0/4u9/I6PXAu8
F+tfRYYem31dvI6gQKqyQeY3piwqiPXFTAVNtqEkQ16NGPUv26eoWVJ8Zj/GaC70P5GgPdLRL3KQ
vaJZIx4CwZMWMpwIy+pmsoPXf8vzsZeoQO5hswpPsvxoiXHPz18CKc5Fki/ZPrM/P/TkJ41F/5b7
soSJ3vJpoq6nvvpHjVO3gZ/BtunYUaw4aOqtbF3xx9j4PrPMMiiVGfllqBMZKwMuij91edGmQBH7
tr67CXpvo1i2CTeWZ/bWKmpLbjI7bN8lcurqFvVvMfsNE9Be86Xcm/Is5+DscofLpVX7FPUhNA1b
HelOfMkWFkqZ/6ggmmUdx/XncP/ulv8L9yhr1gH4QFQIJMnWFBqx4XRKRXsTCBvBof11ouroeJzK
FrelpsYMsmbiBA6yi6inkz/F0rNcqZ+vziVg1MynM4DNymTvKR1ad4GEypbYEHo++FL4VFMbXXD5
xiX/AG6/oTiqmqd4G758Xls32nKyuMC6k8wL9j/7qZQOUqc961TFCZqL5W0AYfVpl+acj2QC8+xi
eeHyPGq/mL0x8Jk9hx0GyDJsGyg/ZYn578nwqbfzpcuA/KA9PJkFJmjox+IPurZKdZCGBELFUxlR
cFqr6RIIp1Vxw4iLaywN5uYcca5KJ7TNphiYepVP/PvL9YSJ6kkZbbjHUhBpd6r7eSDtdXOqAwOC
MgaUP8uykdIsGf0xltxMYNj5+b8iJY8R7e/mGaeJrpzyjnaShXgJ1GIkTzB/6McDHrr4dttV3jvW
yqpLPNzXFc/Ng8sjM05LiNfaBA8cxUOewc29zMC0DF8Npni5uMnxyMv10buhGVkLB42ov89RNA+4
hn431daMRgZkxOFGd8Xnqw5HvQCEymFfZLN5Ru5G42rtRhWzHr+26MV68ix/93u5wDz17rbrDyN/
5ElSkK091XXs8RJ7C5s743/u/3pYFese4hCDlXqkl/VsPEsYsAZW9hIW5WbE5OXzU2/w5n9GqF8w
lD5xeCPljjiMskhbIqrtW7Mrk4N2rgtvizsZ+f5Uj//o2n6GXdQbhYcRYHxo3HWuljK/QnSj1tBj
6dEZJTZqt45aznm8PIgzbF5ITrA9rOupZAVYigvOLVRlM7ePoeQTbR5vGrsj4DtqsgRe9+rCl7JP
N2Au/PDFBkwck3Tx4p7l0nKfy3edp2dhBoNSPIn3qDXb9yek9mfFTaGFL0rz7uXoqO3noN38OkYh
vP8I/ZLxxICSh3mE66t/2tme+TRkJVX7Xnw0XlSdBjR2q2Zw9saLSa3BKVwrcjZDf1rHpTJOB1qn
VF/JRsxZhYORhBu93Tc9yy3acKAUXWBmBTeRO0i1wGF7HVJ7C6uaPI0ClFEtnZ7WfNn/DW2TNzon
LATWeJT9gVECHmFiUAzJT3/rBdpHPrSt1YbAqQZOY2PuUxOIDR2s5pj7lOWSX/4fsfFx4ZTT5OYJ
0VYaXvdDRQn2IZvGz8emQGb6ufTrXQmcLER75qZLcGv9emZ6qlgtEhNRDNlDD9U6SLoqpgtua8Vo
sRWwlTmigO+rJNFbs2JXER/EpSrHKv2tXBsKV9Idjl8Kvzwf8MoVz1SPLKU+iHs0sp1Ol7LPUfiQ
4JKw4xvfi54gkXyAW2jqAlsghotyDhUYBzDg0GJrT0v5/RCigKHUk5tHSV538DOJvhh0se+9/J7v
IwHKjU0XnDcVlNco0NQP4y/VnDOBbIYbwB7sLSRIsoBUjvCNN5GAkJyZUrsiPIUHhriWMvyIONzQ
VSsq87DPG1fx1W9RkSEdcZsnWBKMnnv6W1j3kUJ6iopNhZ6ipdkbwXe7ErwdeMzs+rdLkVHASoFL
F5yCpQ5U8jmDD2yp0kzBqVDek/Ngkmhd90XtQVtnU4XJnpSBTlEaoBWiR0LcQBdMVYR1/ppYiT0P
NPhn5dzlZBI1cqNdltxlfFkAnxYRaX3Uy1Wk8EZ/TZP5hhSMfhJr0ALwy9MWzkGQGdm7jNoYYCto
jn53eL9/b84JCWyBiw8YL42JFbIvpaiIRNiBw0NQfV/+mXcmINYazbyBsF3Y57/8LXbERaA42nBJ
8ehz6W1ZpQKOsGQS4SrzB0/O/quhvB6PHih7ZpKGqYj9ZdjRcUg92SEbi+cAg0PHMhQA0FKJ3ZMM
fRM3KxYez7iqQSftmm2SES4AYToY5uuHz9OfH+AIsmNMLchAMOI1gwUXLwDZgMmXaD11uSROOtw+
UIeDmFMlesZ9AYSPz/rDGaPrnBuZy6xRmyPWi2Hw1x8l4WWyDinjY9XO28pwqA12v9sKOB6t9Qdo
mhJtGHaVn6QLFNOyxKitPyAUCil/bQfi3/8kGbL+UI1H2V+UunoEL4Y5/zny4jCAn9d0JleLSvhc
YpKRK+2Qsc5S/ZfumHC/f6l3smFh7esQSkdL+sqJPJ5VwqWLqhrbqlBjS3AgwNewqsnvFd7IQdHZ
xLVJRSt5lMwN1EF7al33PvvQXYLsjFIRQvEocfG9f96pK75BUWwaPsktLLaHIT6FILIp2lm4ax0g
7+Ibavi4mrU7My/xcjnEgyIRVkdhLqEKCiN49040gvEZtCSlg+36QfpFSCySBs6HuDHaIyAw/r5L
eXB78b/sVNaQXTT+3dzTuR3q/mnJB8NcylyTFcagx5TeRByPDpA5+NupXPfBzC20BqidOpfsrBL+
d/BUhGneV6XY9AGfSwiUOMWq4XbOuavjzwIig/2KqtbfypUAHhry8mZfo3Ex3WTPcvUIuRRjyV6Z
lwy3zI/A3Kj13ICBJPoIoGMr7EUpF+xJrqwyDeIVMMP3TcoE+qHjkAXysIDuUGqwuAcBBe/p4DfJ
Cp/9tEjJsXwr8N9RxsA3wE/825BNed3STce+3sR2/jUNzgIJZI+U1FGlXdhtjkM1d0drMU7m2u41
Rz9XCc0l8NJ5bOAApreJiH+ig4TG83N5d8287s/NOqKiff+9qkwy+cag/1WXGs16yQ1UtL5CJVtw
pLK3SQE+qxD4NBFu3ZCAN/6VvePLo+tz8wLiO0wPY+wP+kkvR5v8r3HF2gucUATJhTufryOuDrDF
dH8ffUyVwkgJLf8jehY66lOlaZkPDOkTCHYnf5vwRQT8PjTpDJSQ7WRWtwlkiEeltBPQpqk+XxkQ
ZbclLuFy3DSSPRFca8HDDbh0qcJxF4rCY5JHsbJtDFdJ8SW8umaYHLPDLTqVVAdWuClTn9dmAwXI
xpQtum0fgj9n8AwxAcK2VhG1x+ihYV64LLLLYKv3kJOru/TdVnGjWtdKkRPRyArNKGceVSzCXxbA
sXjHp8yX0PpaKjCJ3lUiyXF2dDx3UhXUxY04zPm0FkPUHPfCK/KMnQunBSf+kQLE2x1nzvgzePoU
FggLH1YxusHIJQQsMSux0w7s4ONsLA3krhro+x/zsS47I1xcvwgim8qLDXON6PahJh0ApPtnKmrD
KN5zDuPO5WeN+YHLe1gLkgRIhEs91dboEFKK93Dsm8U2fW6XS5135m55XFZXyrnlAo+VMtu8hlxh
z0ZUOmz2nFGNVrfEKA0SqoWzON2B26YHc+xj2rh7+AVF5yC7tm6A3V2EZQwLELpsBbhfLYMamy5A
gtvtWpqd8hMynsSEBUon7hRqFQeXabfFkluC9RDgNuqigK4vgPBk1kZEK9d45b5xrb1Ei8MKObMp
0xEZCtFa9e3jpOWiKOekywo2vHYr83X22sGDbs72aj+ywRYOuj6MVL5IosDpEYJld1U1nXmRN6fM
nLwIEAvOabsA6SvH0pfxGtcqvyuO1DOKykOjs4KJR14gcB+TBAakTLzAPAF2T+VGGPJx3GRLmKaR
zjxbw9Tz31QOT08E7VZmRYkwCkvAstZ0Ihgn9+bcJip0hJz2abMgvMx8+JeTYMXl+Ql8S1jg1+LV
LM1q4KqiIribplJoZ8KNEXvPKz/55teKqPnuxlKCbmBctUWGxE/xnKiMUmW1qhNJppvwmeVDay7+
dSquDFzgLdxI9XOr/NLLVWiGVo2qtyILoVS+js7M8nkMu31lQT3i7OyBc7ydt8K8bA1rdntBXoB1
fkXaX6UdWlT8GSx8vsjt8/xm3X0AChC9vKk6MBZWzRRvaR9IY4Xrw7gLAvbtzQmDzTa7it7N49Yy
DQE08mIi3qedHKRu7b4hv9Sc8RPijNxgigq31SetMYvJKz96uJ2ZFplTGDQJM3DzNrrDLPM6T+ww
1hPWZ3VY7VtPp18+rF4c7RDe8vC2m/Z5uuXCykqX2PI4DRP+Ck5xJxx1VLkgRidam5WuKqyc5AwO
7mnJqPw/S1SnrN8OgXKKKxy+seFuFBs/GcWmS6XCYHaHTkrw/SoxWTgmrl422B7+4C+2s0K08naD
MIT89FFvh3axJCxebZKSIKI0Ir3zmgF/006Ow4ihzjkh+lY6xOhJDQMW80H6fpQ+pI0/jINMn1Zw
zdeZMDwah8uKsGz964+PjZ435oe5u7XEnkhy4D5E5nZXkSlHlKLnFiUEKS5DBlfKSs34/PHx5hNQ
j783VgT89objPjx3+umy/hS3RcqlW/jhPblpbNDf/tgzdKLZL9yt4ipTzYQmbpfkWMhCWb0vOREb
t6NRLzrR/62RMUFr5Mtyofs2xH8dUSq2oVlSnUC9uDYeyx/ENDTYDrOCcoxSBIobj5e6AWGn8XfH
B10xvJaLG9oc8RAadXoF36fRxN+m1W2pvOx5IsN4j7KWtCQ+dh4KvNPd+froyOx50/0ZSBXdzV8C
Efam7d+s2fMKRbceyxhh5NmyR2aFtD+EM6ABLwoq+sAjwFu1SOgfwj6YAdfYN7dsoUYj8w65jP2v
HgGsg5e6D8koHeKPKZK31ed7lCzb2JK4YVVVLndJdZrq/FA5dAlrFbObVZz9DxigLfruIJwA2AYo
Pwfw7GXXjX4QJYQXkO2vEHJg7m0rkoHKkFLsi8PYPxU+8B8sgheZg75eYT1H5APXQQ8L1XUh44oo
PybI/tBEKTQ8s8hZVipDG9c2EZ14DC5UpLqPUrA/GsmLhwcpsdlC3SeEpDi2c72/IfVvwl7HL3J+
RwRZ+QeDd3XGZSRfVpZM0WfsYY1SjsW/+SJTCoi7LgGT84xSvUfveVrn7HdxkgwziZLMMS52F93j
BEabctxGG39Gz0Wyy1Ik4l1o9y4W6AyxyzgvRXLxZ6trmXkxCB3DnTgcOMCbsr6+kgO78BPlRUiQ
xtBkclR9gHvo1Ea0QANZyOpCVZ4uRJRXwtqEF9jmdoiLHe6d5yMvUiGtubnAXVtAj7ncx/YtE3Rr
7Ynyc2qPJMdJdTwzTzVJZkSY/5MD2wgT/wSAbjKlzziciznqUMOwHacWEAhQQwfhq7CfEUbIwhKB
SyMogFN+dpcN71+YzqSYI5Foq72Es0aCIOFHA8/CK4KHha3DV42v+hqUXeFHLSs7O32oG4LTCgBk
FXMJetbg5MQF1MxHXl0ptMuyUSyOOhHc0aCkuBAINU+/BEjwbC2it6cFvc0OEjiigfmQv53kMaqz
lky8UxQ+WlxhswqanLkmUa2KH61UAR9GUoefvPik69RdG+5h/LfuVfYWeH4n2kBPim+NFpWBtIvB
jbl6dB9OX28YgBuc7znVx3hARusWnLvgtQXmMLyR5qZNS2dJVFT7nOb8H5C5CTf3/XmpU+wt8raq
H6AYLOuZBVmK1CRhpOm8m/jY1YJyCZgXd6lHnyemJKewaCTwk0VdOPoOR5HG39jHuwgmw1GwaQoJ
xktWBGOxLxIxvOVdYICi0Wrx/YPdE67BsRDoA7JEUNx58BXOewu1RQs2I14muBa169fc+eaAI9YF
a10C2qkDBETMzTyxyI/ZHxaZQRFLr6BJRcuNDmdAmCgrY2OYc6Gf3gNsdbJ/aaa2YV17+JZIV9NJ
i7D+bl2rXxJngALcAocWQ9xEn3nCN8z1pvVUCX78c9ZB5dgjjQM3qGh7ND5M9Tckk4LWzVTMyCJe
pymVoU5EjgZYcjNwQkvBRZtnQ97ujiI95DtwGSImCiW2fCbeSTZGxC1pWRV992+B2U1bOBcLN/9E
NwqwFIoHL9xOYU47j6B3bYijZgrzXPQm1gEF82opN5e8yoUJ6gasuRVpQRF284yxJcNWTzgkP7b9
TLN3Ng5qYVuIJsoUMaFsXlyqma1lc5qq2KcjrS5xuiqBUxSNtk8pcuNhaZBvNc948Fc8Um3rBice
P/b/FAFPMXZzvv/auyIyKSHe0Hbr2NIu475xAnebVUtA93ldReUGZQD67UzHbZdwhLNlwEZvZ2jE
meL0WhgJuF7O6Dp4YX+qnGPVBDj3UfI76A3bhyr9BH3NejZPSlL20i0oA3fNbG8atDx0hVvoCqnA
i14VD5Gc9SgkNzAgX4zwKQ12Mjy8i0WKwZEDJ6NgH1fS0MJIpBWlyoaIpd5rrv/9vDopBDdyi4mL
hc9ymitk47IdmPnL3jQmoU/Lw5PIFUOrhxLBziA/+XQbuiJBD3obyXPFV6ltoh25wvcSymuou11U
6MGkvhvIVOOEFimQvwvfPlluDAaoO/2EbZQuiZ+2tTOOgKnmHJiVrZp6CQuZq6SMWwQD8mhBAxKQ
xmcwp92cP2l0mo8tPgs7q4GSXGwS98yeU+Lps/4iaLlAMgGkREwOW+yxCmmut8kuHe6xHhCwzbGW
/UBXFSnv6eplA5U0StzWUzgxI9FNz0l/4CRt3JrP1FjnSpaM6m3ry7h1cmwVghdR+3J9g3nozm7n
bktTKBoznM7Q7WVQgjt31nIVi2f0zEkeAIDwxTgA6Vu86eyhCHpSRJI13A9/uU/qjfbDq0kWDu+u
UblzCyZG2yxCZ4Uqs0kznGkQCgvTWr/ZYPWEepuGX+ybfVgPKIbb+ZRbF9ctjhE2SOh8tdojTiJ5
ZJ1zPCRmlOdyN0fmQMRHzKwSokqTEyfsvmwveocRnNyxPPFmRmHslCrgcHO4zIAtI7My2s1LWVgn
blYoFHR8MP9mntM1DQ4pMFAxaRW8vEYvg1IU8xfX+pzxL3YjXLWePmb0/FdhdpWqf8JzvZ/xkktH
XaVw1/zjVcz2uVfVu3VXQcVTKD3lopcowRo9raYdzh0+cnxkPlllgsn8F+nuiYRWHzMe8JIrOnhN
qfxOyoa2hzZYaxv75Ncwzeb+ceB7incLUnfAShySLtI4e28RfsLXZU2BcRVdl0fAfWejMDlIB3Lp
m8WoEAfvEPd7zoKBc3VH5VmW5Xu2LwCS7m2Kb+1/Hd+nyzG1P68+oVLk6tK4NfFO4dXWJnobnKCj
frR8weof7VN7OPyhgRcOV3yrvYg8voYvNLcAV1SSwU7tRXiD6MH6KGGubIg4p0VdcYuZFYv8UFGg
d+6RwetI1vc+Xg1wh6AvIg3awmSGhl1k22Qa3ySrzVSAyxIR9DhYm0bNvsd3k1vFJ1eqCXAxVPbm
NlXJ6NnVAUdlUIDfo9WtKL2Km72Z1oEM3N4ib4+vqhEzx9Nki06L0EIsHSjOAPTqp0k+rDwFJYjg
RrBE3dBUe7edDyukkqTSavq6uUikfjaERo5jiIdTq2vaqNo6J+8S5nigfGHq4Od8uBCKwy3Ziqe6
d3NIpjpBzyGqWyWI10zU/gvAbVTmdhkvU220pdT3JCD9bHddTlKiTWq9qJJBJc4Bc9F+V/Jx8xKD
l/jPx196HvfS2395y8s+fJFMhaBrZS9GB+9LgVB7Dk+b8PCiY8mHIB8RgbFW6ooj3TdOIcoawyJs
NFJFqs8RxBBherpBJzlEflASint9urC4ooFRe006ftkx5cajNZPpMiUaJ5LLk1tNwfdveC7+/py5
2iLnaDlOkRZqRZokB0wLPowcgGu4DCzArudZlkY/XMOxTqa0x9tP1krnfGepnoMzoAXFMntkO7FV
zypxF6hycTt/Xn1y9cmELsoqk4FNmpElWSxagjtJa5gsyabwxXiLNlYzhIh0w8bmLvunroGaPFj3
H+lOA7SFY5otyhCKVRA2KaupRoiIwOMFabRr8QSRtedmOhGqfLtrtUDR+rBkuz8BRhLVbRntD1A7
AkFtjlzTbGTrDFGaH2ZLKh1iCn87NKpTpQzmq22n6UuwqFNhNH3BQbFV8bJvaEJb81R3UUfAKVbv
WZUnwn0wVEaHjVu3ZqoVBMRJg1fiS6Y/ewRnMILr1Qse+cXv62SvL/AkHY5fYJ9hpYZSXORKFmHI
WeQaTGIiHdOhz15cuTdybxUHGDz/ZiSDs9Owtq/pz3BmEY/cCZa7y0CRd3rxdgdzq4bNAOBpF8pL
7ULuR9nubHYHpdYn68zW1AaJVJpdH6YaRlPjyiIhzTkoLZrWp0Y/FUFEodYD0Sg2+wntsTHGavFl
3R8ICH6OL7YEkd7DuBhZBSlfXO74DBEfK/4OZK8XSzBj6JaSyLEcxrCRRNx2YU54QqnfbYn3xCNq
WUtWm3QB6LH1NHRDcj6j5yrnTgAnDq4jVWAoBiC7zIKRn/8WmzrhIk7QIkIdBDz0+8NxCSMNWW+d
/WNDDm4OEUrrVUAjzy6+ie7LHgMsKPUlLT+Nx59sB81RjIMn6Dl44wPBJb150R/hHthDAMs9Fg+c
sQHUnS0HPsH2pALPSrxFcqR88rqZksy7MavA3oHTUh+shv4roqIMSBgRK9AAhRdLmnIi82c6nFP8
hIUj4IAHZKJC+unYE2EWPNCn3DCS8gBCJ/2WC6I+MdVh8ISsZhE7zvQBhyulT4p7msfuR/WI1mAw
dOcs/QiTtn7XcpY/yQiZJ8H0yIvlcXtM4KzdwGIts4clySuzK218YRibd+6TreKc5rwh8Cqs2NJq
S4kY/sTOBFDG5a+C00ngSl8OR45lA8jcINRLyRgdTGFBLd0N8PMqn6qPNgPUeIs8E7QTNyK3EjgR
sVBdUhJgx3BCyN9JuXzFQfv35eL1Z29FNU+CsrfIRuQWhUvAS3r6Nu2dfgAoQeCqcNJTPgLI62rV
Sy97fwrTarf9NRhWS5NLk9YRqxSccTGZnNMXgkkJi8YT6iANfKSDN+hZsL4lAwUnYf4iOg3TSA9S
ALhTO44tIxMlebUZulN6//Pm8ydsNrfcbeT7fFK5efIknjj/2BRm/EN+yK+XTgM3GsNPYSZJGKxp
8T9jYc2e1y6arQgTGaHbMHy6GGIUNfP7Z9XurTcB0rzztrz0btCwBvkKkxS612bb5LIvTyNLAf72
mRwVaXpF6wwtfm3hoi56UOcShFJ2tTKhVWtjiS8G4gV1til/mSw1qhenq65UWVEMJVIHr4CBZw1/
Pd5PsFf61j4KH/7pjfVG49FIXdBaSlPwb5dtMWphCZXreQQkUMnvl1dSe1r9j7RlAQV/+1KwPMXX
h0tqoci8g2aWRW0UGZp1WZAZu+wVGSc82Ga+bQctTJLUwSdDemlsZOmyE8Sn7p9fo/dgJP/9V+pZ
hMBJ16H2+PGv8FUf8tYRBKZHjU/rvq5aAlXcZaOjND9YmhEBe3vx7G9b5k0+9xDZqZ/suNAlwIZm
3EoTWDA0hY3HeY328SWuqXSL2R5dCXgu3J9yBxbFNxFYWSsUXUrJ3jb3a4hqSxo9h/xEIn1fA2DM
Uc0AujWGdtHEJohp/U6A2ShlMEJU2Oo0FiTUAbOrsv+bq0WF4RsSk32opNdiOW7zBwbq7/sIbDgD
U4bbJgkFh6YpR1Ot9/lwbnwawTI7J8I3KHttU1CvjYSkihWdRbIsKycc2XDXYfBaCWaVK9CqpCPF
l0nVfaLwU3v90wA6wUcadgjYEsyHhvZ26XstbA+1jluMoXR3hY+Ufjzqu/V5rc+resGwIUv2UfGZ
2ScogDq1EViEuDv8Mxw6hcWUwt6RyxfSWuibKaJRNZlpoRwtFhdcE8w609xfeaTcEWnmn8juypcs
AqEdvYG+ukliZ73H0WJLov9HbQ9j/iHEsUGVu5+V1wya+HOzlxqZmEB/JFDhrAtfFD1fh87hXuVU
tUSKLH90A0x7gha/rEzq3wKb88vUU6/gJDO6NxEaQTVT2JGuJLRPE9X9P1ul2sMqci1nGVBueLjh
AlwpkcFrc0UftcewcwmWZCq6cXCxrHtUVXL3pphjmd4B/dpYziZFDr0YI/WVvUhi9i/7YolidU2L
/JGEgXyKwFuKuMuA9E+or03TvQ9ThIUPOH22Dakh+3Vl7HyYGPmEOJuuqR4FSC5Nj1BbnF28UnZP
7AbZpTwCZT//PZozU5MIoEVHTyUilPxYc5ZXJF5tTeBM668v8gBLLV1QCT3VeeqfTQCSjQLl4Ofk
neODBoJMYyzOaD0L72fudAr2cnJZnRuf+4CSBFStmGV9kCV3/0bg+fvlaSzfaelxCSBdgUBizY3Y
CRqF/rO97vf8MTBPn+pk8RzZhaMs2SZxOQVlSVPbTJ8Y1lpFS3xrHuVUlpq9bVnLG4W4jck4prQl
9jenwyFydS+64nlO+5ZYGp+EYd2selQuAX24MFOP1y1Yup7YYtyyNElcO3XKmfb6TPR42muPrd9v
FsLEX2eHufjfDjUAW5mFLJrJV8g+x5b8WO0bU76xmM2bfcm6lpGWUKF50xffV7WBoctbDAQav0+q
kWYZxK33RwYY8BvWbSv3kErNdi9cRyJfhUqinXxixh5vrmG/U8OAX4bappYfOdVdzLYlmfiN4IXG
N6XuyeL5TI8/IeAL1h6nFpmddic6QBDJxccvPWjnrYUBZDsqgZMm5EvUu9Lk1LLIO6Og5Q2qoFCe
6uK14fFwMXeftc8DuAYcnOiwn+2SG8G4ruzgn+3PYatYfKbdyoNiSR53V6wteTHHEstE20XWVbQM
MMOUnHxfVoiu9/LAVfYyorf6d5DbSlsKB3fM82MXH9wroFLaZu79Rph8hHEoKez2ll4aEojqFkjD
99HXPcxY/4Q3nanZI4fDj8PrQC//uEckt/RLbl/geauznwpVi2GBUSNMIrFERPVGkZEeMJruINt1
zmiGYk598ZxzkKXWP4heDHnAyNsOYsMOSVUk/ut2/L5afPGKnLFwR/U0iAmqLLr5hOt1qccSfE2n
g+OUjKKItWhPybItTpYaKsqdjAE5wg6SkIc6OgObqStPBRmcdAjI7poCwZaM3QokuGaCQyianoji
v9ANDeWwHWyHO+bF6En3j/QlLD7U32bsp4/NY8aGmBb6gptTFmXjK3CMwGCYkxyp+9EHg5jDDu5K
VVMQA/rF1WfZnO0yeBss2NTx9z6090TtbUwZp88pmmLl07Wm+9D9fKZwFmplqbmjvORuhnjiJAXj
4yVnrF2yJuiyT+ZYgMdklbaYUzLNIMcOBM/7p8tL0QjZ1JkVBt/LL8WDQgogprRS2mmIi4nThQmO
4duDS2HPWC6op+3/gYLg1H9inuEmA1UoYLyFHhjDNCUyvWeZRa1zQfM3fFWNQUDZuYv1O9unJFTU
tzYsuj/BJp+Gk8UgrjRvcFfbpsX2rGO/rcO2JuIIg42GfGwSiWG8EsOf+qt/5YjjHyb2AgYtNoaa
7YXsYhoi0KgfO/JRn5lRihjOqku81oNz7gLA9puiecigA8tRzlsnaotELOJzxKBDqRxwuRe4Ucm4
4ExLKhBpymJvrsaNspkCJ6mNCTRiowO9LOxKP28qztHRKneoj4G0cdQqoTYHrLkW2+ctnCQx4Qsf
loDeYySJq1M3b+MVNkU2D8mdDcTr+A7cH6Ts9BUmNYMTD4ymST7Mps8vI5lg5oXRTr8iuqmIbOlz
b0k33OvOhUjTT40giTBPb8rsxx2lkXqaznMakxeoHBkTQId5XnWdCqeWcBehPxiid7Rs874rOhsR
XHX3pVQ3PQ7CnRe4Ko6vFer7slwtoGuZqtE21Iw3es0XSbcx96wzmnsZQIApVAR8gq5A/nmn3Jy2
SsOuNY/oVo4vfOxbOzfxdzFv0zomz9sS/afmMjjVGALzfnuGNHHU3wdMOhJ07JYULFJOjORHJ1Mb
f31zHhIrbCDBaBeK0+cW58YCwwQP+4Z7Vo2TqiTE6JTX/rNUjtCF1EKpXc8QCRhSK6nh6UBjxR53
40GKNuPfZHobiSeQJS8SY0fjMwMDDNXlitv4XYfoKJfV+cnEE6zmfRjZvHyBf118Uk362cXdMyh8
6tAkII/RZHEtH+P+WJmxmoTUOQ579LrddtCsAWYZhK0pMz54Lp9qCDdghiF36P2PGd11/Ej/XTTd
Ve0+SEppcwfMNEocdYCVtL5byyl3MBebUsC+GG9vGFy9ppcx7Z48mLdmAgOgi5lLDa7dYFrr24eH
Vu/J8qzEW6iY89Fyeak4CwNE/rQz3cL3VSy55ubrfP5HHfj85wPBhx8yjRYjgE5pCVULilPek0o5
SP5ZAj5QXEWopELA2KVfhLUUZi/ih89KO6ThJGq6voAByEgd8xcIHjpKDdrwqL4Keo2icTznCIVG
CO+wgBbhWtst58UGd9W/5cLN5IXt/xgMsY2JdtRvggui8AR05dNoOvbOE5HXwUX+ZYizZTxUmJgY
/W/nXJvy00V9l5KM1SMhGM8ftQjfRauiQkOlcBW9k6OLPxfajDm7Rmw66Vh52/6ZIxbwa56ZHIgg
rloZgjHweoOM2PnukWzSATx3VowuOlMTJTVgrTQlK69s8md3dhqa+FY/XpM7PwpWmCGcgx5fPk3i
h6ozzVYJxyyu4xeSeoqs5jXhB+RKIEmlmgVorogKPkZjdJX0ie7ImfiERzgFFSe+xBXxyZZF8kE/
z4jmi8vuCzYhe5ZA3v0hrxoQzbohIezvjwJrwFcXOWTOvnfnZpXKGZTs2VYq4uwH/PpqEm41/A36
f+GCX+sIEzdkeqFA8G0WUGQZ8/lqJygb+lmnPilyw2HP9ZC6PqcW3GoR3iQiRVG5PE5oxHQ2JXVY
xgFAMG+APDu4omsW9x5FD0EAmYfU8InVQfL/lDCTfEsK1NPRnKl9r+CfEHJr+ue+y+/PmoLx8kfX
hXgMqrZlyXUqw3hE+4vGBo3mwZ1ifvBys/GxLmHAhTR/1ufgOb9vm2SaO3zXjhG/RfbiHkhiNE1I
2mXu4yiKfGdOwxW2DvjFHYXx4Ho7V7ZMh/jrAzCqXkfr7KOUfSTyui7qeJQ/v9qo6TJZ9hkjP3Jr
ufBIu8du6j8y/quxHIATxMF+tUsa1qFgW4T7lBbLzzixLMZDsuBZilZX2uwKG8a+kkoasv8zM+SM
v0HRiBIqe06Fsca4lj618v6YSz6LmIOqBHG4IQ9rQRky6rO/RQtYsWlb2yX89VroSdKUtoFUqDO0
btzIkOvH1oDezz2f0p4Czj0x/JD6DZ1Kp3S9I8v83RegY33QbGO+vwu2810LSip2I2rE70ZpjiAs
YgOPMfg/wWdVXZZscot2h36pAxHkqYye6fmSjaggzHsJaI1s1q4/HhHeTA4z6GOHpugUtpE0XRzI
0ENLQYiDrB5dRap4U7upgojcTYYCQTtkU3+Rh88/heGI4aseDSh5+SeORQhZ5OuneTH705YKgmkS
K7Wp+vWgD0dbrIqq787EAebpYGgpVvsvpeR0qnkjqoE+hRgynA5DyDF6T8uTusYXegNlyWuispvz
8OEqdTxjIqL0hpd4y/9utxWVcAx5ND8IXxCIGRJTO5LNrx4QnRcmOK/GUTtHrTudedzV3bAsiac0
dEOQHYvGm4Vzcs4Q0UIYh8uiJ38AbOYrYvJ2VQi3DezX+ZQGJu2tj5meBXiHyllLbdNJqIsDcfkn
DRETtpzS+SQNH6uT/EFHEo4ckBVIKSrC5ByEotYtYDeQUbh0KuRHPR+PWjiY9jHm80g59v3CSpAU
aTaqc5FYQCFpxZN2qWZK2Ihmk5zT6CY1FYQLjOgIdzx4qI+rthKO73k20/FNRQidUDi7kMG2cBOE
seLpslMzUAHceqqlgxz014aG9aVLi/WS55e/aQ0DsH5QNW8jCY49SzG9mjWKM7cI0HSn7x3jka3z
2VhdxZSgHBUgHTH+L25DaNPdSSqdDVUT0aLJRBWBsMGhB+vaUqjMV6eTNLZMZxOb22MW2ewuIHTt
mRvfDrSPs8gNECP3zkTcaaAnSKh3jfDkx9SKEsT4s19q8IdpVGWToM26UQdityzBBsQf+zbP3ysc
UMyEpADv1HiXtkmsuFEnf/EUcExqNaipdfGDjmkFTMKL3FuqQd4eV5s4Myy+67KmMAHXeRZnrDQw
PWwV6in95YwenX75UTcTieZTkOj60cfCgmJczTH3huh8dmXn4jZlX3L5zisNwm01UfkwBvBpdaNv
uG0jyK7pdPKTqLQfPkmM8eEcOuBLqff0W7YtUtQf3RyvTLWNuPYqwo9TybADzFdMlG1TZ9DvYL2g
ifBHthFVDPrY4RgF9dzzX1be1GDUIAu7PvDIj1KSKKIgsWH56mIkQE/DdmJnLivqGw/D3L5m6KXq
JPTHO80bMi8RueGQ0APqY82TdVn4SoZO/fZhOmzPh3Ohsm57v9hk/zrZyDaYnYvRTffPds5yGAaV
efqSEFkdyRTCiUUZkgTeglepc/qp5gH1OUpxry2lfkn1/cbl/QVfMYj71wVLbcCDG7xl+WqPTZWA
5+s7jk8RCAykGcN+rEtwgEz2bKZA0nKM5rdPCf0osnuNc7w1pAO6DhKv5zKW8A5IMu57s9j40s0x
0/IeEPDPy3Ycqg/kvtyAYVmUD6RhBgin9jVityFOjcRvX5ZibbhTxeZSDooL+blgregpwetclqGd
wEnUwWajFjyUjoDIKeIhVxLG2LEocKIvfGDJutgOkgdcwnIdFxM0+LNJhgN4jTUWJWeymKEah81/
3OmIBYlSNOsy55p53fSYmWrx6EG2h6FhNpCz7THpS0Z/bqrj0SCOtC0l8IhiKRA94N87Kd3dLUxI
UqnGg6nDw1X7HXSbDfoA+Tx/XgfWYTGEDN0aGQvjSDMgCGfMpY5NohG+DUbUvSjtI9xC9ElnSHsQ
6HzfHUaHTUip8t6o5YK+AKRbyNsIws/Hl48bNQEH3ck/Ea7wLt/V71pESx7dpyZiH22EVj3kuG4o
rqbVub8EnxdXViV/sC8m9IoAV1YR+KlYdk3WK0Li5y7uJA1Eb9u2rMXiD+yBK9IOxVa7gQPq987O
/p1agn4o/9aoxC/GR06vFdsfnVXXSvqAMtu+4xAgFWd/777XIsWWt4EYiz2BnlmQYbDGmNd3xksB
DOFINcCc9CMqyMcEnyQ7E3H2cYV0fR77q8gs3fc9eTQ6JO69lKonqstlKxmnqNA2gK6FW9mUeuqt
zsW1nVeRnggLEtK0C268N6YYpGt833st4iSifEKL3gHQYUbSgJ9opUSoZw6y3QwvKOtBwj+G9RrH
3EOl/PIPyqLkCm+AFC+hYwLGDu1Xhuw4reViDIFEjmEzpH9Q/D6TRBQIDMVR0O9o27Mwsmk5s678
NgLcv4Gh5e1XN/G59KnfCowYDC9zWBKc/In2ixsCOOuxRmdtrmJNg8QM3/aB5jjquJYs+HBEBU7d
TgZyG/k2l5gUXwCqbQDJdZw0xSzMLGaLQwX6Jde7ynOV+LLrkkOx6qXb7xjGqs1TbkMjeZmYaXZS
7ld7+6ItQ00A3MFlr9m3dNqzIgY0tAPi27GzTLc7OEyAvqBQh9APl/5lHcGeq7qpnCAhAka2xfXn
On2AE1v+bcyoidkOIX2tVTjVNSVcSW28Lng2etiBdJhhewnHEG1mEV7rPLsrWZxHXw2EXHv+snsZ
CRSlZEbG+oiBtX/SLzx4udL0C9W7YMKPT9ekZYvxjM61qnrgb5EVW21mb81H3Eor3Dm8iX2PTW7L
KZunjUA5SBFqXE62IRQ+S5DXxFeRG4slGAXyhDDKK48IJ4r8Pizw0ELOoXCM/oA+AXsAFsqDduAR
ciQBeDL0OyYs8hS7hxY2pniGNUnmXu3BTKO1e7ahMnJoQRYc9cnZnM9iOS5vRKOx9rlY/n4h7xLk
E/sobTm4b/4BaDjsCz4Iz/DLZNNvmOwVjGGEaEez8qETHCIAtfLtUxj3lXNOL1nPmfI9XB7KtLHi
kR8GOa9JmY/gtROJieQKsOvj5r/qLDt781MxO9wxcguhcsRvl3nAL5m67Ro+MG7tSOkhTBa4HXqM
jZJKDVCfUhkTpwo5QcbAY/dFQ+H3xD3U6qULIG7lcEzeI3Pi5n0+VArnTvxCj4PVxqUaUwHuz/ba
AheoKbPlEA5EF4re///jRUt3d9JWS6ecxoYp5bRuxPaPFEKe4GhiEoJoNjPwLPe4C0zA0pE7TLof
TTkhgHbUxZXS47KqQ/NB2ot2OO7h2J53Icyb1JNZXN/mHnJA+FJah/emSYjpIqzhAZrFlHRp3sgN
0Kn7uUF0hZunpjylvPjwgrOKXG5fd2tM8MLNyOctCjVE+ozpPP+SrRUQ/r5OnUlhcuJWUpy5FUL+
wM2LKuxHKP4JZGySwwEYF+ETV2f9CV01SXKTNwk3xlyF35zRZQCqGWskG+A2ypPSCBxLIGSEQ17n
28DlrPqgo+FlotJlJf83peDSn8ie7EMiTWKEwJPByUOb3L1G7Huo4bVXByFK7/F54AjgE0kz8JOk
y8taT6Z+opcBJkZLz5KirkczgMsQzJ/9Rmhw0HzOXwXVzUgP7BzF4AqoElDgF+c9d96zWDe7exM3
Kd7VLkk9QdNYnDs1HYAkOFSwjnxPkBOFT94Vi8iQDnW7DmPN8uR92LGbdKYm5N70N7MBLNYcCIUc
Dkh97NiJ/AH/FVQXJAaOqMkMcbIyndbsLL06p6DSZmJvA+7tGX2m21eFivzI16b5shXYd2g/pQk0
V0/kCc8xj12yFIJmwv/2iOBr6w2H8IcZG8jmRF5qZt1TSRMJxxFl0ZBt/uV0Ws3h3RcTcY/j/2p6
dbKQyI1kUdN1Y9V5h4F7oiEQmZ/vJ1E8wV25LVxuOZTP+XXc8ChDV2ctdejKk6dWJRuW4rWlgz+z
r+TuYDhkH16SUhRa8nOWs01NNs+9lVE+/pX7fqtt3BRWcj+4Up+SlYzY1uPbw3N7rNtiCl47J8Ll
DHVYcRpQp230Kk0RQEbMYJ5UbUFXK1yN1af/Y8kaxV+rBXX0owCOkxpRK/ELwLcwKh2kvG1RxzN3
ynelMpPq4YCDPaxzMWKJGFJn27HgJ+SlDjcALBiwXUBWkpZ4/hDRD3eZxBW0nnUdjbOv0vHJJ5GI
ImFTnkHJh6LaMZ9THcyPEvoYaUWc17pPU9rxglGRwEv3/rk3fksJRyxg5LcgIfYYDy8Tyoft/TW5
EBf48DQtoTe/Z01Hhz5fFbbSBqiIJnvluP+ruGCecm3gTIv8b11xJxlWPRv9X5r4ZVIxZnIDvt7e
nvdwfBRBIzhzV8gWxW75DyVGKQpIuZy4UhfmYBQzlbByT97f7HJehgjuUOF+T6Fmj0uYaKodGdhW
IRp3Engxz5suQvOhsBlpIwmeRzDn3PcOsUKhyKfHOi7GvsrFRgrQAMINEC2IwEJ2JSZRkDzl8qiY
al36XKIUqCR5ysAg6wMlRnklK0HEi3WPmAGKZMPDFjRXr7f9/rhmz7Ja+M2O7lmJmEGAHLjYjz/Y
2ntj+zXNsTQaYleT3GadcqRxTSqDl8Bmw/Gs9QfoJDz+7aeN1Y3NzYFjtAO2NGNY/aU/pYmldwYl
X7aDqFoZ8G8gYPIBqYMbovOLhbxL96XTcOv620YlpsSkUFwylWQx/SAD62q4pkayK55PefOoZ8b8
RSynjnOrmDtC+SuT4nMNnlaTbUeD+Ad7YbYc19z3kO542L0VzhDEjBz7GOvFOlMVqeCyOG7rBETh
iiUuxwo5szR21f6lp4KZXqEIZBKJrw57rH3SHs9TsmVQ4qDSFBdz2fEYtDstc8WVXTTLQ8NHIkVZ
UnfsPICcb+NqSx0Ty2fi+/X0UGT0gqbBaZpDwmjoq1OkU7RgB8xQqL2byZRV5REfgXW9zmy2mQ87
d+AtUocTE8dUUQZG8Ho3GlmQBnqew2kC5NWcRUqF2Wp3YQqqvKHv1NEjBi3Trj6DFHAJVicdrNUF
cUJjs/h5FEh4wM1onjIqBsomlUputP/Q4v0KEqrRna4gxCsq/T5UV7Bk18E1Gt7cPOUECrjnFHB4
ObuVZuViphZ8PaUSKufBATo45RuuwtuDfPzTSrEbFOXm7hIe4UTt9m2Xq6jfzDGPGMQwzqLRGts5
FTszdYnQtLR7YOoypvwmLRMBIBqxAeUyfTUWD69ismjzu/lC0+IPcPgKcF26IrCCGRv0sc7sLXUm
9FxZHl6HrXg9XRYmS0z1vS5pOg5JpzaaliFZmHeVKOTulkdHPcT+fwoJuugjiUkdoVrC6LXxxAUx
FB5KNsIAFVDJBxiAyD7lYf35iFcdJcQrKciOCvE7t6gNpDfLyJhgZU1mxRwXAO5CFXRNIcQG8UgR
DY4NOxC6Wk8IZSB1UHlMg5nGSOERzeWIjBDkF4JkQyn1/z5UIYgZalta2pFeSCEXQPIxxw/eYlfp
4vGwIYxSb9kQBeMOlda575M8DMCqw+JLh2L+5T1g/oIoMXGObOkIdCd8AX0+rbNwJKIUkwYOLLPH
bfB15goYmC6bT9nMsNqKehAUTX+Q5cWUUk/B1RcdgZMmygje3W50DB2sIX7JgyMKQg8qFiNexHrx
r6drALgihTu8hJXF8I3e7N4QmPgOuh3S+Orhhkhhv0iyix8SaoBZTmJmcGnSs4blnkn3hmrXGsUz
/4vKqJyfCy8rKXMGj5TpKioJUSDi7AGMbIGC3D8xeNLiqAxED+7MtBHBg+X//5lmEI36+neg6hqL
F7nee2elwNXdgL+NTo+hkwaPspiGvY83FQuuguWDe6x3W5wrN9JxIF3ZhRr0GmwHs4jXnvnVqT7F
GKiYupqqqFW/UqgZuDGkxmt9SeTokHaQuwA/m5TJx1pfHULDbStQ00fn88uywWxwXCxAAWZK4OCl
r6+b/0ItWsZrUGC3tX/fWAVKNtpziHHpi+2BBL+32oKwg5rik4uaKkuVCg+zIhMyHl7b4HCPRUVA
bLJHA8agnC7A6qkTkzRtShyMr5pJhfHSe0oDp86dmHIRWL/sfqdQy8Ut/jYPWzEWRukp+4Ch1VIu
l6TiqoD3GQi/av6xwn5kXZblpHFCgkGls+2gh9DqkJow+jOo85fXz2HsE8J/hEcqpVlolbIvfXKp
DsIsrZe7aQhdMMBV7jlcauFtVPVNvLqqyK83uX78FbN8HKEXsjWOq3YujwJLpPtnHYi46oDqKZQv
wKQha9BhLvYHZESWyzf/1Q1/WLHzopaeEBqoXF5IBhiLH8ClVS7H/bGMYvKpQyexmgsJOPuabANQ
4iVWhEQeH4hOBr9bJmr1oh6cbsSV3v6macvt4oix0ohR+0ZT3TWHRtNXfiyzHKH6CZXGl4+QOmc2
2QdJHY5NLwd6npUlxVENJDTI5JB4HM08dM5keFp4C2Q+Hh8KITGbPi6sw4Wvrnwwh60LMcf6HYAJ
5ICYoQLHkC3BsSPMwXGEky6p86uu3+rHZh+uqnaKwO56rNKC1dHCcQ3uOAUOxZMXWil0ojiRgwO/
RkdDaDNFxAhKHuhzYmonf9ekI9wt2eFdwcGXWIfa2/37UkFRuD2DzDHnqGMerVIgxu6mIJ3EsutO
WhHWQlliVkR8FTjTK1aocR10pl/tJWjaNabQFdG7vCe33OsbZ5S7nRhxFj0cR1SNjfXeGKLbvXPr
3Z/tDn+f5C94WwDjfBCJzLcakdRSA2dymu/o95g2XldQmkV9Wn628r8wH3lvd9SNoLz/LmOp89s+
LD4DLU450r/gWqTzb7xus3v4wUa00Ju21TymBaTkxugQDgx6szXMq4vFMJOlsFk0GvxYfh15lv8+
rDGzelIlOgNfIlAu2kDFZprCSXCinnaoFD04F6RgXC6969SyJavYe/zMhsU0L5ipdOUtR4EQU8cu
ikbMVpFTq9lh/Vx0TmbyY/v0rYTuAxrPugq8KupLKmxLm6+cOOhxo7D9aKli4wiAB9+YSITViUkV
svoAiGsmhDXBem5OXMRPN3KewOCKdUwge+hOpHDiCu2LtVedC9uNfRBjYobFo1R2M2ahzJLUjUL8
OSgZ8TofJsTbgFxTTTmikjsVv3P8LZu3X4ZuWJwm4m/KBmHVBC8lKFC1e1wTI7Ovux0EAusQfMau
vQS1gUD6aXhedjDttkb2L6xoyPU0CdBWVeG+xJ+hX1WfIOScozLGXcnxwIYfsNziVibVgcLGl6uM
LXakUKMTXO/FsH4qCQlj3a+z0Gnc66RjT3oh6BmWfu7IyhuIbvIrIU8+K42zYeVaaQAEJw+y/tM7
MjxhDJl1QxZwcZNwExbErpJ1wBxmZ01Pr4b/ysUHPbm5VFL4uL2nRnuWoNFbpWlSBZXberXMlSjI
li7lDPt2vdbk26NaqgcNZbgOMC22gHNAO1p/yW648BPfSu1Q12UX8OePDxX74XOo+e4vbXTjQGsl
kOoynRWhZA7S5gLzHTI9PKIt8A9blqQfb82p6+Nr/XSZxm0NAqbh3gXORZhO2Q9SGy4qDo/VvOGh
9N2Gi7XT+dTGUTJa4v0Al9OE/bYqo/sdXcYSFRUhj5EXnGjPNfNcZHZ3OK+slpN64PZNvmLcQdEm
L59tuQjcRBOsEY/zSj8L50aJ2unkmQtUdEazPpa6ThMxtICE251xLE0fYokyYIWNWb90tNSfpEKV
auAolPobj/hG9mMmIt37z6+LVJqEahM3KNBkrq1hUmPtmOZRRY0UMnyYXdqh39pRjYTQFrqOpNER
vvltQyYiwaL+jimrc0pahJYAiJaxmu9Q7UNTHTE9DxS7mRL+CeRgueOJfjWjvZ78ohz4NJN36t9b
yDE36Rfyeifv/H0VsoNdvgd2AB/v1Dm46obYj1RHsNQS0IYMj/Pbhjp3jawrZJUKwb5YbWSmYu6w
qMVPjncdTun80gxjzlejPFYEaAoqAzk4dY0+4eILDz9xRS5w9kSr9qamVqxBIaGiyEE+2lBs608T
DUjpu3IQ4q2Gafi0ua2HN2rqaHDg58SHTffsZCNx7BlIBJciclIk2ZLjIdWfvwjWdI/JMCTKDTW8
VTLB1J2H9JeJFx0UP/IU0ceWOQQL4j1t/gykBNGafH6oxBPIgS+XN7qxr90i7SKILioWdZ0QivE4
SQA3tu6WnUO5Rj4NC3e/PqIPGcveWDVXvt5Yf0w390lhunngfS1Qg3uC/WlPIYtFzY4FEezHM0Gn
tPqb65W5p1pbuJDZJjn+mH18IjDZzJ7DNDQSN21RE2CfZQ3GMeGQ5ASd/vy0+XECDww+nFuKy6VB
c8aymUjHwmpOG6CUsciGfkI4Z6Wu0FDmTXxC/Z5PxHXJ1yzQCbN1UveK1qxzKuGjX2SwybTMxRSQ
KqRVc3+1x9RVESVXHcwVmwO/t/5XS12AjSMoFdRhqWRLMvyldGk7tpMu76Pzs/k3CGVV+jdBCoKB
n9z36V7CfdG2Vqmc9SVMMRWALfFZZg1NKjCRfTPPdXf409Tj9a/jlzAMKVjfStOzf0EBRS8FvnOR
Pofeu+dkJE7+u4RREGVe7zfLscZGxYiDg9yokTuqZkYrOXXCN9hvutiJ6hDWE11lwokGCfx8LeF8
jV7YAevLz7kemWEG/tEwaDOaKCwJsvg9bpVuMkGa5IadxZuWFfEP7tf8MTLgvuaoOTRCP4/xO/8R
Kf02FM9rrbQ4MPv/RlkzbIh4nzS9lvxntKmJrcMOEXQcPt4xEqcHBdY5vy3P5da0jygpAiVFq/sd
9i7QmDXwBw4wqz2vCEZpQpL2saAXg5yEAk46FYch4xeosH29+uuN2bHSuGeWO2dM9kp7oEIJaOFL
6xxLYrY9m4oCpdikR7CMcLaDS0VcxciZVDaoQKBhJlOjkWpnpQ+4BmEIZ8PdC5SB3jh28zflldnV
Q3H9V6GK8JVnoXAgCfq2BoDxourN0RbTokwuWTF8cQJMtlhDdmZUeLhcFAYtIzGK6NMSf7povWfV
CXXKBmFpCyuKFi8NKbrBoHhxYkl4dCI/tj8qhPbKysO8fkGajOWwxLofv5+LlTyWjE5D2iQHa9qW
o03dcB4nZcpYK9Sjw6Uywsu/xZ0B6FVCllOSZdtn0FRnQtdp7vH9irfP/NZZmTyJldkCUXrEJCQT
UjBnXAGi0xgAzOO0GvHPfDK4ru06g6nzU3UumTXFndD11fN87KZSyLrCLOBpINGSUjqJ3QQGAnGD
Jwnmnv+N4CUyGP7VMEsjzzQIrfjIwIBpR6PuzLB9dEPdwvK9/DMeOvY6v1PbTT94WxIw09y0MhZj
80dUDUk06b2qt2kkvHWmSnsew/VyVYXb6FqDEnWTG6zSC0GCoBM2duOrCcKuJgq12T7JnuIYb424
Ef93XuXE2QV4JUhIjUky8yjA+kYV1owKZCE3lQ53fpZUKHsyUZjJ4HNHSxiAqlkpLyjLgs3WNAKM
la1eaz3Ir2piFCEKQsxtL5u0ySmGrrM7M/W2+Iyq+BZayVlF7RlkfZ2XlF6zlctMni5ZDBodz26l
G93XlEi+crsn3CsXTQ/49sw5xKfQlMFoab4r1JuLQDq6k/YjUQJIcdGm+6pGmxkHjnb1MqVW6UJA
IDUkfBNE6yOPM9jgBuIFzeowLQmVY3QNBHGGF9QfVIgLdSdUMhexUPSzPW73OpfptIVORLxpipF/
46fQ4ywQhdlRu9lVUanVjD9D8/IqW6gyhB/kgz1ufk9bfKwJoroOJDaYhnQTa7rQh++y75dHmA//
EwZ9+PEE4mDyniE/+hOwVbLhTbIw0PxZ9DSF9NP1fZQ3KZZiUST6YtM8wqqq794y8e2ZGFmcNREV
eh5a9q6hXaGzlH9lYmi8k/zmVJfZ4SZ+vKx4KhvPMxJlXSThBGo8QDrdj84Wc5YyUf6htOAhhCo8
+Qp8Hb80tEfvFF6rPyGaLpPByBAIUqhXK2sGcSjQVVjIYOtax8V3i9KlcyfEuXoEp12ZQ0eEuSqF
XBKLCodw92p+2zC3fmcjqAIyVSHeL3I9k17gdmhyut8WgNxPkmWZHXoSrcwkec0sydTypOzrdKTe
iyLI4JyddaW1LxxzKkaSiBQXmZNLSdgDdEZlpsC0wGa2OwoX9aJiyQycuNUEdCak6UgQlsXtL8ld
Zz79l6rOrDIUoW/5gERb9M6GOQdo+qDSQuOO3FVpZ92F/XD/zLgdDy07egY2MzkXGRQN20GoyZAu
/nzALxW/go2XDwl3ZoGLfhbxT4WO/z7Wb3Q5qpbt5ZAudLfWh3q8NHg2zWQTzHX6dkbJp9WW0r/b
HXdYQpWEEeTYkv3JBvA+GbPduZ15ecf0J+aZNdyjJdV9zMfFNeyXZMgUmn/r1MyKJ2FNMprxtEYt
F/FOvCxXwZr8wEiBhFjGZHUwL7KnyFHHqASkDa1W2u3ovSBpfWFV8pe5qjsu6T7CBXLte7DC1bx9
TxeqyA5G4z7cTWRZBr+NHBEDfX63QHSfDTQxwKhA47K3wGX1gFApEgW9srDgjx581BphkI6ozPTW
HnL3p0IufD7c3lAzvDc4IDvV79V0iNGBMMPbniq5sKvlr8th7D4O5Sl0qOOj7PN6+ggogJgA6tXt
H+2Ho9/P8nJNFwgf9ka4/Sc2pqjbUoAWrjkIBeiE8goDjncMN1sc8Zott5hSJx06XaX1iI5lAfBP
mmDju2lR9BgiUMW9IlpezVOACfFF2/GNZ59g3DupkwDeUQt+8D/TmPXlrqUL4DZz/OZTAOlzl0El
Qbe38pVEX+as+tI0XLEkJq+vCQ9UbSOXvFnyH/SVWmb/kCnBFHmV8ix6DGPLMiHRavrPWeNxtCEE
7WcD3fUO4mRVOGL/SMVlXkh/jZWjZYtVi408k447+obRBM2Q8nVWcwgtNQZ1FEGaKgu79KGuspaq
3MNrvXL5PosAIsKtL/F305muKN36d+B8/PaE6Vs9WbDMZo45snME1V8D8K/SC5tP57wLaIa5h6Gc
V2q+OJQ7DXJFMrExUwvWKvkOGMaAcQ9bLniUoE4X5bemw0VJmZ/zA317+s4w4gKcZcAQ56u/kJZT
cHBtyFDw4WDhHH4aQby2NUGshpP6N2FZkj6gwfVHbiq1aH+pW7Ok7o8iz8SSioikRROfIen+yzYD
C6+Q1YfSb8+pAEFbGSa3bPd5RVqJu//xqbkaDkLzzj7KgVdkcPgFkzzI9Lvw0xGCxz+iuECaZX2R
4eeC//YKx6VCQrxEsedZia/pzuw4fPRqzhYoOu0Cpux2BxVi0JBLqVP5zhHtcluIZ1DbeVwM+dJg
2Ur8WW0q5+GUDEReEq69x+1ilOvTNKyzZI7PPy67Ez1h2Gcm1u6Ng6TmY3YaOcs7N1q3nR4DOQHQ
Nldt9m0mbrDGJweC4yfeqBqp1L4BXu1k99ir3a4L8TBbWwbbmXoXI9ifTBKg8BzR3Di6utz+jgcL
ZgBOhbSSlRRckyRTrFpEKRDeDPIpl+CKMILhNC5cXf/BlRMuEfUd6LG8yDyDH9DSRv936zZnG7Ir
p5pM6ZGyQm2/6Z8Og0N17eVN5z2D2wbI00mkefRFyfhtLA4J74L/U0k3IZjY0bSLQGDa25rvEC04
nwgguvOLnBgvUSoil8ET7m/NJ99qnIl5U7L5q+3MdtdFIO6cD4Qrbno6svc2hhp5CNjPCY15I63J
LI2zB8dfyLcRocVBd12Xbt8VHQ8//4VMNXHNLRGg4NdS9RmQhpAQE/JI0ZKDPsUcemB0ixbyCx2H
ErBFE833EGNYRIsfq/HOY+ZM/JFN7sdK1dWB+BaIuf6I0dZomj3ePKM1t1bGmU0KiVbs6IBe+Mjg
odnYqs9g1C3rscOIKGJI2dXdTSCxqfYc6CyGZJPTKhRCCk2B9DUavlHrTNeGkkecs/FIbkxSZdK7
4hOgI/28ppko0/sUlMfzV27DAK4j3Mb4fykba6YidT0dyLp8EJG3ZQGGdj2Qh4BqjRzj5tRpyLhR
zXIbMBJMJOcqXa1NU3wNpuDlfY/Lh7voaIEVuL19e7AnGdTW8mNRnd+s8XjwUn/KEHEtF/mYZKBP
BUvEw8z4NsAYZReaqxuqtscIZ0ghUlusNK8vt+sdz67hdtx8ExztZy9LUf+KmhNuG+ZE4WcdIYSv
2GJ5vYSRsydUw8goOr2yLqAXFeZos67/ZXh+ylSEsV3pxEWurhM3KwDPmoV0qICtpYGYiev5Euzs
3uFGYBLUT+FdlWbyiLakGXUeGA9E4I+ZW+3uh8eZwR1nrxyzpqRs4W8PlTP/Nz/DCEz9aAaysxa8
V31jM4sChxP6XGuBbNgfb1n8fiu/Z433ZOTYPCP5VUOEY6Kfm0G1/PFKKn+IOuQgCEE8WaryjRdC
WgCYturdMtB59wmOwx3HY3XZrEV2H6JCVf+pOqwgRgMgQJqVygl4PC6Oh25WkOR0DKA80dE+d88g
XXeJYLddIwNUWstJX7hdr+wL9v7O74qIQmGkjjg7wqGTs1U5QhUGLovLsoxKoponRJmofdGAuD9V
c6ttVEo529NCwV3vw7wyhsmZ0MpM/Oe5wiRfiM7fXSI+bS5PxMjT54JDlXWfZEn1iUmTKWAAY+Jb
Giavou68x8j5zlb/Ha1o66cgzl/QXOpynG/qx+aUwIhqgwydQtGdeSAM5G3COXM1daXB6yjuXI8p
Tb8isC+ap8+ICNEfn1nB50G+RyI9dmdfVF1Ou2SWWJ6b/MjJ/aRkKUmEcbn5GQ5V7AEpw/T7EoMO
Bp6WHDYspNNPOyS2Rjya/Cqza+wAKyejsQL1iaBAZTHLw7uf7Oo29PcmH9E4zOiXTptE8GweOEYn
2hyV5ZXmul5quWXXzTe1OBeSiG5uJozJMGRF989LIxLm9ytOgcvE+wbr61Ttoc9nu8kcIcIEVRhS
0NpvUe9L0t9SYKIP8k8HXiD8kPLU7UZ//joJJdaEfFLa6Y1WaXU15+bqu08P93apXfGqXg+Qd7Bh
vZhKUfvOLq3C3Me8OX3/3JlBjQPMxPBNh41Cw7qZavk95tBkWwwGXALGO2W0tW3Iruh23RG7NPr6
OZDVJQYuymhGLxjTSLf1A6ISWNHs1QsF+9yRxn7VJL1NyGyuz5d0Zl6eqyNXSrma1ah9l7x6wvh3
I4/5oG3oCtJqIl54a1Pis65ZLWfW+lCaqF9P7g1kxWWg96gHf0q+6hgoZ6kud7Vi7ZLIffPkZTlO
H8Upu+DzkUc62uk4MXkNw69zefI5Kdu7K35zoAl+n23rqoujD9ZFo7A775LZK6Ip0OEM4TjHebFH
p3gyPtoFyjykCxCiFAnsOw0oZtZtMv5Tf2l/oDjG/Y5u7XXaGJkxHnMUJLfpUPnJb1rBtDBBFC8A
4r6Qou0NSUggX7HkubDUDFuro+lLP+ULuAXPg+QcwL53pacTOwhWQqEtaxZKAPZm+twu6V3D+O2u
t6F2AlW/dqXUVRxdaMOQtVa1DUjSlS9xelts16lTPO/DNcz6jw5Oq1Xy2uiOayWAhLeMRDWYUTc3
JmH4n41y1/cf/2TQo+JveObGd8BNCOfFneli0HqGGoGLQTLhhWgoQQuQxJvIT5jLlz3Rc5Ge19kc
2M1KE2P2s2zIJrddyoGXhVL/BwnUBMilU2ddCj152XRG4mPHRFZ71QXpJkowNZXqECAUHQ1KRlbl
I/+P9pUceLWxtf6TPSu83MpPwLVv9AstYRuymrxZXsFlSAsUNpNGd6tCbdtEt4jb5/C6+s8dczMb
F0DKeYqFCnbeDlDFRaNw3iOfr3sdYYVerCk8HZLts7Fu/W1+4Vw/lgkuStmtWF+beNcL1qYsS88H
1sgam9/5BJUQmVfNDwHpNnXQG/NSc4y12/yMhLrWzwkGmyxWwhWV0joz/2I9RSavb6Nfi5JBEonh
roZZkrbqy5ZCzTOFjOy7qCP80jM6tq96xPJRa/vGU9eKSW0gvh5nUzflI64D1MTq0vnw+/cuYyrF
NZrQoHdHPtsMguK/M8OX7+gu3auYYKn+Ea5IV2pbKHg8dHVPcE4Ilw20rxZ+oaa6QTa8+dAXMJw/
CToBsLf7uEOdf7A7AcKyMndlzRdAqM19faaBLsNGsDmTvrC6tySsZ/ueQaU9FXPC7aK262nSYSlC
HBk1XsQ2gyWEqXyMi9vwLyocX9r2oc4woFX4FBO42JkGOVo1wDFsrW6GgA6JwLjn8kf6cRXDdLBB
jsT/hDQrzDMfcGM8BPN49eLzh6Pg18gzSzVGmWpDUjHPMt2569eYDY+mNJbE+6o3u9wxq3dq5wdD
1yGt4TWeaDS8z8ye7Vudk6BDaMRFszGbEmF5FtoVc8J0atg67TxAwlzjXluFRhuDfjTVouMnVRit
U+fonr9PkxTXoO26x3Y1se/vrlmrGZieLwQtO/Mgd7fBZ/eai3tbGrcYSNHYyPAADqyD+nFIkMED
zxfpLpDWtM66DtDdgA20eXhUrykuI1AaX5RZxdhsVItNbsGLhocrq6pNPaE+fcr+aYE3/81KsFEq
JEmMXkDXjtTboQMdhZzv8qotqiQTWUW30adStYbwSzMKChrWfm1jQ9FpwA/SsgoFrLRuHIydd4j8
dkxsmC3xU3Gj+XdT9a7V6I6fi61qT9Zu6PWauycsDkSoabvKFdkzoZzslWIl6h3FSQL6TFiPB3U4
9DsheGHAFEgQB86luhCUugq+N2GHuxjIiH2m2fHqiuf6KYw39CL134C1zKHAeVENnuQqstZZETVI
tznrOJDDX862PMWMUsfrLxP6ExjRBCGOqT3Okf6aR56MdnEkwNkmuh2+Fpag4Sn49SQpcwRzr/1m
HnHNiG5KwY0767/e8hOn0bUqkEKNZzZtK0TkB0rcCM+JbWBVvaDmPKzwOjpDwFtiwk/qYDEfD6fE
Xdd7zL/BamylZ+nNZjatM00Og+xSfVSmHQApDjFC8I5myj1fVXWw8Ttbc1kIe2GIqFR9wWQLj4oY
9d42ds3pX5z4sJ3fr0HxRnmeGZ5YqCMLrWMGYBqSyGB3KXGhsbeCPDOBRoUYG0P5iAQl/5u0oxB6
lvrXu9cF5nSWJe2dYLjZhaj4h0Hxt3zqpXNNGnzZ/IluUSnu7VrZfR3/zxkeL5Xl7XAUM5fckdRo
wa4WgS1h3mwmJjiNPOjOV9KF0Cq0MrpyDVFM9GbU/IR6EtNfUZrNa4gpVp7o/oIck6VIJfsnb6ri
iQjXo2OiWdOrCMp07E7FGOkiKyz77fSy+kgBBhXRwHJ/L8EuQVv7yz4/7SFygYwYxI2t0vJwEQNZ
jagXVbORWMl3/G+5jTmLQIJA0eh++0pc5h2Tqy8y1UOskaAmkx7mv5DrRKNgRdyxZdDvITZBoYMB
y4dslOQOIcoSvXtD+XrigjxILfSotwtmLemrB7FLfEashPXxqW+Q5oK5fgBf7/DGrXjk8pruIqz4
c5AlHsuvJKKAuDbk9yl3KcGsYIZgzTv9d6WshcjwMOdyXrTbXCW+cIgxo4KleSCDzx/7eF1FA06x
qIM2xNAjEdzcviloyyykq+nqi1UjtmO4I/LkXzaF6GEt+ClPzwi3pFRsv3Ec9FOzyqFNfYKEeF0+
o7N0XgR20Us7m8mHgmVqS3iqVnspeEDQx2SuSyiS0vEEksEsSkxMztKiRp6OM2F2Rt8+GAMWHVll
EDlAk7Mjr+VCPWXcMHXmMGEFc7nmIuDakAy97B4Ox0Sgpui1AZmk6a10+FUbR8VVYKbU7yepyP42
k/84qCBg1BcSo+eTu7BNGLmXH8y5Rt/E0I1lyFRZuWQKGU0WnG5VXHW5/A55Ol5ZryPimv9/85H1
sgZQ2IRlvaLOni6H8dtKco+GQDEG2ySX2BmUs4200OljDs4RUhJqKKyZypDvz50pd2E6n49rgNeI
XyCdHrr7gax2WQuwsho2eqy6FPLa3N1NyCtFX7s8sJZcpfx+vf46AwHNQ27AXVZQcVUcHo0z5KfV
a5d18Z1gP4ZvIWrgVCP6abXuT9lZoaGGBfNtA3pqbW+t1WQfkUiuK6SibT9MvxaeNlAob3PWGO4S
Q6c0w8er6dsIOWzkkxYE3VhbAzcj41avKpmMi66asJlebrTIdYGd9lsSm0dwL62itrsznmp/dNV5
v99Nr1zSZ/B/bvGdoquOJEFzGY1G/b3nfYKN41SgvoCZZU9YXBI4EbrB7UvPG8vKK0GAFRGXBaFu
Wp6aQn2nByKqwl6Uy3FQ4dEKS305fVt+2+PpIfwmdusjkQwEILPMju2zWdP5uleWs9Oz9p7D1Onf
l0k1poqpypeV2B17snPBHjIMBsJtCg9exSel4mgO1Cq+nmsb1z1maiL/z8AJ8bDR8l6eouMAYecx
rgBK+lCyRVEQWuVGrIqp4stRsJComzVG8AIM7iU7roocpgIv372MgPWSLDoBVAsXxwDJdks56Asy
77BDkkrCQrkHYvFcbHoa0eNEfeJBjLoVIC2j1muQ3kQcpepw0gyrvruZ158ELDLkI8nDWi1fdxXm
v5TIB0sOCRfddJnh0qehMy4mbrzXxLHaTxmIUuLqEOl9XY9b1hhljsT464a/0y4fR0NNLmKSNxmN
6n14RXS9qZrF0IyPrdLBIzxClpfneXSAiASW0EiGXwDJOs4HHTRuWbW4AN2VBwFpWtetvf0PXpt0
pcr7snUNFm3rLvmf9vdhQ0CPeCWyho9iQ2yUpz+PYLpRfGlVS54qMCrsCZdLfExuU7IZcD6SsL5I
goM8X76syzLIi8MyE1fDPP3hjEPXQ2ww4QkOqUlwLA3CU/SDz/Rn8M0j5XtasJIZgfy7exqByNPt
VrpPidOFoJl/hu7K3e2hen4oWfoGcEWeNw04JI2NLVYmqLxJYi++nAXSrZDKO+oys04zoi97J2db
2thLHaV5P0dvcKybi0TNSrTkRB/c1zoOx8tUmXrXOJH+GHyQurkVl6bl0u97/9tglEbaUNX0Ckuj
5Jl4AcMPXkv07ItsD+ecQIOOObxnkjbqkcMFKtkg2mIPvbAScxjzHRyScOc/nkcJfE8L+Poq5uAh
6u4/HYANPCtBcbCqdRE8XiNbjEXjXQxF4qazzQ36x5pHV9ZFKcYR0psb/qrlqnOyfh8K0A21BrVl
N2jkWvOI5ka1B3ixNVXAt9F3hhL5XMggtW02TFMpfcJ1UHG/QIm6UhlbCqafO8u2xvPlIh2Wz9CK
MVwOiiLEgUTiSbSHQUtvJ9NRVJpJvddZx5+aEvKMKeR6ipls05HvuPPHF+1Op1IVYI3fTRTk2L8v
haTTsRkxhRxV6xCbcrN3dgOYknSLSm3rObW0yMEC0T2AOV3CTfxMocju8lVT2i2Z050mttuGLWj8
GCgrS9mGWeIjtdUts0nUKMaKkHSWLpCdUAL7zxe9T6gkVM1VQe8yfo4Y9j/sdIKIUkdfEWclhPh+
ljN80ERZLtoQiuI5U9B9/RPyrINWf0HulilRO/VK1+2fZwL2msBSDcTGznT8BL2yfBARZpch7WDO
lA7hiCJZuOmCEO8dMGB6KXa4+2mzK92diQAAHdIVuuhLo6AClPjmVS+U8qXAOoFxNztieuWdbzNu
suVLF57qKYeyGSZaV+ZH0RSlhFdmjfhe3wT+ksSXZGs6lcATfunOg6cxa7jp7Psc3oHafD9nrqzK
O824bRJuuhvQpRl6T5wyFsfFZn2S/VXpTskMtEIwpyXmR96mpuqlgXHDB4RM2nO9CVm0FRS0mGoE
aMmR3MaHbHWXyDoXGIKcLh5jwJlolqvi7hZ5pxD5i2o4pIuVC6nb2XmYIt82oIa5a2JedPlyeeO4
K0N/5Qnl+4qBYDRlj3JwLutNKbFawXcnlxg4OyirdRX2K7An2qmRr6XX8WbTSVlgPQHxUEn0Kh5H
lDrG5eXDlT+s7R7f8zk3uhLkVnLiO2onARSECTeOD6dHnCX1twaLG6v1j6h7dogImrtWXooSJ7X3
y35kWU/rwBL0L09fw9qbOLIX4xCdgOc/FajNrdZ7qHIm19eyL3R9o195ydYDyNtFJJTxusj85cJL
B6J1DPhsrjRv3fKb0M+HVy1mbcDIJiZIU+FbMZ08/8Tufg6W/+su7DhSZhJ6WUyHTnwPhJi1RRFX
QnfsYVcJbefiMjFNBnpSZmtJkWx7qUbMOXO6IYgoUC+4K6rU6N0esJOMrEPWBSI/7LPkyB/3C/VZ
LmskmqYwzi4wIwLM3qX9bym5r5PqSEHIFFDz1nuoodneHDZUtuyoewNC7HUP8FhLg3BBZvvcGi85
wWinnNSSE0PHMcO4n0W5bYh+2q3TZwzTyCCIdq92bekMA9jBQ6Uu0lXxNsOoiFGYMKldrw0/hLiv
pU1/Rcs9lphnRGmxpoi+3bi3ftMcb+0yXuAzZsbkOHHWJwXuk6ecDiaChpEK3Y16/fMlt727/jb8
9jcw+QOZCB6WcLwMbLuR139qdr6bB9hTtp2Obq6WQnJkK5OJHzgikie5rphzlF5Sj4OUlHyY6l9c
jeF126dYDItl2QGZ2lPEFMlUPQpfoRNGcMtk3XDxPqsCIv1YHjs4YCGBI6vcGUVIlfSd+OddgHGt
DDUxwki/2kRHKrn7mTxDnBwdsGdEG/CgWsLE9t4u/PO5V6LaEjhS4TORkXKWt1z7bFUBdpR5v0la
HicKg1Er+hR5xLzWzlk0O83TErTftipxssc/TOsxmAqu3yY0N4U/5tr1msr7CN7WdfCN8pDvo0uh
IlMeRvfA9CoxeYz7yYFqcwI0GdgvgIUA/Y5T7gpgwiyE1ai1/1gNOjcVn2YR8h7Wv1ocJoSxi2fL
x73W5npEu3GYbvJoeBWG60ZhAvgufYGD5sM/LWdpfHtjgfCfdoMA3r0UI5zAS7kxCd1Ao7WUVzUj
sw/8ywubeYQ6t+p/0Mlcx0ywun2XgUhTF2s+oeN150XkSi4JcdL2G2YKoMyX4uCJcOAHOCmZOPp7
vJW6Wb4hmCnM3IgiSdAJ8JwAmc7l+oYVO9PI0IfxeTX3bGfQLYb28bfAbtQB9jIU1uHRSxdxwrnb
/lL/q3l+7qMbG27x+eEpFNTAFC9Jwo5hLE8tgWcRsyGv2yOg+iccP737r9iTVMZEVXIT643rJrYp
x0q2KJ8/O0WWb3pmgJDjhaTqdAc7rbk3zDfPXa5/hn1sU73zMNG+6X5iWh3IopDdwv3TRHm6s5b1
rRoE6xmdSmYlIFdlp6ZjA1TUxVmSJtzYj+gSFYmTU2EYhwUrWzdIXEf/8t6J910M41cvpoFfuZvj
qPRfh+6HU3YE/CmCukw+bhK2ySbsndWsL3hjA4c13X6q41jJAC0zZVktbXLwwLJqPkjUOqSlAdQN
QZswbxu04/n/ydEH+SaSOfCvF7t6vEVd94UdEveln9JVO4Us2x0pl2e9RI8EsuPyBjQs9zMITtAy
//3kI5e4uoYZXU0HaKeo1DD7E1aEv5PW8xOZlqO43XydCu0XO6NfJJDI8LwGi4rx/S4BluelQO2i
qkXwJd46NyRhpaI0H+ljGGXSPP0twxcxf7lT4WPbBJgDgSIDI4KnDICc6D2kHFHyCOcyqxqufv8R
Xk9G9O/p9L0tKHy3Yk36AwPBuxqV9HLzdDiHZx33BbklhHDYTUCZdA3jPwbl2X7nOzXO3p/TgNR1
cCk6a7pv+HgwNvltKZSMQCGMIUVZwGqqAODgpeGgMfizjnpBQS5c0SM6NsMk+L0yLQPxrFRaS79A
xfr2prxME1S9aGwQI6hqKrOtUdsZJbtJ6KaG1LZT9bhQugxjOuxn10+SchrcwByW63UXSG1mhoF9
0btZuR/cy+0jJwb/JoEV2nyMvMaPK0dOWeGNKR6wtz6R1XH93mg68yXYSHb9OOdsEEcBOesybx+s
5eiXYW1RSO2abfHhtBIGsQu55jAdYkFqyoDBiFFh2ktgy+5gnGsOsctI+NYeHH2zGumu93AW14Dd
FB5N707PJBh5n8c9xnOTBAwoZSLglG82/ZZM0md6jMWk61hhf0d+W+pL8RyQ36pFsY9RMoKEwuGK
kveEZituOvYRPABM6S322zv+qPFm+EIzPEV1aLkkeGPjcN557BBsl3jff7uVzPcZTss9XPGjqdVx
CpOaOfdj64nVlhmKzpxOTttNP0i0KlBpx2lW4sEDA7vu4B+aTgjP6qmKgl780IIf8k3fV4KVpRwd
qw9RqN8hXL2BDOdN0LDSKk52IMugw724esmzYqxv5GjYQ7ysfLQHy933IoC7s4/T8JHJVXe7tTkE
tgUtRRZK+Hs9FNxE6V+gmXtHxnlsjrgFHIWmCrWzSZ32H0rDO+rhS1uhqzuSdoWIwHyg7v7AavmN
QhkWq8Q5Zv05HTEfD0IHZXEDfxg7CpIAeNV6H/MpTW6kXS7YEeJq955DD1CivUlAOnniSxxkCWtG
2usPFgkZa1FNkvNt1QJFIIsgGwq/4n15Dn8pG7npVCTpzeK5MucXwCq5FthFzLN7LK0Iqmn1sJOH
FD4x2zIiOBawTuPjtpFoKfa29+XfqTMVCYxwboArbXI8zIZUO7UxYFgoG8HDQkxf5IPN+7uc38/x
kyiv6Cvm3F3VfqNaATTIwXmKjLrPqTWwgZQJFYlr+ECtYDJBAOTUEXQdPZJAl1LfhtdLwGBn/0PD
/zx9EnAdmPlz+Ge0bvMfrAugT/IOn3phS1gAeshkFG7ZGZm8G57k2CpCd5HJt6EKk0sIHt0uZ9Nc
ectmKKG/+0LZMBPo3CRnb7qf/9S4uV1LODL7+KOjVsX4JuKTMSPrjvzBC7g5fAWcauW6pVU68Duo
Jq3tDIEw7sBVX8xhpJnQM7Y5T53ZWVbEaG5d4TYKCaWOg8KDt+6I2fM+pYEb8HIZyMWTJuEf25AT
kYsrxYZ/WCZ+WnDkED9jhFj6uH3oYgBIQuYHDGt7aHag/DB8kIEEk7DF+07jHXrg9jXKrVpm7WoS
pXmuMKm2/sFHrpW/1O1Z2q7WvBOYbsZg31X6R2n+4GfTcZPvwgxgDXpfUm4qtit9Rm6F6ttzcXJt
/wFyG6VhJgmWTcge6g7p0eKhG3KLevV+dqCTAi78x+sEpQPkPKVOrdy/uAEURE/sSgyrazx/dU/y
JhfSEum8PRNAh468fgFYohvNdkT3VoSNBhx106pRTy/40tVAVQKovtQ7r363P1Z3L/4KxmC7DXz1
hbA0L/wR60rtIm2t7pur2mZlW1Dmbaufxm2eptmzM3ovQEIsHafg1gwlDqnIHoGYE+y/xvthKU3t
oIefFPC05YzvfkT4Dlg4BahZM1ZxErvDT516eSeuAOC8rkMa+InCtfCEHdnWtJd8Ae6xK6f5GjGa
UiI/RvcDBAFGS1lOAWjqRfJaAR6kogF/neB3tD8knnGO32nuMflxkuqKyzE2rKOovGN8P+UbMlKM
WLjYEo+ntI/DIqCBY3ZRM/QLgCb4GYt5UV0nXbOx8ddxlfUKvOppScFFjTqSSPIHIGSLcGMhRSpS
B5eeX6Jir5la6tF0/tWgRLjTmJNxW24SzvN7IlVNkRufGnk7kUy200d6tSyfQ9bBze3wR+fClK7S
eWRfotEvXu5Cz17eBnfAKSt/jPI2kxf874Gbpi7yYCLuCljBJGsZmgRDXhTr6cfbrswyFbj0CFYp
Mn/tbAUQWUdk0mHZeg56squHli7en2upfzLdoHEOX3hCzzTNy+vm2VMWI7Ilspn+cIL/yq5Hz8k4
wUBaXoDk01pvJ4SxY/Ji9pZAI1imobOGuLARQ8P4GIxH1Fr4jkdM7Z8T/zkqZ96AVhzQJBKrCcW3
U5IreDirQF2sf9AEtOjeUSh337cIwmFPCd6adipLHgKRIZM5lsOkFd9nvHh/rVMNe5s5BeXqGzQP
JhXuomsLW0DAHEgVqirL4ndfRJL+oNi5C7cTcFJ7vuzXVX0HvudvNCEIGkKNwHHruVaahRyKh8ie
vr91lD2szrxfwMYYPUKKqaP3N+siBvlQQTxrovUgvjJA4eo0c4ZR2CrZrOS/jdArQRpaBwPS6N9u
U+/7LUZiki8NVTLdMV1FXyjQRcu3+9nbyEXmNuQwAb0oQ+xOKIJBa6bwqjgBaCTNBvtpqrinsm1n
QY0uvLXiLcZd8Z+eWMp3YZfogJbsqQ/rhAW/1ij0H284y9+dbg8gnwQ5JnePudk5PdDjFIoUXqzB
nP5XT9RbnP8vdro05NVJGJiLyNqRCHwsuWbWh5eTyOxRr6BhDVRY09r7+opp7QUEdG2RQj/horZ2
2RT40LxKdDj/C7mOTy5XzDR97f0k8glS1fvlimaJbxvXd+K4iF+BX68ZIDxvQzUVw3pNN5X8LbRa
0bDNSuKsR3YPjXWWYmvxP8GZk+9RESCCRkZ2uyIxeYr/zpSvrrei4ibxx8k3i9fmt+285W0K+cmT
i3sw6bT6h0UAAHgYjxSXE68TOqzbz/tlvwDTKbUkPAh/EdH/JmtjVOeG944jHUOvVsMkIVT7IXON
GeBO6rkv35Cvl28rmlfPXx4Q0rR+VZSvHMv0c3cgMqo1nXlFLdDPdJST8VQSSJ1wwloFfXqzV0TN
8DRrWEgxRittkhT/cUmg/klI8adw+16UxYaxJWAZ1ZEvTYCmxh9lX7x/JoZalHE9UUdlXtssnFt5
/vj4imROHrPZU20ykPDJbdr/coUO0pAJzfq4xvxhdwrHVjU6hpNx5pS+cdQFfV/qP5bOamKmx0fm
LLImnHjExRg22YORh/18aYtMCafUapdkaJVHcv5fMHhmQnUCuypB74vqyrfVIwZ5Z7Oxtyyqj/Px
+TITNjwuI3HS/ZX09SYXBSs8i+c3t+FkuGvr4EyqXcJPCVjoNZerdlprb3l2LGjTLHZM7z9dgGGF
QRxBARKw5SjCFc+kc8zOg+Hye2wOBftCCUuWpAscLB6ZuZPXYPxj05xC+4Fjwv6K3+iltSFAGZGV
+NGs0Nf7Rzv1SOPw5thSfPQpB6AZ7UKUYOgIPsSqjCEt5HLvlhVRdurmuvojK+6W8DhrS6dV/PFg
L2eBpBc69voBTTRl4e+e00OMhGSsdpROK5czy4ci1tX1nbnvaH3VIwf37RjtadekFbIg29RTIQmT
TMgkEKklm/uRrkyz//PRebf/MONlkkxo940BEwFydvgE5W9xxTJPDnlCVAE0Q0sSMX6gQFUwph7e
AGdokARlG9tIkiz8UI6Hdo0+HDp1ZpmnP1rSdrtrsWwwsP/mOHzw4Y9PzbS2TbapYQ2rAwg3PW7D
dSQ0QTAg/HRQoLlkGLxINBq8LZL9nz/CnDfpBCBBrZsGP/+VsQOtqPwsahkUqWkLgu1MNLnDfgqG
a8PGgvKjK8wS36hSHxF+UuaLrr9dAXdyyz5bwOJzFsTPBX/jGKCJZdxzZqHbYgP/R8ANi+HHY9Jy
kMK7NJP3WoSj71x8hcanoDDdc0dBbkh3FzCix9mg/+/Dls42aT2QeGwLk33QwMqL+AxKSgLKkIS+
3Z+cpByc4AAV2mYtoK0k+Jq9q4x5AzC8wNyD/HMP7Yhi8wrueiK/ct68aQr7fhi1bA0v6yuEWsyJ
4d1bMw2cgAmSIF/3TKzKpoH9IJKFGr4869kI75Mq3vefZ41S4l5vlNpiYT2sVWI6R/Eokz1m2qMn
S9tkBgwkYMSh+nJJ/0+eHZh6REEvuti1hd4pgytGAQCZBIN5z4W2RS9wIEt4z21K7LQp2I3zOHQv
tDkU+k/bRFFMqJAptNyW2cKycnJRKWyxc1GqAp4Zlp4JZhOCDDCmyl9hvo2TXTW0Dby9gyqXsca8
fGSv+MvQp9TvWKk+UY0P31O4ECgEuJcruvNqCb0xxoTumxlfWNC12bPuEJJnhkF7xt9txfDTc7B/
SUrcJ7vbJ9B+SDL3rhSco0u0ZeJvGdfLhFFOty573IqAzWIvw7SJrJdADT/xGxQTL+W0w+jJfiQT
TVIOb4s6bmiCvmDcRN1hHnjswMZU8qItzsByvfu/V0aarQXb/p37iz0B+7SgFfaJoTbDPirseGK5
RiZ/M44nzY5On1uOSPmExGRmBaLlDuj3pVTl9XeakmO11B+xfzNwE9bAgjKVwo7SZkUeha3WDjFe
3deJ8L24lNe8NOldhJ8qy73JsfIKHLDL6vrv6cubF3I0Vpyu7rOBoFmw6Uyu6tHXokX8bEhbBcOA
4bT7UqKuyhTlJPXKSisMhYZZN5WGFtMm/ZLXki65YAMlj4eRgbSmwY84t0KNxHfOdrNkTtEdO8C2
K3ek4CwKgFl3k6nHqKsu7J8CX/nsHZQZYdQg+5cfDVFtcIS0mrFmUzGffzX/tXd//Md29/GytlzZ
LmqpPxwFnevkV7G7hASSujcQ5S+HmZr7rKkfm0aup7sH6xsTxRGpdXNinpQaXoK2lML5rNRlnf5b
7RsfztCSSBENckyiOX6v40gSTOEjmcajlpLPALYushdimtuzwS9lFPpT/LqNww+Ndim6cJB3wBma
gBTh9ADt6oGvdXsJUWYVznMxA8grwtZwoaPyH1elgLtaTP+dQvMNJkJMUtmXYhJXYuhq3nuj8FM7
HojmMSnr6Itq/nvJ7ntnv2hM0wg0BkJMRlMaWgv1WI8FRvQXaQLAdr3bxhpP7/SJtL9uFvWYiQKj
j81WluBdjY4M3DErNtWhJd2NKeQmKGAfQLPh842AyqKOyzCmQKJQwaPZbhWexHAAzrk1+ZdJqr3k
0OMEk2LB0nKNLNYKM0X6/qesDEN8s2c7+RGJlaIhhwndhMfTx1ur1tOSw1S6DcJ5FsKf7acL+5cB
5eeVIqDFkVXKwPDa5PgVtNxkIMsS0VbYFlpT9rWf8dJ65cauuAYbNVzFMcoGNjhXNXp80hNCESsk
g0qQ5XNhs7DoW1jdZs2mIIe+5KdcKjSC5wq7LbBEIVCAJvppM10Puc070o5B9wMCdW5V4hMrQQWr
mdLRN3z7XQUUzCDsDJgY6CEsywbK12EKRSZgiJBvjcZcT6ey47D59rXTy8IsLsS3gtRPLJ85Sflq
cQZ0FMSUEPZe3o2qJOmtO8aQACDydIz/CbXtl2gJLOOk7cziXuUvQ8y7Yys8q8C7XfUjZQJBk7Mk
K6AbsnCfn3Eo+Tz8nisYdhDtmuBZYK2DxAAaqHxvPwQjhRo3Sm/5b+j6/VpVZOfnKPglVIBEsohm
NGsCoxyZyfXab8plL1zXafdicD2UZ9zwb46OR2CSVzbsz6ohOipSBTpKQ+uwdB0sGTCvpl2LgxEj
DIyE5Q78MigAI/KyJO6BQAzJWFVQpOyDhtZuUVVAiPv4ZeEnVT1TpnXC+j+5JGpqiMEjgaqFB64x
if+d9hWCMzapCmuj4TX9rktWkO6aVbKeoqeR0vnKQFdfbS3yl+S+3kPmQvBN5FpWVLdlfdzqSnQt
oGkK5/vsj7MeVq3kFVuVSk3kJjt66kXdj6tsIo5W48EctbZNCtYT1ZOHyRtRH/l7Jaud4ytqQ/UW
r7d8u5KCdVHf8ijYjG3Y/o6levdeaXz141wTSOnZwga5KiR9VCqTbb9ibM8wkiNeaMeRBdbjYLI8
qDMvm/qwbwuZUaYowoHyuRX+EQ4j3y2gxam/mmXwEjNxmktIZU7F6zDX0BAzpxnXbHia5VrXt4VQ
OEMcXRyJHK2Uks6E23ozU/RtKAcNFpNnbiaqbQsGlJ1OuXayRA4YoZDIujYct2shjN9UYVLbHg9O
z/pkFnXueqlHPA2RQr1p3NyseWwaucbEWgf5Df92Io2eXXBKIV876oEoV5qLaAfdBf2WedAsAkJZ
Esd+pT7/uXV5ImIbWBSyZHy7/dTNhlj61NxSi56Iq/cqJO711IImqoWzW33X4kF18EJOGlXBB72n
vys0t5eDypBBBApC0UgZjGRrL9AVOLCnj8ScUo3INT+jrSnXjeMomy12+Afb3g3JD6p2+XT1i5s8
N4K+UYnThdloBJh1rMuV8LTsjlXFH11Bvb1yM6WhvTUuCGUrF8OS9pKAdhPMZcWms4rhLYl/M9QA
XpSrdYphtDqkpIb/AuBl/WWxUWAn6UIiJa8skHJApwTKqGmjveQJCyExd5DSxycEzb9U7KXqssk+
7xNQFAutXatMjU4xsUTqHCh9YkwNo6FrOS6J1uKlLpF6JOtDa/W3xV+tJCa64M4NGzVd2s8vFGpv
tk+mKawJjtR2gqUS37xheB683e6CPnxiNcJ1vWzaH1va9XDIBiY00/+ER56ThpeDpWqLk9cUA3C9
KC8SuVkKLjQAzXmToZZUF5AL987nyBMKaTEA0k1qTxLauQsxuHcOcPIvU8HkS6UFO9XGguGOuOSI
vCZFoGB8Cemu8Qf/OlXENDSWeq4I735L/6bAxo7i0KMtW9BBxhB1ECj9ifN5ixXhJaCYKb6eOzkb
+x9Zr8qqkqv26mZuhW/ZafJwKF2OCninY5qofLfEZWrigpsovvjaHsbpu8uN7mxhVj6isW4yX5QZ
SJ4o3a++69BJypVbjwOmZmWuXoKnZMZR0ZiyNMHq1QQDKuY9P54UTFe4eiy7yY4bQniOvd8AExYa
JMl72IR8Q5OH4V8nnx+mja/3q8hF+4r+MdfgySYghwlUcXKQdf726cIEM1UBhqYhLB+wP4ATqU4p
YVPOFFq9937NEPbHAiwZLl5+L9r0otC/YcXRJuyRcCVo9wnzziEETnOGNu+4bV7aYMkbVcoGHSq1
VW9Ke9Cokx6t/Avp8uKp5oJZbSW0dTs684ia519IAPsJvhQkvsW5SMfm5Av57it3gmLNkE6P2JGA
HzvrG5oARy8s4URGek83W0s9U2/Ba6jxzGXGum1VXi55G0lR4A/sEXRSg76No5XUtvdGP5MM75U5
gP+hTGKX8EFi10vPZbUUGu2ahzmxVe5cE3gbzXIUYfX8KsitOAy3QKVpVsXGfHpuea4gk+SGaKZ9
L74t4fDx3NLlyHG4SKuk2Z8CDVySmIxFRwC/5W57IZKiVJNk73Ft1MX3FjkH6Ovd3CSZH/ycg/YC
aEMsQkAGUcnVic2G1dtMlZi4aKDamXJ3p75Kk1M3eGJY2IiBPfZLW/URnIu5WwmXpwTUJ97Shi3R
UdnyuG95a8oTseNLkYaOLvJeey72GR2jIG0cP4I+73raiZ8LzL3D9kPK3IylQO5/t6hFVimS/fnG
M4pEj/OE7EM4aZxEUNn0vIpVwfLWJnqqu/zfXIGBxvCHIrvZW5llGE8g6zll9zEKh1T/rOayk+g4
X9NgLHvGlXmBYTBfzErBoJ8z8RbYckEsBAlYL2UGwK2ar0pL1R5SNJ9G4123yXu/xFMANfBp+cL/
r58OfR1mlm5QmcuUTHmA/xz/LT4U6YHMIPgCKedZkwFXlvp3D+2iyW/Er5mmg8l16BazIy27LYNJ
qf3GVB8kN16abU2L8l8TjlU3MjNx2zONkM4mx4UFv9cRBfX79DbiOBxc0hG6J0fD+cvNYfFmKP2A
7DTD6Zzso7Lkm+raLC99aU1xy4MEwcc819Qop+luFufQNhBNU94K2ssDYEA+LAv+gR2VIQRMKsfr
pcYkZLgsKAh2w2/QVrZcL5rFDbogU1/tH5nWKO6r/b65Sf2JHlRPrspcam/wjQZVNGEaEfCA2Mgn
Z1DVD2HJv2oEUUHgzk5QJkLfGZPmQoSLEsL8y9/5BQq45gK1qLxMZdVonuC0MgBK8Gmke2ubNz7i
LvDloxIWN4KeNW0jmy2t9gjtjZWG+5CSxhdgTvR+EMaPA26E46rmoFeXPO6NuqlKGh6c6Da8enTO
GkWwZRycKuVV74SqxAwDgBN7cQM86sA2fg3rcubawZEp1lD45c9c1gp3VeI7o4ozJCU4odGs+oJM
1y7fZhIH3naPBpnzYBDiE+b2cf8xjZkBT2AOoy8HHuzGz9HTTsJz4ADYkudT1ywUN63kF/FJ6o2H
ywwjJkCyCbmZnK7tDJx4qyruuPF0ONwlt9u75OjPjCq/gNuzLLCRhNLgbAsaqAE4ZIMDMl0uRigO
1Q3penVcf1D9nOioSnMMvDLkQgp6jkoy72WCGR7k4MCk+dYah/Sm2jC0FbT8tFloWmM0+7pXucxj
grh3Y/+FvZEN6A5qJE91Be3xJBI4P4DIv6tOGjUNxoKQflzyTdcmYfTLGAZs/5UO6MHiEn8o1i/9
px6HF+r/22auJWdhkrL6OYJxZpjpnL/6sQIUa5cPdMnOernyeQ3t6McAN3ngprGkquGDAeXtQcQE
oYAQA/X2Kj0yHOKLV3StCpIGaiZ2+5imilEWvHh4uSt/4NPZ77u096Y5aW96wmvK0wptRTbwIUk6
BF0QxdQRJFY2c+Tlek35jctFiWcMU3Yqw2WZpSJxu3FKKol+iiuwKWSkX/JiYjR/nhsg/gN+f4TP
4blYDxnQEsNbH06wbSmKDeQtRgFd8Y0QoEDoBANwYpYnYPuo5RAaJTT32CaL6cy3rMXQpX9CyMeJ
euebCuaaBPaotACjRfabROFbufXj8n+EhMsSm46A1q5hteiU4cTsLh+wt7W1/Y0c4ympjrsdapw/
4YBzHBJOIaGi9y9igOE2GEDSSyFn8p7iZGRJl9IpbLd9GWpx9Jd3MMcxqTo3zH6s7+3W62PGlhbR
OdobP+4A4oAL6wto5OQZgGXGF81UWvaQSU3Sd8Lvf6H7gLje69NVWHSMyMUm6QvQeTds+SBZyTAo
0qmj+SlJl3AIN8ZdMI7gISvksKi70pQqRWium6E6lRIRvxUtV9muRjt9DQoksWdunOp4uUdn/DmJ
6mBnLTRPI2wO4ourR7gi6V66JvEducgoyA6t9xTZWl0WoKACTP0aBbzFJHlj+GA4PMDUgWK7penv
zKSbVt+/rECLbhoormAjm2wEOS8bWfQPxZm7i1Rh7TDyNtFJuQu/vl6O8M8AsvPLlvChxNEZ6vMW
mkP6emX2Z+mYahtT+hjT1x7kRGYrzMm44UWkl/fA3CKvHa5kJwnJTAHD2uTZl+ivtQtKqM0zKS3z
gOb6a1nTcHdSjotF0SAWvtSQ8fhQvhKtsKam5FclO1zBaZPINofgFRD7Wj6+6ns4ntuScB7G+UC+
mEXo4YsKbZvYAFuCSZICHNge7UyPo0rtjMc7JYjw3sjqrX4XWlza2G8rlu5mv2bAFRX0BFRFAPOP
f1rHJsGzji/s6pdjjP0bqWwi/p817h3pWjXxVDIsh3zlQPuF+Z974teiApfqIphgW6qkB6u8bSR6
ls/TiGk8LT6glmnOw6z01unRXlxDclVHyvXCa8UI1bawLptIW95wBOLlciA5EACptbP69XwHhKXz
kRoW4mnNCA6NTmMLAjxWXBlTzB4QD2NhMcsFWG00kWTSwBgbS8IMDqpgskHz8Pi+/hTlWBCTyAYW
KjZ5KYSFL8V+L1AK/ytBVPVmnSNMsp1iVyhna57n/m2wRpvLDkexOiCtLJY5H0cRC6uosDexkfm0
jZ8sf2NMyvKawljei/VmbpGqrnOgujCrv9mFJ5k4yABeJ86lKEcyBwqd9FU5lw/qGVRrHd/waPRP
odKAfm7xlxPSyOLD0Ajq+8jRXK7QSOyTtx6Xpc+6Jj4jZ11ZYp95BLGMw9Rv59vUI/6NKoz9ku8z
I9AA5dLtJ/PcTMB10p1tXnnIPMvZDDyNuc6V8mCP38DM37u63q1T10vyhYHuzKVcs+OYlw06umAo
DYvT4xgxdVguhyPsWxjltORFk2SmWXEsr2DPlXzbPQ9oQi/A84RyDkfgnByiP3ee+fD1Gyt0FqHr
GevMdYT6/lyngreBORMJTOtcjRlNdOPwmb6dbvFMnvpIHXXGCQwbZOaek5i3+mbf0grdyh9m2Ifq
MFYgGdR8RWGmZ0pmVjPXC0P3F22kNsfAjgy0WlliMuqVcxEv0p6tN2QVUCVVS5TtUrfcdDy3oCbR
LtGcKASusmKGnbdC++EtW5C4lrFTThhMyJb7cfAwvko+5V6jHdJdSCcvY+TJMRaWEUI8DloW3sfX
KYIx8rVe5SKDevqgjIJNwRubBG9Qd4UHpo75GEc/YJBTHCF7nIzYZTkwq85kYSXIJKpaUewx/0YL
YURVyzLSf3gpliOajmNG/C5Uczh8eeNjIc2JwraI40PZbQ2z/u/HCqt0yAqoArLcYbBPi06lmyeQ
oTb1FrFiZCnY60ZJmft3OH0lA2uP/4OkJY+HEQO4+c4WkhYPAUVtDMGi3JFsEWUHhur07XaJArf4
Cdnv16l0GGd3tV1H7NeTcOTGnCr/JPZSxyi9kN4qSaaVVOGpQEwGK88pLOPc8BFV5OEmJ5tRW5ko
/ikG6Pm3S44AY/SdyRosuL+kapqmsAufflIO69lkmfXmIJHlicRy7eCZpKfsn5/GwB0RJMPnhBtu
Z4wXAM1TZJygD4BNU+H9gQEj+X5J3Y8YRa3NJAoMCVPNOn+UVwiN/Uub1wS83IdtKnuERNB8eHiU
azvkgcGUMZFtfEM/NcXYAntGWwp3+zlNd57ARPzbS4AdR0oBEKWFg+N76ipHOeAxEzv82XClGkoU
RgcPxPbvQwOD48fMGlC/J1gzL4PvWTdkRKM8GCzR2HiR5WiWdxbFLCitLYEDc+yRbHkfSVZIQJHE
xrMAlaTVR4AfdBASGlT7gF1XVe2gptDkoT2bQtyX5YLybsmLQlRO7qdSWDZrqPhrMsYGG0xjIiaG
ljNR5WY3/1E9Z51GNgq9g54kGw31HdTtX2L+vsIU/FoKIO4azC8PmJbQC+fQUtY3U117afYIXu43
GfoCuphMqJb2XsUWyIgMi45AkLEC2YjCvlvqDg8x0rYgPga8NbU6VYLME6KbzB/eje3tam5te5Ou
GJTzhT0gWEvcJpcTs1qu2iXCQORLLuxK7PfCEZyc+C6Yh43tLYT7lWV9y0wln7YXis47RlJUEYf8
2sGGpCzhhYIbisOW7iiuU9UnnCBvAPyBrn/aznfMF3FSnEQzXb6qxqyrtD3nEPL6Tu8mVcvKpOTJ
wLoEW4h6hHAJ5KFNGUhdoigZsHbn5Lne2XZD60TmyK4B87/gcXHderqs6syDeX0cyxrjrv+Ktfmb
DrOSIfZPQX6cMMS04eueu7JlYhapXlnRgi3VqksoNMGBJdbG6BDKj+L3eAclPI61y9PUmpnOPAtO
Nn5vYYsNWl2TBk8wtY3zrdCj7Gg8az+tNjLkaj6NZ68rFzwUNaUOjxmwyShoOAltsxpzJA8/OE8A
VUefazb4c3pmZpQHzTNahKB2xD2fc2mYxnTd9GbbT7oNUX2MBKPwCklMT/ocwCwvlXFSWD4XDvWH
iiEe9xa7g1KNHfXRKjgtOYUx5WQ5wO8fueljEyw0WwAGTY3ZUaPjGUXV8pTVGD1tPqqApImBeKvk
k2woQHwVac1L/R0B38C2Vi8rAyUqjxoxLtUqcVmH64iKc8xHbiCC+sMwd2EHCWQu9gf6x7bB1CMO
T+g18QOSxXpegpGuytJ6upCt2aOIoHpJ18BcuYxVlx3sTL3ncJQm+nwpnHE/BVPvrURKXQRU4y27
3EmrwTEetUsTGKUHAet1/qfgEvMtHH3p9OST/FPCct1C47v6+bHZqOAJFyftd+gTwPlXiDOg5df0
GFuHwfmaxya6O+MktaaR101NwjxAfDVCKwPNXDQHC7n6s/6QO7RA4mMcIMdIamfOXHZ0xG1HbpU9
JN4f448hdrRnCgLCx22jJIkUD9JtS823GzgXUSp1is6AgG7cpTkNa6j8O8MK3LRy49WJiDWH0edc
FFHBV2jOybarzYJ35zYKgM/HnYGnP3RxpK2iDKVEJ4ni7kL86CaLgFNCnndXYos8Haz/JaUuwQ/H
LJ74TVSl7YGQSqk6AHYmrzwYM4rNKSSzCkvtDcKB6kQoqQJ+KPaOatq8TUiRsNhNrE//OOHxfxYL
elNhsfqVPATOIwTXIEVvoLocz8VJk+ali8Rtrcxny7uP9Y6YH8/+zY1R+TK3ECIywkhk4qrvgj1d
BZDx98anotc3iLCoAMB1ggb97KZyngEdQe7/fUeI9o0J734ekjFchX6jOnoVIuXJL+IARJ+gyYa5
p0kujQ4EqvEP6J5TuOHfnsSeSYdrrmNP8MBUvT09K7VNnnBfpM9+/CIVaxujwtzmPgvXnoTdi9OT
Bpb/k3LL3VmHXPoB3387p83awYqZHVyG+POinBdiMCKWOr8WqfgIi68HpDqkT0nAfeudIAidTTZA
dZRM+NBCo2hD7Km5qMQBvL1+MUWk+X1twHGS9avowULMqsMwqiL0FbOw8IqK+jhKzFo9VyvTEYpF
/CfptcJDTcw4jHq8qIpRx6UYWJVxZcvWyHOIYV8yITAXL/MmJYCEzzeU219iMPZEf3ADBFyYXj/o
P1m+RyTLxp7Euza2Qp7yf0GEE0Dphfh9lhdiHZvpLzMyUxgLbKTVkhhpSm4SS+kZ8przISxCTJDi
smDdSI1WYuPEn+0/RqUstRuNg+o0EwW2SPiKbhELV1mrY7MYw8GW7UYXESlsmrclt9ODxCMO421L
Czl83r1FPoQ4bB6XgBnD2qzogV5DUGWAUkHYf/hEVGhi3f6wqhfVhAvl9CUVh2mCXtcNwLzaR3kT
GZr8jkl5DfYEeetwVB9oeE8id5llT2pixYMqtr8qLO1SPsw/g+J9b8/shtRb7IPNyW7z1lODFsqF
nQFCTv1Cx1t3IComo6bBa1DLO1Uo8lFoiCRFUghU3uyT7iZtPy8YsoP6cDQsm9itD7yLJOcPoPvf
X0wxCy88aIfFwZbNFH8eKDhVZ9HxezjJhsi5UinjUmL32cDl7pkqj8eqjBnx7BJyTPSvMuHe1h7m
whD/oyXJtx9TKmEMvg5e4CfGD1GfmEUhlSrIk/ZtX1B+kME9/h059Uu9c3zDllzeX/JKpWHZ/wcM
YX5vStJpvpz3D+s1q/eTz6f5doE5s55hyGv1pQnGOwzLq3nPLco06lajCTaBaUaZq+ysXYjQ96XS
e0WCF7RDz2IB6VwLrH1zLlpO2FjTfKF/cXUqV4XFAKA5wb7v7ca5/r1STucYX3vW1k0qhmNuQOnE
Hhh12rNPU1jMPolOPsX+f8AUsG7n0LezHOG6+ctkRurBLY2mOR8C1lt4Ki3BgPIMMW9Vr8kvGi3d
CWoAERKxKnBxMQj2fLFlGn+15uFglLzkc+Rm4pVA3F2Qz+4da75GmQz/0g9tilQCEyEfddDzbZI1
SxVO/TU7vM02rV6t0s2vRPeiMNj9HIEQBt13+0Lw3HNQPhYWWIndlEAB2vgzMY3ECXiDnuEIX/T0
GIr6E3/+XULOSqL1lj5Eo9vKbkEeSuNsqFUF5dfjIqcGLU7/Q1Lo3PuPM17Hhh/ZHOXKtbfX78wO
ZhuAWJf39KoiEFgps50IlO1FiZtdNqrdV8Hu8Sm/vq+bCkxmKoze5keRmAVzwp2bsBV6tezo4hzZ
C22f8LtYVod0608Jb7btrUV5N0DOK8U1Rega7B66g91aGw6J5FUfOVOWSG/ehYTYO99+pu3YuVbn
Zx0iSHRdEl+WcryG/FX1Z+XMLhgOrRuA1j3ZFJ7/K5TLdF3XsRECmGFlPHxO3Iup04KrGSiZ2B0z
120q+H0pHuu1YDOlGhw2OSsXHueDeC9oN3FgKEiQT4VtHjuFRJx7ZdbsSB3Y8dPSFkTSgZPqez2t
Yrgu5/lU3JFAC1sTKuFooFWTFA+n358JX2UeSVmlJozNajJ8G+hwOfSG2kQrHZffOli5pa6cuoHd
hG3iqlxAvzHqjlsk6kzL/29a0yPJb8F4cOI0GC+tlIb6w7kQGl8Aj+YVn3ZLIP2a2pG0RGHdCHTU
YdEFdtZF7U9viyLfjHUyXos+sPuIvgr6dTnW9MBcKFprW+kp+5xkXM1ziDqRPcAZCR3cqSplIBE8
AkISnztWo+nDNw6yXPzAkbzNIGI11Q/LuZdkgCZgimeweZne0PonAaKGfrhtW6jlV67RaHT4sV8P
srwXMHDfAuZ9IZPAReGsXurfU4uAoAiqqIHSzdJ0CK00ZuwWuWg/3jEBWFz//9idhfH3m7j8Z/8H
KSYYoi6Wzl64SxOGLoAEt4qi5RSbSp92WmwDScbtbRWW+nIyyta78kZfqB8HFWcZhiZJB0gYU9/Y
eF5SQ16L7lyBAGmxaPSFkB/bGzXIa1mdbEltGYF7LZfELC1+5sT0cgXcMqrMIOgqzw1l2qMUwUMW
VSAzzGMIIPCKwHT9C64SoiCwD/urHuooimod/2DXplANiq2H7RXUfyx6TgfyhJhq9uxTAcY9mj68
aP5u8e6An9LAPZnHNClokBYGD4qubW+KzCXqyT8nfMDeDgT1KzZ7HdWpZsSYKNrwlFhKlMOxykHi
llnNrZR0HejrsBo2b26jIjS0GFSQg7ha4XXVNnBQqfHjTHgN5U4psl6p+pPjQVibi61cl39JuY9V
2MjHYi/i/5Mqp8li4iFMMZzKt+UgyrZCdp5iFE/FpP9OuKMXLWLEW/U52uy+f0S4yjw2yerHM3ua
9pMt1s93fVSpGa0qld0iOQpIgUTNhSQ3yNvFG0oGMmeDm3mpRsgTsEOvEuxl3/i9Aa+SFUm+N1qg
kZBiUdnnC5kZQOzfDbeMnDMi31rXDMYfM+TIIdqc1XuQyRSjOL9Efgt0HBV7bSkrrFdCmHfLL9z3
N1wbNWdvlyJCbZB8zL2Or72ZgxBFS2XUVsaO+ZmWOShQjYgtO1ebbfpOdxZ5QtgrFMOHAyvAyyMY
EYYBzwM0X6bWQD7xZGZV4xeqv7/6C0jIOU+B4YZ/NIy91Q/MVY4OxlQ4hkLWwB78ZvXUQKIq87sw
lDw84a5GZfSSwV1UUw88MgdAPvZbWX0SrVyBwZaqeDISokc7vrP2Bq564Mg3PzONgZXRcTgyxYVE
auvvkf8esr3ACb3bNXmNSMxLlIUuWcm4va1uDIUUzLCKnwcy6vYdfqXupdekH32KonINItxXzqry
vi/ugIztbP6fgJauxSXA7dbEt4lZzY197nFakatGUDxRWSgh1FvMD38UyNgj7yso8FA8uZHh8f9B
lrwmi4bjjSwA8/tco4MZsjf6/TOUmzL8/R4SeTTlNS8ffBQyXRmdi16u2KOJ9coq+RgUDmuS/+B3
1fZmDD8D5KDiS6dCjU+CquBc7bXLpBxb2uO9TtGqEXsxNcOmqJ0Q8lJcR/82RfjEek49od4Wu/fG
I0gu/6rG/YDL0qjAexEkYrWhy1smFBQ/8aidkfGA0YHKm7lHVVwFqZh25kSfTNJC66RKTFUrz0rs
i9ors9HhkV3rLngI0K/fr7SK5iHler2NlED9zxLetM/9U9q9O7KalQHnsijZosAPLpyvPLNdLpBV
qccYnDQS8yzHfuqH5IsEhfKkalzpeR+adbi4cQCz48Pbpo7kgqq5lwLwXkp4ez78eLPsMXL7xHqi
b4euOU4pf1Ej8v1DjdLOc7zhgVOkz7/P9ir6mlygTNBWSmCHzbcEoVY1QjoRS1W9WSIGaJto8UFF
jZjc0aVNqo80y5vc0KLE9WyJ4VAcKzuSLAigj9CtezZrAOUJ5jVCg/Nr01imHzefylYi0TeXgsY/
NsMyOeygIOZezkaSlUVyrxxGvfBMomhE0IwSuLGcm1OhdSDzdM8z4CUyqYTLqelp/u5B8N14KMbM
yORNQGcDIdF12gNW+hm2WfnZCOOwQKVn3NwQyyAFN+54gZhB8cDJoaShHjeH/Yx2bxqtgR5TU8wy
pP0m/jQhY8LgrcSaBlQXCMbJEMx2c9ym95C5urPc8IO6Hcj9bB0Oa5lHavmiV/XBEIimXq7magc8
1SmDUafR8mshhLv00Q4udNu5XPwEjE7CjIbz/T8sOdgCqQNWfweaX0Gu6iTxMhf+BsdCEpJgtaq2
O2qChE56GeeimxY8J0qxjdbQdIwE9iUr8OY/dbc1ckNZsol+rCISPZY7UYhqNCZjfxioqzTvqmiG
4cv3kyRZBsyFn6i2LsEM8oyoTfUNaMtCqpr8DKIEgKtBRzTap/ROmtTBdGTq+Dt8f1Zhcoh4uxe8
iatU7UDv+2fWKN8VacM4ucCP8f1UY6N9K59BD4AZAq3wOTL5wsHHkB9KzbfcXXDa0ptnZXb/8r4e
LWvwapUAe9kuhMNrKORB59Zmtsrqk9edRNsKcem5+PbLq9XctVXYeXF8UGw7etthbfPBT+VrrTu7
F6pzVlfxlJdp7wIJCUMBpFkfyq5UH8hagSgQkvUTO8hIVCmZPexu+PsN8TMIHASYJRdaoLxunrM7
pD0TUzfvTQWYNb7aeCdb5HPTzizmCFN7+Rv0bz9NqbJNYISJmMHo+G67SJ1aeDCybrPajJVVo9dp
VwKtvoXQhOkVoz2DbLPLe8TPPz7CjQj+0djkhkC97Ka4VN0Fdtmnh3NfnwGBxBnzzopHkP4yGRbS
BSiHY7eW2FFcripYrw1ncRcI5P/5nKo64OJIeie6cutn6c2qkrgx/jmGqJ6zfmfl3gGh0r+utBTx
d9H53ZlbIYnDH2q6YeRNypUVyHQci5ShS9Eb+48JcwFzrE/HWU+R3TrHDmIq+5d9V4frUYDaT8/6
oMXc+kgvhsYk8x0z8yPKYkLFR2LiEVhAMQWeQeQjiJUWqVbvonbIHxa7jF7JxnyJhST3ynIzIy+x
A6xe4C1PFNOhR/MZT3GlfQa0T6qcZh10yW7BNNdT43ihLlT+iTERp60ObWJ7pLjPuAZ/b2GXmjAO
BxQkLIbSO3OWTXQrKjuVfmZc0H6E84nrId3LnAvVxYSjDFB1bOGfRrNBeLgTqpaSccmpM/sn8R2B
9kAhnDcs58jGg8Her2uqCRnHvT3VidUhaNP4IP00N++ZcesU7CFoXZqdimmXYdEPyii+C7Jp5Gog
DcguhjlHMoLqJ8t/uW+PN7eZXh4pMpzAvcOUdYbSez7A8H03g/22iqIS2C4nXpbCZ3B4HetgdLTc
3CjwxsYIZdcUvrownISJUZCyCuBFKqG+YEx3w+u4dZmqcrs9DRNe31VEGjZi9h63nhAvBCCD7G/J
VH4jh+JMpN0OetzL34UkBg14CtrIbxpvStpClz+ROd5fZYwjtCCc/xWLzRr7dA9y9P128fMudjAZ
Te9G1Q6X6qKeB4Td+jVjHZUpwxlKIlbDKIzcCs4yrj+xTd6mj2+pq1KecUZ16ylW6t7qRlC2kyrd
lQL3YSF04eE2j/KDHGV06igo8KU980O9BtRA/HWkpKDxRvoo/HInmexMDtmTGYD7deQDmLQTw04d
NAcah+pDq/2FQy1zdF6I/NnUF1fhl5iKsKMpfqnttLmxo0g6GzVq7lrDUVOJomrwILT2d7GXSE56
V0uRvNlsqw1Phwc+fKKVyX2z2YwHuqAZ3hEFQYULt7ijWPazHHfOS5EKRCXUbUB0IJE0ZV5CLc8s
AsoVA2b3tzBAu2O3/k1E5DW3lpxs4rwsjQOnQu85AG39rJ23xE+4wOBwV3bjOAzuRZT62/t6sR53
I5uEml2fQ6WQERryahY2SCIxK9fQCxSgS75hr/22sFJMZpY9kkF6NCaeMwLfgfflagj3DG/yZPNZ
IrBQChOfgzWbDz9TO553tag+FESfLTYGEqA+kaA5QllSMLMTJ2VH+r+s2pezrg8mGtCIaK33WMph
i426qp3N1qGasAG3yJQi/595SLBmrti3W4X0J5neNn919mVWvStOhkuayK3GA4spNyKDvEX3GtOb
sIJgom4Sd7Zu/AAahyeHs+MzvJsphqAUqfkPLom/2hfKhYxSc2c6wstTkonbCQUyBKOUEarVsOT4
DOX5TAIl8OBd3PetasDz7bY/emG8VMW9JOZLVYrmTpTyblL3dEfeOITingoupLijVYlFI2WWVSRx
oxHUnHOzES8gW+XTTKjgGgVG4N08dcia5Xf6EUjEXTKvibGmLkQUlsGtXXHxO6yigxZ2rmsxUzV8
8SSxsetCIxjKx2ovcBq1zKvsxI72XXqs3cYbsH+9HhlOTXWcJ6BqKm8p/vcq2TTX/ZN3nrDoUEYd
UkMADIhF2eV6z3zdOCT8BDBw4Wq0gzW8ZA3CmXmQICrju1z/U5sXScunzz23BHCtE09yXkRwqjQI
TWGf9mQthjZ8n6uradWc5f61p9E3/ttZhlyfxUYrnQImiMtG66MmkERvjm0h0eNdA2pNWZUGIEzx
NObLIqtjERkcC4ZefbchyUi0OPQ7xMKmQ8bbscHH38VJuBb/7a92Uh9Adbf1+v4ttCvVjqQaFhwZ
DKGGUxXHLTqcYKWKxfVORF7ymwM68MwEPzfLtxR2flcC4BIECCn4PKp3ob5rsYCVPcDX9hnBHHkq
4O5Xx5av+tT16oI2v5aWYz/DTzA82qd4iV9ev1zDoIFWX77yIlycPoyotGMFnrThukUjjwqJ8EJI
vBga5OEJf82ai6B6XlEfJPXB5YCHvqBw7p4ri3Xe3Qp3vh3fpYbq9qLilUwcf18OBPeFpVVfx4Xl
6By/PZFe4NHZms7bcmZLAna5xp2BoXQuweQMIbM3pzMBUvsYfUUTwJ6zmbUylQHAb8oVTcxgyg+M
Sw4o9zJ4h93hIBGs35f/+196AqK6vY2bn7pfGELJfy/N5aQ20bLRfuAXQy9ZqZin3uMr17TMfi4k
tZIdZPXEvpZU5OA+4PudeTsTMXhjpcg/CBwNaG3CsOhobJl2cRsHcpNGSev2V0/2d1f1uB9n7XTs
ddD2WmlgohJp2ZdTMrk+VDUWkg5nVy8PKVlYXYojuFPTOL9fvx0kSx/p4z9xcKIUJ+0K05v4+f9r
pUoN1Bgu0qyRTCCJps4OUWnQuth20T/QkW3iKuRkoRo6PO4Rz3esNoiKef2vlV0KwxXSmXeZPOkt
sJ4eUF8ZgQynMtPppMOpWaYlScIcQGdbqS+yBn+k6uy/WFhEgULM9nzhWdgmi1VW5leM39Ie0Iq4
6l3gtOjGgEHtS7u5u2l406aYZxizhYBaw+fxcsVps5T+mysv9Lst4WZW6k/OB8mR77wicmw8Xdy3
4waf5Aub7zCuQtOOXMEI9IkzlNX8V83nY6bFBvejftM3adj0uX8RMs1LCIN+KA6+cKSxE6u2U8Rn
QL+L7TPFpt/uHzl2T/nfVS4QDM0b1j3gY0ErxuhjR2FWuC/Y6/KuQMpvb9Fxs1o4ImnQj+zuciUX
uy1Oll4/9Rthck0bfBIGArZIcQQ9yFOvahZkG78i/ErMAi//gBh67tSrpTtFz9Xjm7b//vEDTKnV
XP4zMzIaq8OODqCGqGbRm5V90mLBL5IF7EXFDtzd35PCe0q6RPRx9933XMOS97f5BUR8Sepcet4L
/R0MpYeTw2Yf5/bObZDr+GzLGr3lo4niA1QJVzfiUIVHHk2riuFJt2LkRorIbDGzSJ18dhMb0fkO
ME9ZDCEqs/3J3HCbJEkxIUZ6NH4k7djsLIM778b+4kuTP/lh8/XmcqvTxf8tIqVpVnIzTCqN7cq5
03rM+ncGk/OWAMrB0FKdQ03a2Hs2FgXjgwwi2YTIYZ5cYDkrcFI8BDtUhZiSX8I48L27hI4cpmYz
weN6Fy5bUN+atJ8s05YGJyOPLfl6U8yP7bFj4IOQ6CkJb6IvLZMhwQNilTGRcrdPkO2RPGPFHfKD
K6kuIsqZYtSC4mZuRrDYiIjLSeePJcg1Dfk0FedU8gSu5/RvUjFuFtLhGG+heozr72/fV20HKNWy
m8bFb55U984DLfXwtZ5D0M4gwlOBUgU33werZ+c3X3rJC6vPXg0Hg1jxkns2KXpaCuhZQtKDeMsi
niMKPWgZzuTfUUvIAiKTiPS4R0cWieX0OyIIGDh2fHaFt02cVoAc2bFtgVMLLtsfUOC7d2BPz3V0
gFDdiXNhfrco99V2Bm34f7fBFbWX5HK/ka0C70l6XkJ9Szhos2vzMMiY9+Hz/pZr72XBlceBkGeW
g+j97uVmCtG6Gmh1TGgxcnKrP8L4BvfkWw3gtax3/KpAT7+LwaixzS8trufG0BN7eSZWlhMADauL
BxVr/roZQ3xC61L1VrmrJaSfmHLPG/wOVTvc5POIl+RGtBS7SB2Ctvpq8bLS3dNbPWvHF3THmMKi
rFf3A59q9QK9OA3LVS9c7Ajellr925G4agqTdfoQKYAGdxSqpIgLncZYbzzYBxvyffy8AGczUypJ
DdmQt6ymvJsCYOwVUdgwKeOwtLLzG+3R813l6CcSmFS2tp2q783Xww1fde3vitpMtJNZhT6RT3fF
Nk0URjv3TOczBEN64xLC2C1hGpFIr2Jh0uHmU1bTAbcBqcZCBwWZWP60MZnHRDKivDqYWsyxHuan
X7Bu8xJuO65J/rjEOstpjfV+r1Q//FaIphmKah0A4y7ev2KR22shO9584C+XavQokPz/soemCsat
cUpkU3W3lHiMKVWvlQnu5ghNtIo6FNt6kWARDLNI0nSzPZea095We31sQgttNTSgl9lLg6n/GKFG
lFk8Q7jGk6492PvvUvwhof40AcksSK4ZOlCg38c3qB9AFa6PulV0NUuJmzVZpZGI0GzaAq8p+9qx
RV2xMgJUpxWzInRy5yxR1LU2AlBYVxuMNCr9ajMZhyinJoQDyz3KpZOQHguqfgtf+ExdJER3K/en
YMoJN7R4ZO7IVjZfhmoicSVmJCswj7i78NWz2fTeesp2S/tcvviq310gtJNgo5xkqHlfcwPGKkYW
D1DRaYFs1Bo2s+N0nKBN5oIQ7ZUwvrpBlKPpVADjbUJ1rlVoMOMUsKaSK4XLJJpL9jMKOoAfR7PY
cpUi5VkFIiy9g0s+YSXpSIPB4UIlAK3qA2C7+fZ2pyMhI1xKz0wsKgGnibIfneT1FuM5zU4VlFuT
UceJXZjuHE89JipWN2iT6fn0XIu5sk96s9b5CXDDMuFZ+w4+B/2EjWyz/rSP7bfKesXluHxz6Q2W
hAZ2PhJNOOsh6m3SOOWDwtWhL8IIV5JQ6awjmzcx2LajGoYDVpHth0VgSNAwZBDLdIJIjJKyTf1u
tAzYxrwzp7fLP8qiNsePOCtv7oFCWV0XdLLR7wzJpZCQITadAmyr7pnUSlaeoCNxv0IIlE98hm+H
Ac/WPDewOt2Z4hDdYfv5sexwOdSl0gxmqB/xC2xaeN5OyYRuLLHHCktk1K8Za6LTiGo45tKbyjRN
w1shQZ6w69iZoe6ZwneS+OOfOphloah3mhkXt3E/T43S7r91ZBJ3YXemSfYrJpflZX4DlWy16+DB
mvCx9DEYRdzWFw3hyUnOdDDcbwfc/yBnC+Re83gDRqcsSqi5XfPndC72CcagHoGn6Bs7fBP88Rlq
dERe9W/YScwwMnanyOIso4cx0/cl+goiP75u4wXkn7aR5B5yPD2V7AMXliLeZmE71Zuj5QgPoNXT
JXBifnkeCqiU6QW9IdChYFsaAys3LEMDmoFfWpojvrrUs3d50jRTHSgeRaGic8yZLNuhUTPj3tFP
iUTBaE9QYKLJ0juC0hy9DdQ0PJxwwmbIIxie22hOA7L6zeLg3JHdckofqSbuQMq43i/2kdf2d5OO
JdbUFzEySsvWHBJZ/xwWafs1hF72Fg70yrZUnu269Zz/4iQhy6hV8FkW1aLc9rOo12UzrFkXyvrX
tbvoIwOMjuivPumY520dS8tLXB4BpKZe47+zkd7bDiMcGpZYEamNW7ZnffgxrunPXh5s08HVug0r
zqWpY+no/9lY28bnevwV/OJu/xAswdhgr9WCCvXo+mBEDzy66GQhXby5n/AlhRbJ3TakOT1/VmQ/
kTgl3PxZmMoFKJVU5agYMFC+x6LKo/26k5Mpcwg2NcqBinxsHgki+sxw0gLdz+9UdQ2lWz/utjqV
ys3hpbX5Yyl42GhJifnbHEYbEunYoh2tAYYdzMH9eapYFg2U7VK6ImIevcR0TbPXH7xQYsZmZW9q
8xkQxLdnKxmbM0AtIbtuUbM0oxV3U7R/WJHHsK2BKvR8f92ZEBYMIw8+6wzOfedWUTfTxu0Uj9Pl
2RFBBeLTGZHum3ZMESUMnv2U74fOpL18oG2Xht0JPp/W4BjKHw62tt9BafzbwWcgGPohu7MCWwYJ
4sOwyVmOwfNTPq7dLxnhWOQ7e5ZIC5NESmyvJ3wZgV9ZtlmQwNCZHhCs5lGYblAYBEiBLjuK8oUl
ptHmUxHNPIcMsG4DWfzYGz5qpoFjYHE+n0rl8UqpJ+nGdOPJriWlHJ3rWwDDe5sz5I0N+HHZzqhs
gnWLayMI6g5Bowzmwgu64iQ5Uq4DjrpbuLA7rWm4a4bv5GbskmWbznFVfnwsuid3A2kXqldNR0cM
/kZNAE/2OwgaBr5KGk8FrgycfeHmrtX0IIufUPAJ7V+92Hv4J91tW69RsUSdzGnp0bhkvrDodqfU
m1XoBcyPZd8emVsAuK2tzQqwlqiVREeDVFO47xGBERolxuH0jMMCJ5qN9si5dRdDnItya7C2dnga
D2XCazOIayELTqL3Chr0snZhsHkEdkVTY5BMuYY6XBiiq0Nj/YDIDP1TxDg++Bt5cqq6Tc+QpI+f
TLvx1xqH5JB9O/V+ZhTObzSW94zXvs7qREEydeQTRfo9+63TsJI5bNYGB1a0so5bUAVBokMHelbm
quJIaYd/ZxMqhCmrSPDBpAf//e0me4uryHL82ffEBMSq4pyZ4MmvSms+DgmOSPrJ7tPA7ElMGIEe
+2yDRga3cBsM0rUqqpAmGTuEBxpA/P01jqf502lwiRRLQIy8jwLKniuTeLdLnhnFRzdqkIDwO8Mz
9VyEEXlJMQ3yDS/ZhAzwcm9pRgzljKk/hCEpleqcsEk4H9LAoIWxPyBRTTs/8ftEuCMb/9WyQUmY
H/HCG/Dj2PkhWCTTZ2nWKw4BlnSkuTE4N56EP2GU0uHNdTl4Z+jKP1x+AbxHUzY2GkbHxdCEdHuB
avK+4gB62UE8gxgu9PEw4YtbgkqRdA75WuaevG1l8cOl5AU9wPKmu+vhk3vL0jN+SMAkzVQ3Uo0E
eIBOAUKnyInQAI/335J7E2ypYUV8QloJkH1OJbFPj99CtzltBL2v/FzuYnSWfR6/C2Dp5pupUv0w
rzO8qHaFeHYSIzNmbGgNXY+tGV42E6Hg0PWEAym6H+GLsQF7l4eBaa4qpbQLrbWhIaZDQE6LlULE
CJTk8tvRigxC4dkmU0K6JQDGAyw8b3eOGWkELJFsXUS5qB5hvz6Jkuc3nwPmWos0XmtrN/PjPxwu
pNcesNSLohOZORC9USFe3AEpb2c8vGp4zr6u4jh1D6DcNttzaO5GmadFs8QGit3GxR4EDj3oQtpm
4mVCE0fIEC5IG7cIZn4HhJjU0tWMsh/Y/AqnfzfpKk4L2JgO6tpEnXflfFrps5x1OV/a/GQK8Bsb
flDPrYw//zmey2qPo4GCwGfAbwuq7UmaQP+BcZfvAvIwHQf4CwQisF0VOhgPogMQUq8datqZcCQF
wgXcRpkFhekJTn2hl03JUWxqwR2QrsNZS4Tv3Y1dpro/xjTraws/eUgtfWJo7mg/QrV1tjTzM/jF
uwCyNDh30g42cZj1iyyGvcEo4Y5ZSeok9QdlRDk5bcu8e9WmJuZeDMKPkKCyIS8TipuizfJ8gooE
xSmnu/pA3TUzsoT/DOJN6+U29Rv3DUFFujuEFBK6zMrE7V/Id/T9FGSkh28AMN3NX7FXMXji+VWT
u0oezNfQX+ZUwaKIzrgpn231ivLcAkR43/6TRD4rU8hHHJh6vSlVCAJqZpMge4ybxkSOfQfyE1FH
z6yeoHHKTbI61hlYowsKcR8R1k8bYGwheyidtK/owAWLE4AtIeTMV9qH1Ainz3N6Y4gaWAudiTSI
Efb5Tb1zZq3s2DtgnbRN95sh3gDh3fm4/H1nV7UDnB7WohuclfBwxjJ4H1/ot6kMXRSkLzEOsokj
r4I7ggTrKPpOn2Id5f115p71xT179vmMYEW5tMCjtmj1Y8A/65uhVuQRKFSm7f/Zm9XtsrUXm68R
gRE+eLyX2l/a1kQJm0vHcJygmm3zAOLYv69orec8fS7SIW+n0pdtinBMreNw3SO6QMFNiZMLHsnC
4Pio3dIJfZDjfjeFE52HBTJNe1GX/LqXdOutUQte5MWOWvdz8KlHkq44ucZHagdkXOWfkt5z7OXp
YdD+hiK+otnySgmkLdZZyrK0I53HkoR4XkyHK0jVJOZ8YdAQy7ioGp4hKxyiUbrUzGFSEM0MpMns
xrT7PqXAlP19mV/aGZHnEXwzehVd18lzDccOAAlqWA+jDvHOSeZuPu1MEQ1sKJLsJYbP/GaWZjlo
20rwq4RnkgQ/rQAIBq1NJhE0zAmlPdiemMEmu/e0yJ6GPTW4ANGlmuOrWgeWlKpLY4py9Cc5DnWd
mieFNztsZOw1TNy2JzkDPzf6oU3458SXfNrBP/TG0vllHNqEMWWhAn/4/LanSvGhSHX7pAcImA6T
7lTMKJnSDHofgfDYu4TFKbdN1h1ZGX0TKOeOVdfGiodGTMLGUk4rNRNLifYexHCwMtmEjJE2of82
dEjqpgt2qRCc7KrnYsAbSYw6IYBqenXGmdKlmOUkKjAxRey0wO98C/hdikvnfKV4o5iUfVEfkb8o
PwRLKeJBXbEgF6D6mUNbq+ti5YZQszpPPVWHzFyyDo+B7utZr7tRDQYQXXAftm4LfPuxBAhrE2oX
cm1YMH58qEWwJpKRD2VkYIpJecuTzRg+6b1qVB1a7HPJzxDwthoTkOI13McncikP2DAShZDodx10
BXrUChncdgAbF1ukoC22fbU98pEf349cjS6VlKopHrsGUdXJk4mHC+3qdiV1zRBVCBVjJRFgjcWj
a9106Mhqt1zUtpAN4NFyQQtwKENPm1PilmCXDeaeaXTFoKGYZTEPhBH1RihyWqYzdiCzrDpyiad3
LsEEGYdaSwpLfKuN5h10bVYnzhK12TxEpP6kZrqTiymZ+5BMOvAUFfJnm1xiDWHMhRlPwBAWtQh+
6af+SmYHEMF6r//yzzhk+dtmgOwOWGZghfPSPxR50UmTlHhTHuanmXn+VFGTKdWVr7vZfBB4stTa
izH21lQPj58AqYwsdE5y9PFpHGnrPGaxCMh9jvH51zFYPOGDtUpTVh6VqT2LwQX0NW+L0zau58RL
WNELHysgXFj+/MA961m9fnTREJZeCEcMCiXeTr0QFa7PSLSg0fWcmbqkHX/qSWQ7sr9WBqW10uOP
l9uBPiYBSHuYWUm2Wii1o2DAEUzYWeqfvwjX/YaiFWbtffw89E3CxskGhNCN69gl0LRPsZKM0PGq
Wa2QHcFu465gxeE4S38Da31G0gmndBNHrpI6ZkwzHUq17a8vakFOiVbDwbSUUXpf38XMpvM5PkWE
DNlm2NbW02fI1uoSNX0KrPNP+PMzCQkvaGH3B92PJUp/dIKcqZ//QftDl6XASuBeu+4BVZ16E2Dc
tqrNUh98OfSLfB6WEwpX11pr9dJhxqNbiczPp5Bj42OnOls11+xFizcb+kOPExuyWUX381lHPxzj
mr4o5k10GsFCqb4xcQpn0UjkM/amrIdTTMio+xcjNIZlGp056VC/dh5LE9d/IiYjy0agww6JzApQ
O+u9/9QceAtYcXMLlGF+t993DK6kp/N1DC5kOkD2BjAsSrcaQF9xwYkKCAqMWPe3mSMe5m3SUgA1
mn4lGC/EOfKbz97G2e1HPI00/mUEkkVe2suvLCES3FFLmb2id/qQGxHT9au6JYqp6/btpRhDKMrA
V21j1Twluk61vH0UCJ6PZceBNdRyy+Hui6hO0uVlGo8fJW+RCiNpSjeE2lTdlHxfCJjgNUerscpq
hSyHXMaxavDoaS5UZT9aHLurKQ2IF2C2lQSS6tejPo0iMv3+vetwgiq2YYrbRl0p7usnF958qwvy
RnL0UkZaai9JWENxKUy7WHvdbLxRybVVVl9xPe5t/iLt513HrO9b1PBkj8h5xbtTVsy/LLZelloW
XdBiRPaWW6toCO3Yzs6SrJD1DebLw+jobTMsUaCepvxVjsXAUUogsVZpzEK1/QfqsHV4ENbNY+wz
JjY/tbN5I0rDNOTI8yd/v1kF4DZ0+ULpzIKAFdwWjWR/14EA05MvPa76sHa65gZGHk0iHjmsi7mc
PQHziKWccP9JqByk7Ma0FtqeZ2akWFe2/Y+yqR5LLxYhkrTkylasnn5jcmq9t6vrisR/ZYTRJ2Vu
T2IAcISaF1hYfg7X6z1qyqp5G3TqOpvgOPEAqCbp/fR99WyR+zRCiEPKUis8wO+dJg53ZoiNBCK7
utDmVScBh2kdlR9ut6azLItyGXbKiI/zii2DctzTksYsb+9t3v2ak/B7rrW2ZSCinCBnYdyH7rMP
ctP+sBrqVHTOUX8CR21x93Aguu6NKIstmoND0CGCObqRO/qSoeWikD27WuoKwOXzYb+QTug1ijps
prTG9v0ELAepW9d/CPvFaWiaJAtlWQ4qOHIbbwUXBLW8wCz5nX1BQndbGF+8an8G4xh2tzyVCfbh
qGW4m17xorpjziugfymjkqbH+nHyD7loCjEqHkv7XmcFRh8WD+n1zcB2upjVYjfj21CFF2651izE
acwpE9GIfmnFYOSPy6lklho4zwGi1eyOpx02XV4dkdH/te8nQr50KGZuKQhvU05ti6snIaf8qYBy
BPRzHjmUsJlqOK8vFZBgV0Sdlq6cbfddBBShM3rA01x+h9Ql4iDglmix2JPtuKOWuQ4YutGW/YMR
MdRktF00giQs6ZItGHRvcVtk15mjiJSQFYMMdjK3UjiBW50m0iUxM91aRG/h3UHp8AYmQN9Bnmcl
/N3CoqAfVf4SDkClD3Qz66KMD1h41OVz0gV/xRYxN/szmMVgbR3KPTDIQtM9xmx2JYUp7WRKmBWk
irfzU6jCkAzcY3o9g9dcq3yhB2rK7LOaGJE99CiwLMy5CHIvDSBxmjlV9bZ8LNLTudPtDK7nwhh1
7E/5iCoffm2CKsHuFfQavCOjftxE0lt6r0bHLt4MAlJRkIW6i95YjJGAzd3ziH6A46zPqI4bUqDD
zhHxkyfeakhyV1C5P3iVaD9NRvuSFt0ELIo697gd/ywc5oLRFoCs02MTrIpGh9X4hxt6CWizqWza
3pmsc1LnFQ4M0FdtE4aVOXNN56BIk+vqaPKv78WSAfQrKAsEK8CtxJbSqk8pyq4GDhsWe76WmoKi
zSCijBV/dguR60JSgoR4PsQG00l79S/GjzLhE2akf6LOFcxx7B1d4OzwRz3W/PKwp06bkLDzEVbJ
jlviTch+nsC7wWl6YM9FYQniV+Utn93XHl5mCBCbeZz+MouwX7fSFwss+rLJVcfveRH8PblmiaGQ
+gtml6UwZsBsA4rsU0tynrvOYvZmAnOCuOD1XHGnPBqibknohaql/mQGdmLm8+11z7eddydxVZ52
/Yq8JNY5xTRDveOEsMEGhv0DGqiTxEiEsGEMwpYHqLPLQefjMPv6vaFHG4dfSgGvKK63VMoKmErS
hUu7mT8ndOUKXc2GkLtOppY3b5qPRdTM6Nw1YS95hDrCWCKpDFZjRyZlBCartUHiwD2XZMTE1+KH
NrfQq67FuHoSRAvzdc3m36yFN2R3KC3epB9uAB35Fa7Uwt6JQu1D+Dq1PykvDu1ehq3iQrCJ0rpe
I7WsU0nDd+CV91opUU9z/zwku3U6wyUeDplqXLEH7WS2loBds7t4q8CqpqgWaTcGx2DWsV5UdyVA
Uj6W02YA/N0amWUdsF9136CUGnNFNa8rnuLnYeUkFYzxoBXZ0iDOrNTIcUSOtgrWGLhxEjCSeNA8
tiMOwpoffcc3ocpXvQlfM26Xz2frpfVz46moOVLzntm6u0fSxWlUktHP2GXW9fNP3K8IUA0XfVZV
+VrsYscx8QPe9wmI0OkU9GFDXNSx0JxRxtXIliQoF4Matvlk4txQzILCczKG2h7kYn8jJmQFzoAO
qlYacmOeCo2RbSZCamv/FeAsIhMf1TQXUxKpXMLr8nnH7Etml/Hkn79SItXrBbaplB9dPreXlBcr
49Lca1hYS4xwPLrQAnz63Wmuw6/bWiQ6mS0eRkiHPtyFdxKSwde+M5pMZHTycyO7WA1/Dxo3Clh8
MWYiSqiNVXaS3zHj3FfU0Nosr16VRC5nbvDuVTviYPylKHaa4rWJvXoxOFP8b7hOVDUH3D69u4Z9
vgD2jhDo/mko2yP4pHyasoeYqQOiCWfbmLIilLR0JbCAj9GX01CgsdiqbDzI0E+7vVCQHYbt6l5R
rB14w4PXwnHtGeEbb2vF24xSx1SKA8Baeb01OmDFjeq9XZutomfxf/aBe58regBSO5SNvmdHVk3J
PIpMejP3linkCfGSKT0Tsco/kXVIIbiQo1ftkJB9gPw301Iu9yoM0knpYctcfblJdFHd2quorfU8
WxNuJZjvxUpbWl1VxNurMBXp34QyrUMqxlLGX36F+XZTBhaane2rxGWDYNNneXnbSB8IBdXyU+Jg
/XyNejXHRfFGk9PNAF42mxdv1pbR9/MEjmWdqwXk9AegRaNk70TWyqGCqn2m3BcvHrJMbOy30dz9
P0RaPehpn6gFgnAmvF5AhCCYqPWN87oT0HzbVSYstnZJrH9JEirFgsemW2qx0jM323jCeFnQwNBt
UY8wjI9E4My2/SgKytge8WYWCJDwoPzx1TuxQBdODKkCyI88AqekxClUpJuoVOOYe+5TKheOqp8z
DPc+kPx8B0M4a+TCXTth2bmL/a9yfyKDBI1Omh4irB0ZXZvmaqeZltif2XQU1Yg0xWfc3quYQmEN
Yrnp08HvefAZ1Y3VcbC6OP8xNttF3wu+HlUcn0Wn6FJStk7hhkcIKS8vKWjEsQPZc/gWhkhZ97/0
96JiA8d/qHimZPCKj1qGlnNjAo4GQfGf2PW3EdZaDWyVzAZOJYg9Nj03hdHOUaoorPwphzrkHJvO
DJdeWuOGEErFQx8FfEUYeQt1jc7NZ8autn5KNw8I/SJY7spdsywr2ffc8bApIZOPC/t4zm2BGmuf
Knnn15owO022S0utRAo8o1zHTPzg9T/Fk9sc6AQA4D7URYdn/vgKqJL09fhM0+B27zJ2SYy+F4Y0
wrnT1QR5yFDYgkAUbsOv596eBQc2z6L0/22RRkZdnK7amnRM4hWyKqZjde++H9znheeTuGFXdEgr
vE5BzoQYarqHEUY4eQAKL4e+HtYM2LLmRgHaDYCwxY47TVIIiJyTw1xygOvKHiR+rnMh1KrdAalG
x8ttfmJ2mNg7F2RoZ0O/Sh5EhpUyvSuyySE7ks+bl8uVJAN/RfArPyvGm8JDFiV2U09p8YvRO1el
N4427CN6iQZiz8Wi0bbmLMlzLu0XniDNJYcxWdHg37tXYFHUJrx7gzdg4lyncmpaHFIdEtpJft6w
nmdfC/y+WDYPfezl2BpGipmFMNNRiqlkdiLj+FwwAblTJFA+8fwDaETXtqqNC7qtKglcNnGjRgwU
D5hXxDqtiLTNnDaN7qvvA7RcB1rckZiEksksPbUe7fwk5qFbDamI4E18r+yZtJWu5hNmfTuTYCVC
Z2auuMCtiutx0FScHcdmM73WpL5pqv1OZSkSPBpPySwDCl92wU6+pVY7OHTO94zpLigkgQKucu8X
vcwb9ZGN1BeZ56Rwojgx1EqmWKb844pvI4UrvP6OdKUPgBYz6Mz1yFTC58UFvMFOLTJ/UGnOtmXL
npu9BAX/QCJUESL/jp7+ThVo05Sq8YkCn2jOUER+G2W3/MuVWtIijKB91wRv4vDnuwzhD6edUoZX
u5Md3T3eOS5gCDig1deE7a/O3PfEeupikU3PyWY9+wXHBgNwedQ7JxfpFYV53lQSKnoYPKRFNhxb
Q/NwV40+R2DdiUTW+IIAov0/WWVGDzOZCC+HHaAcEkBUuQbJeODLH2R++bavXlR0piFj7BiIb56r
qMxZHUtMAM5/LEytTNtiO+3lSIT+FKS088f+wkKNIGixiPp4JFsjLdoflchan/PH5OQBE6FsRW2M
bET44K3ym4b0wcS6cm96IHmaAiTvrz71EElDD/yVOhaPgsB12Wgz9vPCaGmoH62idr3ywyT+8E/F
QctzBW10xUCzP+3qeFZSM2v7+6cSpRiJGPWbEJrZapdg/qGcfZFLd9BeZbRSwJoA+aX1KOV7gy7O
8hob6eooQU1JVY4VqS+xyOnorQAtCeH7sI/ymFG2RAhQmR906o44rkCfG0+T5KO9JtMjkVorr9HJ
/jcQwHrCDXPK2ElSa+3jJpSYZT39xMrstNG6EYDbSUQOjMhcMuEuBxXdhH5FcrJf2S+4S/BkfKcf
XaRRPUWxfUHq4ampgX2m1YYzO0JP3ZowDl23HnSTulR4yG1G04YohFl+lo6W/J9QfmMKmiFvDBxI
Y/4h0GAMGQXY7UNTOk8CCdKBUuoqC2J0WOSGm4koOACJSt/15pxlUHm/c2jjR9YG+XyKo8IzQGku
+U9g2574kBjYk4RqN0mqNd4JVlX99JvIl3g8hQzG3x5dyxtdZphaWWxV6L8CBu9jzyYY9RlqJBdr
flLESCj4NpoPHwFaLK75qw0cvHJ0p1A1BEhtxtquj2c/zuLpY2mBYT0YoR3FtTKZl6XW0crT8LoW
xu1nHPH3jXshEzpec0cxLvNLP9bzCIQOCsIOPZU5NC2ot/w77pxIkfLaBgjku0mew7P+ouR+ZAka
5MJj2M4TYPoiz9oynjqOn9Pg1/chbrChQNMeku0UWbRh/RnTK/EnWuiXUM8bBjt7lwhBbvxjnTm4
pujAuobXEBfTsMSLON3oiGkvX4PO8K4sP2DZ6qakthSd6h09dF9L3iKgwoDHGURSKOh297Exd0Gq
ZA8PBnaC1ePTxUcbdzjVMuM1uB5B+rPf7I7EEeJZAEch/N5WL+Y/waC6e0b7wJe1pv/NZkjsYpoW
fIK1uw4wDPeDmzUVkkeFO2CJcq7aBgIFfCoVVdNvLm8fu9cnPrTFqUFPLyQWc8Cm3zDNiIxSVF3O
/kBl7ULvO6PHMkST++8sr3zg4W/1PYVi+qCWEFBIIKPrvy4NCwSKujPnMcOdmOYxhYiAY6Yl8Dhu
L6UNfizQrcWFhoL4FqKn+zm3GSBRvUDDySUPkk5bl2NBnGaEdQxtbYeONfOi7tbFLeyEq8m8ru5K
ZxM3w8hT0Qie5j+1QkUILcVgVzbe0eDarUgoQU6cbQ6H1hMm8i7zwYTU2bpJI1WrIwmSCEAS5jpg
7tqirLNsxNxAFsp7I5qlKQTXYeJq0RFOqf8m1OuvyTU8fRtCrz1/eZYfjtV1RkVoUw+/S5c3yXlg
JqgGt1rhlQqGRxNreLJTde55GfjoTLZfQqjsB/jpfi7I9q9JVRZcpcFIoZ9nHVBbfQeWa3f4dWBj
FARJYOaWiAVWNenQaqQJT6UTH8QKyfVL50Wrn8yt3lgmItCc2XZfkD6z/Sybf4XFCPwBb6QpUlc4
MldWHtW1P1U9GYmHwaCB38sgNzJeuJpuXbgA9Wa41SwFhGTAWRAenwx6bG+xRVfWeOSa1rZ/Pr4B
GtbIrIA4DQ9EcY19fDmToFQCS4DOEiOHhQQ9klmSGcu6mWn6oW3iKrfhaSCHNdNeYa7hxDM3p2eS
1Awcyn+Sm3Fyf1jEq4NlyJRDkk9EY1RIsjisY4n23y2bvIuAsWkhBUC5gD1D1EpJfdlfM2ft12D8
iNTDrvE3aqpew6zIBdSF22bj56jnkDeHH0J14jTtjDjvtu9Mmxnnk5nZJdUutUigwpEkJ9XS9G/1
mpyY12vf18xzjRmfISDlj9dXiPWaS4+3AP/gMg1ZrzSMIpAfPRnDLo9QXSNY10HB54Ry36B7i6Rg
qJfS0Ylo++BzswIaf6fsXbBY89yMsv2zBw7UktPUbqmJf1yfwrOrgjG5bllLiY9w/p8qKqY7kcA1
o4TxxDdF5yp6JfL6mtotogBn5IZloucF8dvzc9GiDpomP+YEpXROWFBf1J4gERNN+6jXBqYHZqNh
1I4j5V/hvJV+PO1e2O0PM0Ai01zClUBV/oZFkSfW+57h5mXxPnjBuw4r4Gkv+uB8wF2y6/Zw0+nQ
yq5GUzaBy//UeaTKjgDHM8JyRnvcn62edTGfH5eaaybH6kVgiCuxm7NaNV2Kfiof+3HSJMNXRY4A
8EHt9QVh8SpMbMUYlrm+zMeRi/M6sKzNiKZx2/qia2HxhvgkQByJ3aLIlHJymcJk922s3izMaEgy
NjyHH9qprlkCkSOTYWHP+9WniXSn3BnhzGnf3xUhPRJBVyPySTE8t4FKKPBrdzO7FIr/DwnIqqM/
TKMczqm1tBranPJTwdC0peJmtvvEUrQ13oPoEPBlPIWUw5YapXOIJemlCptcMCV4WYMY6EG9WhzJ
QAWLwtQlRU6yQ7Dm1HIhrWSnqzpJkX/TwCg5wzN07XHkIjPh0W9FwcpdgFjLQW3PeCO9852OS6hr
uwYJXqnfKpk3EiF3oqdDr6yytzoENlJuCifSnjKRfxecZxg9XDysUMheUZ2l7Tj8jJeA4VIOgoME
flLEkY7i0u+vs+iwtvrCB7NlYqKK4Gv6ZQyEFy3cV1E/x2fnKFWkAcHYDVleswsNqTCJoXCs3rmg
BwpyD8QvYODur481VrcQJQZLrwbAElAgjVcFiQMC/kPSK9gPOiTLnDTKAq+R3jbFX9IvgYqO7J4h
LEu8VBGSvi77619bZrRiH9FgCzChePf6nPkiTd0dm/tZv5uysXsvOgnrCwMn49L7P6YrA0B951x6
gFP630zpCmklBD3Dg/DYdCwksbU38kl0e6YekQ8cHkcTghQGxCvaMZPnjo8K1wkOdDj+C+1HRDoc
qbpfgwA3gZ643tT8E6VvRKhFzrbegMiR2NjpgARLW+9kcYFz8Zkr2TT3bKLtUTV/3/V0RhJid8cO
Cb1P8q8NEGbuTTomfl5378uzipZML53uff+a+5wBeOO0ACNAuAqjszIFlMgI5MfPjC5vtqidmcWu
WxUUgucBylOq9Bnp5Xqhf11PupZDS94UxfoF3cs42UQiDrZy7kjxhTrgqb1WaURaSBe1/73iaG/0
0iU6krblOwMbfcjsGNHYXYAoeFNld/CRWidX5JP22IdjLYZ0huZbyaK2ennzCIBN1QltTFIQdcKR
KeXgie30ffKAt38EX/ckZNfnCIRBqnh9+/56Ph+GMZIXCf08OLCpj1AwLthA0EnryzMWak81hngI
EsuQKSsL7wrXcuQjYA4nRoQlARscstoVR9GnJCqkxkjxDS/qE8a9cjFd3tqGRiUWB3GiqdYIrGDF
JaO7WBtqGaLsigZLPnkmBxfxh8wKd4doXv/Tx86QASeveEBLwsAcsUPuTKfhqV8GLbUIS+zheqw/
IMm5oyCqnepAi+s1TyAlkk0SloBVeIg0uCsfOEjGKhA+FV0ItVRTiuTkEnfrb+aDrDFx0d5wENk2
XGkduWdxgeiopp9JTT8RYHoooW1Vm5+fTevKSzz2TYeL9d0hBx7himhWhJli2nywgYcOoI+2TEkB
zv678x0W8AM82k5CK3mN/lShWkv688oJZjEdTxPEbasON7K09UOT1XzrWKgdD8+l4rHgDzd6FLZx
9ni8d66CQvH9CXMxihh0w4HrA0VQpslflnAjhDL4T4okA8BRjO+ilP5WMFvaEz1xmhRB9ydPKt46
m0J2ZurtIzYJ5S3GeIXBtz8ijJK0nZBP5m1ozM4zsI+B3vM7bYEg+2uhXE26QOEckmC5Wd/dGqeI
8NWjFWuEP3Bfq06O2uq5p12CMS5KYjt48VxBAbXLDNyi1cP63SVO0LauFlri2Btx1cgryf94lUJz
/eZfF1HnISrESU7t+27bycrDPidhuSPOsGwEQiS/RL2Ce873vofDUeQID7iURHGoypBuQwYxmBeg
yABs331cWr/FxvwvfSDB3XXuacYe2Ch3pmzepm0WmIsKEe+SkS+JL/Gz+EHj1Tys2ebhOnuBMsS7
hK9sQWmytogJUXxX0hIM+ruYTvsugMT4j17H4t9RbgH5xuyZN71wplQzcugzQBEvzkkvTb6cB6Jw
gyUMnFe/8GXbL8y7BVwhgkXcvW9Z9+NOmngN+JI5hn03yAXVxBN7cftfpbwvx1lacAOpGZmb7raX
NXHsu4ByyPDNHFTC50+WUE1XoCggNb1vXHA/9cGvVtd0RUDs9uCcCnZYbWAEl3zq4g6gCwzUqZ4y
OYboRfkuO8aS0kjw6bWr0U8Rtb1jN7AkM8tmR+LI132aUfuofkKYj3aF3EEoWR70OEc3OvfVXN8E
ivruWbLmmAaKIM3v/2v2MvvR1aoUWUmLfU1YJQ71bGY1R6zDIejrJa7+C+dxpLIc/Sg6X3SApERF
XDpn1Z//g/6f7FHbBwlpy5s0iGzTniqctyaqZi7DO9eeLaOnpi5kLiDSAQ5yvJxgc5ff3g142EyM
XpL8YLre/bUzbCsVrti7TB2tCAtbcooqTAFB6XbT/0vWKuf9jjhBlgU3HJPFoLgYua+fC54m0HfI
6Lq7GcoQU8VYA1kvQhK2RMF3OzVqsFFJ736oZf7ikRKtxNXHMERX2XVTh7pyi/tMANgq52Mx66gX
pjwXNjq5DhHWPF1vKm2Qh2pN4fD8ZFgl8pKgnFkxDy/xDsuFd33FoCjUSpZvThbXc8l1W1hiI69B
bXZV2rZf9Hv7FGTnwHJfP+5YTiHySyx0/lCX5IRsgg97Arx8IjXeKFfE3EEU0ahOce6yxUwryq6C
qHOu62sLNCRC+vlHPotIdspMoWqDLmCp2NdZM78LuI9GyZSbNEdXxV7CVMrfwq4i3TciGGAehss1
0dj4fA/lF7F8MOPdn2F2Y2RA2jS64XDSqVjirgObX55vNGeRTrKYwh70hCGRLIhk6hL7Rek3d97+
3SUvjMcyQFiexkv72tq32S4HD4kcNjCClT14hhd4UWbOqtYXEeUUDh8WYgBS7zu5ONe6zbkidj9O
eFaRuh6cNkOtpxu7zGPQFAtXaemUhcpSXALU5fi89Uh4sZ3zLNrJwf7YqTu7HX65lQ2ZTdIcYOgU
r0UhRFwkpKaHEnJFU6vPonH53Tvq5IdEOa9dy0CkGAcwPzqSCHTSVssQYUnDDCY2hvOKp5KLazGV
bypyR+nmEYMMABwlGgf1WQhSLfDBsJcZ+gXOfuiFQspK/c38U1x9Y+6sONzBrW2vrqYSQjDlMX7M
5ANvLCkNmJvQpXc6vaX+3eqGg5TwKIxkdzHZ+xHKKD6fTjH1lQ2umxv/MnGYn/5C6i/90ECUNCvt
aTFvpn8jLRhC7xkZ1imMR/XrGmjt95Ghg/SYtlK+9JpCSjGuvtZoTIMH6BCyIEav4hwkbz3IXx0A
1UW/INIytENlGBQLHuyJyOMz4qcepBVh7Jdpe8lmsFTNX7eqcWrTKO2VNnRmtBwgMSG1Pp4deHWZ
q3owEwL2FhsMyzj3MheH/PnoGHxvVRCkH/2HlkOtMNdKsgyxzp6tuWRZ66131tMR9mHTRP7qe3ml
iT03b3mzYR1FPnmHIHs+dM+/Ta9F5ai2c+wKBB5UpiotL1h3Th+skaMEj6IoW2VFNm6XsXVZ/TG2
lWYkK3gDY5w6Ph6PUuUK1sTwoFlWmZA2uwwR2D4u5VeLvWmBcXmRUavAc1TQLrlsH2ijT62SskAq
e7X3jgv8g/ieT6Jufb/RrJkK6z8/C/WvgpjEoMmOfmE3zrYUJmw4HbhUXiTjGcX4sCCHW8ELfinb
tXZgn7FrpizAXJ8qFsOnY/neBGxl4W1FaOA2FFI3UN0FDt+aiSDN3Ys9wYDEdYpzVL1S+GSJvxZz
Hz0eD7aEO/FG+86/H9laeElDibxIQEhFfnOI0YYRs1/YDjGl5bzwwRk3DTdclwaZP4LiZJagePNJ
KDDWf3VC7T1uqVEhYgMEfuXGeI7LJkgLD7/Ljf0FN5T+YgsUeA2HMOdQMlEYBMQgjYTkpEEkaGjb
9PRMP/ifqubUJaCLBEJWOcPWlYgq67UBbiVpJY4Lf8k/8t7yKLzcMAIN3zy9o0jwfrytfjzpY0lE
8ZwNbZfFRjfZ2unRFQmHekOuAMCqHEOLdNLlXnpPApNTiUD8fn6e1xhrJYrrPv6wpggeuFK45mn9
LbGef+gStCX0jCcuZu3Beu8oZg78SdMshgbCju2Vi0aSmwkB6LEE8p9QOwPpfAuiRhUKzU3h85mj
Ktb3lYD0RHlfckHY3E4cbdkd622P3YRghHzD+MJmaka81aTg4tMFRug/uejecGbq2oX7y87UAJ0J
/cPvdP3VcTgjJilU4x/2czScYGX8pwahwTAcKWfzSwKKaWAXeVHQRITqU9PlpjwSrkOeL/ByDbpX
Z55210JnRWVELYHNYqXsnDfTYoJvm0uIQMVmNGCIkaLDSETSzjxTvuP9SaWiFDqma49peyHm9F7e
ClMJwGgi5HRHOct8/HasJms1m2OqR7RasKkwGwK1pFcp6n6xwo4cFXVZ5Nr79e1n3irrh77jPF7X
+C30P1NomjnRsfu6u2vYeGpMio+wpu/9vgRVSx/oPKFXeS7ORSklph5GSUF01qiw4+6jjTrmcqjp
p4sQM4wSa70aJhl/Y7csh0Rdqn9FesUPcFUghxhkr4Ou5PXkjxs5mKhjBMhS1HVhUBWtWg0nffeM
R4AZuHgSp5R+HDXYsWj1SK5STHPqf+oUvYko7JcbPBcy3SQmh6TCYwrY5NHQnUBLTXb0fTtflGy3
A16WbzqsKgSVgUnSASuQWyheZhLZT27xqJvnI1jI021Q+hR+x7PJ1k04NEqo7Fmdor/lUoP3rUFc
4C36AzBvSn1hGezZuaI0SYSew3OaYWIG8nfywuPk2KhSbbpL2APixN0HWz6e6Jnz7hrBKbgARc1A
FsQw637TSNAaGJVT1GKE61ta2zuvZG0LyoIbE0PEfI/+DpdUXQKjoH0HyFv2Ef+z8a4zqMNE60XH
2t7MyCo/R56bCW83KlDT6RjWwUWoxYHKurfLrjupO3rxumfQFGUx2iL9x7ZNUEZZncS30d7vO6qQ
q7D3dY4lrqhiBOw+wDI4kjhtTLRax3qf5IJisN6Z0d4faOAK8UEcXutovQEhJfEzLcOnY9bgImhB
nXw7HlyzWZUOPM02hjX9e5MNMNZjVY39BmRhOTAHPcAfpIXW8clbUt+cQswrWxnu1rI/VCGt2oxp
Z+mRl/ayF3bC+2TrPpD5TueVc+8hAabOv2MgKwe9RYkq7AdErPq71nWm3stsADTbp5LCHshqh1T0
HBiU1AXWeAp6IW5JNGjvbgj2CJ7nOVCmu/P6/w9l6bmRsudgV94uL2B96kQp2oSaRxdR5b1GuVyS
YIMAD72CZSvq6oCTHTTArMo7ZtPHfeKKXzlvyNUpjxWAMrqofng0H9YYYDVjlh19wQbEiZ1vmto4
GG9mD1fNStbyT5EYJS5OZ6570f6DlSADPgEZ7Xyc1rvto6JQeFxwd9BEf4cmk/c3CfRuOV/FiBkK
l7PGWLPqQg4m9BsgFxOMH8zLLouyKNa224lh57TAKBJJfa8lRQtPCWiFTqGjtY3UdEP82zW9ctA9
pxg/nBaAeAYXTgHAmOf34birHL2EFqLLU7HjIhS3n3jCs0VHpQXqcp3D4fY4sLC/CyVucYBLCmgd
kcS5tkkiEUsXes9e7lRCl02nfoVzcVlg5diXGKXsogj0kARRS+KjW6tkOvEqYQomJMTiARZqzA1w
iMPud4+p0YuhssLLDDTQrKXLLB90HeW4FR+in1hg2DMYqfk96H2gcbuygFdVdbeNu45Th5Ilg+Ta
2PNtjID/ilbxY5TsU0c4108B7srjhPwuwiuhupqcfA7xMdZzMD6mRjAr7vZDLIdRIyKcphFRVMHa
SoxnQRJi0eqhf2sLWu9cCOC0zgUphW3SIbQrfNgBpE7rgAo2a97eYlBu6PpTV/HPGfVW+7AM5Svq
wxf2w2Cobb3LP+95I1feEpasS4Vbp4zjBUUJMKM4IsV4lILFhX21GMJjhIhgRrU6VVIQzldNA74q
Q9hXxYfz0zyBKckCxKp4CQnqkVoS3/ilX3LDys3mdKEGczRABAJ23DBkbu+wqPoiooFeYyDCBTEb
EIqJuVlyvhVVjGULnBQ3sOIOATMqM5In02pe3/gPEuW93x3NsMpmTsJrkmpSeb7trMtMjvMwlA1r
eYHYJLK9Ae+IDfLS8hcsJ2NPmW5Q58R1yEfH/iXaHepQXpEitMV0gNco9pIwi1ZTOR6RcoThOju9
1hlu9Ah1TrsW7LZmBnsQgVn6+Hmj827Ypfa3Bwsy2C5HflnY1WqAtTS8k9pOCQ0ohAwRjFTrp/Pu
5l0EYbdwCl6HOTIQT1c1lkxtGmJr6DqMBNLCZgNpwdbigAFm+4qRbXaaafMNw7ywU8tuj3f9R7BR
Dr/BKCvPb8ZGDeoVpR+9Gc5bxIpiJZiN4128zDG1PkyPFrpEKVF5eV6Z8kYVlC1jLXQKPQvSv5ll
5O67cy9qYscKmz73Vq+ETqFltsmP3nQFPS8mzTT05KmlRkpb+1Z9m9m+jmEcOjJMH+8gRB2ksZnx
4v/ffMjU8SjkzmYVpYNj97dIV+2QSRxg2uViFfUFBtpp+igffU2DeIodY22lenB98si2TT69x7RM
BKGVwImI7AdvPFb08TD2wvCDmLn9o7AhYDyWKaojfjnQuOLb2XVvAsk4w46CtFlMUVBTcq1iHEVm
s27GTBYDbfHiaT/ToTXo6Z7yzVRgu+O8G5dlhJ1il2/AXHpEA/4bqBNyzJQICAdHFIp5QD+Dghtw
AZ+h5aBPaB4BwrDNVc2AM4v5v6rn7lAHSE+Ma6EQ2xJTRIRbIzi7DW82JBhvrzuxvykaH6qIrjjy
RmdEQpToasrC0QOoeg+4nynVtq3iY16nMmtxnQoMvJnxkKk/cps55lhxP0jv2Z9c6Y0s20HoRLzh
AzQj/1FheeuqNmIg/rtT3EBZcjoG9DoVLtUgakxMezc1s1b9V0EOST6ebG22CvxHCOwzLc4rXjpz
ZH8xPgik39SsMOyFWnBF7e/e7iXyvgCT0KcGnrC/+uTYEJX8Qat4K6beCN9mITqmHQoD14mtog+3
mW8AsB/vBsiPbMExHzDOZNQvrsx0LMcjQvHiVEyPLLl/DzbvqqY/r7FZE+Wmtd/hydTtMP03tHxQ
xEJejwq/oY4qWoLuUNcc3wXAXbrrXXZHWAWbcKuEwVsEzUxEckpBPrXREpwL2FyBJCgclMDbVn/1
4gx9MsHMGyPqSPtb0R4jfszSSUtC9Cv/wPgRDA1fOFC8IV5BLV8Ejqkrg83tbIGZ3+UTKuI8QzBk
ICeLXFgtmwV5BrVLxxnvoOl9y3AniZE5r891KNc4wGF1Qxa7ABQwJJq879uudjBW02iA3TBOOsXV
g/C+xBxco7iQc9nJ/zHGP42U4isXN+Jobr8aI7kIm/10tX6wOnpEbeJ47he/QtnFApHHL3L6+kbq
KIts6z0yV8WKy09rce9rCnwsRvajPjV5ap/iV7lwZZN2h6tJ8A4nkdES14TXBG3mEE/Fea2snrdn
CfUzerwPwv59gG2/1fXylOTtCMZL6hRuR+2mL1yUcGJtFuFNK/hUOJVYOF8KF9TsL86WzaVUogTK
mDOpKC1aehD6xmPlKYbCYT0spN2Kpy+r2zstA/DgM/hgsUnVc2cvyWnLJiIO+X+bzpP0nVRjdvYB
B8WDsbR9XlVnEYvdy7sZEixOYejcpQroxkvUjCgxXwcnfhvCxKdGzLmO0HUO0vvz6kX+m9EJoErT
CkGpVVdjsF/hamYdusG2v+/0r2wXhdHePI6nmYEVBea8izJA5MOFsipnlEzjtuOm0s6T8+Xq91QQ
QWi+Nq2mo7Drs9e7z3nED/3+68TEecD9nrpbtO5E9pHy9x5ADH/p8pCD1M9+9/x5j9ISakcUGqSC
VJWnuTGGlHalo5VBOytEkqGwuIdKL2aY8ANSUBiJv47jzRR3/gYf7yjZDanp1y+tAlYisoQMDw2I
MHxZDbksK/sxwrfIHTAwiC7AkR/JGADfeFCfsu1LDEZUdHReNvsKZJ4CDG9d7ZpnSoZlqsqJ41xB
N2K7GkQpk+tI/YNYM98kzlC5pB8EYBhQQ9VYZ72g7sXJJ3eWtVuwgYopsnZHsd/bdgUslZRYxzSt
24hTU1YN/yrNkS2UqbKHWAcmD9ifsLZtdPJ/al9gCBM00dcFoe8tVOGFdddMdSqcZDdMHLEvMzlZ
4lVJHioG+L9LxeEYmAdOOxmpKAmqhA+8VXt65PikY0yVg3qAKWm9mm1g/8JAi+ARfuVTHVIm7mWX
6PChfs7Y1oGfyHHAW+nF1h5cSx9KsVLcem0eP7Za1yrrJn7LwFoH7YM745bF0wjGwX9Unv7XlGI2
272TLY5V6XPV6Vu/6/nWOSZhxHi6E0Fqb1d0y9aZHNexgapjO/WbE5pU5c7BcUl2mxHZaokQJuB6
iLV7K+b5/YRt1U3PCB2WF7GJujsmTocGnjd3tLGDdQMKYt0g3neWoJqxkPyO3Pv2r3MX91kCrp/V
OkSWE/7QtMl5lGBUmBvoU2anjp9OOUe3oC686T921rGZOq7G1rjxJmbURIMY9xiZVKmWIS/46J3j
CQokiI93bL9su+/jK9FWek5Vs50IgGaGZpSXGrexrUKgjBpMphXqsMnpGit5LRl7MJfHUm+UX5sZ
1o4SXk+BTXm5RBTKW3fsOR5gJ33I+c2d3wV/oOAgK6iYiaCEcRk79xP9Fiuh65fQmAWd26k/UAPC
K4dYqs8rRap5759ygZADQKSm1zmXKQDoAPVTZEB39EKTj5wzgnCfOwpez/Bo6FS1CyiC/BoFdzdV
robBMqhdWeH0yDVCCotfcSUjMynWWc1Z7kfFgmi4/3LaUXjPvdIUSeWcVAAPytu6FyoIVFsTwqb6
oyAZoL6RsYkkWF5lOy7Gm7CS6mfxCvQw2SDKu0Q3Odm+4Ft5VIraMKIXE0ME4Hu9wQscbrEC0xA4
SNaCuRSzGut867AU4HZJMLqaG8373eCM0zd0xHrooA1S7O6Tpm4sQeWP6R2I9KTwDwfaynqxrUVs
ZyMv7XQKcx6nNNuSDQvuA0q9dxSi2t1YEBxcYI5K4M3rNBpv83eGa9r1fzqM0Jf8O+HkETlrWTAt
GM+kT4KdtP5YTW8em0ifROlAy6SEbNVhkKXoPIFaxeLL31qxFSwSbAZ089E6oElLNkltHMTozVL/
IlD3o0Nb5vQcr99YCllC4VlfXKK0iWIrqq1DeN8Nbx9dCYdcPXmfOrsyj1fJ1vwIwEpRNPCmm3cS
Dk+AcU9OpPQk6n+Mp0Pci0TZYlarBw7zorwoBJYI1y6Sn0kbdhsUhsfnmTfn9oLe7pDq0cNV3gaB
gw9CMTyRIW5b8lFNeNJIPI2PfIGindLbGZuMiT4csBLhjgN5iNqY4JCbeDjaGQpC01Y68i2D25TR
GjqFP+ZQ4ZoK5p4ml5GGhNu8YgUms609bKnUTpYjvfDdGb1dZGkY3avqN132XGQsBEGS3a3YYmIi
huYY56itkm5uA/YFlo5ERVqmfDJtYm3PYBdm3BK4Pvfesgkr/0cJoqabl4hpu4PfaVWez+c+ebZI
VJLaoFT31o6G0uq6FFcJiFLuGe1S+3ZKlUxghSDqI0B4b6gYakvOO2OXfYpTxfLEXxtDqa0hHK9A
tFqo2nz2JUgVLDgsvwFSFkJ3f646YXeNtbgz4M4/rzCeMS6xN3rGPaHq3FknUY8elj98FsBSRdbi
Kcb1aWZHQN2uCpNWYUsA6W/GmZ4YOu++m0KtPHuzW4ZmM01Vrajf6mXra1t8b5zq93SWFHyVHR2m
6WAs4i+dE4nhqNfyzVpdt8A+9N/9B+S9kTRkil2HkGv3z/b8bARrdTjhXNABgAXo1Tl834IKgwWr
3jK21oepBtbiYXsDgaj2cB7szfTg2LyPlevaUwQZMmnYhBl1QsQVCtp2Gw/fjTLUFRbHvBprlYLw
ctt3VWnS5TEcGtGz1DcaaPCxapsgzkHsXTsckc8mF5Ip0c+DAtYna4c3pXTa7WQ7ny4Wnmi3gez9
ASjGp+OtAOiTRa9QqFOE/GGdFIE0nxriYHxG66X5/pLfFWa0KQO3ttidgXTFB09y9eAAZ87q7gDH
aMC1FEn5OQfcJSHSoGRr7u5WOiWbTMx17PxwX/zImOhGZ0kw1Hw3VVdLUeXX7cxIg937cNPatTVt
+oWmpKERXNUtpEsMF3mFydgbIJFtkGEyR0f5X/vFyhUk5UX4xAlKQr1w/LAjh0iMxQBFKshxHA7j
b36Qgmr4S8zTdLmGNKr6kcMmke3oeWpuOZxXtjG1QEijW+EUYkhxSzXpvrMOsvZ2lDjvMWD81RUS
u9AcdVG65Y8o8PvtFnejDgCVrJW1RgiozEFXpvKSEEdKd9g//4Y/q26RPisusZzXFw2ZHX6BbGf+
aXrdRGtxjJSpNZs19myIHxngA8oT70OGgLhCXiPwe//eLXGTZEagUY6CqZVRg+D6sq9iZkrE96HS
CiP7B7cdY/2q5BnxQFyoNDU/FFTHRUBdr+jqJdIt6uoIT0D2FvJmJXiS4BvL41HGurrhOtadeCYs
eN8Jgs3zKLOg68BGUSU0cPa6SVSKuZfYm61uLdlEnrln5HjjgW91THAsbv+wnErg7Vk5NkE2pSH7
FaO9YGjNfeeEWpUecDshh9eyi8Z32HMCsvtPdU2cGRGba9tCJuHgU3V4WmOjR3ScER3jDq+Kyb+p
xokAUP386evmmTy7cZQtsfeuW/KsCNkoOP6N6LJa8GgU8hBWW8CIDwuHFY9TZp2ctU9FIISUsfT3
2fADsrwVSWchVGxGtTyOWxIkZv0gkWkBM18+9YsZaTRaZJBs5qp6hRzZ31GEOzZnFqyYsLjCYepu
/Qqz0Ah4Y647ffFnH4m/1j2C3kYidjjngIZNerPJnFEsIexObWEjAm5hZB7M7BFGIHRTfcJ5PL+K
3WpzJyIvfU0C2hnOWjoTN/x0WKxrlmMGGCD1pcW6h3aqVzR2S4azqFj8ZARIRaRaJHiAhDTkr3Zs
C+Pie7n8j+G/r3qiOQ7duvAyJnIPm4yJZQm5sWL5uJSg7UschL0sLv5TGx4qdJyRnn5nQHsvF/N3
qtMRBkzzKLrI/iKDFq+hGCASGl6hYD0Px5ZfYFZClFZO5cQzkU1maErbKcrfRzHS3EsZ+42j3ISC
ov1wvzUBReTl43rWuiKiwzHHp+5lRDpyzTYCEIhgZAT36iqTaRgTk1iVcAXDATccFz2eGxZHW3aZ
A19SXwzPu97YKyCpKUqZ+SKpmki+2yDX1dNWXxhXAk/BDkhcduds7NnpUTACYa0oKbIdBq3ww0fg
ilHGTDocByCSlIIk9Xl8c2ckt9Y0W40ecuPHzbrbnmJKYTmvviZ4VQterUXFpGiw4BEIy0oAS94k
e4ECt2Ni+tGt/F0fpBIvaCk1642fHl1mohEyH4l/q5hs3yGGALppxpNUCavMV8zadz/Z3s2KoVje
OaX+t4Bc5uoOpjhIt+Tb9+aMlbEjcWkoSTp/8mIml+VlGroqgKx/FEl/d1XN6Hu3xJieBEa6IhiS
MRn/eGXo6iW9dYauVPP3M21DcEaLqicBVKkL2T6fix+T3DrTdiaz6c61wbDEPxDQJdZewceEFGUa
VfM8bD35dYkLAfGgVUWeqyZGU24/HFhwxy2Sqqs0qWYg4H3ERQ4WleypGN2iEL2S6Q8BofCezU3N
oe+vTTe2IK2TQboxLDrXf8Hzo0BbLbacPparRu0uKP6BLgz8YSIC2Rkf0R9xqjqONXXGljNmUyhR
mBKzU1ypVc22CfY9UwHTA57WO7MJ70Qh/LOrNbQFm53XO3bqT0ksaKPBQS9n9icrcJX6nqbSySEt
9aoepTSjI/W5RnJViy+VveJM2w9QrLfN8MZsxODcooIDgC5y6vTzf33it++hwyvxY73MiLlLd+N0
IFDaOiskBGp757kkrz42R6att9hsq8o9BaO/t+yr8JLuWsqBfcTvVfvO/ZtcdQClqrb0pxWZgsBx
TMA3tmygKymr/Q5vWApMbNTNalwoXxlLJwLDIA6NQpGPVfopBSgmkyJLWZ1nZk2IUZMZp2RDVkx3
zDahpCK8Aj+DxgN4+nTxVlPVGGJqr6r/niddGdjqQ1630YQl9QLjfdq6ZEz3VsREoU3fkqSM14Qu
5nS+e4rApZZCZ2Y5PfufUdhStqxLmrkxdEkbdO3b8uuj/fwg7mjo1yiPVNWLYox45UnY5v4p3AyX
/hHLQbWL41HJIMP2ETYGuRsSiN/RooYg5W38HGqLx5aHZhqyNAn+16L+WUO9uMC6+XQjxPRMu1wT
orZAaD1mbWzhc9OI7Q/w5xzn8n16QCHOtI0k8EB5eomF32upAcl+8njGbiXl5L2wilRklkhoxViy
eZhiR25XmlrbU2iRoxNntx3HC/lFnimwfz/ka6OZA93JbdN8PAl3PrB7BfzbyxOlTxEvncGCxC63
CIkdx1Xfvp9RluIN1gfe/CpxsFkfq7SLsLv+tBw/1WtROKFCp6G82AmoVAKM+NPU+9eZGHoUSXk5
DujmsAQBvfsFFvmh60pZANv8NzRvg2b7WKoYNPD2VcgNr5CqUznbiGp7DbqHl42LufnIIiDmJ3DN
wZKRuDD8WglJNhU2Xm8oHhIdrPsRI4O3UsGn6SqfVd29H4w0S7kJfVDj/pdZcXqJBQ4l40qBPPT5
S70I+axpKN6Am88vR27uinRWgYDKLhd1kyjUD378TpHr40+HwDj7gb9AkpMqKUELgahzCUOBQm/K
661r0pb0b8P+yyDmYPdpzOlct60VRpqPBW6KFQxKzEZtj1ByhJGcaStqsLPh7JKOylG2BQtLdG9u
TnMHffuzvMLgkTyaHYg8+M71b3eD+hUaZNWQne83gs+BS+J3VqUZmrP1LtsSMCcE8unOd5e31k8v
/AOExAQ5SjdxkTZaDe2pnT2bs9VQI41CT6rRLXvxxuvEytPaJ5LahiOqvMSR0dCAWJIUnpv3qYER
LTw071yQVuVPwBKp2peVEQL0yd8JEHETaLlKEJG7t1ZWWHWPNcBgrGLNMKno3YEbbMdeL3LyGwRr
CAwmdUkAWkyVT4yoKAAgqZbs7uF2N4hWgCKcq2oFFkpgCAH2lRNYYAwO8e3tuEyCvy6RAkwLQG8Z
KZd7Nv7q23l9dLp5rpG6JtXBXhcypqyMERcoW2ILPPn3Z3vqR5v4e/4cxvX0y416MqfqOBJykpid
r+whs2LI7fbskQfJHu66vW2MGP4Fs1KNwWC+Yc4vpEYNQZqlC9wxKkOuOQ0VBcIG0XXiDJXeohhs
RGCxe1Wb5bkBPFcvj677/hB5xjya3c0CP/aZmZnKxfY7jlH70tA/k3k4yAkEAdVH0DO2HQm+4DQa
7vBrK3YyGz9+8ZMqxNbKb7Y74F1frYgC2l1fN1Ld8diLb21cKagbQo5KjjgpltpoTeE6xzlmwmGp
hreFJ2PorNVpeHUdJaLhZm8sVMQjt0BQ/eeza7t4OO79dZ+vnj+Cv9cZLVC6aUJ+CtfxCnXDI7Wf
4zCu7H81cyqfc/uf6bj41j62G2wxPsmUe8FLv7rqTh+2I5lfTdZ0Sd/TB15MKDhz9X7PtIeveD/e
SsSUgDWknUusq3DnPasqdFkv5KCo8eHQ8cKcWRkHHxUiMTiNcCdBcFd6M86LZPjoQoeGuzZBfIt9
0FmBkinrHHzl/oKHAAxmAK9+DPNJdDS/eZohQdMs9O0mlrLNDggMfixMQoVtLbAe+guH4rcMsPav
l685Hi7Y/Yh2rvxLZ3ltBWVYaV1z8Ly8a7bi///pLyJC5h6tOmx/AdAPQdyryQja9o5ae4bsnXBW
OChLxe7lqSC6bwFq7bq/z1qA0RD0PqsyR/u7hNTjeCaf1krcWfONUxo3XVYqzKPFT+XyBnXjd2R+
KxLwHn3Qo9MpII9OMuH6DeL32M+lE38rskmW1fF2+A2z0Npp75FX6pA9l0+BaDbb5T7Dhh0kdTlM
seEp5XOeth6/IXcSQ/4qqMbKpY2XNQOjuBrVwJpi4CM8PwBb8F11GU0j1JN0iBdigOxlT+9JB9hE
SiDS1qXYz8WustBrjDHdcCGA7OH8Y1p0dIkJZFEq0pcDKzM+uDa/PTLm5VFm052boLzMVAjw1nR1
wAhiQrCAlE/Lc6dRCN5Qrw9krQSzvTJDNvcPyYlyFtxuRJb9hqLMtKXOLy8cycTpKHazXCF7OqUd
yqu+vZhzBPDwy7TdY14xikaPa1GAzz5dr+tF793LIH62sjJf6FpCFwb3g96mmbJMJelF27OR83We
9OtqTRHiM+k5V0Rlc1Cz0ybt67CHFYwxky7BSgMG2JIrSGUj7GyarRcz0O8EoTyPHph2psZo1mtH
VfrFsQ7OU3wBexHVP8Y2ejeOJS4nnuv6rdIq2H0Hvrf0wSw4OF6S662Q92ta7j36QIEuVOLLIOfd
Ab/6EAuOHIYy0g1BfRszrGIhYUhL1XPGd4ymktyrKaPE9vBpG9bhGWgDhAg085ClUsDkXrfE2Zlq
785NPVt0eJHGSEbYwGtF5uoE8kKqDVAjKinF78jVqA7AsrUEyxRL/7nAj7snXBEk2qovNV7xCpBF
qnxGeh5UpEWzDGg1FUWirGi5eSy1ZAfSMaheqwNmtmU2oIzCSnR3w4d3kgFzuOoF0V/gKR2eweuC
WuMtBqAsPKiF2n7v+h/N7cfPfdP3gn3RovumlFwcR4Yb7PHQWgajwkMJY//Qmu2PIbZwnjP80+wL
h4gNnusOsIWQ2JZLfWW5qsS2NR1m0a76ZgJHA2H6y7Xxy5HNDco8Tm8erwmhACalMfSCxXFwZtTz
KqbeXu9wIGett7zslqoiF6d198DwIt6bHMNA0gSvot6TZFpKmYvc//nl4DZ0JbOKvEwoZN9woDxm
xM7OZdTrFukoN84USbpupfgRWhk60JsU6y2RAmAjtZx9SKVOQ3zFodHAURMQIQgL57SubA1fEt2L
5wxjuiRUkGgor77NsE4OlHXtAznyPFh+4tkOXk3UtOakv+7YhgKftbO2swr5Wd9KodVvMxUqj/CC
GE+rkxJ4+uycAldDqn4RD/OFQ4mmGFe6ii/21/WdNuI+DADmQrO0OKgpYoSAXss9sJJmNQ+GRwhc
fKIHRvFi4UmcbQJ37Umw061kFtvXCggN/OHtfajPayCMjhVAwV0/6ptQweQXoBiFy37uun+/EQub
Jcn5rCREaRJ/ubdcNVPCzLDnxsv1tVVUGq6u6fcYqyCp4g+QvTIf3xsFAxUZLWGi9ZYihM5Zs9AD
uLEnr8qsC9iHEtGl7eNjDUCxIAO+Js+8FcouyxffQddm7SssY7CawJa9cMxFvV0xWzSlPNfiJFir
NxnH2LZjZ1l+D5BXoiV9ZNBgUi3OP7v9/BD/9MBUAsWz2j4ONWKcLwCYxq6zKUs5TqVU7h2BCNqh
hn6oa41PICh9LE3Ec1GmBHrC8LQGyDbQ+KjUSkoh5XB/5pVhYczZbJnSBH51ereT0FSNUlRkmVeh
BA7lKSVTq1FXA/yX2hztgsv8B1qWcY1SQufBpwR+15KNunjRNJFmhEPL8z4l+9NF0F5ToA5aSLu/
9r46PbwUQqeFnR762dF/gln3f2U+rwdbWnKwohjImb8pPvP9O4JtS9i/M8OW97pMUUJbrapW9g8w
+AoODYIGSK+LXdFaG8072pDvJ1xAbYCmn68m+MkLoWrobTFdEn4XUqbkVHQ5EMq3MLPP7p2ba4Fq
0C1yjPAzAlEqkDYhXSwVCjKcC+JVNM5bYkB3UgSo6Q9qFM1OOFHgtznmDmaMjhz6Ij2To8cvYo61
0V6Y0f4bhwFYWpgjaKJ++aum17PRpySAv/FIewOzRPByMpDZXwNsj329QN5cJIOWlExssvuIusST
pIMHXxxK6ycJjLa0up3K8ave/5Smdqh0dKoyweAWvpPjj3kud+Ac83uMo62jsQzgijiebbLdIgG0
S6I9TG38cY24ldf5kdJBqTnXvyjr4je2oXIjD/RgJuAIGFLc1ZsBMaKarFnz1xfi5yqsrViyS8IC
FeqmlPrsa2XMJJqpR6BG1CRCnXUjjsPLhTaMkxR9Canie8wtf/GU5plXN0JIoOz4o7HVLgogfE16
QotuACB6nUpCE1JhpOE9KbzsPxUVFGqnYk/ldzbp5nyQ3rd8Xbl0sLlb8L1lRSSUTodKkdb0mxKz
l5vHoBzQmIuhSEoIh+kuwgWFs22QiowfJfqm0OeNcMpCKBSt0spzJKlFpObLSc53/U4E7bmN+6/A
2HOLT4Bl0Yf/hnPI2Gkv9a1IBjl7Di6JWQGR0TDXZlwYLu6ZNK0yAaasWCt1pAhO3jGo4OBChiGj
8CfMur9nQDEmZODkg5mA6YqUwiP3A0bulfEgeAH0nZjQWKC4wBmRjFTrxTh/nnkb+o/hcpaHqFio
JKrguEDFuwLP84/EFNJpvYEcEe0VfgVAAmhAhtiyn+bXhHDaZqgeRxhgLmBCOdjk/HkZ1nTg0lw2
mO+FtBPOYWtDecey5Jy+TuBEaKyol9sLgL2bTeEMuKKBycBPeEZ5aZ7FMRbyKOjz+sNTTRLqBgNp
l4vWtjz+HuCMbCy8c0K3C1GhgaFQ3yraRXCQ7DM5i5QRXwX1cxB009vSfcyNeqWqlseK/9JE5+NG
e1PlI1SQYQPvujY7/6RD/gPUOQIiFB1YtuXQKvZ58ZiwbdoenzaNXsdFbVuqN5NncU0LPfB0N7Tf
mUwmcLkkTZ6FKAbiAMtUzisDIb3crOezozUjs3ATNS0raAmrA9HGILeqcUm68o4tqclrPDtnR416
xuO8C9eJXmrQYmQm+1piBq2KvkdqNkRXNafL+AbXQ5I5i737buIrxSFXXEsq72u2cgVqUmzs4UKq
DJQQbFNkxFYi1m/u1rBJdIoP+L7zbZOjYqKll7/2yWb5peWqG6TVe9embHw9FtsYLX4D0XDe2lpp
WyxuYYApHr/45SACoVRlr1n+P8O0WwS1YLpAo47qFWlwxx52wgt0imcQUT4SIhH+6r82WxzjUkjH
977AnuOESD+kKNjg3vRBHhRo377e3LlYlSx5L5SSoXo3iALlPSB0AG8Erk/CHCsyqbR6iz0p3Rt1
yCrqAJYy70OSdrHqjEkaiYJTR8vzUaD2Jf8Zju0UXOYuQL3oRsNxMWL4dLkV1XDC5Rm+OOXJ+qMz
apTY7cJ1a6J/qwlAgK+QBRwFFTaVrgvEMErecHW/bs0suWARzOYKjzFXTO6UDF109c7JoQgsGFql
HYlfkc7Oq4Hdj0j4s8In5+4DPKsA2ig8xdPpHIQMDIkmcrrb/oaHFa5JhRiDjX1wIgmqk4TTVLLW
ZtRY0OmerFDewSl49M1bTUYP8M2LiolEC6dsSFNFCyCtOPcT1OQuICwXlDaTJUygxmX8k/9tWEk8
JWH50/Pgb4EMD4lquUo5fTYdp53n5eTj3wqGoBrkVH/oV/9sLVXJP3EB/vEmIxfnctZOkWaClpUQ
tfRwY8WfJdzHMWsnVnX10oSjfNT2vk3J5opmCjRttxLVqvXN71yNxE/oG2JFZ1CxfyceIBzEn/vk
wSbYuMXZx0WtIhB1HSa1ApZedyOmEWB9M0sRxirf2xgAlMSciqybXI0rFyWDYGznMV3sErunFFTk
77oje1F3SOQsMSvRX61tPn4veGmb9upx0skdPxFmd8R0xwkNilD4HA9o3d0lgQB2Cjq+adUjk1KM
yNKlkfb35n7KebDjcashEuyLs6zESQuXHBWoqt0VbBaRlYTJc2kvLzfxzS4BYYl9Yl0W+Z0I4xA8
7//8vam9BY9WZ1JW3HM6EBW+PEyLDnRNxyT5P7dZjwWYfYpqV7JwkOgLX51NIGk4mAWoKfmMA/e5
JitPu4UzGJJNOr1QLC1nj4n9nXh/IgsUyVkOSYzR4QwyigI/5DHGQe61d4sXoLdvXVSYcny3AqON
DVerF+LB/pn5Jo1MGAgLqBCS2nWT5tIveHJKsrb6KGADrSH6REBtFq9tPbY/7TY0bK9noj7MO40E
V2dIEi3qi9CdxHV0UBqp0gNckOYXhyHw+/4XmZ1IwmT/GiCVixVJEfzFCrfO3CSVMs1iMGrT0M6T
f5XLOKKT0nkFvUbbqP2lCGeZSMzAPTRAKSi1nFi92c/1M9veZia7+jexLdp8qkROAnqdTpiJVGR/
/XB25xyIdfb7TWBOnjS0qVAcbAGqKu69ANHNjiyEpd/ikoxIsVOAHJyeyFagOQUeasm/k/hho+La
etEZGjz9WmSyS+tP0DgrXc4vojnpYZ+cjunCWCWKtvdRodllRjgaxvbAJW8REK8yU+Mjde5dPc5g
WihXfJsAlaf8BtmE50w5ChNlQZKpGXYYVRmf5lp0ocW5MbHKtrwwSxZJIKCQkQEgDyDyRWJZuGoe
QWchzzJ28NG9KWIG9WE9wEFldbB5vUGj1VZ1b1l66/WN2i08S4IA8uQdi0+OvJ9AVJcEmmKjW0H2
VU7zu7GiUihFKwtk5zEoOAEORfTiT3XVSjO9c9AxH3f5StQZytA4xcEWj7cMdTuKAGFhyQiYk622
G6vPfrP9LnEcp/O4T3LHzVLDKjebGgM/+IrQ5xiSdXq3FP5Hfq/aJeTjphF5X1H0Hx/HHeLoZqvG
P/B9UYF3uE6dl+nGOLvI5OwTLiTddWqLOYFd1VNH3nciludror5jiH422ya9vWbF7tNtaBtX6xYo
coDWcBXf5bAiJbMs6H6+OW/OjoFT/XZQyG7v5A0cb51vDMOhoK5k2cHh+o4XK58pv8Zxp6EdBPUY
any5gFghpPFjyB6HPBBnVsxz9Gxm7lRHkVExG841OxjeUjE6RZZ3EEFAXO56Q9Kifspd8+iXa5Q/
/44/dtbjthVIjpbHa//kx1ZJaxAt9MAqk1Bp+d+KjzUkKPNpXRfTHpdcFZEnWAA2/VKCrufqpc6+
SLNzfgrpw5V36TC3z7rZ06SosKs4QvoK4vZhQHB93Pas2z+049adRyOieUpUXT7Pj1l1ljbSnCCT
fJfNlIHPPlhsHCfmq3+IhC9gYjnVl0q4aUe8MTiulDtfoVH8h1asFhBtECQAjejT5YLznAp3semm
ccM3O3u2kvY51dyfUhgknFUx+zZIK8W574aSq/8a/caBhoGqSa45wQwKSnc6Fc3ICqcG9tlbhKKa
lkxp0GgCvSLatOtmTyNwTbGZbld+63U33rqN5QmBV/F7ft2UgSAKQcIqOIj/1uNvSyqGHTtUVv3n
Wh0zQcHg8w09uZM/tBzwDS1pB60UaopQe0CkeYt9wJ3P2ZQp5rIlo6ISKQiw9A+f5krBRCHDNTNr
s9h08AwLzUrofcN5Jg5OlK9As1k8yFvpgwkjYKLBzhBbWCbkd6Li9bFXkMxqkg8R6Bj11IiHA7xu
+9lT7Oaz6jnn9w4rMeO6a0uud/+ZmE/QOmgAGOS1v/Ah6EHTBYH5/7kpLV+LTkMr75WtbVEyR/d0
drokBhWAXb2TGrlZFbP7II7oo2HXcOSQ5zkESiGMVGlx/B3seRxYl4ycsDdDYhx64st3qytfSpw1
jEVHv49CaUUv05Wz1BXRfSbW2uU0RHpsoBW3VN5X/5tF3tyG42RLqCA4a70w1jtPuiy6C9jGXLsQ
6XMzv+4ZFGIv4DBZ5mGbRp1GsjCWwyog0bJlG1nhGtg6+hc7QV2kUf9ZQ7af/pn3jt/lMIGZX8bj
p5X1/CuQylW4hGWRuMK4muvJYetXsvjjDOz4P1ts2zAHw5ZuKpAhFXfvaWieHDxiI3ilRDIGt47q
4O4wHPLQtmxb5058QWKP9YdXI271JNnsmtCrJiwRX6SEGafhfCpmARhEHDmFcb0G8MX8gWfzIiId
gNlHXhUP/I9cvQOwm1R0gndwVLFcUpf9C83Azza3msmEbUO1S8n5NmEGbmo97UvhJdOh0vw+JfSW
cjcTD6pbZWt3t7BWOlPDubIUiVLrEu32Q+DyoznhwixDz5QuyI8Kb2eGJkr8MAQ38skJohB7EeLH
Z+Su53usQef5JqJ52ozId8HxYPgoK7DfuS43oFFBGCVKUwGqDynhdMAXq+A1cCK22V51NxfO38T7
dWsjmfHFl/sYEB6TDWGCf/tsmKEg9De3LGFPM4d9YLckA12/MFGoUetFWNxqGbfw9DeshfA83yhr
IAGRg4FZtmQdoHj1aqmrAtgROtSqWDZOrqfXllBl9VVl7jzL8eQfg9hEdAP1KdaIPXrNUKa+7y40
o+UzsqtnKByx7WB3hEb0HADIzCrSKrlo5phCHuxCgpUYmiq1nWxiwdY4WV2cexF65f+nKfB7uWgE
K7jqSzgPeAdWoRgGHxYJ0c7z+sFb24S5eYy6WnOUQf5+PglBtQquqkoUUn3p1nsBbCDp/CWg02Sp
I54LfIdesqwqWYmyjnGA/ozfTISl0kgtHbXIUxk6lL0BveWR166NMg+0mY8FK1+8wVjA3/BqkG0C
Roh/GWhpiSMvkUv25AwWaDPQEesVW8233KGRt013bxrAwvpx30p4dz5eQxv66QUBVSmRCRtw5LC+
O0unPFaenT690AQB2GJzGey/zuVcRGSaoKGKIMOXJg681k7nzh/b67G3i3ZRilKr9NOoukUJ6Rf2
8Ahiwit8RwDfwfM5hO1OPf279+GyDnQ7EoVcc+WVTWC6GfpsvJKPcf0HUwui1+84qTRrm2HKdAMK
4EP5pVyyL9wP+m2wJB5KopiSYvi//1YlT3/LenKxsdPAm6ZWgPIwCtwVn4J7TXfdW7WbWqTr0VhW
Rtar7jx6SxzTNuOxUdsaafTi3DPeeGv6tTMpndJA5SWpwoTH3R+9ijPdqIHTe/qxnwdAIMxm/NrE
lCroXfBXLBCz7oC2XLp66NaqX4ygAxtdLyocq5qPI0166fDGJIJyLILYoNqornX+EI4o6ZcvNr/0
9PD7jndgqouUdOm4XY83AtvGhiuPdo0TY/ltZzN2C+SdlaTg39QZwHs83hhfe5Q0u+96zLkEvX6J
mMKoqOUY5FtmXjU8YvN9qHAX9ajcG3S2YGlVjZrAlmN+mgQeVW2ewK/65vjLWj5XosQNYQj3kyBU
dIXQQ/js0AO/HcIWkClgJ6a68blSe5NKLSWgrrqkoap2GIvd4HtqsgLd6vY+hrlcUwUXW0UUnDkY
q9anjXYxfSi9SBq+a5xNobM6j73/gD7hjf3bKgLDEZbn9MD5RTuelGixPF9rGnyTCOU3HWTDAApE
elSJLNlHVgMGcQTOCuQFSY9KYHQsAK3iOU5Umy/170rPV4lDjTrl/D5ZH7cg7uEGoTCG/Q63HTng
h6fKKb5i7loQ5dG55PLS1XeTebAAJ0NAvTK+5hWFBjgob6xwUpXwGTFgBf3vYcue9XbcwNCRdluQ
7LUVyxz93bqLyPI7vq1rb1p0cpZG98ZpWqa4C+SjX6zn1wO4airb6pp8J3Oo8l180rtPFkhhIAmF
VGdP0GEOSrBNehWA4DNUkvepvxrVIhG6aW2ZCSahmwQNmC8Eh31vEmwwCkLFFOus1wloyfNJ/LTg
7QrXhe8B6qFNy3eQqLi0qVrDfcSsHt5X3VRgzzbaNOh47q4ekDGbVYPHFX6EHS4at3EE7yq+lW6f
dv8qY85dmj2YOh+yJwbjaQJ+EQbuSwondW9+aOg97G74rqFXyAggCVOZy63SPCVORX+jv1J+floO
AfW1Xd8TbDFbY0hEpOT7mSJFPSpdOGMpGVUAyUm13CipzxPKu+E52pfrWz7C9i/S3D8fBSNRYVb4
YdaqGw2yRTp26wx6fjtWV5xNQkezV23g3ooFGOS+gB7PAJzmcv2W1w5pMFc9WzxQEgYwPKxas4Oa
ENLBmqy1qs/Yp6XoSyAD/i0jHbDINIPqOEtKhH76DFqMQgVxWveEwvGiMXO/PA5XNSq8DLnymYfF
JSkSDhlxpezgACfwtc/ti72moYaQ+FnUIy5h1wxdJDwJRX3VTT+kVrvN8/gdrMGMQSmDOTBzm4Ay
IF5HFBE71uiuaAMgn742dQntDXYwguz1OuBmquyc+/3o6Q5j1lKpUhjbBCULeYKj3R2DtElXzUZO
Ykqoj8PBcml2gSdaWQ+jfSBtlbQS+/V0gdcltL/Q+CrmsBArsDbsjJwABVCtlqwTZEB3ii6FBzib
PqZqFWBAtXABU5Lmyfx+OKuE8p+HjEdooKoiq975um32SwARYO3xQp7EbHb3vp51OWzSMYuXklDe
1xWJ1a3lePy2F+KLkGduNWOJVc7cHk5e+Any9arZQhWgkY3p5SXCV/sciRvq4Gxg/SzpxtQ7Y13l
uQ2PnSqGQYWbNon5qqpvl/+veAwPhDJ1h4BxEb65xJesn7qRpxbR2STX4XshzFgWdD/W6LxxAPfS
M9qN/UDhFXg5sgjLMdSDkwd8aKuhSNgavrzzD87Gm8wWbiOpDhI3sKFnw+bgt/TWNQ660BX73UtO
i/TMJ9WV2363oGXHMmiS3uzjisLns2ytwNdHSsJZctjvdWdiKM8afpPQGQijN7K3jA/msLCiK1gI
hanGSibMRfxCsc1LlB1Nx02ASfMkHwm7DcKQUyvYUX2WKehV24Awbnl3kJgUm7+VKp5CUfoDr8vx
dSjui2sNNmnHl6B481E/45NcZEbIUvFO35ln8d4fT/NHr1jToW5ou0exQvFh3wBMiLf1gYikUTeK
hovc3lEMx7f2BxAGI/LjO6k9eIvUXWUD9KqnPhYH2+/C2AiyGQb3ljJcr0r07yF9WbzmkzKQBtdv
WFh3CweBsrneuTCQ2YOaLoryC17mgLVlkNf2JyFU8TfMO0UKcBxNP7QmnqOocDTI8oQbTbuWhl9d
VATg/IfYWmoD2QPCyHmqKSphdLQQPpmdUk9Xl+QdSpr9XuQkNU9aruz0KeQIMY5fqJHIhw0pr/bY
Uo94i7aHV4Z4FYfRzYe2nuXaPuNLhe87D/pAhgOm/aGyK/BLj1EL/HVH9lzsjIsdA6wgvQlQ9jQO
U9PxTcR5shxtUbKWrEVKmWsKV14z8pgMMi0FLg4e/wpni1prS7BPrh0zr4hnJahEi0zI/yuUiH9C
TtgI4RBudHE0qrLowPkokWtZtkahN6e971yQx9XhtuCZE2yZLyflffDGwiDH73wJbx8lUSaxc/Gf
DTSE2NFL+EY2wRsk2faXTImCTaB+88sh5ad7VyLYK2CDPnZnbBoYW0n4jU8Z/DeDIoV4b6RvqU2e
H1RdSjOXRlnLByYKXsas/IYPTSXPOb3kwctt9y6lMOeXrR3AmZGIRCsRfBHQjOKNB5oH1F96nnUo
lfNsug5xoW4+dJ0ckDVCu2uHkOmWS1BAMMTaJUqNFWRQV3NtkomSbGBOBY13Y3HNzhNtLn3D/Sr3
aZr+TZn7f88pKgEPAiWChUlCtlEGCz+S61LgG3wbrSJG+7xbr/3fwRbE8r1L9KKdDuNh5JOIBrvN
n9B22wFP181AAWDCxsKgR0rg5Ca0tzkY7o9zRBCUM3TWkElDO2dGfQSoXboqZWU8xP6uzr+dExKA
6B4LMu60hGF+yAdtSc7QVc1k9ZqWJRyYuoTsTT3F8y1u/hmCdLBfqqAllblLRYEuS9wpNw4+Z+FT
a0YsIUX5//dzk+emkRCqAkDnXDhl5VnCKxbixWGgouDN7+uHIwgnAPsAJgyVvh8DLp6mXcfE/QmG
Xi7FFf8xkc0AuFHNeq5pZvnfW3jUEsjTb1BIIHKTof7wJlxD/bFwEAa+mAR4Q+5pvR8XBIe8OHyh
YlYwDYD/ceM4w+6mcNhqgRU4OF2qSCLYA5Wo60Zf9Mekjf93kh+Al9wTMHGPf/sA+uNN2ogfp5Hz
hM680+mZEYGXmTI784eT24N97J/BOcWNFzXm9ZIWDGO3+P504+IzbFQ9+caZSvAyuXctjsa8QluC
gdmN/1NY2+Y5u5VQY6dft5oNA3F/ndjvuIUrx+Ep71t5t6QSsZ4S3h1Z9oLjM6AK0h8KwjL8UiRZ
saWUdxzwx3JHfABmlk6EL3YgfqUbpCKzh7SMdRCX7lnHZDtBMgEiH5is85F0gllX2CniSi/HREbG
Dkz712N3Jeg8BP+VZt3iP5qpNmzdlIhZEk2SVG5mDT4lc27mvDYQe1nHcrKX7dz7wcIJ/T7e///7
1KSCgd/m5J/VrMQb7FmE4MtVxY3L5as1KI3tfOKs5w36b9T5ZQ65I1Pz50VUIoYwJv4wAqDgLZMO
PuhjOD3Oa+G9wfIwn7mpHH38fHFL2s2urqmP/HdZ8fX+IsSTioqvcms9YxtVT20I/DPzuSfHxLU0
THxk7m4i/CfRTps5j6YhiYB9z0dqD3bYOu2MWz4hlALfB4XhuJq5qWPbSX7UIZeDu72cxXZZqV1R
wnIrYjCh+Mw3T5daX3pdNg0j3jdGMQROkHnROI1M6ICP6CCcju7aZblppnLS0RgpYut8ApVSkt3R
+uZ26uF39oSTAOIjr1JoIEA7vgM8DMOUvc17bYkRNB3gHgIInK+x8dUDM9unqzZReXOTPYDnl5p2
7H1RzKzzXa08x3PWxoqbmYbSgr7Vk/JCu0o26OEvHHA5+Pmg//oZywb2/Q31SByu8XAIOtfB8J/I
D3nS50efXmEOYsMJLbXv4XE5qaPnX41DlsGLbCvoi32dPkNtSLmUqJA/jea1kfASTK2zJ3FAbX6e
yhk0y0obzXJYS6tH5WrPSGmYtAwXanLJBkW1e2ROQFtSUGmU8xDMwpQFZ7BZssU5FsPF6dy0zPCH
lzPQC2jAmhDLotqcUc1BX+5l6i4Ij8dajc0K2OmJFGiiS0GUOwgFq43dSApyXIyFnBqYE1GZePRD
ObdScCwOBt5XmANEOdjxVGAcISKzgcieHZGIb1JYNXCCKfWnEQyu9YM7UdNtK820kiWXgM5P7LaY
i/R2AL1PyQ8Rqg8YaWFO5D8xzV7m9dM4/hBVWI2aKpepO4pm+i+iKTdmkjeyBT3amiHlC/L8u4v6
cyGAZQ0iFsijq5b/s5YbJ15WkfMu74Ayjr5iWbq+gJ4fXKtheuj2cB5krEjoEQSz/QoVT0qhqcIt
HKIuU8dbcta4nas60BmLYHPzL1Fw/XbnW2LcAY/v/AkJasWXaNNavju1x8/+QsBxPhUoJEk79xPn
FlYygLIRPgGSYrnc+GqlxIca7bWy12Uvtbv2yKdyEzC64cvJ36wByZGpQPvhxodVA19tnbvXaTBa
6Z8qTSCfk5Zgdj6eUshUWr/CR1Lm3dxO1yjCtD/ICskY3Cy0lW/8RHdBsybhZC4QUuNQWiaKe8BM
Q5RUIGjQlNnx2Ryb8sS5Ec/um0SR6OyaGfMIVbSTc5Qhqq01Z7eJ885f5RKcST3eEaGGK0g6WAZf
C9wDU8S9Q1IjYdi2VGNRYwzF1xZGigplHrBOFCWimltX5aXFVaMJ11YrDigAOnkX7LAozXpMk5PR
9CVgFb4cAgy4xIksee3Ey+9KZjNJ/xQxcyISuUpGCwIbMnkIfJzAZ/znun01ububXCqRhJJ4Cnb1
wggHvoZRADt6vtgR5wN6JTaLBr9pBopwScvOTHRKHiSsvNIkO+aZK6k2SIEvDJIuMy27kUUIcgAQ
GfMxsMY2nmEvNObfu3CC90CaUfMXMy59fx6xXXEsUWYniAa9uWlsT7Xjq3MsJEc9OSJFdYSenuRX
7DWv2XZE6QwkVDlkf76QDUZbTORnETCRy6MKGLYzBlh3wX1gHsSl9o/vt7FZOdEhIZKPjRFE0YXv
wjSzr2XgDC16xkzJBUki0dtPWYX/JWfVseEf8Ph/Prh10nKMARJbxR518cIWNnk1gE3a90pYp9Te
X4q96fz4eaBJPRbb1SD3Pjp97bgmfY1vFeN9BBDI0aKSE/rVXdTNnJvLyPMYLhPXqo8MCNIuQMAt
jMipN/aTuchYqLuH7uqkV2mq5hgxaQZLTXSd3LdmSBRlP+D8qFbsZiqwgRfpmaI7Mr3zcq4JbJDC
PIav7A0SSfZf/PWLh1lKNujWsW2LPRt9xyJSk/TzZYjMsuU2qJbgZJ+Oa2yoZzGUl7T/pnlP2+j9
WafhhIRww9pGvdr0IfMysdSfmkmCD23LKbTKjYSHXzA8E4DaFNJGNdWcLIFPVctu03LtA1phNPaC
F9ig5M5xtFB3rb4a8/Oemco6HCxAKrSVjU9wuhOO7cdN++ESLA49j4LcYofMbYrQT2WUo9Tj3NJF
jiTosuL5ImEJxNmWlBY2uq0SOzgUPerGVY/Vtm5gp6d17uKyM8S2RgvUPTTp6UQBK9GmSjO/x1ZP
23kld/JYS8PEAWMbJTN9mdL+/4oRMETQQ2TFeUFX2zOF9i5vtatHzPfkF1qidPsJCLHMFZuMH1gH
sMX0GdzLAt45B0qppZcKcdiNu3qvP+R1jfdyaN2A4pnH4HEDdymg8wYvKiEdHO968JLs1oZqIM8o
pC1GF3VIChP9LNaoyfOR0pOZrme4VTrBZjMAvs9b5hZ/pXajJ+lOhoid3HU+1nkKxUwIlgcnN6JN
Q5XnA36fqXyazKO01fgA7n53KtafeYnhc3Z1Y0vyxCPTvmZa79QJ0vOvVXhenACcchz5XXa1EH5b
pQQW8csUGLp18YVKfLvTTtPGSMoTFiiglVBLxVkkeED+WG+BpTgeziesMYIhPZpE1xJIKB8uVmEW
rdEu0S0VVxIkIofuhr5ayG4BN/B1Eq8yniJuMRWTNuXBlwCpnmJwFKjNNGtMKiFmivjYfhNICYfq
TBCiV0tUryNlCeGEOczsWZdgAuNmOH3DmXk3+Od+zNu7a4lO+TmuA8bUkOlzo6wgIrLLMzOcR2Eq
QahA+uN550gZplEe/REe/2KpilgXR/SKx0STTu7UBXJZxIp83LS8Kz1QeszsTHOkOY01608T6shI
ETzMCgk7Riey/GdXuWSGK1vWFYUSRn5FosB+cltiOr+rZ0aHekYuQSPJAbHfzBmFnpDwtyzSuvNL
UHOLnA8DOrL/lZch10SK8pZ9bH4Rv6XoA1zHdAKKnAdE5lgcKc1zxm2O1UEkHRLAC5mXgEsmyjmg
4VcpwaKxO6J+GxEZoUkr4qv+vDkOEeZATlyMIEjJ80yXji5cMLNMg7qsnYdzuCXSzU6G7kq75OV/
d7EURQbeiWpdO4u8KHSCUNjIkdbrDWJiHjZrbrxjfCexjbIAJGhETHm8/GouYot0r+PH6F8UcqsR
3rtZYH3SczR2ERswPgfWkT1E9QWgWxfkLJYqvpEjfHK/x3R0Sjdi/jFOD98vgBv/sGfn/VkkRR8a
sNaEuv1Cf1c12x8+DrblLiCaxgbKSW9zupSiisKZBM453bEW7y2HrDE90afqZyFwn47kJSBIjNiY
pBjsyoK/kmSQMr4Qm5cL2uzZkt+5vqUF+ymzMp1T4pzmPbG2TFQRgx2cv3bwmhgC3KnqZwcot/pn
qy80eeeJY+vBzLO90slfzLjboDYgz2afIwgh/FTykpBLZbUiILT43LLJe5OTUlDIJV59hqcRBXaK
xDkD2z8MXX5D9E2I6u9foyCmzZGPnSwESanRx6Fxur/AcT8LGtrwDu/RuDvVCtbZn3B0hYwNucm1
FxEAC0NvK9j9oI8Jtjby5ihVd0v2xYqEQKI5dVU/2GdBPnBRKV1oL9U/kq6fc0Mpssaqr8qCkIH8
OUk796YZFoKIscnxjD3MQtRL0hDHhfSFXcdS/JEkp14YMrJMjh93EEoprmrhUl1NAl5naOGQxOXu
sROMnu9qA4EKcnZw7JW3FiGgDK0tursAxsbMJ39Y/dP4CGBvEpcGHI3gWVn/wYGx0BYkdCmy1XPl
BHx4ZqS5GYY5LP6JtWF0wlKDkqPaOITR2S7wo4NqsXTj2Dv+nkg7O9mgljbQsvTTlFon60fupinJ
bMs245ZnmiZcQeUDX6npCwFbZK0XWjUFFugzs9yNgopvG1vv+J5meFGHYHDw0371NdbRfAw88hD1
d0CDLDtAACY/okpnf6WX3yBVw7gF3RU+TX17mzZhntsEtQcurNS4ihLjwwsBmDvoSfft2Ydpap30
2QBZFYkRMOlRuOspk871CuNDcqXlC+RfNBKpgvA1jyzdIXysjXWpSnsb7X1zYGx1ypy95L/nA+Df
evKecZ+5b612NDBqcdoeS1Fkf8Kn0LiYV9qChILgoRh8Eiq3OLc1/QcqBC8WGYojZTeVM2UD3bPr
bXTleAsfyHed8k/9+fz6zhg2DiYx6jYeVv4Vd16KSXfQt3U1XdhPR3LPX2sAXi++//3IedXzMCcV
LJbSYAuAX0QLOcOTSMMyKPEQQsizBuMYSWkXB8b2IAAVC3jiWrzPXgYOYguFeUc404GYJ1fRGaRQ
ae2Pra5aJITfZr+vA0Nx/AdxIS9S7s8j/3ToU0IzVO4FtkRAmtcWCQ61T05zFjpyJtCWjYcDJpDW
tvZsxyf57Qk6vCKwI72yMERRTqeIPa5Y1ZTYF3YWzIZLE7mC0tSGnwDMswXbJlGi1W4P7teLNJUj
QKZtP8LX0rcxkfDiaLCKCAapc162qmGjAui0xzyfZJVU8sZOa3U6pAZUW296sKkoExIXZHljYGIP
c4paD6C9GcQl7+79pOnydU2NiH73Isqi1oZ86g3KE3W0trL6Z6gtTvnpAdj9kYHAkKIeLnrZSWvn
tD3w3kWjae9LW9r7SyOqJwQf2U2aV9gpXoYZBxnWui+NzXu6u2HToNBEUiXLJPJC1l55EmPeQHR4
fOyrG3uz2YhT86/GblPX6dVuM4fsPTHX38NW4mZtYGBYleSrDLZsGnXwjwoUYvwpyAtHorLMW0nc
wtyw/Suk07yEDmCMG7erZ7YtSpHvqpsZsGperQP56Q1L8oFdulQKFZxU46xc859ECGjtLmD7G0eH
0D9dLeKGc0oWnkm4032y3rr/ESTpjCxy1su6lL9CbS5mizgx+TrWRyhd5aEMDKmCzBy1SJ9ePj4M
7e+0ILkEHFi06vzKb+AGyuIY2X4MWJ35rBzSZqhwz4tnd0TGhRTlTu5kcf0UTcufm95tzeCxb/FN
bdLJO1a5Fd7jR1cBKKhwuNMb+20nWf2BnrvF4CF7JdAOcUgRp14/2lwg4m5bo9660hkMIuTsM/jB
DauNR0oKtR+u/Fn1EHpl6Pwg5cFX4NFUKeCwfbWmvHXsZf4lLUiAHS/dnA8CwXTDdjxRmfjqE/pL
ca5oKd7/CpoS+Uu1FisO/jSAymvuw3joaRgmdCa3Nbzgqn5dIZzqxRUba6EVsLr7ak0FRg+ST04L
DsBLFfasxJTXtYzeD4OLT2H0nsj4cJ29wvxZK7RDh0q9xsFCV17/6nqzPXT043PkJqg8qJ1WXP72
wXd1mtmfaL38AFmW283mptCUACFuVYSwFx/BlTZarL5x+SFxpK6vH9Oot0ic7Pv1oblf8pbTgawD
t84BTT8HAsK26cesELxKaqv1RCq0lnQxJyNwBOvBVjxh/6RtUuhssG8at9aCNCFc7H+WUUcF5eeX
P8sS3iuyPQ09ilBnmUAyHpKLd4ZVZUenUoJc4Xcy+rpR00itNNjl7HM55/wlRwHX/P1BSoczLcHI
K8fiZabOTKDkc7P4lVtdWO9hpH4/XweQpTa1JXBj5o2in1o4R5qxekhkJb3h4ZZwOnTuZ98v2G+s
+mPKjpRnXxKIaZ8KdAi9jDBEE6lGaOB1/XxbKtf1H3i6he/WM+WPSD0Lwtj6zu4Cy1HbfKmsAq4l
fSVQmJmfVDoCmdH2YfWCPZZlI7TxFVX1Fmzepz/CxK/C0RuCyw3Ta57onIXk2zgZG363U509Ig0m
XY27+tEnLMVD1LVXBQntbIsRHI7Oa/N8uKTKluDMNkBtUjRsBtsI9x0291T/uEVU0vUjnpuWUukl
E/fHzs0NDS2kR5rEtq2lTEKulJSvHDih+4Jqd0ATLYQv9AiBzAe7jQsbdIUkyu0DH7/0SQ/k/Ibe
D/Kfan0A+VFYUG+XdS8GQpLbq1JZ++LU7zXKeVUcmOhyhQ2xaR6lX9tGJBgdDM9OpQ6v/WEsrPV/
sstOjzUNeoQz0qwW+3sQ1d4uFAf/9rB6apX1BUEGwW68RJT+fS69Nxj9lThAnwpgOYYzqRtwV4ik
eV00H6pNou7jSl1+5WsNrNPj/bN4T+vMWb4RVucngyW33LYrSzHWjNmeqfQgNDdKCAEmYR8CAvAp
gpcXukMCzgBQsIyW2ghbPEA039F7DMhN/YD7DeOx6LP4x7xIh3VcfdhDSWjSax9Pb6YTWkAm0TMK
2w7ne63jgG/S+ewxHw5ARZ9UpOGtzfejloBqg3546c2D+1uFywjttzrzKDtf9vOQYakUfL9ATRlv
QPrYPLnuU7ZdTO6rG2/oHdJfAXh/xA0PqtdyDfqzoNF0Zi5FC7VzhoLYonpNFhSMVFo7KFzshNU6
mXJQ6FTKxwhvTwmlKoeZ8NM3kCqD9YdbsRcPUIxcCTb9/BTmGVC6QukcDgChI4zCOkz22xvOxdW9
b19JNrCfzuiHN7rLZf146s7XguzmAahPyssnQneHicfUPFpB+xyfPFy16dQqWPClSjvjJCvZnOxy
ueeh6aQcoUXWHFswVMetH+Tpj2Zh1+8BETa/1EJgr9grrmKyGQDh6bxm68BMTek22l2N7reA4ZS7
yWpl7Fp4++yQGaKSwhAyOcVMXtxeeXuuyyFUgHtPaI8MkhaoZDj2tDY/FjRnnPyrqgfAzqeRYjX3
u215SzDuP/fQsSz55wFGXCQj9Dw425Ma6BwetmGC0ML4t7btt4sri2ksjL4LF1c0T2MfSsCcXGhM
6bD76eePNgJzwDTZjM0SVpmyninW41YoGgdzu0Eyg0MH5Pyfkq58k8yJAr//DlrgW0nkhCk+hN/j
lN5ekaXsWt15d5W/z/UHlQpxplUI5Cd4UT0nwtT8EwXfLpb171Zxm1+C0yRLVV9ypWIAcME0y83l
mZkVDMSLWownzlTeNGDWsJIau1av0CFW4bektoDPAQj+1OdI2eOYgURTPHPW0VqPDQCsGelJqQSP
HBSkwTGuTPI2hK/OpnGYbBFFQqbbyHzKGuCRSbT8dUx93+elnCsGlUTnk2a/ZRFxyYueZtOec5r3
3UEq6XuVGZkUPioYL9ngbBmKCKeLMUcmYWwAOLPXY8DWbmygO/9i4Rk1XEO7AuzM0Wd1WfDE9GqJ
0QNPt5OlYoXrdjDJsX8pSl4M0tjvVxF3YqfjMf6lUOVPDy7qKD/hbnhCTTorsDUSAiYyzhSnb+7V
mmTLdkqtk2xVH5Gw0o2Wp7OCegw3hMLOP1hXAL+ClKfu9nrhUlIbakj4s9PXIxauervjxRIAAbkR
U6wJjjahJGywhkJSptu2whkPw2QiSPaTUNlJGoVEDtbjUGoO5Uf5eLze2vyVGlgOW7f4bHUfLgBg
BVr9zm1dy3OGs9oFqefVIzpQ/qgt1yUdq7Z+6p1A1Qv7EG9UHfKOyqFW3WOVheWlpLb0uvq75fHY
Ks1NipJPYjkOtRroLXdqQy8r37/qiOnz+XEv6d/SoXDTWWhDamjNhHNxR3yIlHbWEnDskX3vcmAe
7Rd5frRXz/bhuezXyCtvag5tBxWhgCX4xlMkzyREZFQ0LkZ7tGyij+i9rWzi/ZbpeqKTUdlOig2V
g3YTk5olHFOwzHSAQ/feAbLmxhAj9A50gQR2IDIPKCMzai8UdGcT5/BYVADFXoyYxShXsEAy105S
L4L13c0Y2Sbjf1v2ElVBcA/K0EAsYK0TKz0JWgldj5sJf8dGJnXydBbJwX921Z80QB6CXXxxjz7p
5xEYq1QZ2TN9YcXSfkeflVAqSaTYHhLE869U/Z4VQJujlTqJy58r0Jy6tLPDKlGm1kqKVbDQKNNl
Aoc9LVwHUzlqYAQDcn8rDYy8z15/twSxNg90KeQ+hMhko8bXv1vMmuhwykq2EumRsDI+SteenLrE
YFxboWiFg+qYj7ceFw3PrsFjI4TjovWSMkqAUtCYu9kKYbr9oDTag45a5/ORxp8Wv1sWpaybLbVA
reCG9XUZVUKS0mjkbBNNM90TMer73VloEvMiXTK4pPgUjna3pAy9ocMJAYCHrLN9cpikUbYrnTPt
cixMxI7BwYNjv8ykw1Ayh/MPN44PgHszLjkRs7O4GCqzQ4/qnwGDK1MDql4wrsTMVZOkzFpYSXgy
DeiWAKKTSUdV00pc/hfa1r1Ru2Fqu5XHc/4v4LrUnMCaK/2H5e6bq6zoZkcsnRId/rAEFVakGThC
X73zyghu+hD9CmXtNnJQO4Z0XeKuVuxPxn7o1bweP3db3dhHU9yWVD2B4iTetjW29t/xvC7YoLET
4yAFhLypKM8/g05jS0039smYHPMX+On6sswlA2d6i5CA+OH4HlZuXCMiPZPl6GO8uinPnhxMSGyr
q/yPkkTbricE22iwvIxNb+xxMmb6raOrmtEug+wrSxd5aaqlY5r3ZQ/9N7LkUeJpLgstdb6FrITd
JYmgRMnzZzmIm3mNxNgNkKitsYrIEtBmcyRlrfxBrYi1tujRw05/Ms2WCSy+T0FJOSwGRA/q9md/
vyWnafjx7/rzDx1I9sS9RoxqkUxPc61jtPiWelj+/GSbmP75G7wM5sjb6hqM1UglnEG+/IkFqdQN
k5T5d1R6iwLS4lN28gvvDJ/TPyyrtGUtuAhuRuhw9P62vejtRNMp2vCxR6JiqIxGNAp3DKiIB5dK
nrAZnfREqhrMN66sK8ium/tGi5WWDPRlzOiU4htTU16ppBcsipDcFmw0S61bw2F5xEiH2wOMWROD
6hMEsa3YHjtF+o2Hq47j8tbzMKOrOIQXIHGe+D3RBcVV2ryqmtmSGjoaG7lBi6abUh5cfBwVEyx8
KvY8TWroTYyIV6uEES3Dbh8t81s2W2aaWCQ+k+aJ4tfa5hkd3ZwYOod2YKSUV7YOwbGY4BgZIEHZ
c2q+G93eMNLGOJWZi5FUXQUgH8IsdU7X6b+d9et2jsXpP3ruTkbzDDzMSOwGY07xdiZ4SXBx8Q++
UaKZ/W8zbjCOKRKMNWjOV/ErqrYO3wu61Ymi4n5Lez3n6w5JQij0XQzjI6KE853+ULYc0KLnP4JX
uV7JVDs0fHSA7n4sz94Axxy39FuQBTtzHXbpnUtBocw2NZHsGQpFiJ4zHYCPljxnhN8AykcpZab4
wPOA+d9HS4KYIfMGsGby0OnmpBuwA2P3NxKQFutZKEO8wkR3113PfLicGLgz4ZPi6oTWTq3EgzzC
2fYvtFHHzUJNazuRjfcJjPAL1RJEk+oIjNYKt4fzpwGkA8asG03TLUBAFpJ5sICFaWOdPjQomB0q
2srE6zXf7KHtgP6AITtinakXkB+4ErPHMh0ccr01nW5BJSeir2utKUaIZeygX7uaBZeLXf9yW9Mu
zpdoUQk50h2QM+D1YZuUMjmHWOVi77QDqNSjCHlFkl1uZ7ZL5QK+YohGikcT5IXgxxaWTc54jOpQ
1r/UvruootNhmRLAZ+sDaezjQa1u1fciFNymlz8EG+8VThNqWQXwT6dq37BTq5OLx9+8Uw9d45L1
H7YAoNx7qKDTX6neV2nmNPUWRZH6GPA0FwylvQ3bCN4lIWu66helh12EXl2Dc6eMl+95DvZ0H3rM
s/45d+fWrOeIYXjkFbbYtDHEnn/y7Yip6TioWV81ZLxDYoiEaVPDdNGgUIMpvYghwkkkK5vSbk+G
lfqG3brkkEc+DeY5b+2bXQX7Nj/tOUGK7RCyi8oDAfA61E+8QYbkjXbwrd8svgfDlCicxXmacq8l
tyQ7yqXwzHQecV5kquc92wXhdWIavUfMUubKMwS+y7cH6Icpm/Clkx37kGH7h0LWqcEpuIWnvN3Y
4Z+kbVRtJ/wJGpyXs7X2lEKvEhMmxrXE9++FCZlRDn6tofS1ShgLt0eDyFu2kT5kRYkbOKjN9hAr
vWuUrqq6IAPCCMGWzVguLjiSHckhwqrwsZz5SsP3fQWWDoveKAJH2SUFiO7JBRHHIZPhdaRulqir
wcIFAI1J+ypDGEM6iiDpKo7awHhmvXvl2/X3kzNUt2msHi1jExkwq5ViJriK0kxG5qJv1yKD0z6R
clK1pvLguVCu+bFpxHGjiHg7z/PzgXbKGAI4YVr2+drbt7lIK/kClRDP+UEesJ8NySzicJHWcJH5
dPhJevS7XV2MstGcIzbegQ8Z5FB5ZgWty/Sd+kJarBNJ74mh4NQQJ+8PuQwuFDtQRTqv8KBVF3GY
W0W6zi7xQn2BQAUXHHh7UZ0GER+U1d4DVPX3frYy+eomtYM38TwtLJjZo/ZfMw2Y7veKVcKou852
M4U0d/Nd1UjUDWDfqi6KnpoTw39tyNlaCNrguzbVtK1wneIjctBVCOhecfrvX2KGrEAdp8qXQEfg
MnyDF7GttikRnQOoL1VwRhBtPK242avnrLp78NGi2Aqu2LTtNAhdBl3hIvKAumi5v9FJrj099rkw
nK8If+aWhnMs9gmVz//SpPzHQ9KxD8PK4MM3Uo74j7tQI2Pd11655tCpDyqdnR4cmQ80J9qNLWED
vdO56ETVOuAWIDWh/jBlf9S4jASbU2T8rwMr2cBeolNMGFTryLsRu6FO/UtFxPuNUANzbT3OjgDf
xBWMAGODJjzHZ4j8yba4mxcC6okxrl4q+R661DVsX3ZH9Iqgwi08YfyWDYAJkn2lK2McrqasbQ8P
9NsdESTMoiilUsnaM+n2lfx5zAPcBCOZ4s2FwEtJc9H/pwEsMXlbtydRsHTomb0jEiTl/2UV7ZrM
fyOSbFfzdUUwlqDLT8AzvzyOd3lXysEz5whAz9xODJzTVFEqMMWKsRjTQ8q1/EGIVbI/xnqynSZa
VlWn3uxPh4ZmzApk+yq3e9p/CPyV4d+CeQCRvOYzpVhwKUzUEpkeOivz5OUFlrYQrB76qRDPgYlb
m7IRWwmBYQBZSSzpHxUNcgCDrdf62Zp/RIcaSUfjLVwYwaXO/N+g37W1kHHovKR6JzQ++oTUdVyB
U3jnX1U6JsM11ggnHgRKqKT5ewg73aSjYDoJd6Ah0xPYOSpop/lvkNiP7jxkYocMpcauQrYSP4KX
S3gz9yle2lEW2hlfTOpxrGuuKZ3d0IU+kEFzo1w79rGeWIwPnZKD4ctZCCpgNF+vxzL+s68D6qEN
dwDTLsn0G2r0WFg37gnPsrFrY3oNMxvT+mYKeJPLLbUOmAyr7ibL95R8rZdPIlZd47Bk3OnD9vc3
Rnwh6GkrDh7LqjeBTjOj8ELQ00BD48ufHoNDPweMF3v9+U9/agLTQ/SuM54d0BMpfBruL0Aee0s/
PmHs01KD+0Vkl7jTkQyd4+O+pfyHYELDYKhewr9xOu3M4D4yqGVpIb519q0iZbaMgEbFWMqFqTSm
XXrn18yp5D7vish39EdQ/sm0tMKvRARhxEWaVuKPX0ItO+p6A7mV0X06KXXChY9vARhYG5/9LlF5
hsn/K08YqsrU1ZnC0a1lzV8FJqwr0QM4Lw/+5pa20+SqEnOAONY49il+z9dYMWoCHkLxBHQQVTRT
ph03HUu2/q1Py3U8VMq3YzxzjMa5sgxVs8jwyT18RoyTnvGLJbMD6pGG1EFWWdRjc/01F2xH4j1b
4YOfaYsqU/wYanWKnu+ZLqjC10Br5K+lG/junUK564l2JI664RBvzJmBjEi7lYEzymaZDk8N3AsM
zOByRErIa6kTRhGk/C3xEYftFi6k9d0DO3AVbYLb8ra0AO27wNZDrTzBzqmgEgOsld8LxxsQPVqH
IH1ky6r4G0hUELnYPwgnmyteC/PYgRUEMxnCBp0oMQqbU+ZOITQMltxwiHzkV1GQtaj9u3NuDm9Q
TH6WMAnVLXSuDa9GVvOjhrzb1EDus5jfRjnov8MRB8BHs5dIzMtVGBfyFGLt+IM/OSbYpbCwZg/9
LAyDjY72IsN97rpm1upI8E2Fr+AHpX2jnBvGq35j49TQn2bzAMLbjabk0TzTjdQIIzLcqz65iKMV
Sw5/eU7p8YHsToW6fFQqWpqHtIwKrcy/6rE2HtWthLvevFR6v1qsdqPbVDX2kjrZMPfen8N5Fcvg
DTDG+Ii/uge7nS4V25ss0eIfH7oonqJ2F0jynb9owJKpXPp+JOblsB06HxsuOW7YrvJ33skgAWIC
KZhRpEZsj88TTmsTcedGK5Iv4rNsSaGPPAUKH4fsopQBhyz0xiVuPwE/0eHhL/Cq57PRpT9OB+s3
8dA8kfpbKOv3eEYm08JYAmvD+SsutB1UedWx40eHh7Xm7SF9neBCQij+Qub/2QJxk23FsOI5E7Uq
XVri+VIpEsUpO5ceMR2ZLpZaP2PAqV4p2z/cmv9PdoP0OfPRU3jC8ZirPECh7jLgvLZyO1NVOzmR
9NTOzdlcDQhC2AxIH3GVdTe0WVn67KnfCM503anzRqYZcMcM7sXZ4D96gdBDQ70AByeU+kcM/Yzd
ZAgZwvB5kUf3XvzbhDghkaZ08LkKSyx1ciTCCcPXiQaz9ityVQd7mODKDyzkJ13P8hyeuUnSRAF6
R1vcHx+iWL13GJy4IuWFHyum6yXFbWkPOClSofpNe3Kd+Zto1JVFD/A93quJrmrzlZYO1/PAZ6Wt
15FFjfyW+yTyE9wdEurmL33QQyoOlJ1o38jigH/tRNFYhY8A7S0iAayTIu2+wGDnYq/JZ6LTc3P7
2iJUbxzUtxtybouuArKz5OuYOKIZRwgAqiWHFJd0hcn5yAAk1Ze06SdfUku/8oDrcupMmAYAHMy3
4UrsljSxf8osJYAIivfo1xVr5iCrrzb8Ln6FO+8leu/QGUciJy/L/bakdZPgmE21zfc4lpjSIvV9
GdoXyNzpd61b25DJ6qOrGouzn8Z7FIIknj+Ez2lwoaeYrFPsx9mpwcWkEfjxO+vP5J3E0mSoEmxX
Pi4mTCiUg7d7zh+taLP/d3v0zkP0E9zOfDOKPXJCXcnH5tmc2jE5FTQQF8WbfVUND1TV/lNyQHvv
fVvA7em4jW/jXmHGspWg47bKRaYa9e/E5QlbNJOaoDjZe6UjdPPoGCE9dkzmuUKgsOkMfh+zjikU
VhLBQDvO2baop0yTleikFrMP0kD31Y6vt2G6xKPTvU3YA/ZJWT5CtxE6pc6SvvZlxS2yOAZKcM6U
lYhaoH+UIXJO4y6J29Ho/qTUG/zVcbQR/kqY147XoQTVmD6WPdVJrUQecw7AWkVNafzPAD+1XG3Z
4FXQoPHBRX8l5AlB8CZE5ZwjLnlaPkpCUpjJuLdJ5WaGcRlJqTEG3dy7/g/RM0ZNoCo+PC417KpB
6Brst4zyOJd2drw2gMRV+Dm0YI1ez2tN85bcX4mzTcIgxObStosctLQaiqLP8aXK+F10fpDyAif4
N/d7v3ZKDD+i6lQzlY56QSBFkmcyRikTqbnlTFvV4osBeLGzLnbxsmMzsNDFrH+JHO0jPyI05hDm
4DdIZGSPiG0LRx6tJJrkb8b2yJI4eb6vh/OZqMp8DOlIdPH433dClF6N0CwyjgGc11Q1vu+O4ILZ
9x0S8f+scphTMYWF7OgyWSBYPpteY8eoR7NPhJaityYG8Ci6p2uzyH1JN0/Es0cIDcggUj90C0RN
t5BIInJJkv7QqwsuUGQYz3QtIxbzTJ73BfKThY4QQcmqnc56M38DZf05u3Eg5RiK+YT7BVCUZWlg
sQu3E3ogZvzk4js5/cDSSF8ltv66aoJqjFhCa9UvAPRqk833T2bl+TY0lQ2zaZ34IE4CJHLioPn3
0rKhYxSNhJmixLRABSyU7mwCPD+3femVwvf9GCTDvnNbUw6JKvSmOHQk9PpU/fdA9pu8EA7iQkAO
vFVBAaU74xgrJxqIhqb8xpbkiHTQRe9mp+oqOjcCEnBhRHJhiPNsEjKPMyAV/wRjIERAHmrSsY7J
Uziu8g6BTgbXKFCR+bxJUEoaaHblRD+HtuWEs5bJB2KGX0dWj1+Vx1lOd4IluL/MB+1AVkX4ShSk
zrIsHJHtWdwTWPkrIf71jdAEXx5XHRmgBjbgDfz22EOZUQWDSQ7Dw4aGnjt0KcnDJzmJ9vHxS3CG
19qeEmKQ0buVICPO3hYX8yTapTZBU841hzEexMNOrmRKY26SBC0vmWdc5lPBN3DHP4x5bn79DdGe
Ex5ejkHTI4r+LmpxIdxPmjettmzW89r9anOYFYFQ70PTntkc2eGz+sLSfgck2i3qicXyBNpGLSwy
ZT8r7bFRgBqKWDMl2fdFVFVdJoHztLRffNM5uP/awgxdJmndA+bn3aMczkbiUinW+5pk0UaBln7M
6SaccuhKVORBdmOYqm2xMse2tTLLqVnR02gP6++Rbqn6YHTM7r1KHHhdsCDWtaieThIXwyrhG0wP
3tUix19Tu5Ym0cqWur1NNtfgY3UJDJcFGN1hpSRhOp2JSL561M/UyMATpyHpLIpPLyUHynGoMi9s
1E5TBcIQg0Hs/GmivnYqENlob1HGFh4luUUthy49gioreTdgZdxGF3SIuxS/H+k+XJj6EpVBEGSH
JoxsQsD8f2QFhGbgxVOSj4z+jKrXnJbmr8wUbqOw5htx5ITgsUTWRa5lLZCcNFADM3/jR3LpEVjd
GsJm/fkhiUGlJEjQyxMb1m5qaMt8AWvHy7nY0q4RA8E54yefApib+tTKl7iCOpfWpbat/hQ4l/kG
8M3t6QUEDOJVMG2L41srDDlgo9T0wRVALOgw0CJTrFKLd8fRdp1Q2OYy8ilskCriVrumLOi9+kTL
DbgmOfTYdc6kXRcLelcewPFQzKjWNcaCfA1t+swm/ehlrxwxWLZ1031Hlzt+5A4kCQnYd49gn4C0
+tdJcw3Job4Joo4TglBJBXiTdJLy0yaKBqNMgDhC4GnO7UPYV5IXDNekX6kIt7HcRzSY6mgfI5On
uFSjb71P2qQV8iMeDirk+uWAfstPd4B7qiPIwJLJeltIqRaWUL0W/y4l/PJcxphA+uc+HRnjDxnJ
uscBV8BzXzvWFBkW/mNBXx4McCjZ1gkA2ggvwe5cgK80DO1IzuSVxXgglFA8x0JVpBkY1T402zzz
zMJpv+qz6x50vC3sfcnHBvQ8xygXAZ4lZ0pGp5hMTQwjghyqcC7bnolGRCsJd/rGagYHfpSNcKWq
VnshDJr5WGfmTc4jaef4yofe01H/LV6ryiUc2Fab9h1CrH5QaAozp21Qf0+LfW9kJ6LP5BkLKdbT
++T8L1ruqpQ3AyHt9xF16uOuzSO6n7b2v71B0oYujrV77sxsr3SCGgGoTUIgUenj8t5Pi3sgD2tG
Xr6kE42Rw23qB2SInVWswdZNP3lH6npLlUEaO0dFYuVTld/lKnb57sLjiTv6NQ7Xe22BWiNJkIzB
mavZGfQxNklf5rWKTXWgSgwoQW6bEdDYs+zYIf4Ohow6byHg3QxPto5ggABPe8OaBgv/RI58CHBj
HYBoTqPL/4GMuW+oshqTUESirjVJT2eWMn10comqV6NKTnuyEL3FL8Ihl2JQ3DJOlvCWc+m2Zqee
3Y4coyYtXETJFHoOW7kno7ELvnbn7TutVzuF7FOcg9v60ST1tSrNwiKQzXURBhibAbtHRK8WPWgx
jZWLzwdtvb2mSS72EZ1ZFKm26/fiZ6+kPvRENVY4U2KcyfkqwwoMfrhDzGc902MVuIp1pBz4L35b
Av5KQE2b40gF4ikGL6Zb4q28fuU2p3KS5g5WFSWTacS97qjYxcrPcc/PutDLJyPz46CS4wrqabEx
LNLJtxgOml3K6188yNWsKSHC08qZ5qPnBp2DFT1csVMinDMyoCD6XEEN6+r7bSRP9W3LpggHeSo/
YUonQVgmx1FeY8DPhBguqxp+nIDEFWMk1/hfEMKvunpWwel+D0ntSkRmLs2QEDbha6a9J4To2oxF
Sb5izSwMGT8YF+A7aNzXY2T1GtdPu5Kxx56jMrvGk9s7Vubo1Hs96crDp5kFlydNEwu6I8YrVu37
lKyiLF2eWnIiMfeIDVcy/LjxXOyzQaFm6456/vMyJO2Sqo+SeMRcLeH/7UuVrlGWIulCKoaklRKM
isdjUFCN6bfV3LtfVVE1rWOzpPDTCLqWacjTc7kMf9mjBhThYnxzB1RmrGkhWPH8B6QQ3pMLwirz
sU3Q7Xhy9ZShZ4Xwt4kFHV4jx9AyxQ/3MCSoya4F2FMOp0Bv/1+3IgxfhqjMzC8kXii6KQf/eY3Z
qoRatbUVlb5pzAZCogkzcoeIsqUxRxAehB4lP6LvlmUMEM8EP9qOPZXrjHeopmiHkGm7M82WAYO3
N4NlTIdlMz5AAHKxkZ8PZAlLmM0utWyBL1WlSD/AbU9xobF0IfzFoJDA5eWB84+/Z6zXJiGgAP9p
nuUltnvIcV8asa1GXokWnHlgu/PWOnfEV6N0q8ar51xU3TAMKyCu2jjLtPGUCMtftGqj2AtuCJsc
NvqNIkefoP6cxo+S4TbLUFFgfc/OtW1qXlIZH2BRHYWum0gLPXWezzNv2AJvmwcUYNSSNcZf7ZXX
Wnnle42fqnrz9zmIJfqGQdgRzuVEu9rS2n6viPbCAMFH/xO+Q8h8dIqbFmISpmbFwfgdaigDrugL
2aKKe9XYCfc7yotXZslQBQDaukQbiuPtbwGJgjM9XSQIBUlxfAElN2A3ZZBBWC+VYibrisO3Smuf
3GeXiCQGhS8ipqsIXcjfMSwZ3uWtZmBU0JyHX9ce0SqhF3Kp28KD+0FEZXUlkLMZTjVOBqQPNYJu
vBy2QS20Combr7KRAIm2riX/AomWu779wH6VBNUU1NZ2RAT7o9VW4xBqlkXqN4eQ5GjMWrmryC5u
9f85WEUkrNvjeR8ESVaxMaKqxZW6ltJGipfGAZWDiRPPShKBu2xYsEJZzBAKc/BD7BvWZFTkKKEh
iXMIMd7PgTh5kZWjzwx/8ua6XpOsxylJYitZqmjAPZsmmot3cusCW2Bs7ZFg2VZyeljBVXUKq1l5
NZL7xLnJZm8c708vkGnjnc5oIWyJ3b1FumznI+ys9OMtSvvRVBdfPGr1yqxwm0IU9s+ek0FcdCBi
Vs3xYDdXDG+GZ36U/E0yUKfJ/oV3bWhArik72kZ66UFRJNXuxuSs4RASMkaT+Cczx+TwxhHTxbvh
H3caTiX8C1YupXJ5NHjYb+dNl+TkeQqXw0ICyCmFUrVSsCV5igE/LFcueHECDIpY6wx6w69rDcK3
jTlmdW3tGKYVjUPeBiuFhepZJsGyHnb8VROv7tQgG/wMTrMyTatCkvJ4QHJM8lhEIaPfd4qTSjXW
ynkgNOJGxJLt9KjtN4fjM7ZAP8+A24AflVrqx/m9A+GrpZSHhzKoRRo9YHG5JCgkC7CCQVxeHAI8
CsMccMMER18mysZGLl8OdvwRDM6eQJe559WWlK9tJT08px2qAZHQpmLeIsOmRKo5mIJLyKuzgHP/
kfvSfRZgIiIvafSfDECfuEWtG3ehUaZCR8J4MA2DqQ+hcnn9HDo79HqVSfcXFSnONmE5T7hMsuB4
iBugjhJIVQkDS3iSx1y53QJtr8yx3CGRXvociX1IzTYrSUS9QcP/k3Bt332LSjrV+K0Wu7NIswfr
dpF+V57VahQQpID0+of+qlnjgGIbToTIo2RYYSZdCiv3XMsHIx90NTOb3qZZDbwNHzeApmb5Hfwk
sFxCCnpuL88tBzYmWE6YGsoAQZcNfpaZtEzjHlgiwPcLRXbaEceqLMX1Uzbdo63pj5K74+Gwg+yJ
bi15g1xCVTCbmfzrMneERGaCQz7kp30c4iaxe1GCMFNyHNK4syWQBJnmWj+pxZyAuhP1hzpo8Hc9
aGRBbzrsZVnlBNTw07KX31Cqg/gtQZh57LaWYBc5IaktR04CJ8lQEDewBUxEYHNo3HVyQvH1Qg6g
9/7pyFQxsxEa2XtB0UzjFXmzWpHFF7r+S8Hj/0navI7sS4nUT2bnXsQwWUmQ99OsOjEABzPIa/L5
yazAtkOYpccJ2COowgdiEjiFAkFzD92r7vkPTlH6Nc0mnRY3BUl3EB3byol/IwAPJEHT+4cc9faY
lhofh6MgKBQVkH2Ahs5LR0GFBLFuIZnGlkzF9sf4SseWXBopomM3X9U2wNv39BkdgAWZUIVVoJJa
KTmHJknJBvBswkPrL3X1378xHhEpW5YmbrZBpINc4hT1IYGkoteHcqt4lU6nB8F6NhNAIQrFmm7t
yC9EgRP6exGDpS2f+TbYhkxyky9ltKm8TlcQRKiD4L2gX9XJIgEqpnjlw6lwTTxlaVdXeDNxl25t
j3evXRPnDkUONNH2RUAJ8qzl5qDSdmyxdrwImlV/hPCifF303MirSI/HKDikSKYUvem8axlrUCU9
0DZyGSBJpX4ArqEie2qgWV7Mt1zjQMS+IDu+t/K3ck7TKzsF0LLysIsxkBeinXPOxkw4WrCtgRrO
crzwIuZyGEkZPaq7o95jfs5yjbrwK825jl9INKQ/cEDsdkWEoB1jiRmJdydkSBXaj3BA7I2VSSH1
kbSEulCVrk248Qi/s1RaIQgsOhdeQc1osnyigHetM2knU04GER4sV4/LRj3OewyZHzC8lb8qc4BO
kpJnR/LPYKypaR6ftnoaDhp1SpTR8SBsPFzFEMc6XWGoD0/prXnaJ9Zt074HeGjPRl6wthEeVP4s
F5ytS0stUchZYSE6/GqM9ioEkc576p2dOFd915nxRlhZLKnkW9etnsn4FRAij5v731qwN3lFU7dT
WZKjlijCJ9LtbzkdyBXfdlPBOfw5/McNd2QCjzvDNqcrOlcYrKnLs8t4CPf5vc0cgz7A7ectBjMQ
R1QigcE9BxCHwHzTcKWE56Wn5+q1mLNLOzBqEWIGE0DXi7TBIB4lpeCqOHQNTTA949hm+HB7Zi0S
ZalktQOgoqY+lgoR9w3/Cr82YkV1tuSYZPoL5edeCi6WMixw9cUmyHpa5vZoBMLqWujbLtv/1urT
DrDxLAkLnVFG+yP+rQj4JRV1lbqYnMhOCVZn8m0Qp0igwzvep+7Ct6sg3J4RQERpl99pLRK0ueVb
1mJy8a1EJFds1jJf/AkV7VuyCJuDe1GnpxUVCQNMwhl9bsuKEJeETjDh56RssgrTFIuu/inLkQX4
rekqpemj4GYw/DBuyRhZf1OKuqcpsYIMWSfmFBdD1Es1hBigGx3dfbIAZI1Bu09wV/A6uhSEqqUx
IKg0owAN+Nn3k1RaUTBtKez3f7cYLIsXJT6VmmMxMaAL1vBl4HxqvqYjiekyemxBPEU1s2BmiJr5
rE0CGcmubr7vDJ2mmj/shFcLhdSHev2uDhJjg5JsVw5XkRqmHDDWj6tjPGTM7wF/lpsQOqDyissH
/llgZ8Xlrn3p05mG5BNBC+rON2z5PAxIfRFrz8lvlI4mQabFeev94JIELNg3XNZW8kXCI6K0BMPN
g7A75LCV/3r8W/4T/u/6q6hL4e7RmcnVzAq/Wkvdz7hdPb9fcjLGCjBNwgMJmFj0jqoO6yQyZpY7
mE2Wtbzg46pTgEWjjbT5wYucenbFf27+YFaT4Lssl+LiHg44k+5O0xVEmYHP8qypoCGQsFBVzaRj
BDeIBnDxKT0PMboMTWgsY0bbR7jbs+NiLBP3X5iIr0PJ8xEyHZwK+/WHjzTjKj676KdP0IL+t9fv
O3PEtXWamfuToDYF6jI4tAsVCrMAt5HIgsNNx17/UugroOVneITjtd17qJLALwvRaqKv4i5eva7P
J5N46OUrETPbBFz4m9JILN2LweeJG8eckyfh8mVzViqgBmg8wUIrl9ndxa0mJ+I0bOSXDd4RAEYD
gEQu0BSh2wjB7z11KupmuCPsiEE89lI5g4siN/qyhL3HmOwVG3mmiSZyMKc8b8/BX40+kvUu3y8A
5eIk95KCYi4vAfRG44J46qvjaygxz98FNHojs0uJBl+dcZSmWZvLLcQ+MhI4itOE60LFRuBcjFhh
ME+bZcFmA38N+g8vfdLAC8I+QIqcRSvwnkB6TNkCyb0fH9AoEkGL4ZWzCLSb/VxKg6erCGnrtFA4
QN370ACoDUBciU7SQVEFJMXnD3C1UpEnFyRqlfeNeOUVMr5JlM5bM2ZgODIxYmKMI8qoCK/BWNUm
Vi7ySVgBWolfzIcgabNsMrqQGkHd9jbHxPv0DNP86m2hTw0gczHIHcATj0jpGJSJ26x4y0ZpCAaC
koWmW+qhwBl1IZIyhAt7LzTiJlZJJpVQ2EiZu97FdHEDR6m5Jpj9PXhfCM799AZuxyjXU43HlpIE
qrEmf1CRhicHqwFmbK125zgjjQ4+5rzrtYbjWZWlZAS+cLkkU+qgX5wcLQJjwBzLtRrX3HWT1kpC
7iBy5wIOtBTNatA95c0GT6oaDY2sEJ6yog9jjZ37cNw1jBbsHzWK8PC1VpQ+M9wvJjjf4ZxOeI0e
HVdZPUbYjonap8BglNR1xehB74aewMg5Lad7T66ZcMyTC5uDAKaTm8tVuJR6X8vxLVMgIQPfIQ/4
m+ErE3ZslOw+keSntdf4dK+DzpV08/5QE2Ux6ZbQnIe2wa2/nUJ+O5QDy7fYUR15XZu8CT5QJlnp
rIOfkw4/764mcPgMwYvFOM/3Pg4HxordaVCYRNn+JigEbHi+QA7CsIbRyb/tqurwJLqpeFV9vQuM
ybdEA4JHaCmh8bOwwottuRlShHp/EhFR2JNCmyiJFquj5wrfOZuqqNK3K8qV/Qv1oP78HJ4xchf8
KjPhsF+PSch3W5LtuYsrhcMRu5mEfZiB4RDmYgMLztELFXJ1lf2d+zOj0ECbJa2nXvwD5rK3Vfso
3zXmg3BbQpiZlFQkL07SYTQrOXGiMXCXO8RDyW8eabkB3gkIrW+lRW2TLOMnSB11s3qC0SU84OEd
Sq3OV1pKAdjSJ5FEl+x9b3yHcwyW24WiNcAeFCAT4l1GrMZ9aKkSgDc9i7m14yrh9beE4J0qWvVr
GBgnXQRm/IgV0iPWmBCfkvM9nOVUmNLrCajVxW8b/WRbMD4vAGnTDwRuhAYo+sI9U0OFMhnZ0sZH
vISkfng7ge3m+5BmTDZ8ZE+glthJTco3maJwB7onY5I7IJzM1SNH2uKgFbr47tnt6B43ruB/G5DE
35JRWkjlhZk/gT1xyrmt/2oOt+uu97zIObwDrE3OQ0vu0mVGz5arjVNZMr1q5LJyw3/Wz2pS2QYC
JhZByWIp70toOHMTQ9KccIijKV2KckiJ7EtsKIwYZwfRaicnomv+JAZXvmBRmOUp3FhfUmZMt3yh
emea63phwCYghU5PV+EFROdhDA7ikfUZOE47E0AiD33DEBFxIKwBk/8YhLyBgXi9WMpvSV/fgheu
NKTGC8HUAsmUtFrt4NN5ACgkB7JmTzYPlr0hgXuipzUfmLPsjV5uHhVvEKSRZLRDCqTf4PxjcI9A
BFEsPYMvJjnXKwAaOmorDhRNoBEtBoMN+ElgXh6Z4MPE3xSIfPOi8ppZLPJXfuNlhbjoOFA73cmd
RSlkb9pLR3Q5sb/nrOTLCc2sV5YWKG/UNX0Y5gVYtfqSADM9NfbmeWfe/NNaBZNDPJlEmV1BrQS4
GVdWIReeqBwCMsYd2idp5P9BHZAuM38QpWY3CevZ6kW3NOANuHUXkCuVsWCZve9JFnjApMUxJRYn
Hvsa2cC4XhqKdKbSUH0fFzjvJzfNFxCC6fVsBepHERdpwcOS68Li1SMT34W13apJOX+zNCmyZh9m
CDAapytQ/5zEcNc5rLYUHJJReqeBH2IOnSwoEphmDAZvQMzRyEz6loWG8RN7mgeLRlVJjL97EKJh
R9E+UvjnG/kFFpNSK0O//lIbPGB7fC6/V8unC7Z55jGciryH/VkDUv4k3C1anRHws/ldjTsaDd7N
SBoA5/4vpx7jhGIM78VW8ccqLOrzy2ppYc/NMfOs0xLSww9EP65FvLXqXw3BBKFJNMDIoVeWYe6Y
evnCaHvkcTVIm1vmYUp2z8zPLLqHK/z54QOFVMD7MaVz0U/FKMKmCvdLcpH3AK4nguohqpZ2CvEI
qTz3OpDu6u5U8Bt7D4epPJJpOhg0VyGFjp5p6pkaVvMA3D81zC7gz+i14zcXRi1SfwWuleppAfv1
3zhXq0L/3/SRU7LMmMlSjyX0f5PCr7+s4KoZVksIdYyFwSuac3xZGlqvBvnQ4HN/S+WNBDRQ7Kbx
IQO+PK24KAhfpoFXwRh0TorATBxFa0dKTlRao2MN0Ui8DxNpfr24HVS0OZm5FtMW4VO1oWq0SJTx
x3KStWXe2m2swF+VSslfHvBXv8YTdyCPd01yoYSSEKVGziUsZ/9scoNsRWU5Mw6C/p5MoXbZ+sPm
FlgK1ec8dXa3UWd66Kgm14adNbu65ZQmQfdhC29rfL0gvBAd6tkSqadpLQbzvTCY6UqfJtyKNLtR
giwBWHiyrzZxCUc98WhjSvFChWCm5fRX4P1CDAjYWaT57M6M1ry7JYpAox/Vjvh89HEiD2xex7PM
WMOZpI7bSglJBcEpvzpFLR6ecbpgiywJE/PR1GZo7QRYD1ZPUAlU91A+8JLA/SaW0NVJq3y7Yw3b
Cc9pSy8dcbwEqoWjlK7g/5lrqJQxK5johldkFcHNBkApfGqdPrA3l0hSNxeAS5x/Vb3LAQnTeLEX
eoXfL6kiHxXSay0d7zAesNSd+djPIPjgKu39Lwyj+j5ow+IcW4JpplzJmYemvCvc1n8gKrrsruhJ
lUSeHBQnjFGxh3TF9t5dfFoWiQIsxJ6/e8sVRh3QpzoP0yKMHdu1OaatS4dwXkqg3FgA9rs28tK8
muN4IZ7uJOk7aYOsHyibfqE5a0CrVLpRRio0ODvYMuJKvI2Stlnz0PaIkbWivtREvAgnxGRQYclT
dpFqhwTtJx35ggIcRet6ocpO/OFP7ZcL8vvoMR/h/NfK8R5bXYuVLVwwAb0S3kjInP3KhebORJ4p
zHp8CyqTwba4/hjQIPfVMmyyyrhz40Hf9vSVWR29/P4Wy8b46BzuyhW1vJhHrueF+73v1395g41O
4aSY7DmztyAH0FB4uzkPsqMt3J12b7wMQnl+1rjuVo3ZTre4dtWFQYQySvDIa7LL/b3xe+Y9X2fT
ipAbRTwHFCbA2QFxZq+TnghDqSGlKXrQy5tZYBhz+mICo5NZeJgJnRaTQa4bhvwa//Ma1XySthAI
ZgP6HEHt2zEdtEenY2pqWCgY9Ea5uKz63oZodQbCGtXfASW0Ohdg2/BWFGd4f6bplpazI2v+YQ4V
l8EBFfEq8I2SXFEcvD1ZKMgWPshdjF+NTLt5jUQR1ah8tdy4dH1NcXWEOtznTKDeyYsE2HJBLhgt
Cmfr1mNa8gCLsBD9jGtW1qyKuGD08Zrjc3lsCk0Lz45SaNbvkZZP12Puecb8iB06JzFlp2T/0a50
pwDSwLDWDNt0E7IocWcUZV2iE1MmRLo1oUM5DeA5bsXyC8WxSJvlLocMCyrY7+mAUDQG67eoOwH8
QAd8RHPFLlZVBHOpVW1F6yQ8+npP80d0lwxVXEfqZn97HaXHy+bYxxU1veyfn5mKzU6QUL3AxTGp
AEJA23K0+z2miKjTAbv/HVYHVHCZH4cj0+c70f1upfKv52ERGsHsVRxFKb2d55jDAFThgHpIQy+o
eEAaIY70nj6on8foJ06SAExkIABZerqgEOtPaAZFrHF8Md43BR8C8P/gSm1VYGlSEcGNnluQzCJJ
7qx1YO6m4wRrPNFseGgmau1KR6WXe3vWszVMPbG4So9F2XXsCe+38oChv8R/JR2m5EiCCip8S9MA
FXxkFn2qFJeQ6w+bk4JzQY5yat1eO68zfEY6IavGz7MoXigvQYnaAmi9xckGCMxN8zDkOzbHgzJZ
ShMrMb0ii+ELLh1fqewZZL1QHUN/SAWIJXn2/7jeF0O4NqI9QSAvlesMvkS1HLf2D1DA2h9SfauK
/ULYmZ2Ft9i8x2yLQHRBHL6K3RNvAK1XFT+1VntNda742i9EEyV7/DAuIZqr8mRkXDjN7gIg5XE+
D3yO3/heXLn4GzzfA561l+e/bEuv6tpLV6hPkQ9ENfSvQKZeY33CzDS1fyO+Dp42twYCx9XwsbNJ
H1D2XyGN4PfAgp5Kn0BGzDLd/a/rU1sHEoaQ7PavE8A+/9Ffc7TupgbVevKZg8fbxMU7jmeJZNqO
F67IzU4TYCC7am8BAC7q+1bcFzoANKpWh9kagtUh3wVb0VjmCtj/SASJowQKodvDlbo5NkLV0aK9
2+QJg6WMjf2z10vEvaPUtLkP7wdN5zt0z3Pd2jdgiFSMc/r8EaIooehG3lVPCI3Hq5LWAe0phAji
QTVvTLdjqxsoCKgt55XFa1agJEqU2cfu6l1ARuxnfpn3BRxJe7sJ8/840xFenqDhQewfjqe6u8UR
0NbbKPwJrc+H8ugdNbSyMghcHieLyCfl4zm85+oEUTfxAnZv8rFL1yqJEEl/YxasBnCI60VZ6Hk1
fDZXlEhZERGs5lO83p+3qnI7BUcO8CNcWVWzb3yqwSGPXKi2e8XA5plYdPorsWAdDibWcquvEiS+
Ok5Y6n3M5qFO6FHGCJtcRVV7aTBIVXQIHi0dHV1czkYzpLp4bWHOQy/w8AOYjyUYZsn3L/lXBGjx
Gh3xRk8QSzV2LhoyPjDZFXWmIhjqyHhnf8vH/gh7a77pceomlrcY2uKhuWYPpJuNTJO1vthVKbsF
2OzCFxvTp4MJWlQ+vXWoj56E0WTOfDYK61yy0hWKBdGDBdELwxcJahVC1n9gCDgjmKgzSU77jYlX
Vt4KaSXawBAQCpGUWLcE4faIRvTBkH79McyloiUrBNjN+ufJegQm9t52KxloC3jAFpCR3sEdcy1m
sxjcovP5ywhwal6U41kuDGm+RMG9fJLs9A/YLp5U51ULe0qJZLLfuxsFFKHQwUISLWIXGrThWc0l
opypYZxUmmAWYNZrLV8PLTPZsUF1WDw8G1dK+Y4AFL9EKM8GvjLlgF//5pMk1VZxpu5MePGqFB8I
HSvyIfy4Qmxol+cTGzOwHBLsrAi/AM9OATn4ZrFeKV+KO7FUtTIMFwSpTVYJ9pmopE7zU6LfheAw
V14U4aSXVe9O9L6b5yjpXuVrpobEI1hD2KVzOHnyLeurkGMSUp9suzVGIMYPacbwICbirTn0Rv9s
EjtTHOoKKZNK0RXtD33CmPLoE7DScccclKZG8z/DetPhbHEggf6/PiA4dPCNfDUdoyr3c/coL0Hk
gaQVMqtP/VqAbmrCm0ZxPw3s3jghe9ZT4ztlR4DSEKDCesknZyWf/NcrTSH3DeY+5t9yTVBdCgiI
FvA/+F8pguCu5X/jHaV5UqBd2hu7x87mY0RCbAVXh5HFq/yipHRn9CWLZ1y8yu1WKjtggNoDGqSO
wtGx0caom4Kz0fQBUB0UfLiWPiszurz7pmlbZWQojltV7pWlfI6C3wiaVSzAjP0r266JWcwYPHmZ
r+IH97q0MvkajLX5xvvJE9/V8qb9OLD+mtkrJawVTPig1afqxyHWVrstOBLIB8vtSl349vTnHiXg
KKzrDAEUu+3mjgHglBncpbNFHWS3QVgTMpB7TyYczdQPAgAY0dflx9LAi5nGvJGCnNeHGbozq7GC
7XEk7iBo19qSNCIiGxYou51edF9SZbW0dEuRzRqAY2rWNqng/A48uaZEaeqAAUHc1uOIdoXHllML
G7N+aCzShqDM2/TyGu5VXM6D+YaO4s41Ue6TITmeVWdwEUYY49l5YPP58Tj5FKIoSwyg4QEjv2Ss
D40wkpAUbeIaHc1JwJvsJX/OzShLEJb0NNKcy+3NGoHgekW23QyfHycL3BIQqKB/p55rVWi1UWqZ
CyDJeEMeqKyOraMEsQ5ETF/4AQ3rcOkXHQpwbtYQhc9TDD+4jV1v8D2a1240yDo7EM52h7Dwngka
u5OSJoVH8d+wKUjm5GNsjg32vNnyuURpduM+LoJqXvL/PxoRPAr9LxnzwBFxgzacQyrav5zyAerr
YaTYpwyscPxEyGY7sZFt0ZjC8u73dwFvEkmazB/kjAAfBI8Y6cH53/7NVHtvZ0HfflHdRJD7j3Jw
LbilcMeemCIhwjQUBXPs39eQGQeHlV6PYpYceivBgxPGORQ4vbMyyl10leH60Vh45tDaRJpcUK3z
lQ/eMhDfl5Fue5zYQqiGddTAHE0XfVQA31rWUqCYkBH6lQi3YSWC/k+eV1nHuNKaBQ00Tm82QHno
DLQehAcrKZZdM1C9tILjYBwMJ++UHnWkQLZYup8cL7XHWciIDjsDd7u8ZWkt6bzCjci2NRo8LspM
+HnyxW0ATOAdIMGvCMfuZTw78lYRvqS9aLGhVrRYN9KZk6MB4GIW5z3pkLa5PWBf492Ofd3AV1as
f0dK8nk/blod30bYA+OOCK6YbNxKD7V/1wKQSUDvwRNivbDkJT38esER+DgTguxrLUZk7RVMV+5W
4jMk/qdRfjgslL1QaX5udetWuzE2SUCLTJrHncrOY4AvzEy5gTOxo31cbnlWFihl2fPnm3QcxoGU
raMIHvw5yGEmG5WC1UZTUQa0J+rPoqgeZC4J3svKP67kvvzwKqzONHzWwGCuUY0DK6P01iD3Y7FU
4kpn0+NzAa48qwc1upZTPbciuxdjanqCRIi9OyJtZO8ZNmAJnqlAIN3/YPslCHiATItIcqbdjKqp
zTk3h/3tncIkBEuUJOOwJ4A7kogqq3KiKD/Wb38dGgIbF/tkRJjbasKs+XWvMipXQ3YwhjY9+Kbj
1gm/Y+hKykHZctIn4NTeCxGFm8Bpcm8UWOODDn8v8CQlFZWsOPJanx/OVxCHBEU2qHkynEUhx28X
pMrNZvTIve2+h3Ynpgp2uJcL3F5giOwVds4j1a4fIfH6Z0sis2wAznAgehW0KcLcuBcNNPmbX918
UrqcF4qjdxgnBKMNPIQEklYqW7P1yjCRYDGY5zf1O++Fk7BTN2FbukjJI2E1TfPG95E7PWVRLAkf
XbYoKziGrvtFXTuurhyXawK+kI9i/4Z7hwfdFKONI8kiWhcxypbn1cu8BiKZ+fvmi4DsPax4flEd
COj3HgDDjn7piX+sKa4Un2zCWZSVzdCS0bwWZFb84IE8Fuys0UWPZ6K+iRen4gSld5schWWnviIC
gKXGlKhBfKltDzteqBEOblYDZnQx97PCB2hlAE6+I4AeG+114eeFI1XEpNVcGqZ4P/qTzpTjkf0t
dbd+OPvmu8C+U4r8++pSYoiTwlMWYbmX96pbI9vMJX/ogKAAu3nU/wsPhz7ZC3gfAW8AHkullff2
X5VfEtVmZVLv8mFBBKySl1/quxhjnd7mJt+6zXQxCsoqxHR0FtIIxbcZU+cjKMaZjVKKPs5TCBTp
Fd95VDb+ntkIaffFTDB92tykC1+txEJAEVvEzFlc/YK9p744soW35Up1c5LIzsRqnHaTv2CLFDbn
OUrijmXkA/RadeMtRErBg7LmPEljGUAsCMWUWgGc9xenOK1kbb6K++kdYaB/WMLw632SIN6myNky
0olMaBYFrLyOktEyqXO0NFkr9tlPaHJUOgvgRDDU3/WqZbL7tJKyQFKN51v6dqmy5NJ+jJpnXD+H
yHzPi16PbZbm0Zw0ysVyhGjD38a5z6UFp2Zb7I3A9AxpwSw9nD9BjAniyP/2wghJaYYlh2eOS0nf
9qD5w1gAfcdhcl72SsqhlQ7NYC01tYs1kyhiCWHYN3+M3t5fI2PLc8LJIeAK+ZECdAsAKshod6r4
oAORm4Lul0CQNRIg0rvn2oZjA3PEvyLfEmI1oP2NLK0g0iosTb5LEReawuSzvnKRiCPgFOrbqVoi
VZLYpf8FSN7geRVAToaUM6iPL+oHVtZHTmLn0BSogtGEGdlbjTGPrJZsCZ5lphT2HUZ98rYm5d8+
l5btACINDmwQhQB0LMk/HmXE3Q9mnGm1bv6125RHycWdIt931hbNPWLmKjgnXXiblDjHorR+ZQfq
8jA6jBO3BPyL4IkMi5oGefAnOW13mddsX5yfr6HbP1nGiRRxsu0ncJEz3U1cFf7wEt5FztX80n7R
diPSmz/ncL3kbQMe7wlb4Zkvs3oLDE7WXaXmd/tejAEHHro4Z1LXsDgX3Hd310tfUqP9/LZ/xHeW
vgB6wb1zvi1atn1jFDek2W9qLOhjPJVHmOBoPVWwEq+hGIqYpCUUkb8EdQmNp85ClW01f0sdlFH9
E9N+g4Je1N4BzcDWd9dtNhzvSlh85QRAGQuBr/pIM51cglnOB8oHRJO6zdpItrzNHME8xAk1bTe7
GQtmE9p4xr2U8LY9S079P1KkBROF/d+Bi5wZNk4fnHEgqABrztrSQwNW6FecBDTuiJtHMNrOAq5E
eEQmiYjT3VwAFsNUib0T4ay1X36BXNoxur4jFr4OW42FLaA1EN/kqUhR+KiMmDWy52j1wdqYHNpK
cY+a0hjHhDP8tYkL/ed4xeVweJtyN2qOKgpClWKAw3zF3BmGIstPte5obJQpzUExZqrWw4KRs0Ur
NXtcv50gDsgVAGfM3bo5h3qUKKc3fWDEMeQEtONKupOzhK1D9Obg7lhIfPV9XCrktMXPe503Hqu0
fkDNfT631YWHppxH1bCma2uuKvwDvp8on7uzP+P0OW0E+/4E7X85bneEtFilwKTnXG31MoAW9eBD
nxeXFzEEbq/nHPLWQxBXtrLN95guj1Cyo4N1G2c7tDNICB3kc7vS9rsyndjPOrt/49Z7IF8xbNSe
ooOeIr6bKKLPMH5BGKabPB5RRhAc7CQBjxIIAixBcALj1kxFSktOIw4UO12aKULDqhAxDjCejRMs
i7dCr4B/SSJ6vU5UykB6UVSDtZg/AYWCP6U457oMadBKvate1lIZYuqkeFxMQBfGcQ7si0iyPcCD
FRFZHQCeypNn3GGWwjYx6K+a4OPnnIv420Y9PkY8DRAiDLKkc7QwnqcDGf8N/O/bksSDuWsYlwP7
P6PUq2zAqXdR+3cK7q8C+wVpMbiG7OGECwTAZ0ubC4MczHzly+2BwrplPq8DpJqM79eFMQM0mhLl
8dgKdIiWSw1lqXUnbJoad/7LOlKAvYq1SyuCJ9Va5aQnrWLO6tEqIGiMy3inlwPxGo3HPg5MVE/D
+/2uTE9G0WIcaU9l6Vs70qg15MHSSeyTAFNRaiP7hn0DaEGITqUh2Yz+Xyu2UKaLdXkbtBw+W4un
TPZ4mwpW2nJaF/8rkvUyd2t3ZDERaZHpgETof4ViHfEPRMgMZJ374w6CCqBLFS6x1JzBqmBhj1e1
wtbU85g3M36u5Ck5kstVjUE00zGZ544QeqoiPnjeyRXHjUb2egPOSZVGgIuZa/UOP61qmjKu40m1
Ru+Zxz7/WZzU2R+TXl3UGF8n9TcnC+83VxaISUtf6zJe5HRDkP3c3iRnPfPuDCao9La/YTI7TFXq
QwQUOljy1l1oZsbFedPc3199xmjSmTp8mO/5J+7cX4EqriHA++KHSGY0bi+rP9MQHPIRahsbBOir
80/cNbc59nzzQWGicCEwSeS9rrxOn9ZrP5x97o0u07WvELotDebyd/oi28Y4HfZ6r6Lxv/JtyFoR
lOp3XXrwmLv1uSEboKnkNL9WPS67L6C4B4uYdngghUoWGBqPbzCF7Df2hf1muysk0cUKprDzRkM1
9ckquy67Vm7LYTYlmLmzxv0kZ5D2kcCdGJ+DE6OAFS3OpnB4rgHAWpTvmnTBCFQ6kx7RZJR+Y4us
9wm2Kk3kGb6cqYEAw+eFZixAG6FQr1zQwJKB2hdtdFdggbHh1ZrNAQfxJlDb+K8l0ZyQ1n8wEBlW
ArAgaoJvbTL/Y8tYMwDxldu1X084Z8TLzHzOkvzp1J3fGz+fw0/wdrvrUP9h9XrNVcduOVIyfN6y
L1ITN18o9eoDSCXVuvZ6/60zfTQckuVa8UJf65XToG0pavWeUJBPgQXOjSR44q22oXktKH133VeO
641oZzR3e/HLCXCXqVMlnbosWkw9+ghoOAR3lIPy1Ddrtbm88GyyhruCSW4OXMzEx/Rjtcm47oG0
ms8SaXwz5ymV2KdRS5zEEbUL1kFE0Lz/XgK02k4YT7NQAe/dwNp/+s9uzbgiShMkfp9dBderb2iF
kaqMRDNfcxSPNB592hcSOq2kDHnaGBk8h1nzYUen+s5TkvErwgOBw8kM5GOmeFfHVt+PoBbVzg1b
I9nYMynhuIe/Ljs/Ux0OsyrS1LKonVIM/z2wKIIVeyWZlhtzgcMJvY90phicbjKEnLY1gy9uLOVH
Hy2MWBHslYpn+lq2mLSQ3O8h63RdA+Jx0SObP8fWh+amBnWo9UJyQywLWg0nayvCD1LdAsFlu1oV
hOE0FlolosIgbu7c6pybTwbgCH8Oh2dngzkuyuC96AniknkyXSsjv9jK1Tffcwk7i8Ows5Ivc8oB
2wog7zo8Xw9GWrtD/NbANFfE8SodeI0gvi8redDnTQVrrth8dgGCSZIiV+5Vqo0Ntoyd1ogLBprk
Ahr9sjN2yP9XkmlPgPepMqCrjM+s1Mq0JcqFRgO7GSRcM7anYxrCGBr6VSisWTW5J0EsUijCaMkM
iCENTdRvc87cuH0h5o0EF5gqWyjIvPPIxZkmqmQLiOtOu3SCdO2T8DiuKYBcRzGTYoLqV5baCheg
iy+guCHCpKJ5TiMAYdWjCH0MjJurHmbzRHBuCnGZPohN3GhfKLwcVotf42eIQ/1/6s4I65jP6+zM
qkHThabWiZ6YLht5tdaeb9/qKCn83XfML/Hkt3Ih8aQT+M3KOzEY05yJo40NTeUKyBCZggiv3WZf
qWZ+xDMWkQbtVDS29b2+AtUiWta5/WGSAQc34i0LkJWtJwATEMPSgOBHIiIjOoLghr1s7xtV9daU
NzbpyIFN97k0Oa5FhvV0DmxtI4N1umJO5IN7q+XuZDoo1+mnHBz79ru+st15CHle5Ev0vnCs9gP1
PQ6UKErujRD5n1otL+uRB1d+ho3M7sX76WPukOz8beQuWMZL1uKJ/H+blUs1m2JZ1WJux1MVJAq7
G8uxPe0z1ECSxnhWYQkCG42yzqm3/5V8FZZFsktPI9Eh8RcGvzyiAgF6i3JPEXTkb9Jg0ABt9PvY
vupgoscScbklax7lGJd5SueKsSj5kzCv/O4Dy3b2AGcJRY3RBV/faNkTiApDzeEVgdQfPs6IoZ6S
1yJjaub8NO/v2xwwdsj5YrWXwR4E8F4mpdxCE/GiQMRreRBb5iqKzUHI81axi7s/xf31XBAFWG6N
UBl2izlkOGYdTk2V20kc8SU0e9Xt5GQ4iUxBBQ/S7W2Chhn5zbgYoprxm/mZClMz/dDTMrUGioBv
WU5fonKNfbN08RYx7+Q6UJllVQs0g8s/mmE+2Lj1SARG2W40ertU7oTcrqv2S2/1PzxWaNl30eLo
mifB0GSPb0zW3gwZg4/vs1vCvxtYXM616KC2sltifVYgXusNX6Sha5g2FovZ81YegERTPm3aHqo+
daT37f3E4FppjaP+Rkpk9LzQhJ/8AvgjGC1DDP56Tt8ufrbD6G5SnetI6pFyrMJhlV2FghpiQNtR
0AWlnEtDHvmOevuA8vOOIEAnwmRrAOPtDsTc0b/fBoRJozo7gd7L47jDQOcf3/5iUVxkTlsyH/2o
qpciHvm1qcUSkrgQKdOGZgIrzJnTG1qZp5rwdRgyE4TW7l+ZpQLW5utTBQRCDdc9QnCzlj8gtcLq
pTHnHDKSO/paPYFQnPwKAJwUXFjYt9Yl/LbZmQaCFImNiZ5gtcId8lrXm7Esx7RjgXI1Al1YslMK
SwASEamoxHLvRIptUO7dO3s5FqZENPqSG9PyGHRopyPsW26b8gjCCp51ZddaLH8U3dt+K6KLOtSp
t9iO16kpgk2TKcvQ02mF11wcQrsSiHg/FY9owncDz2eMcH5LJkZfobU40pAg5gX9bB9kDskcviZw
WT9t6yEAiq2zMbme3ILsKuTR4XgVo/FhAeFl76B7iEsLLAW5dOOR+C+MS7MAug7RO3kjq/GiugNu
KA5Ck5Rs3I5U1nWu7dAGaBDkPRrxv2142lFSzlRZu9c+LKkkacF1jwVRkeDAr/GGtQjLQwDIDXYt
Be0cdk1DrgzcLAZwBgYycCsth/6P80ooLySrQCrsZnW5YK5O50XPyVib4nZtznwM6dJ7d23ia6++
pyEk60fh1HVnGR7RuZUGhFpjNroYRQHcQynutXv/wRW9g4m/QTtjaWEH0hrJOKydZDBKOd5wbaTa
IeSkMV0HbxDkrUG9bDiiDLZLSLL/LA4YEPzHg4g1WWy0CrUETrRd0U6vUWToTgiVA/aL+hVXh/h1
XpdWmoioYFZG2WWGsIPjv7t1FbajafBJi+ksNP71dViSFUb9jaUz1my4LKquEwoAnB9JpL/FUNTK
z33zgSO7Esuf6XYg08fO8LIzIn+qU86b556NZmcIgx3plLzgk7Do0lzEStmcEbVcA+5LW1QtGaiI
s4PsILA7F1Fq5zxCsxVfZdgaccOMftdUVWjqIBCA5cOGW7ZDEhsMr2ZwbnQtotUYcNlOOPFoVpa9
sLSW9uU0nldZQCXFe8hGiH/4vayy3CE0Sltlw1LTQd8WhWOp6NMYx/ywH/S2XkXbmSPMkBycHZO2
CZ6juwYA7HUy7mLFWDFdQocAn9vSWsXDRoEeaD270Bnx4Y5T8NlkJcaALiXHZ0dzm1yGEfJep63M
3jGP6GvYZYL8TkOi0+NIcOmV76krMYozMEcMEprF6jc6F9ImGB1n+YMKUUNOnwE4psklWaNWAjKk
7i6CJ8mN1ggPYWnXHPuYIWe7dd1JTa54joDCPzxV1WyecyT59CMqZSkbMg2+HT0DrQ/7oUcNU3Su
5fcfesGokLOBk+We97hZ52GcpxBdKQHv5lBFJVBFrf8IsQ3BrQMl7UDHS937ISxH3XLyldnUoevv
rRhP9YM3kHXeDL693uq4xlYGEV3UAWBburoBSoP8VlvYwkBGuhgNR0BZQ22HAvq5NjZ8NsnDkR0F
wSd/LQaQedC6Js/gpUi751Vx43Q8tOaI2CminOpm2wwivIX1WmcVfYN2N4bP9an0jKnUZIIoA6gT
+WYHfA8tHb8v/LB16Qkdm4geAtjQtFdgQkH+lFCxSIgSleXKT9h/rdgGdXBkbe6mv0KueFJ1v6mz
GGo6etNuadY00CDpXWU7MFrBa0SyMZcMKesiK+YV86/P6GGCSzkOIDKPGtdjgs0kgE2mEp3pg2Ep
bP8PfBz4LF2PPsL2pU1g0MK+73S31IrAGO9+fvf3ozqW30BI9FSFhjASOplkx3XRWxLuPoZ54KF8
uCHH96bAoJq4EVyONQh/HuANXi1AjSlxinHvb9JoV3LNmILeTcse2dkoBg5S5U8WGcrJOGf/bN27
PVJmYM0mFd9wW0d3bSSDsu6F6FzcOnNDBLBiN1OWhWngIumDfiQ/6h2JosGk6SrlFf8dFsiClr3l
KGE33v3U/j5hIea/eIu06H/JXvL9b8Eo1k0UYkGzlWmpmBsPPYUcfqIKV5EJttZpg/0IoLjMwvam
Mtk4+JCN6SnZq5KGcWQ60+TJ0xJsTMrRboWowxnlrV0jD1ybtWwUWs7lji3fHX/q4tQchngPP0Zc
W4PdNDEHPr21/FKD+0KvETmQrgEOVtYAvOGFYTjWKoVMKV06elMqWdHztRKcSTMVhMVT4eBbk0p+
shHqQ/UX06Ze5JUIseZ4cBOeDtj/2xkP+RpAu9KjRW+oWuboY4jd4Mh4n20dCGYuAZwG90sP9i9Z
inxZMfBb7m1WPMWIy0Ef9Xw/mUs9CKC+FbfqG42G9JyQyiUlj3mc3yBPh2Bak51qlgQP+4U9TsxA
IoDCbsH5+4EktfPky6T6uBWgK6GbR+A9t3ixsqX3kuX3k2xrZPugMw8UHyTyF7k9qYYKhCtk9uMZ
hVx+N1OPy+n1wFodyKQBxQuwxw7wrS/9OL1N/3kzoq9XmucWom5PE/QVZrDX1UxLZjK683s9WJQK
84ZnNmL+9YQi3fWp2kbaPmO/KBBQtXk3xuO8sWVsop06rWxGrl8cN1usWTvg5Yg5XjRmO/CjCByk
v3SdNiUMzdHPZImYX/AoTeJEuewGH6+IUX2CZhQJjNc2Nt+jhHEgrNrh1F0VcSC7MpJpkhz0exo8
dSGNNIMUzCzuEH/mNTooWLvGn+acxPejvq7LRBksF6Mgun+BNuJHI2b5DXBD+pW2gZAjFJbKkasA
zlGjqaTqpubUKED9q/RPGPLQYJhpk4ZHPqQ33Su6ygeVxmPKyNnHbXez+TkEzApU3tRZFeEBCBAl
V7KXRYdHAzc2C3wdQ58HzJsCFYcRoOpoI94yN+E0wijHuV/NgcwnX1bj2pSzyMpuSQ55fvdMgrGB
s/TgkBQeKGZjNQhID1+GykKFLH2mNWuMwXqj92p/IMN/6cZXuqHOh2Ch6nXRKr2k5jZyYGpfVoU8
8Zfe9y+GAHVlRFfcL1YF2uRh4HwDQbTW1wvPg6ln7Vrmw8KbhCIa3JgWN/EX7728J5kekRCGGWgN
aTr7IzsCaF0xZ/gjjK+qS0mWkEkZ9lF3hgI9QFjGy3/yxlkYY2amsgUExcznBV/haffF2yxhtG3t
eigKtupha5uUvk54ghI1QCHlVhUVePJxMg5yXwPLMTRWy93MD4rcfFeuWRbvcGwtZXf4y28p0jNr
B7KRKETaYm+FPXb8C4IHQ4mTIp0VcNw72ok4IJY773Ubmy08/pPE1Ea1UUvLeXvu1xiHWJUWgrMr
Q2/FBoX4k86XhZfgffteiUkBZSym6xDahnT5p16eymf03C4ARkLJwyPK7vM1yFO80N7gPeDToAsS
AzqwNV3E8dCt/3d1F/c24leQJMBmEN+zIDpMT9Gkcp7LLhPgXWlAcC2Pp5G9/M5ud0rkqVlDGaLx
SeK29koUB+O2aN+TBu7doVQc6DlafK/hLvLAFdYNIPYoSTaxmZ4m9w6Gn+UvIlDHt1Ha3M+d9dAk
hYIxd2vGg0gpRNWfFOMrVwIPbF+a94ACjlmZhNHy96AVzrgfyo7IP07lEZ3uKC0nrgu/SZEdo4YT
EeTCWO4P0fC+oPcQMat35RYa9YuA/SyRbSpc3dp7hU9v2wc9As3a1mtOR4dOF1lNELUsxB0ZVQd3
n4Q+3IMtdS0ponlu4RGbkEluV/vnTFJ+TytDJ3o4mMUx/z7nbgtPotI/I8JJfz3/4XEkmEdLc92M
Gv7ekYMYn3s7ERvRpXnBZ18Kt0Rsy1ttEYIkb1FFkvb+q8X93/5tGhLs+HqsQOk7HNxuFed49gi4
3GtMUn9aZeJgBld+8WjEGCbhTuVSaWNNFbVcbjG6opUllSb3L1zYye1j71eltgPI0u+XrvEZEvYG
ACtUo0aGgRxuU2Tv7TDz0UaCQYkXRfIlEH78lOXDV3iSIuDgDQXLbGlRxcmhMxKflwPb9ADu+zSb
FsOG0ZX/dmk0RRxvsI2eXPQ/EnuJ0caysuafQUB2twSfpg0qP5RDjzOjwQRYkzkzeOq/jMV0gFaB
P1QlBVOjYR5mWBw2xmu+8pYWQDjs+x0BqRAdOg8CjTHkOJQsnozb2CXl4yBfi4w3tYEx47PmUkAo
RONUYxZ4KnDProV+mcCi0Oz6Qjo3ISfOiHUuf69s5u8I/qJd8g6Dv1t36zVovtGEQnxyVS5lkUH1
pmX7EZFZlIGBeGiM6qlNbKS0JKwjxkjCM0W7Lt3aY5pWgsMvllcT0RUDC/9ibIBuTUuZkpjRKu78
885EfAEisXMnIKJ7NQBKng2GNJkyd2mZxTQi66z1nFd/YtacK9BMKuggJi90/3KFA2MrCKMQ1LwO
cTmEatFM/6agwu5yibwH7lGZPFcvytJDY/qYwRZ6Op+hAJ5SQHlFF5l8WogBbWtxWF8avyHeJYsK
XbaUaNqaosGCjxndQJ44os8Hc8Tf8m8mTXd6DJshfuxshYfD5vDoV1RZvvYQsbqiuidxpRJqEFX1
vzwjRvZsZZ1rVeJGx+FYNcE2H9Pmq3jUBXbpHC9Aho3moOHdaQLOfp+rlUQ3JtEvRm/BC42MXUJw
vShxTdAb/6F2SVCaMBkEN4+2rytLng3nv8Ugon3tiVqoATSWpZu2fdi5E6FwRGhb9tCaKkKearOl
Zv6lX7coE/tmIHioNu+WQdNfR/SC1d8tpgyPlRHyPB5ULTCV7W9iBke9QzpeixDqOLYrZMAbFse2
AhjM3JCwy9nFDLmvEDLoxlfIT8KX8Vh7sdcSWXGVuSwfMTyOzr7cEbnZ3srYGxUuRgnyyQH2xAkI
oCJgCvx8bGybIKPWsEtV2+/0DCUaR4xk0Jw2DC6dQCX3le51HhXVdmoLMcvJ8tlRAjjVdTnlMFXl
kJ6WAyw1Z/vvOLJvHUh5saQ5/eZI42dxvYB/tA5QMZD2zh2vk+pLWLCTr/sirL/ukcb2Gqb9kiOz
GeKnZSO+eIwwFiohLC7Yu9kR/scWmZOU4CSFRlT+8vpZff8iXmDOS2Ncxzr7XzWGVwsYXXCbopkX
d6aKcw5lH2+F/uzRklGEf0mL6xEXnzkGRVVo6r1YPMHENca2PspalNVD2P18zUyX5uWR3OPobXHW
XGQob+vfX9mi6xLbOkV3xwP20nFVa7CtOrKG0zYjGLgMnoSSMjb5Pm8z8YB058kXCuFel61SsRmu
cA9Fn+d65zwUQPCQRmommQ7w/xX+mYsYqK0XGLcIKlz4XsOR34JMiW4bSrMkL63MGUFVZFaCQ+lK
X0NxVEWjINTrkTbfDAg+hKFl16yx4CUCQLzAyw0xkwllc6axohRrq9Xhal2DjXDZjaRyn0CMECQK
IrD+qh2FMU8f3unj3P2jSWEtFO9qJFDjMOBbqHg8iNa2LPG3hwwUT+p30ht7YsMVFjMgG5d7az8D
0BNi4Z0JP9kPHty2heFZrztpl+2QNr9UzVrzb19qI/RVsA1g1E4T1DLHcyVoG6/Rq/USsdzzzhxV
7sIGdxXIT2iU6f5ME3GOfowHiDAU9vw3Rn8NRhnJyyygK0zE1ng7LzWYRsO77HX6TsfT7/B43gU0
zn3a/9aOJX/TM57mNkyuOX68scwrr+RjVkiOC3E1MRnhmo5uaiLaxakiVdCN5b5t8q2NgNeINABn
tTUXD98heq5jnmN/CyLrMTLMvlTFnO+LvE4kthITeJAUPU97h5BSQDJApdvJo3haTBvDH2RG3MjE
7FsNsTGmXjSaVo1P0LBYpyVpFoicJiK4dzGGiL+X8nN5Z/4FgyCivwDAsyIG61ddtiwWgYDs/VVg
Bh7EoiyvTaGAgzL5LPiEJkOudOwNmLsLWHiew7R6ohX3EDhG3C9EGsuuENUwcJQYzHu32G3bFiHp
RbkI8/C1KWB4FP73I0KAMjQDkitZSWRzZ3xmAT0Ofb+hPNOzml8N7VU0G+pqwzWg6CPdpvQYSuyX
A+krQVfM7tVB9GtDbuvK3TA9kWLkskTYWkX1astj5xiXaVtnz77xMFAKnrF6N9k4en1HbQ3AMb/+
BQQ7s5Vqkp1vW3z4367QjCty5r/b0B5oj5+ch9+DrOfIUYtbc6PqBrA+c7DtDy6EV8No4ryXMRHi
QJVq+B8sAxYhR/G6jO840yg/w9GprJCoz5xJR0Ls84zJMYF4ZRwJtxrz2lzNLNLIpUdCQ15xd/wb
KICqBKsP9FtoTCVOINTISN23QeiFQiXHXlLElELUQ/rENe/HlweG1mvnsd1BkCMQNBsJyV+85C89
9dBpD4O+uKS9oAvbsdflgiclQap4vB5lEmVUL4cCJJV7kSvPMDyFGErrOsTyrchrvVK8ac/sb67u
rV6f+xb+TGinxToePokLgQ8kvZAUX9IfjN/Hfmi4jkchNWXc+2tku1424tzGp0QJCjlGDRL2C63z
4GWF4cHACt+6FGlgS5FUM/imMseFm0LlgGWh8E+lLdlpnc9k7lE2/rIcJSO7RRoNX7Lu+EuQJZj+
3Prlo/iM/ijGarDlwBf2ucQAcwY2/BWVnST0c/tzjaTDdGnoZj59i8zSv24wN9DjDtJAdAFFQ8mg
ENRAVnwBI3As3zeNe7yiJdf5qxrmqD2e0SAzJFjfQbbzd/6mQLI59LDjZO1287RVfgmpjfxhDyPO
rnor7vb3lnk1sDrlwaLMX6QdNx8hn7BiIP2nsMQTt/BeR1bqmIP/jfHHXKp4c7BlN+JLZyIxBYMc
w6fPYf3EmUOT9Y+D5UNQFmq1xKcH/A0dowNzxqKLMqptogG24OufQEEajpD7GWyvuB5yrCoVdOru
wOyxo3NwvPd1H9tQ5mff3/x4I9uwlOupLDFlzDHXZTMmjRbVb2V25oR5HLoMFZvCbFC9RBUohWwh
qwg0dcoPmKHlPGQR3dbFHbvq6JTA67kDwJLV+YiJUtDNLhUE2zIGhKOd8qz2fX1x5VuV/7S0myld
zsvD7gvZkaH2ScT8kCFs1zp97ZVgoxb0mZuS0G+oeL9BqXWxra9NT6oV19qNxG1PO5YhqyPpO90z
1lQ3UW2iUFA46CcLwsT8X2oHU3hgwqGGOShD88B05WvGkF27aSJbO7BUqOjtcM4I/Jel13wY+r8u
h/tpYbZeSr3EnIG7RPtqiM6SLN5nrvz74hkxi11gtqqSgNbivSdoM7adhn6LcD7n0w1IeMFHCKxo
9e6dwD5KNOXq6/up79qAg8tHyHMFUJZ9RXLsyclwdF3F2fpKEKt9axOz650nUKNK0g6PYAzdfPcU
IAgmljAzJJheDiKwl7RAyEbKC7ybPsSbuDsYBWX0nBisaHoNFVzDF2/p17csR/0geeRPE5JYNnCT
cAh8ps6dYmaK1PAvWdSEB5Q2GBU9xks3oytxPcrYnzlyCck+pJNz4M4YSU716ADh/Tn87t2lg/tT
lFeTqsOgc9XuPLMrNlIo/LZxpS8K0HarTna8s37HVUAj4NyyG+dUAUcywxg3uzgRq0D6r0oaWUZv
IWHUYSx/Ol6puocyDAwSvovfZ38rY+uD4Mft2KsEAeI/n6tpuzDjm3ZEp+pkf+CfRspE/EfAXj6c
OgIPYQ8nvf/y/CJ6UvdD+MRXqhYEkGZ2PNZbGP8gi1VwyjJrE1N/EmKZuEOy03mvB2aZsOGJwh8b
B32wifQzvworgK096hzG5kelGoyYFZce5PM5XOwPq2raC8tvRs29ZKGzYn7NBStfi7HjccrlSjqd
j680H/cqNZIoMwGbnlVW1GzkWc0aZf/3hJ9IjUGfA6i7aAhTUgoWWs9N+6bBQBdW6ZvApIH+pYgv
tC6wnZtJ41so13rZlfNaRp3QcYWskT1TRDeAhSbPxAVc6GIICvHuUQoEDeDF0PxNpygMQX1wn7Vf
8KjBjG4nJ3tQU/3okExlqIP2L3qg1p2yprwke73EpFyZuBWINZKfA6E8ufSKImKfxV9pGYiYtwo6
rzUgX4xCNTyX/3bf4MD5HRqj3FeC6lJARtDCzJTfO0cRGBVmfVuM1zb48xr1KAl3mhYszShB+719
MvtKbqS7u9TcYpE7zOJuQBviD0X4j0kxHAAg4NmOWad/r7377xL4v48Ym4W7PPGUpdHt5atOBDFl
r3j/lGTkMyC93TnVXjaIHO6rUqA+CLlO51F7vNk9Xbttg98UPSefhs7ZTBkAJiJWHnZ109Bd1zCN
cDB41ghaDT+8SMSkLibCKmL32jHtyr8nb36PS65brmjOjcVSnF5uUj6YiDXBUSyTHCan3guuyiwM
fu4PDw7g5EfNxoJONo/BzVzdqkmyDXLNVhwetsBBpZ190NNe8Kq64+XBsJdJY1+lxyeSOHmTzSlx
R3qtBhaXEahGBmqrbUy5BTc50pqYZ5pc+v2aqJZ5FjI3Auch26ETC3ZGrKlVSGaZFuWrC/8iX/2A
KHYVYcl8Cfz6sa+GELfyPZxSNx90hKxh1DuUAfy+GbtVSGZvVqAQ04xb2UmZz7tq2sADCPmI4FBH
9YcMrAq13Qmq2sriUfDw/wXYzPz/MZjapGMU1xH/B3sC7DT24K5FfhxUZoSaOXOjvurKNv7wWoWD
RH8f2XAUbIXXrk8mouUdEDRUDN+5il7+641n6bJjTgKLPcjtAhZ2v/kcmwoosPsS/pFrQ4C4dOL6
YpLdr1tL+RE1VA32JI/651t0h4T5J5OOR21lN7VOe/iS8JJtIwfrhlJLi9TefwFkj4TwAUMQKQqX
JXKqhB6tO59vz+xJqo0/OMQ2FYWtV6BxD65OzqPmVxld2LYibDzBjmeA2AvX90e5oTdrN5W+QJnp
1Kzy3XYLDHxOcqqA9kvf4KSRoyCxv75xkTfM/iuYt49jnUz2JssFDUOcgdY7UCrQiEGe+/BD0Oml
TkEu83gN11q6pqfEqOTfGbvZjePEQ9v7+qI20yVdwBtthGNhZKRXcvet0EJy4gX4IlHj50bnnmfO
b4/51MY1DvusmNTgttjP0swIirRSKa3aXtm/SGUjAOdaFnKVxWXgtkr57RwLAMAU4y/TQw9FfyvL
XbCefco6PSmkMf3nYu7ABK8VMGmkWqqTGAnfbzkEU5Sgg0XKFDtWIgKBp4GNTkNnza4WwRp+vHma
aTxxZBKyNWLNESpeZssupz9YzLxUTgijCGOSCBB6tncDaiHHXTF2Z/RFrgMZrDQ3rQmnLNVL0njx
sdNly0uQEnt0rPNYj6rY8Omehbt6TblPZOp75EThwED+3TNPFQ7qXcynI2brmnsY0kBJ/M89kmTV
MhMzabiDK8koBmKmcTDB3bDvH4gVyBQoebERCfWsufJCUv3UGrGRJyCyj9g6sJi41l2EWsfw54qJ
s6/RM919JTK4YV6M0BTFWX1n8FzRVsK7RvCnbjjJpNIswbKiSWk+giwLU6KgkROPRUPnwvgew3hE
ol2NzojT/99tCtUPVrv0bfqEQpXXlsLI4c4HSMAdaDFSJfo6YcMT/kjB0lOoBonuldNP7nf2WMn5
WWvGW6M1wCLUdlOKOeJqTKQ53djEPuggdIPqT+5UnHbem9WsZWppKlRzvCGLWyxJY/Zxr7FjC1A4
sdwEpsOwKWsKULE0PSCKvaQcFYauNMgRhFn5k9oT9Cw1sUE+4N3AblgHqO5TVnnGxNAkZ0Y426ht
KlF2vJmjW6V48f3U7zWD/hp5TKsdYuIfFeiUNvDwQSUT9kwEIQzf6F179QhjwqBiFDpS8DpOlPkx
ysz+Q0uyJ0W4MhjEKP8Qf4sJwbLhw/NIUry5j92TwbvSy1FfghkIayf8det/6KGSgNhZ5Ivltp0g
Lb5s6IiTaKFXF293fltJQHRxZHj3wNGO491oBhyoK8SR86Y+5Bk+vOjRUM12I0+o0j7mWx+8s3xe
VapM74X5cxBZu7EZfIWS6M0t+McCVXUElxWWZtsQqeUbrMckQyLx0so1AHpIb2yOAKDUwpyIIOVz
/uyi4h+zQ9qcff4OIWz6P6YhhZjV/AcmF6Sa2zsU+9vGakleJNdLVL0xuvHOnBzt1ebqi13Ft1V5
gVjblfPiITQg1NLl5DiGwO9Mms9OBT0wwS2h+5rWBAlzXs7wv9MIWsVMhuJbK+TgROh66ql3gK7N
a+VWaq2AtEj/5a40SwZhAzRrQGQ5dCYd0TS9X6Ke1rX5lw88QEQHs86uu2gAiwGw0+mlm+q6V8oE
UpL/M4AkVsmbwCu2iyI5olwQLJLlcHbrYMutCjkxMz7lzSYM/8F6b2qVd9QwaXNpFBXgiPgThX4k
rjO0rIqCZYAMovNceL8xDjj4PphEo+ZB1JV7NXqSa5fmzVKG6Ne9aP1UhLsnxqjZhjgGOtLoUH3t
y4LOxr6O29z1EiUROWc0+34uOjBs8ci52QwBy2pNf/+FyHX3qQqBrLHiwFpSV+hQbXyHmWf+4yLu
+xV3BA3iwpTaixDv0EmP2yWtVLQlg4VzpuYFA6N+kwD7XKsoeb17Qf1QuzcNEFHugF4b23kz3PUK
zf1Z1PR406THDX+lYaotPR/w5Oh4CgXSrtVzMPLDsFX7j2n2vyO05it8mt62ElizAjGCs/OMvJmq
I0FZsr82fzhoc9yC3LXQuGOauCAxZkSpRHFjw2bAx3W5wvkW/k2Pv9OL0L9J4K4ldMWgPR4rbjCr
KLtQm8Z59orzvrzozcrMm6kspIKTwwPWR6lAgxTpxJsQ/Buuy4b9ShyH647+9d16qwSnIJWANeF0
58fWXR00jYqFMqPv25NNte0exi3mVHTPyBtx6BVwg9h+BysSlh4F1a2xpjc3kM2FYB7DAwHRNWYO
YUeFoyA6YFyMFZaEyi4G4f6iRWaZraZK4RgmlU7KePCnBnrVVxE/JV8SjL0Rpr4S2jCIY3+PvaMc
JeINZszyiTQvPyWu0oL+BZ65NehgBaoLD4MiS9rPGbcOH80KinCCGsAeDdt5qI1e/Eg3Vy2JW4nU
l1csZlrQcXvKzGpwYk47pgbSyt0y+pvXeO5rnn9y20rZFADG5ou+DDQNThIJ+Vs5g14zewrh8vdF
ZsVEXLB9D4HSkK0QN6yMEy3FXYTUITpO3RcaRBCdFEaZ6Sj/Los340lh2mAUbKRw4W4Q7p9tzrgC
mCvVy4HwTrwM2CuwYOJaIneJWKf49idY1s7EDe3It7A825vulx+3mSxINulpbIcLyNI7R8Iu2hnd
3Tj//9F6Xsf6Z9v+PzTEUT0YL7arRF2YxIeWnBBMDCbitGJpoZ85R3yJQTOnvApM+1/ShNfqYT9S
iKNvMXZqFkr0EPHYMeUU4915CoIUxU4kxM5QyagoOGQGGooiUSuTr04XzGdOai1svr3mmevZORM8
QnxXmiXQpSb7k7UVYMyRpiZS7YjtAtnhWguShWrFRydrLx3JxHNbCiyTaRyzUqW372DufKj0rBu/
1sYDB00IIP7lcHyp0Q1mAC79dBoU+t9G5HbM51JTJBmOZhcfcXCGRKnnobPgFAKB1Ra5Li+651mS
WiiOmZxXV3nYE/k0MUbY4NaXmHTOB3FJj2SAEmMcLhv1omloXJrEbf9I6go4VmzDnACutvcGMVfN
Km2EPCCBO3MofLKnRxU+WALTVtjWtCe0lQWjeIsRPmQerqJTR/RDWj95CMan5wqq09LJofAMWn+u
IH5BUmmrJ/jTndVRuuWk/ovavw+TogQKkbHaRvt+fVGORnTyFvZeW5MQ1G5is9w7qOrYI8P9yzAZ
cQriChXpgfvdAOQd1JGIGwb+kk7CLzIgEi+gZ38kV7JH+6J0cE3g7iyWuEAknZgYMwYFp8pn/trC
scWLY4ROExRRA8Mf3RnDGoxv6NzMTcAwqkNfx3FK5XsRWhBP7j39votf8GMulZ43K6jCfIVOU79p
i5gTRyADTCzYWW8/NLsRfy2bP102GkZIE9f9S4JxxP4KehSnGHpFDlEH0eg0ozoXYFkfwapIG+x4
t66ZSraIBpHTZVTsX3uiSOX+IkL3BbChLNPwX2R6evAJQkRAVMCw78qOTeqCfrAiVaLgOhzp5eR0
8zBp+T+QXFOUsmjqM+ktQTg33jjImFb/nvadDZjq8xky0AuRsLEX5HiGFeNT6HD/HnTLnQFu2H+J
v9uoVbN1tjnKrBLc4PMFDXlIWI7jtrFBMr5A8Y13iBFQMp3jft4pw30Dn7x1HtErvlanjYSckUp7
fCzdokSIPAppRuN6W5JksG7VylewxKH6xHvt2EX++VqHHVmtJiCQprgIX2nc06vOqY5ud5A61PY6
LqKAojGTyR7jEm9QtKcjeaWCJky1rXUc8boUvsto+PqMM7FiTqv7H3feQPCka37k8yCaOusAUifv
kKu5nFm9TewJoKvlFXCZKhC41HlFYihgfEbkE26AxFVL3beqThAY1TkNLvOfGcNuTEkQ62+GOGn6
eEKfsTT3n9GNx5wsbshGlqw43/ANkaOCdqf3RjYdiG+U7YZvgKjqIdvZiHroHgo2CszYMZi3xZpg
Bu9ZBDZSAVTco0Z/M07FuhvjfhEQk7uZnLze5Rmw6G4vaMajeT3R3kMKgs1u3b3ZqtihTOctlzuG
tFdYLH1g5Sxi9c/W6bN02fmtzct30c4vv2tl7DhGoDuky8PGHeW16dm0uCCxL0VYwjeXjxk2Resn
S/NzBrmrswVbhjPfP07XkeIG4JVHxcgVtsfpbDpt83pkVB+GZmaVskUGMzPz8QTOZKYvHtYWwcqp
HXCK2Gj/Bhj/rQa2hu8L9lL3OWFe1WlUrw7Yisl3BIhwgiC46hZf8XECQl8BhAj++UCXsvgsm1zv
AzEd313Rr+hIzRYJJp4Arj1WTtUL3+GGie5BePj+akjcpkwCeIfZwjBXLyptxj6DeNYTZ+JhxJ9Y
QvEezxcFgB1zfWAW0IIzZPT5qpRRmHpby0N/RR+vPcsf5L0CQsl5Mkn5k99A/b3pfJBo0zdB5Goz
w0RmcRrH0NZWx51uK4pa1IWzBB5pW39ruJOa4vzFVHL70Wd9a2DAq5ClJUz3G+aqJw6uuls85lCL
iVsUBPbmprNw3AdjUE8zyoRLfy9cSITkhB+i1Upfky0yA2lYYnBbfDoOjyVVNrxk2T354sjRlZzt
VHoL7YwEMm01piBRIMpt874j3wO1uDy+ZSmfg5e9AQGkYR1alM1nlzxGCf4NzROIofDF358p39uD
lTp131biFTSurCoJXgb4uZfr4rTsrTJPjvQr94tjabb5tSgU7OBDaldKU0AZCuWwxExozBiurh1k
wYRUgM8PUNSAdxF6j/AffjCI+duDBI2lBheU72YYvKh4uGTf6imze5usKdbt1R7XTx7Bh/FxsqOd
8aFK1+lnUOl2f/cD/mg0WbYPuPy+gHZD80oKS8cvkp1VMLn6ZbirX4D0KiLHa9j7c5n9zPKwSR4G
u/C17GkFV6Q4q7MbfnbPtHFnXq74ts3uwdhFsiw8xz/t65rAzPwuwia1ETpTXnRUlhOoaWSEttMT
zrnE90kChZ8vXwR4fceIUUK1tmZeIO2ttqT3YahZNtXkytY1ecmfcd0A+vO2KRhCb57EV0+0+9Hz
qBNlkQi5nJ9rVEKMxe2EM5HeNTYCvJ9EXnPwSevRaCicSamG4Hvlv+UfpTPlBkM6I9F327pULR67
Za8Crrb7UO/I1/O2ANKF3f7CDlO+VsHgPHFcY4Rjaqa4EeYI1xjusHlWG4sdVz7BCfjVf1M57bCz
RJ6fQcYNpxBtn/qhcCGTSWWkRsXvKESfTKfk96P+byG2yDm1flBog4RRKqNwW4SuzGvDIofh4eQu
O/dJcZ7FU06WJ4KvctT1z/kO/hTlOwKFwHvcRCBeyvVy7JqfnTUqI1TSzZHTjixr3Axm5o3xNB6Z
+ybrQXU5QK4jGLlJsc/10eQU7Z3EN5SlyuYlHL1HnW8V1VSQb2oWJjwkEXDyyYYCiqkU4fOnyplc
oYhRgyZf/w+sCA52tnzMQ7SrdiZfSL5COJTosu1C/kA+GRACiRET0r4Nuc6DIyNGwKyosMmVfZQz
wg51Xeqx+DytH1h6SsitUeoFYpPM9qIioIYZmzXhFBIT1GNo0gPnWsE3n6ZHc7r2wWxuYnewStwo
WLHx0XOF7Bv41n/QTMDpbzD0YqVRfxsH1vY+YML/MyYf4/xCk/2mrCJA9lejGs4N2/WskjiJ87d9
8a6CDMSlxi/Xjr0CMffje/cE9EKWNMFN3zJA49OkW+Jubks0wxDkowXusQQcAAQiIkU9Km4LDUpW
eVBHzZ0H9Rx5kHeGB82bG4vaWIvTuEeXvtcBYnSCsblftFV0jQSpC9T38REyQjcS4QNZQQ60pfCk
68jEstMpE36C2aSNNtOvoA613Ew5MU7wv322kglddyLa3ZA4UtHWNtaotpeUlGS0HUMx/Ex3SF8V
0Vi8d3gdFSZQ78uCjMGikgqH0o5x+qMZh6h6tBgkydSG+Wmkh8mCGiR56dJrKFTtbllqnzaM2f2E
oK18F35VU18gvU13fMiWRdwbmskFYJxUTrtJRLBIMEcao0n5lyexI1hPGoOIBYpHHAKqgIIQ9HeN
B6TW6iU3aWDr7l5/G3f5agYIfT4LytELpkAWFq9ZuVOjEgKw78iT3Q8KLB1ph5V95M4IGJ2Yo9Ib
GxI78JFSDF4DybtuzF2c5YvIiv64XQ3nl3m3syEc0nGZEA/ceUCz787sSlhLTgDR/oSxnUy0dNfD
k0WWth0OjysC1tveterkUikM5H4zKPcPpxcdqSxxCygW/DYtMmyvWkkc4sINbwjvCAMMEEgkCglb
KQ6le2c76WoWZqimQOqu2pXKqk4xMgVkNOG7AzcczUnpqOfb9RDAWOq267QKi9/aRSTrRq9aMKLQ
ssC8Fl184j9+AcOZRr5BBEj/rLaJRnukI4TVH45yJzrzT8wQlCvPvm/1X7IAE5TGgkiyJcBa3E5/
sBHDiybNGLJhcxl/tIJ0iJNf8rl/zEpnnSo4mgSBsqUK/C8ZNO4RlGKXMGeEofyyKCN3UX/KKOvX
9S7Jzlll9L/4t1BRYCS7Xo6hhACbBUs07Fvw8rZUpUJZddDmBShEkqkkHhlI0f5E4SZG9UDG0m4Y
x0D2MoiXAfPbSe284O7hMAj4+PqXneOUKS8Q4bAeSPlrl6jXV3YnXhINFzRVkVK3CKCKFtJitjIQ
HhvAkUH9L6/cTwujKWX64Ff8xIDZvZMU2VUeKCCIWbwQq2yCFNwpRuv3rImD0f6dyK8rN76CYVqa
rNmfX2twJ/kXt5KVvNFBCIheKt1rHVzWXc+x7AxbzkAqJU0wIcU4Ev4i5LCFLe9wbwR5YzkQ1IQp
QnSDZXaoEUbe9SM5UVRBPppHra++32RhlByviwLfRoDa7/rBxs+eWaSAHAVGAQQBxlWOyCEuKEAK
oxkEmnG87oE23sw4wuZFqlCSYIREp0rRjE1f5zuZnUGAmzrONWA7ESjJEzac6gj1nYsJAIktFeY/
8VCv3W7vKOd7ynM6rjdIn1QhQPrSFdv+iBWJhi9DKY0evMhMDNvfviOPm+Q1edQges0J5fFARp1G
bARwz0OX7seo8d9v0ptj6aWuWlOa3UyREx74IEGfuhKFW9Z2LWqd5JLZx/2OSwrdKoyNKs9IK0S0
mRGqMHNyJYrxskAc0aVRsMHYehVjb3wiJb0lpd3r72LrboMQanlpuWObFsyyXx0vpPRH/GreE9k9
5TKh9CmNjyPjYCJrrMT/gv8lUXHqiiNAf+HlKT6R2juQtUzdbssilC0f/sOf4kNYfja8mStZcHvz
Z977zDbjEfZUTCQJJhTzzxCaOv1tAVe6grarwCpq2w3m/xqI/yJ63DAKUSRCQQSqAZth5Wpmb+fC
kKyIxameF99m7Ny7OpZibcuPJlZPu0aDbzEPWr/u0GPywnw3AtmU0ObE8ddk0onmoqLOp000kfVg
NPInOlw6SP/IXKYtAfPSMqtY6KOQlLmvPBqcyfnA0CMQvgIBHMDubW+63QNZ+wTePHFgeI8zyVUk
p1ciOcpz1dDTa9Gb1bhZ2nJvxInfOexnXCrsK9oD8BEiI1oLVpR1zzYrv5BsOw3tvyaaSraWDBB1
GLj0pJ3JGngMNcqlO4SY79Lut504UrMfqC3LGiGazTMe0QOiovFZm9SVTtRlZ1vkIQn+SanbCqs/
bVbhdhjOCFjsjIk80dL4nfxGV7dkWgS3rsa3cAmJKkQC0uuWO0iIrVvWBC/j7XOd7lYpU6Avh4FK
15HmdTO65lh72zwhlWbs+wEb4tX2Rxz2SYsmo3N1KevlQtl7w+vqV/YBk1NN2w33odzlUKpDM6hT
OoOWfZ9kPdKGNWx44gybQIJl9ybjLwPUKyx66biWcybNFA7bt6oz/MXvMYnYLgQUgHwla7yAzhwu
C/uWNKHEfo/GhR1Ce4DNR6bBzqIno5UIR4t/n9pmojHvtsiZbLWNntKV8pF4oigxpqHOSiGYIv06
OwZoo/p3RCd/t2iFF96HWd2DPKYbxA5cRFDvcPVjfIY2b1z+G1QqvgqVMfI93L4uFiIgAX5TC4BO
U8YmA4dbsC/ldxcG2KgDrdPPdDM9NGWfUoLKzHkTLlSVfJkezhJjOA6XtXHIOjQ+eTtN0yMUak9Q
3pEYGVNgUgv/Cq8r+V26/H7sEphJ05zTfzvEJHYspSPLQ8Bc0WWHodWub07Q320xMPCBkeGfGJgq
tkcT1N4C/o6N5+Sioonv8uKMFrK+EuNyDOhY+iFepD4mHI1DDWL/se4ujs4fDeuypCCpoDiJT/lh
OQrl7d5Q1l9w2jzg5l0iFZjbGe/XZ3IRj7mPt9IrcBM8oWUbW1UNR4t1P8W5ShOcNA8kb3g6jfj1
Eg2efVl2saXycown3tg+44G0DtIc+LRN5Wxd/6nzSJZsNk/MWTk3e8S35jatB3CGXCW+3OuP1nHF
efDdHagyBxa7Tgm+trdog51G/I8iu8o8dr5mbmMTN0Otn8bl7ze/5giO1w08cik6Xh91nTB3hRq5
1I7O6Nj7NU0rCB2iXKNI0xSkFNhfd4aBf5zquRolJQoZyL9tr5ZiAVJFsRwljSSR6+52o7sfFkD3
DUB37RBm/bUbkCQGWbN94Ig9QgaqJ65noUSB1kMhzXsLD5CeFfy9R1OUgLBXvMAeEYDzDzf+/JWZ
gjuFM+9BzrZHu1Vlz9lKmj7SaxQEz8ptDz5qDPZztQ3lYBdB0EfjT/89EY+89fy6riUp0ZDJjEL3
CdQwwm+Gj/I8jC+IRwW9PSIdKm5cj5Ngow7AqDO5Mfp2w8BBkRqBD4TAf6rQM6gp0fWySVGYJbWV
NQkb1NgWgVS0yBNCnxTt92mlxfW3zHsy+EXMyA0HqQva0afKJPzBKhL3rOgRhLa0VdZqVGG0KL4R
MWAdw/uDWIzP0FPyZGPLu/PcADIDhi1AsjThXMWMe7HvLrp+y48AYLK4qIGsDdxcTBGlSp94hurh
PeEqu0zWCiAdorRIcsWo7z0twCtumL3Dd4Dto4w+LqaDOYrVCzbS68rQcKVL1il0LEwZ8K9uush5
qhoMKl1dKK0kkpzmtLCNR3PbJwGA7tr4KbhDoVb4fZP1nEe5iHdjU+dA8y8QqlDbtRzVauiX0O16
shbOSoW+vsOqjdwhXgKi3f7qOLi7L58tkh9tuNG73Fg+moIjnnJM27DOPqpJFuYYa+Vji9XUqa4S
0zu8i4Lhm0FBu+pYxL6satbdWwVBmw9mkJaRZIV9LQZ+QLsXKiqfY2sgjubsal2mjY2JGTCd2qsg
ZeMs1gOAHyaBzf8WsG0TjF5tkqtgZl0dqzA8yZ/qt6fubHCZkKI5taPNXTwiikdLZ2aPDz7FepfB
yYJI9ePpf4gK0gMWgaGXFcAYMET+jB4iBPEOpDyfhoyq27c6OFx+mjMfSm4dzBR+vdg+snE8l6dG
1soaMMKtqUDL+lcyN33107ri8sloKWaa4cR5b/glObVIz8doqdzYJxB9Q1EnwK6oGyI1gOsHYaOo
I7DwuUyN9K7ShIdEpQI8ZtAWtudn5RIjmmX4ARIF5DXtbI3qJ4sNzxFa5MMIoNroPAfSCB55jOey
Thf8E3HfWhW7tnzmtYKtP3r+QGsbNgPmnjy3H87J/86MpsVOoXgvRYTe5HxDZZcKQ42CMI8//n+w
d0E9VezC+Xz936dN2xs6rLtdRS2qKChmkaZoCIK2kEW3rcZU8fhN9w4EdCv1TohlLpkMQcONc1zy
IY0CO1wM7XuPEqumm9WtP379ZqoyqfLTfE8vUhTNUkay7iLcdZ0bjr+7jFuFD1FhHJqyuKoGjrig
z8fF2vEuc1qP7TZ27jQ5Py6Odo0qFXLWFM5Dj4WRKl9MuhCtmOtfezNatOIn3TRrAdWMiNosyYEq
4HYWSDlw/rxPhCZqpTVwST6tOYp1EJwog5i0aBvNozvh5BvuCKNzBxZBFJ6bqKqKdqdl5iJDA2dt
YEXNQsEJJXWeKhD9Cyd4MQA0TGMaPUXHmzhsLsvJ4Rbuhs8g0abJ/c+ik0IDOywcDa8D2mrdP8dk
2B6UD2/ogMstHNynofrdGuFtZMyPfmlhTV54RJXjKQ+MNm20gegY21sUxcg8NDHdeaCbQ5xIdXo4
mSb1MwTgtC3re27OSkQ9n1rBQKEGxwNELRH1SEPbKp43eQB2pqDjTnzlz0ZCQZ/j58NMd4lnkJio
w2LG/PLCRyk+d/k3Xk5TWiEaluiuAZhvq+VujbLcM7kbkTuf8lG17Wwl3FuvX9P299M4P9Teq1rw
N06rUL0ChLP0vd+yZ0okTRX6ZUkG3vC75NiRvn7ozeOrg+ZcKhn6wd0qVkrho6CfbGVBE2+BzYoS
Eza2+bW+4cNgORShQlnTMPbHOnm+rbKGavZv1cZDYs9iuZgt8uUArYe2nW6qJP0SKwMDif/OvfE2
NgT3pHbn+xQ/ULcozymWCoaSdnTCMGD9zpxld3oMOT+c4KQ6eNDasUCOU3Y7OaLcWo6vmrEvw1ju
Ht7rsYXJ4uknMhMLHObeogvPLP8xcv+uU9X6UYBm/vq1Chl2t44p3/sTitXeZHDKPi06dh8AnhEg
fP1MdeYj7rYtBIjTVrFb1TCYTG0ntOpcRZ57p3yJsaxo4EqpWEYLw5kqgn4Ak7yEtOjxERGV4iGL
n3eCPC416bRZihRjIBnhzfMttOYOgKQweEN7crw785Q7bLzfXaolkcOGXQVt3wB05KkcqNfWDGI8
4Yh7JgkVtplBe8f0/WRR/AS3wGDINdmb35F7zRy1PurfVistVOD3E8QjUuVjX+df4khM5aI6/wXb
u0BoM9TnCbzt5Zb9ZUnQKB7lj77bsETy++Gwq1HTZbvMGNafZDvBjVAyg4G/1WZrwMmBxiI/M4+s
6OIpxKTPsqpvhScJsHcurT7kpjJP7bm/BMV3knK340FDOjcqQUv1on+vd5UekWKmJBCHuldlJ8rg
uQ3sFQdWv4OyCp6hfYTE1QIWJaS35vlzHpo7Djqb/0GDECoyvTJoaFeyDqkdtcHWQgYhiUfTbUGC
NCySCbW13rXKnWI/w0mvJG314DBN761Abw5QM0BRgmQcv4yhQRFRu3Bnu7zO5vBpT5hihnbPVq0m
cGPmRsK1c+wQrMCw3tiAgU0JirWbi6H554nL/D8V81mIjhVBAXMyg6KbrffKrjCzoImRJa8KXjCa
yKKI2F/Ncw5KKPWvZ7vWwbKL0DWEbcPKs6W9DvzXcPmKxvy+VawvwDptE2AxfMR8Dqs/hbnzq4OV
5CywLaP07ZVd49nrztC7xOInR5o6GAT6N/t3KrZlhd9Z5WnSJejtbe31aXVwffEmvTIzYJUN+t6i
esLa79/RaLXfXa5ygFz9+FunQs9hMSDsj6QVZSiQpf4nlI+lYntiGTBALd/F7LXh8uda4hEEjgb2
4T7QdJPRMk7K4n9ARjOjDiySqQzzIVNAFkWJnrrhX2+CQgwB5UeELk5tGbGIDCMksOQQtclBlq/B
AR9U4rBQd0/AOTKTpIjbQKIw4mUblfj6nW3d0XpPpVOoFXcB7LSv82WCPSqkFHR+xo6m7b2mVQD+
3eheGDClCYbDUuKquNaN/c71Vs73qn74WvBqrmeLdxpolYvakVODui1f60gKOCS6JSJazBeMeQPs
KWwqePWbMbSBBODNDo96cdtMl6YsiGXUl/WuJKezB0zER3H442g9tOL2fb3Qfd1eq/u95MTcpcR7
2sHF+9/kW66d3IpuBQkTCoGo3isoo8dmK8rv2bI9KCv1r0KWRo2w4DPM8u9cQm/BIlj/4yWM2qwE
PiJ5A4YJly/w5l4MlhpmoH52148OsJSjWgJ+98lgG+ILECKM4FmbgX4CaLQ6ZbspUsuUTHeU/G2s
WrXD7G/3GkTeP6qoRDvpsaxd941YIMiAbFnCeeOGJk3u0/kOGNDQUYg9/0LJT/nzsvhTJ4vojlkW
fq9SKQVbeIZGvgDFoBeSZV7YrvpzmuQbkEAtTiv97C8LZcdl2GIqTv9HH8yhgjDG/n/o+OwMX9J9
/x6nCfnbx7AZ7OTbidWuXLFu2N/yyxKHJfA+TIfVjjU8CSVE5yBJgNmpbeF+AvRk5eULuGSt7sZI
CAowqDQvEhDabILuohOCdNW3bWouKnm40zI2PYRbA2Uf0NOkHtz7yHY1cDLhlGDbCbAQuezuVrDI
O3/A6tR67JCfktvegODU6oRasj0a+KxujvSHcxJaBCezCJKRd1rDszCL7y+49iLHP+d+hJ1D00a5
MJMsKSfpE9FklWRYPLTxT8XtGDWttyr42sfm++vU8T2WtU+Lf053Q/TVPl6vGgk5Gbz+u61Ewvy1
rLXT5l1PSADDmo+zb9ABLj8i1N5BEl/Sgl/T59IF8sgqiar5ni5KUUiZQNPjhvFlVaGzxs6UQdch
PPYceqmSlaNp0W6VzhIJSTfwHFMG3iJCDsuJXZl0VUV+Tj7hNXyHWn8heaJzix0kBJVzes8Fp+CO
E4Cs4d/2Xh17v4xK7+MuVO9lU4ykZOTbFS95jKaauRPs8jYGSjJS4temqEdmn+uOXHdtzuVFOVmg
Xp1ZzDSEUtbEAlsPF8dQddXwy84BdcoBBqSjE2VGWdS+NIHqu5vgMhHxdUod5DU8TdqyxZVy9SIf
kkwpO0grPy9DIA93lH98304riDtG9lXgl0+DAb6Bc9oIRXdfO3+wUZTkaN1evOVgrW2Io1CgK7b2
E6NtKJXip1ZOMqlbAnjagKvcjpOMrg3DjduMcSHhEtKqAqiwXQdy+amuthpQ8vYF3PpISe3RI+Z0
Du/TFTryau5nUyPVyBKZbioJNFOdvL+gU9by8qVaPZEwgTPq/oim+dm/+jlAfAhbphgt8kfZzZCr
TX1Ep8OAP+Qig9+8mwr6mXiLUQJ8/LDYS4MSHPelxxvvqqLUPq6z/BY/AuD9zZnHnOC/T54FeOz0
VVcLq6RgUeP550stteqfgS9qvT926qpVJcOUvUdyn9iuvUL5NOypq01dwOVqo225jlrkeUUDI5u5
9kQJAin1q3aIyYhmD/7z1zTjQhRbLvcb+QBqj5Sa8cWyXWq3HdO1G+3llbFkOPWDrsmcyzGlz0C1
JlkwveIONtnlInG6mMODrWeCvz791z2qMDgepqDy9mtNCQfLTckM+4qbkJuxrS7zWxI3Xjvms3xJ
C3tvVy7xPDnWTFFhL85zTOVmSjUEdWL69312+9cFkbmzmywZzHdw00jw6SNqrLrw2nhrvF31Lje2
e0FNCOQiFTBrDzgc9aeIniHg77eaz5tBKcWRqMdyoe2Z/zCfAscTKnb6wF+4K5qdgV9Go1CWvpPA
6frUZgzin/Mq5R7+gBl/iCVjLoSW7Or/KVoReAVgKtZjwI0mlnyQayzyf8Oxi+5iTDU5Cmu7U2Dm
Pv3LmBhIFM3BxgL5ahICsdCt2M4F1ro2Z7L6uv7C1ECf9wCwtyxG6la075cR9N5dj9qK4ZM9RE3K
9bSsQ8z2KLx4npEolUXbkN1nFBH14ENtPPdSf+0h95hMlB0+DNt3ptnjBrqJtof4MNinYNmLXe09
tlVBYpTG3jKUt4cggFH0EF7US4/AFJk3D2syCthIMXphsfyJ5rJCElucE7KuCWjXw73BH65wRXlO
ltVNJpqHDra+3sb+bjdTsADDuDqulSOR/0AxcErzk2vCOhrfp/CA8DihfigzL/DhSCNyjlxM2VZj
u8Y36l78HhPY8NSXwh8GQEWWPEwCGZ7+psWBRCUjgyYD/dhe/Nws/PdhIWxPEmdJES3q4fxGPU6A
shZ/KglCJGeFvhlw2v83AMW0U8Xcqe9jdvFyCKxfhWKyeDbz6aVUvC5Hxa5SHPzV6TQKdcnRZake
r6k6JILoUcNso3Ti5nmZXVO3+f9UHTSpZONlR1slBJr8iuLEdBrmncX+lw9NwcTby9GY+IBy5yAC
VRqlXEb5DjjkDNO9CAxdJ6d3QboEqbVlXZ4p7+/na+/mogTEzBikhA4UpJW+sUygLlonRRhfZFyy
ixkAB4CpNroR4BBBlVed+A+YWjnT7vc4gUzbukKpky8CXZ2IFDRWyC7eZPc7MTBg47VsZ9CT9/ny
M0ZasuRAf2Csw81dhqccNsCnLdWkihxaYNpaX03xoIMxTaxJZZev4QxF3qwn9vLcmBKkEZpxVqas
QnDkYnYkZFCTvENWycP+4dB8S/CtLfgS1URICpRHQKm17dYvPdO2GsC8YS1V4H+wz0BIVs51YvSx
i5BZQOri9D9dSMUC1pbXoFi1syr2NSlcOZldc5CwJuITBonOSwL9sNzKJ7rFYX/L5LYvNawz+x0m
akJdR7L5QbL96oXGqIYJXFhLL1fMcflTUABQakBFTZr9E1uX2BloqLyC2hyRn1oBfDVQuc5Ipehh
IGkx4HcB0yEDBTKBSTHwQVX3zRFyJTfeFDH0thG3hdo12qHsizVJsru/07cAQolysEUZ72rJO08L
iqxyP07p4lbsOx3z0fp+CIPTeSasNVRroNllidJfOowmL3bI0M0hfjegSoPJYkLcqnSYyKVSZoNU
8VP5KO0Q4e2DkaX/CcwhXrP/sJiHIOErF7KvbrW7/vMR5WVg4f5DhyxqKvEdR0Ic1ITSDwwIG+Mm
q/UbSSynHl8GIXbrZUg9mUOerGN1caGy2WY7qdJu4y0m/Sv4jZY4NFCDTfDc2jiHDZKtOS8Tpsf5
gb1U54YNLYFv8tmOIZovCrW2fIJnwRfosUl1LLHx/+UCTvT0zbsQAvig+GPhWkQ6YpCfr81aukiX
tZzHI5e/AWeTzZsBwWkUTqWCraLQXePrpkS5Q3SVqFkSKrXKoQHfZbHTnxtNawnIl/zuaUgTWb1w
X1E+xJJH08Hqm1lWp2wNTH7DMPnoAKGi5aBr7gsF7x0rjv0WdYI2OCnJ6hZlXmeqG6QuSU0xIjmb
NPHK1bHGTj3MTA05dr+bo7nISGCFPEEo5em91e79x+QFu8e2Yujqq+bPhlx1XMn8GP1T6N+ctMJq
mpJoLqPPjZGs8+zqy2KR4jG0toQEReYmQjIW3q2eOXv3HnxRkJ4u2/rroAO/tsu+8CQdrqDiQYsC
PKZuV3PrsHl6djjC/ps5NpkEy3bq1ZZi1E2iknQgXWgGLxltBHxdXuwZVkIfJQsguKZ0kQJIoecL
niNBCbpmVlBktknmNOGQIn292JMWQ80yI3+OEftF7wkzacSqx69rlBFFqaosybIOEG/xuUMeyX9k
Xbu1sxXapvrLoo8/8woh7WmpiWZToWE+ZxZrexISn4YEvDva3ptlYyT/5yRyVSVcvUV9kQ/9ERAg
0OZlr2HByu1y9NqjsFUISGgbGfduapFBjXmx0tSZiplXdw1Hc6SyEWWdQFHNLOBesLMubYsiGHU8
ii/u1rNQlHln/X+TucmU5AZhZBnNVu62w3rPIQuzAGg39aFMt/f8h4y2Ctg6smwlVI5coVETfDAq
SV9T9q7+rN64uJ2/WCfjaHUIpwJEqOJ7fz0FC4G3aYrx80tuLozGASVpjCmodhT0OwSQdYi7BFf8
sRtS9xuA8NGiedAUvg/x/on744xgg7ZEYWK2uuW5Vm2QjjccbZAgSBjGJE88EBMa/ro6pEfwarWm
C8G7EUxxyw+92JYoT7XQ2bcqRyE83N1OmOKDcAFppN0RMHFFNNKZ5MZACSj/CZ4aI8/rgnYuHYJl
nr+MqPSIxnjoIIwNm1/yaR2BK56KPWmAfkjAvQ/V53Syrk4xZGx+2zb3QT7RvNgbGPzeSNTw4HCl
ZLey0zAZlBiUMU+OyZDkrRI0SSeQIWesbo6A9WoBBWLDUmyTCBgTz7iaAczbO4FAmKa1LYBHiNcM
jl/dFr/6R0LNUIWlvMaHFsy5y7iHkk9QUUs93q1fB7xzsbKJOursX4YS3SnkwXVEQZLkoiiDpkSt
vTcvuWTbOb84+7RpsEbbLB7sJSkncHu4t0mrTr3L3P1+vsQ37ydXfhBOfZiutxka3xSlebpBz3l7
odcAbuiG3sukKK6dRdSfg/X/o/IXA0Awp6JLbCeasJUx8tjDQgJuOaAmsqZKu2+1MR3ijy0cbtSU
5viFpvJvXi/lw72PuJIfIqJU6E+OKxIvEZNmwDaysb4B9ZhdoMDrCKVnrHWp/tkoOacPz4IH6tRU
2DJ63XIfQszdI8bmOkZfponwJgQ+63upUiCUKnbLORfhD4j3eKXw0ABAK/gIvj7CZJ3zlJ9ysQkP
ewOotNtQidFFfq9U2WOJBmBrt3t6HvnoDlsnVqJK9xMRIFH39XQs/ChHuvBl2LhYcgwvGept9ddN
PGMEcb5iMU4TTlgUuCqeuoGXuy1lBvQ9T7AcnLYPRJvLjvXk/b0QRjr55/JxqeqgUpJZpiI+kLOg
alrXVslWeBccM9q2GrrmHQ4hEjpIkoNzYtvwC353zGpPyXB1sCJW3RREHDlXHSUeAnf0MKkfCMN6
t6WVTuSVw6oS9puCWIoKx5Bekmt7YuAeuP+S65cojW4mZvS3KrlVfslohMfM4QG6dX075AeALw31
fwhSSnCfteAtZCHelkmBci9jVTloRKj4M5Cr1+YK9lv+u35/wOndb0smns/g617QEdOStFKQ+cbt
wHOwe36oxEmDNMvoRa7RKtGAwzIhm0LiAHSpiBirvXASCezPdBU5i7XL8O8eK/HqhBF3sq15CIB+
xMgfUebxIC0277P9TWAoDqwCYjMucpzsCzIWIEoSnH9h+ONbM6B0DbhqvYieu1ypgCfnd6ZlW6r7
WoH8kp8dVLB6gCSYvTlyScUREftFa0BClLYtX/Q0tvkwQ/m/kja6upV8DU3wy0ijs6NGypkHDvRm
ts2d+YudZchJs1Ot2BHietos8GFye7VuyplgIkxaUY9YTav7VTw3JdeUENN0PPTBaU+WaC89DBN9
bnqsdi7ad/Nxu9Q1LRHYP1V16lriWRXQNXq2sYOKMQ/boxMO/qgv94RRUsjTRuFrM5DBa5qUF4L3
8TidSQtFG8C9CzgpV79cOBXmFjsU+WD0aLL8FcU5QS2Aa6BuhbfGdiAoa7e7m8YTQgHnlHXqoWHv
hT75AOhVFg+5HKS2odzk/dpzXwpKC7iO/5vIQ4PW8/ZeN5l778QZZxDIxAuAYECqsofFdnBE/JeF
bNitrzYaaPB67AzEY5srG2vezpY4sUOW4qB7cIaanuMaZCQCpdiY47LsD3qghSqJ8SKcu+f+L/Mo
IKsdR3HxmpHI6hWP3NFESVCJJVbaCKLComNtPTyHlwhHOTDmSqA8RB8uctYAF7bEbYBedDWHndJ+
WFujZITEglRb7RETwSmDxZt8a5x0/QjqsyRgyHdnkqLUv+Bg1nJi2mMaiAGlaCC9ya/YdX+X07fh
zgaSsyOHWjqHBvhRURObM6dGKubsIzjyOwzwVVzDt6NrNQfY4TD0OXHV1DMkBsj7UOTmdgJouZvz
nkLqWSZ5KpYUR6PkDNg9KmQj+4bgnWzlLkVwEiX4L+PTSf89reUYXK0qo9w6DqcHRDh4cVSWfyqa
yVBFImTQnpa0To+XN6yIg/S3R/ssvcXsWDlyyV8YQ6Rv6Rjf4pZUsk0uAQbQet78YugcH1zdjuKM
UgNLiQI1igFzQ6ERmwiswV941rllxsCx249ikJBfo96ZWjZeFP+WjpTbLNqELf1NSeoOoPsu+mWb
tZwSknq037JqIkwvHM4mMDGyv68x3ZoBjN6gpUvpr5GvnKyzmYZuUHGa3S3ov2wFDxCqzJxTLXSU
avhRIQVj62R5zhAT+RIvmqOTz06asaMku1GYrNCRQ7KDO0a3OS0W8ChXTP9eB4KCetcki2Xz7zrF
YfyeW1hZLJdi1ff9IP3CVxxGbMnqkNLHuZG+pPq1C91WX5ggBlXsDYLYOnKoS54w3vbpDKYyTcyP
ipQznCWCpzOJ62fxObcVWo/2jAEj3XN9FR2b0d2SbYgDKbFI8XxUd99AjK33ub8M80H2hMwdXiBX
e5gaUCBJZgOjgRzPNi0mlslk/fDp2M+zpxRiUvJCyQ4NQnV0ex7LJV/off9B0TjMYNURfA4I9hes
R7Wtcsb4XBmDTLiURKLPfKOAIVDl4FrK8eVLsv9ibvmPL15IGis5d7VlvK0zebVWiqmHSeVrP0Go
FQb1vX1AfSb6Cka5vD3cy17tzMUpff0gBbkuQMaA8n6MrDZf/Z+7fVK7j8cMXGfxx7NBtj16WsuZ
lTQUKNEDu+jB/IPUhCPdFC5+8C6EgqzvX/YKAlFGOFdw6OjJJ4SXosbiJQlcIJojZZyGeHWQT1lQ
Gzb62pg+a4ahJEvjbUIZ5FfSJtm7zf5svxeduLm0Gh4eCkK0ixRhfLiHcWP1kjNrn72SeOpZFwx3
6KxZOqVMj3lgcXBYrwZCXhr4yunfUrgv/zxelzxVaN3/6Ol+Ws1zdoZgFDiSFXVE5H6CDBxUZs2m
hpu08ogCuBwYiouvqoJSrP4S98V5SNAdCuzORfg8lwEgXSmASr1dZVplABhX+KV72OADuQO1oiti
qAbBvmvzntwqUNZOM/DZnD/VgNIQrx95+tsizpHdCbxifsIPELmyCp/h19htVxFUzUCbL4AB79Xm
sUcPCqPvLU/ezyOzcld5a5Yds8w0G9cWDs5PzUeZ1veRC++Tiidozz4SaP9OGAr8OCUSBTOnUJ+f
F/9xVMex0t6rbzm6tRXpzC5nmXv4KxrGlEO9Nt4/x71pJ2O4ShSfMsgZpOWJQZ3m2eKI2GXuzEHW
1NJHfK/1qlTENMAjNESqWDVwklFs+rsvMPCWXfGNFX267iouASEip6aNdG+Wf6bq0b90DtlyQzBg
ZfcwB1F6/HyWjccw5A/Xc5uBG+VisJtU9ICtTF0sj0hWxqFzX4Wezc3FH5BAdXPP3sIJead2VweN
HRyatToUAUy6cZsPxd3jZ7Rwpcv4PO1fX5bSiuZpnTbw3VRfZIGvz7K7h0JhN0whTxgHgxRs76q8
AYZgRzgTjzOd2KFqDo2VESSdlMpKVuvye9g0Ld2ih5MYQ7yqB/ENIdb7xcD7RyWUfRSGBohzjE3h
58YxGOYlHWPn94JZGB0vcZl9qeS+aYDnofx975ZT4XtV1sJRj6QuzceXEONcPXObZlyInxW7LIeQ
EEBuop0d2yxXwKqcA++mY8IBI/xAbVaARkX7usWRa6/wGYWKye/YzCbgDTQiGg2/Xm39RkeUCy5Q
NOlRd97b7dtkWVPF1is6Cmp1vNRzinGK/1xfJJceZeET6TbY7BSKRoHE+koT1kZTf6KmZ334Lrqo
JKkfmupZE68FLTznHRBRbXM9ToQ5M8VGTIMz8+UXrMXIw6Isnp937+h2kIfG0bfgpmgWPbUeMSwJ
TOZGQNz2K39F5A4geXXRrklUHw03psVtnFaOr2LTAIa2MCUQa07vxItoADvGPhbMp48xx0Dn9v/o
WMv5ys7IXkSqugMDT0uzHgzcP1cQjELpqKP3EVAAbcX+SH/aeXezAPEuK9hirTIig0pg4/bu3jKR
1gkLoVLY8WMIESoYkCYXNC+JZy2okzfbkmuZMbFzbsoJ+vIa+vfP1qWO4KJkoXjamqkfFTvlvOeb
6bkJDXCj1qEkf/Mk1ua9Qzo5DZaCOyyC00n4c8mSFX7xLbFyuOjQI1E4GvvKQ5Bn9MRowcPOfeja
s1IueK5OQa7D2yMRipnlXUY5MMngXQayrCyFrs6ahgvhOwB/I0gJk0knoLicMN7wRetp1a/rN+Ku
2FouY/uI0CXiN3l6BaCnVH9US5im9YCLnTV7qTrcGeZfv27GItD3n4kkthilBhYerZqwBcWdvlc4
KkQyhpgoE1+NE6bVcMJ3YH7T3r4lpH4/Lm7uCpLCH7VqgxlJx2PsaGQJkYcIlB8W1LEFEyHZ4UVK
JaGNjYwwbIeRsUSrIOr6tok0W4BZLGeG9DDeLSPoj6rRDbPcNE3J9nYZoZjjzKIjDLG6TxhDUhMj
KEoITeYQEgWQCkXIUpb6aXQ/Z0WX4oa1+daismp2TXE8aT7HKttyKFUNVnNEqyzKhb38vrNq1Fkd
TtDAXFjf3mUIU0nz7+hZxitQWM22LFuhkKkfIJ1QAUj3z1SzJ3kzKg1Wm69p2yE7pxICq9Sk6fUr
fzEk8dy1UINKpFQHsD7ENLkv0yCAxPAv9HYWipbJDSWF0Ql8Q45ZvjEUblEbqqpOQE8+6S+NxriI
ZbOFqqy/tOOYjkCE8e1edyG8FkvRjoOU9o1b7FaPb4bBKfbLHjCEtflI6yVMR3VPmsbQ/kN2XSNi
nEMJMMT4F6Wq5T9wJUb460ERjFIVZkW2AdjnjjxOP3NsaMuoA8xAkzVlafjTPDNaR6nNhvfObcoA
+8vyR11Hw/YOP/ginKRo9LT0ITJIQUwSPi9n0go4QQ0q074hb1slPj5WsUUk9yzrYGAtxDHVLUlY
3gNsN0cWwLLfm/KY37P/3+kc9TH7ev7+rZ9elsBE353WFRIhOtUiXA65CkdpnPza1Rebl5DSRL+c
GIlBR38PbpgxyN4Ft6ajOQPhA8ZQj9+v8Iqv20tjzryJXkSvcCE9Nl4QT1zhWy+EXPIM0H5IrIO+
w0M1ClkThU9QWPICCvkMjTk7i+QyvMnrjb/uqWSGi14cOpUsm22IGn+FwdQsSwwQS76TWrZ0SG9B
+fQUjaxwczf7lMW1oLUOIqFbIFWT7I72iEFw7hVZwcNLpaJr7nUOU0wpebtQbrvtcxPGC+GQ95DJ
oSIBitUwR+MNMRcnnFCwcYAL6j72cgJsYBvdDMxW8jd3QyDVr5Z5A3C26LCXlOY50jZaFEugWu6d
39e3B5SQ+r+2o/at0KH1Hc55SrsVOfJH3xtW8E4610EypEDTRbaVw+xUPas4NZJeEUyBz0LvokC0
OVdh9gpm8n6utp4iRou2zzPQ3Fy3OsL004LYi0yclqYTBwt0bRAHnYgd/kI2D4A7ricl7SJW9MXA
UdE0WKOH+D44uIza340dLWJcEF4gz7aLxjsUzxg2bniFukPRHPNb/4RnHq/PNetk50iNXjSkgq5x
i4sCZ1RswNNzaQ6ZY5L5/W7isSwrHjJcb7kf4SDE+qNB1MfKvdS7MsnqL1Z0yIfC/+OpX8/wRz4r
J/wOX2Cnskfv2DWtbVg8/u53jECtM5owjy29uVl1PMExON+6k23Cw1cGu3HwDgo2gDjP2sw7Bo4X
EWR5yz9kJPh9S5DsKY99liplC5uhGjwFTiK4JgnFFeZ3I79uvjPS3d0MSOOG2jvEvRAk4qpBOakJ
3/J8+CiqioUTTmc9qXDC1J3cB9ITY6P79CIqwVXkJb9Qyb2tA6GGDsGGQj/Vf5OFZqZ/nf22d1Wr
BBKJ3Nnnim6I6XQplRlblMK2xz4LIlbhDo/ZJKoq1pSZFYDh76zjkvoylPZIOUVtWO25EhH/uvPP
+oMObIoDcH+GwQvcamCC4mNk6RhfW2D/jj8VEXXnUadssGUC+tY7eqD8aNcyWKt+b0wKYfMf8PqD
1la10GGPiJMI5IeV4RY/o+z1YQfRGaoOdO9b1Hxgg2+/amk1Kp+QjfVrp+BnrCZdXbEiJlKvJzkD
51kP9bVYd3hfqomqIUiqbcTcMxxtagPr+uIhnXBVE2Ro5AubTkuj8cMaDKxhVPkmM51ENA0BJqlN
+mrE3uuZOqj7kQES6woptuhUZCLr0NqjrJbkkKH/Brvq6KLsMbwFWS66zrfiipMNt0khh69s4R4a
M/0Scb5ySaSQ8rCpIGtWVtgcVFRj4IMMbsuS+O3XxGQvtWEmuotHX5q/QlUllP0vKl9/m3EzhvbX
K5WwzwJgQ+MSCBPE+qkBSggZyz7mC4vOrDdMi3fspIIEpUDT0Xwg2LCk2t4YMYpP5HIdbXcd6JY1
SHFqV0JIlftPTNLJ4HDzDyNetxbKJ644oSbivAsCc5GIGMj2RMu+3hRD7MwNmtLvenTU//oOkHcH
u/esc0vRVJ1AGl5WCfFUqJ7+a3ehfkpsNotZSGX8+TUCkHbzNEZ7hsYHPXSqUbdJvJ+luCf3KMRW
JCpKltv1sSpHc1asWqHZWJQxxT2OwMNB1fhf3ZReUJZNY08/TjCXCxW/DeroxgX/zTI/2CRzpxlE
YXkStCOyUgxjhykQtaEN/O6t1PLPZ/QAFbZMzcgxtIVZlyRzQkjNQ5rfjGNditvMczX4vc3XzXD4
lr71pljznlbMsKNulI9nRU8io9EzTIk3/su82yZRk8F8R8T4k8DFRbiL3nyttjX0ALYjN2+SwI40
K8zsw+bfKU822wAy/XC+UcE3asVshIljTXbk3uZNRAlTdxzQWCj9Sk91dpzntqtzFI31YzSNCYVx
gRMDPAncW7IwcuEvtX+Rgy0eJvj+7GGcWFpwtJfD6A4AEOud5dIDaJUOh8TSTlD6dM6zvwhsEYFH
SXH/qty9gO8gf0AUqpwn1vLG/oRcGjhPGSTfrinjEH5a2Bs3HgayFm1kS85dwITaN5EX313SAmsX
8Kt5eE1p3zn2+LbLq7yyNdmIk8Fmm75LxBVUrE/rN9wuls9mQSwQsIFmIsYcOL5Lmard25VUI4vJ
y4NeRuZEB0BRLpXxUgBPzQdaLq7TGYV0zyfk/p6XuwIHSSKfsVTjDmHDQrzDh4ZQszfO4hx0vY+5
2cSPWTB/w+HUsb34F82SjIBwR+p3s9Soc/KxaZG0HOoc63AaKSur+J9tDaOmPhK9cOnvMmh9LLKX
b2uM3MvLPHB56qxU+h7bt04D2mQ8ZpfllQlODvReAKL2Ai301G9arIRM68OT64WSKBZSwOM6u+cK
vCYveaOZhVUgIhPPPJ/orI4fFN7HYMb1zskZMxXiG+/sCWIfMti8Qv72uhzcwM3ktKnPwSE76OKC
9M3ywwQdAvb0O4RkE1Enz1+wqpdYBvRi8dKXKPihe3aex4qA8xFROn6F3lbwCOvfOMQwdQmyhvWl
LY3Qa3RhG5iBqw9TNGxC9v3mKZF84ufSTBP/ERDUIxO0PTab6IuDBF4tfyMMLvuN5nHWeVBbBGIZ
vjcT9+BjUfQNknSKJs/ITmAYCV60RPGVvk7wL4EiGLHjkX1mg3pG8lmEGOWH3msfe3TUkSWewPuH
RECDzgihLO3MmktajrM8WSIO64unOJWlccDVss6dJlR+4ynfK5SFoo6JQVLk5se0yN+mbiVZWymn
Jb3uZiaPvzme6wUz0tSH61wrif8haRNyN1SnguykXiG2uIpUjRWj1W3mpD7TOg9pghCgnSs7VUV2
gKPhSghjeZSw6GDUwQXeR8WsfQuqmtAm4I9MVg7TE3Pspl03BjkVDHeTDPJ1a6xfIBRO22piKfpo
rBYzcn64HmaNtsAPeN6CosJ777jU9Vwqb0HE/jxCozYFRqtpTy/coHtiFcwE1NGWuUc/PYMWU9Ck
/Z7B7/dxDtNptCHnt94syHlPlPA9bUN1lXp6wFV7apy2Sutm7BVjvMvqUusY9o0Cr0nWLl/xWn94
+E0KOnqrTdw42DR4Tqm9KNsd7UTuQ9550CP/63tKUL1FvK9Kc+sh/OV0EHgxBTfvJ8Yo+FjOw7Bt
3ijV68uC49wSSmmJhBK4G2C03d8HGcPLCNVh/TxhIXwrmnV6KKFd0aeLZcEK+B6V6mDS5rdgPl26
5emzMfQRttz5OGFdIOIMQaLZbmHLeE3jbkOfj1+d32TSU8oLD9+B3/WK8Cck6z1d2TttDkP+8rk0
Y/+NRgv6Yo7/h+BN9WyK8Oecmeg8bgk9xsnjQP/NOhxFX1vY9Ppk7MuOEcU8rs3QWK6O3V84vu46
BfN5TafYH/6qDR1sTj0dWz7ahmxW86e5NuQLCN0ZMM5U4YWTd9b0UWVNu3hkJU3iyvCc7O1WNCYv
ntjDLoIH1GWm4CiJTPw5CgKjse2JAHY0FORRGPXG+yzcY5ibmxbgfjZkPxZ5MmJAhtnjHAZugKeG
eCnlvVl6EhnmXG7iXfVcFqpMrqbM/fdQLSX+jLnNKZ5maw7+W4+l6zK528ntDELvX+4qw/ekAOkq
deCgWv3a/lVnAssjV9RgyVV+KQ5moirYG4viL8M9JeaPSZqih8LQF7Bjh+mLoqtro+9442O2sNVa
8gkVz/MvdUyswOPL5uUh6zBBAmVHhzEt9vlWjFFdgFMW4f4hxHcGwvp93TFgx65apo9xbetYzyXm
pq5KKkMT4ZPEDBSRyP+bjOWdkhvcYLZGMQD7FMdROfyxcnF4MElQlDdjW3PZl3tY6sbBEj4/CURC
6lXm9GBjAMM6VToUfraH/NabTC9atJBYkkZVjZoKH6q8YDtQ/ux3VxQwzHNvhini7N5A1k+0s5tu
BVl9as7byjp6h9Nn22KBLGLB2z1qitgh5XNh8Sx9vd5J7riQ9y64Nyol1+gKHY5bjcNrYlzPkgAT
j68uVvR2WjnKCjkZZVb+KifjBD333gMlCogPtE9cvyExqZiXArCLkIF/iwPf9OEacf6XNQ1Y3M/X
/O+UkaMoa8x8F5obWWiX+4be7UHnEdWMdx2CVrKGa84EHnuONDr7XJCcbhHkncMC4BSiK9FISPYD
1lawQ+cKzixcX8W7NQwlAgE6B3SCdOhyotzrcFAgwZxqeT/qykF73YWEDx3rN2UlMnonu44OK28S
ZXnqPBcnjblFsaD2J9w4gr7tAfYT4gsFqj167UAmafiBqnMjWIremUQaPBTg3wRbRS9j+H093I0v
YDsanOoRPY7mg+aZTF2orfU37eHzrNe0S8peRlKmGINiwAFsJFdfZ07vMbpogbzD/DgAx/p5FuRv
J1r80baaWtj3XAt+kNlebG+ftr2IFiR/8ettdMih7sNv4mBGeat563jAHDEOJ7PqtglFFaLuQ894
A1ibwXaR2Yw84/OB+JZKemXj4LZquCIE9EyUBudH2POWreH8yDcuC/WubW8C1wM7Iy7cZcFhF4A6
l4gxLawvWUc4fWisjdOFrhj9q2Vbd9J9inYeJ1n1lWbzDdUNrYbX9nbD2GwE3Qx3yxQmVwtNVMw4
DG0wkKLQjSJLCZI7414ixjPh1leNaSzpI8vvudrEVcyZwgNZj8ThQBTpMkXN4nXgqhCVNmFgIwKG
W+gJVB9HmWluwc1tiQmoDEoyyObqs13fQGdzQCOpRS3D+b2c7acPGUV/ZaLxMjCEmMzsb/iZAZy/
nayKYIkXr+xoeFmVkJ4yPCZc6FTY0Tfwp6Q1PVHz8SHgRDLJ6gXO684oJtQam+Q4Zo/CIpNXcT2c
2Tb8/P1XJYKSGaRJDfI80MBAaP2s7vaFMB/qWjJEUEjj7LJj1k7X1lKGbR1FWRYE/xPpoXPgr4W7
w7WAeYmHPn/NMAxEd+2caKojAyt57JofFRaCoVLxGuu613j4ioeqO0/PIYTj2j53mKzG5moIpn43
Gfr33YlXOdg03e3toVe16lHIAxeiPU1P8DvaCkQ6u8+vGAdnJy7Vm5O5oG6rSpTr7dhADvluNz0m
ufCqYbanaWUjPDOctlduvszvpzvDrvgsU8bd3zF4BKOeP3MAgVMhlSG++BmXu7jTDgphxYBl8d/D
M1M34FMsH3fPJf6/uK1p8/ifKtb/remphEPyXLPh76PIeQMqjt5V0P/6CZS5eVv47NDbbRuHcsWJ
kQCdcppvHfZ/56RMa6RfAzBwQpQG8b70jiegzfXVW+uIiUzVia+zw65vFtiEeazXtSg4pZZFd1x9
ZCmbTjVr+uy1X5UAWByJpX8mMZIn7Q6cbyAI2yaznRAkyyYxqLB/mvbkyLloFvdgUciXkubSS+U4
Mu7QyWFaHF/YdKhy0Yl4IhvBZv2GcBhOFSia2cNzO/knffHDbvrfwSgMSvsmGQVrZ98/7f25LTfg
vNNvvzzqR3xjegHEefSr6mnT713e729wcRqAcnefd7qYnU24j+8HcFtFRzYtS9HdpTSzkVp+qPBr
T5GGWw290sFMZIuWeZUf4tfIJAJ0lHW0fCs9/bQXYYM6f8xpGpNDB/Y+63y+HfhJUd6YnyRZsJZA
Kuset4FN+jlRRDESrNxrUYS9/07jH62ICwnVy1noiiFB5N97DqSMmCO9mew1nxqZfYDzvE+QXbrm
zxlIrV50GWYPIV15DDvK7XWiia9D0zjcvUbrSkwIcQmyO2z0U9w4viOViX3MPhJ/VFrXHzcxeii/
b2bkpw4ldSUnUqcy13Rp5IyTcqzTylAWOIEFDzy9xYUJGkqWutleAPviRIZdCbaheVhbblOPCQYb
W2NMsge6/LZJMraIMam/d6vMxP4QXAg85Kz4ZItsY6eE7/hmI2CGZ2Hc1ztkYY2AL2TCQK8DlSla
mZOidz0FeXXhVYN/DTha/9D+z8kG+5xYu3/MadOJUso3+wS4IvlkmnqKnBU/USEpThDTI03rZm1A
QMXv4htLu85CrhIrgb5ta5Da0lck/zkKSZkMJUVIOTLqAXKs0Q0fJ9nCQ0S5FacOvIu960SfraVC
zZMjU819NpqUuIXggKg2e0azuiQGIswjX225uWTXzUpJvIy/YCc3G0A0jbdyxp/BAOZnKMgKhw53
95HwQN2soyMGz2ldCepJnGCqgMAlmz9yorJfOBUPQV7wEwf2OeRjEMkniKuiPHJ1LlW8LI8m5hA8
tnia8fdaw6rR3sPBpQhylJgdy497Hk6YVcRlirVFZiGpKyb4QyVte4q72AfR6TeQYfyJJqBblcoa
ZRikDx1PwqbfRJBY5PCftlC0wxQuMpJH/Rmrnzd6d3hd93Ci8lZcq9fJqY9hXVX7L+qC5p9crtBa
eVvv/GMT/iCm39A6ZzuozbgUvuiJrkBIYcPR1UCe4ye8giKNrxC2UqMM8TvMET0DodbbSxhz9CUG
vMSRWLguAyr3U0qQNZDsqHoHg+bhdtZUZBfru1xGG8dnE+x6U5jowW1JkHksO2o91y42mPQSWvo/
29lR3rR71E4Xu1qoKlUvdSFYFo1aibKa+PndvUR7G/ZppYYqVg135kQAmGB5kJQcX6ndU34xokZb
uE1uFTByRtXFVyw2huWaPs4m5bHkpdztUHuv0iNMy5urAnb7VupEKgLV/EwtDNFn4felpIui7AAh
th/sCbnjnvcGuaqnHIpI38QQgTjyHlQulOV7+P1Gd+Y9wQLfkNj9QCbkiwEh8oUCijAz8uzZ0r43
QPzhtg1fNmJDjl3dw44ZGg4YkdbWhcACW3UgcRyoXGeUgwIG+4uelGRHklwV3tDGXlHeANlM8KHW
eSxN2hT5lvdc8BJy4AOcQcOHVQnCn6R58eCjgpxqk9L8IK2zI7fyQKHE8R20SAbg9XK2q+qtgU6B
ttX+uydASg9qI0F1RcYV7+ulCguddts6MwInYg6w+Kq8x/SAhsAhoqAnKZ4Yt1Pu/8wancQIaB9Q
e6LTAj/D2RCMNSovTaKdzK82wePzYpUBQE4x41Lp3tYIomZRyGwlhxhX6kffQrK1aSe62kSr2bI3
y1EN582b06molyXPe6sMgrzDHksTkDD6x4yhomvJwIV/8RWJwSeqm43bJArgtcpzKdA8xMHqaKWn
uhWJbsqo77HzAt5Vnw7QfesS2f2b/b2HUQ5EC7/iTN+bIAFN/e0S3tRkhDZ+TXuD5LV3MzonoQUQ
ZrmSOky+CAtfeRce9AnAIeqK06eVq9Rl6/55rF8SGGqVDh9q+knERFmP7fJxO8DARUGctw35c/dq
y/gwE+uFRB3xoBl9COg1oYXO7Ono/DTO6CsjvhoLfyxERm06zcQ35FTFTri3eEQXfCrf9cXJCUrZ
eRmihUEFvEITu7cI7oy0Q26sB2E0YKuVr+wV+TeCwQQ7wZFARp1iLl1Hwmw/JvVQCZNmb7hZ1IQf
rK2h6+FlZe5BCnLptGu+Ytuna82xyKW6yE2mkfZ3a6xNXSy5zs0lHHW2q6Gqbf40ua8b2WFSbsip
Wt8IPaF+HRgkXlG5XLP2snVzxJhPFwVwmBTFHW1qzh0m7SA7ChaXPIYFsguhBCEa+5QPNgwcsLLv
iN76kv27+6T8a8KsqFSuMQPIhH80b5p02u99DQ7B4z2mMVzTuuvyR7Ei5WysROHhRmoRp5toNZQW
sjVMVJRKzVpza9JS/gyBAVOt2gTCW5p88aITOss93mX6zVqQT+GAk+MGWyL/d9p7S4JXiSdS9cJD
v3SrX1xv5JrjHetzMYCa0BEvs7FzT9GiVGIh13zBVGpNypvbx6Bjtl4xqYL2qLttRDqnKHeSH9S4
CnKVFerpByqjDzk3n3RWJa2A3qb/N/UT3Czs7ypjE3NOCelENXDCrBTy0BTd5OdzzNqCGiPGW2BF
lCpYkRO5od/KwjXdTMDhNzB3bY45BOnPtk5kuwyomBvBzLBURXc4LmD/xaFEWdIjjTtMoxqBm9n4
NUIRXtGy4N6Y+/D4LN+FDNOffIbFIZSimBPwJCH5UhlJyWNs2a6MlT0nkPbcTd5sr//vNf6yYBrA
pi4iQciiu6hni5Cw4G1Btepx57MpF/vPjijA9GPFYafX8LA6/N0R15Us8mGrq8Ht6mBwmbK1Iysq
NDvXOCvCgDdJuUy4oOH0LXfm8NG9BhC+d5r/pSculPaWr2X6IylIbpI4Kqnf9lYce8VR1eqaMZgw
wfDr2IRgzbV/GrqtjNZW3Aoz6ndhIRgcJG+COob234FPsWoRpqd6LSnll7fQm/tdP08fQ8RFjofa
Iyd4IpFVPNthtQFJhYIeVMz+Fwvr52C3Ggz5U63jidJ2v4CPObAPSLcGz7YcEPexzxhTvkUZTdix
iUowwAVXQwwAsfiA0L3QYfXqelEWsHWIHfP+L3xDApWLxxLNnEisJryp7hXtPljvNg97f+rNW0H9
KvKoI6MwTfX3s2Y906fKA9IwWo1zJlUgQc4VtCVW+8uGbnbU8fW7b//PgNaRR5fiyxLUIzljqvmq
WO0BMytPJqqCx+WnMIlkEJV6iuN++Kqw39zEu4U7mgHiwqXfGaOwC3UqJMQ605Ogaw94xbp7ZA6L
YOz9THNCsy49r1QOkrtG1n1mT4Y8PC3Y0lyScgi2Kmc9KL6X4PmoX9zsSyITT0+IT4+PkB2WcM+5
di5955srGlmoGAiiZEOYFWOF9xFjlaVIII4bS8wCQFYEHz8eQu3SjuiRVXoI2wKoMh6hoLCoJp0Q
h1NvoM718z8xQagDxTPZXUrVELVUnwTUg1nX641J189W1qkjgllGxwsGf2Yb+ec7yZDUGA2qryuN
uxCGerzh72mZS5R44k669CGlbT9JAnT/Wp75BdXJDK3BTRtYx6b65Zppo+LQuJPO29JMOb1vz0Gg
CcqbyiKYxjc+G7I0go+tKy3MRwj0416Aycui5JNJUudnMI0J2/4qLJ8/6wIEzwXmUjOQ+UgGkMzU
ATp/9ccqzOkYH705jGQihSUNar6+Y1LsVZf9pICGiTML4XWGLBs281dvhCHRe25zeW4d7reMCcM5
0kvpcK0csjVUrN4ikuExkNN8Sp5CYeqnlYsBmkTqm0y/O+wi71uwWrlWa0qxHfzaYviPUf5vuV35
IOpKApeVnDoo1exjZUGqIgmjslXZa5ns5+7rfTzjn+w96f3x9uAbalOll9Z3bymS3bTgzZ+VowT4
mQ5ek2/4WrdGKjKC/CfiqsT/NNlaphxAFSd5O5U34H8eC3irJqDS1v0A/FAxrh4CMadVreTzaPJ7
dQDTKROn6Xpe6GCwWlN3YWHg894Z91dOeiA4Rnr3OMgUCwqwg5XQz9vtKoI7tU67V7lrfivff5pd
jKfe+8hm+HfDN57+6+vCuT5dRMGjXd0Zl+WQ8IlCrpOg5wsso2DNM8GdVsX0tgZV1kwgvkrvgmvM
dVR2f+RGi7C+sj3bez8i6702IGB+XftxzxWozZhj7U6uqbixzPlnHssocpI2fvYVK8i/XTwRWySQ
hqkoUjJCma1ex+RPpIjpoeTcmRDznNX91zF998aiGKp8sCoQ7w+VSpuBUcZdg78tojAs+s7NLC1O
CsLXMiKpzPEeutD2+8TYlRbxzMKiHVB84KCCi+qQ0YR6lGsxeFrcota3Gne0wC7ftgSCyrABEuWS
W2hgiN/3Ks3R7aLlWETn/9MzAdDFpUNxN0epv5Hg7Jp7tzCGut7v0ktO+WRddNDBvXZyaIcoViEz
enkgeGVIfRelOC3WIZ5pAnTen3T8MYEqPL3W+p+iYXUl2ok10PD3ne50FW3ex//JdOG0ksrmnDyE
HjDBgoT8OR0P474JhCioykcP8IJKQwkegupdYfG4/YNWUrdjlD0XwSSeMAMnKicaXaLh5YkgKdC3
0ZyNccwSBkgFZAFdceHx0w4CfpKO/3xANdD2e23NSZU6+ncrNjqgX3qnDASAwi34ldb1aXwE0WmU
GsbgDNuADqcjcRA6noCJ5CnkYpDc7HDToIV2GGmIbG6rzFyVokHefHRDhAd4PIFTG9xJzDqVN+ru
Xq9AliYJi07pzpYExglriHvD534GryhMCT0GRdYim6UDNS6+3jI8vK5+u6GmyqHPUTmMvd1eCSxk
QHgqYRgibLaS8Qby4LfR6Ulr//ROYN558QYlPsKh83xEpmv3NHmNdUPXn4DR15gV2TS+7aR0YcbA
9RDRZYVSN8hfi3mQssELxXUSH7zBjRYb5ZIKtE5O3I/3cn7qhTT3NZRPibwmfs/iF1UczJtiFTiu
V+KC63ahHsi9Qmm5z3yowc97qcdMJwn2n1iyoqYEnQPC2P+ma8lU84xYw//HE5zqT/LLYh0cn4R0
QWtZU3URDAr+mup4S8JrGrcFcqGjaQwt9ARGTd0ZYfIXSh++9aG9qv5L3szPbULJOf+RA1E+p/0q
N2vNTKhn20jP5sQZNrwV8t/sVAh188gH2h98IjPXYYsFMxyb3VZ9qMgNv987fRB2MQhd7w81Mocj
FnO4Ewxp5mbowLY8/e0cZMelgv+sdxr/BjCEfkyndcekjOtRtxkTskfUW6OoNH+L4VFH3y2Esjaj
bPyhpi/dOGZB5124YjZ28VvAIfx54aFC1Y/UHHfQ7Dt3nIwVkntc+78S1u7Yi/+6XWmmoZz8JONr
PbhAiBeCivwP0T5xU+Bcz2VO8xDsTcpe0wwiGs+/wC7HKIRrv0ubPEedJ3gjyL/RGH9BhJPWlT7c
aktJVfMTkjXKVCZFQGScM/mMWi466aPyOXwp8FzTZw+wWGNk3VhfwUJwH7TqadK8PnRuT/ABo9M/
KZX6cjF+30TN/HPkKaulVK2R6BOmrRoaaOMv1UN5aJ2Uu00CPjOr3zIiAwS5Ly1xCCk1nCWqxTB/
yJKdofvnc3Y/NC/nfWLKDzvI43rWcVoRp+QSDMjSotWtltqB9ZTPXvLA8m83d0iEn5Msi689iwS+
ORYf1q/6JAZUOsPMZHdQWbcRSbIGglF1kmd/Xqe5RI8zNBZjTu3O81lWe3huLaV+SbzZxPbtlzBk
JpBK9SfcqyvqPGhtISUNtX2yHx82ACxbnUJRasaM0LQ+SUG9f7fb/o5ThHdmSuy7eV5+zZzmENOF
dJO+N3c3Sakq2C/GxLdLZg8mP085znTZWhZ3CXgLLAEwumnzhWNf6yvEk1wX8kdNJll3QADbf5Nn
M4SOY3+4doKsJVGKYT6B8vmmWg8ZGMeuTj/tJv1/GDyBuIU95oTLDeubq9vFShe748OjbuzjEeuC
HlIHiJJn1jqptzGjEphyOwyTOOvC2fbAipGcLyTFRLwz9GQrQlpitB3a0/kW2uE9IDzmmBxKXdcr
0dyQaRmRePzUT+ODwzw6NzZ7F5ScPKxQYoGdtKO0QW/PEPjnPGRKcd1YydYnvagaONuJHsemCKM8
B8E6g8Z4vshPsgWk1EiXcuJQ0IDLdaCMPHg9lBbwv5z63CiZPtrBr7Arqobvtzjmlqd6K6O8xbrn
I6aFUE9g6giicklHEpIPWV+uwyH7g6MV5vAIPHxsoEDXiyxC/1+Wyn80I0FMQf9aFBhZRfViKc6m
MCCu4DZ4FdYa7LvQsXjp9Q+zfppTU4ZEDPVDcmFz+98BOVvrv6t+ryhR0o6ggPH6VuU8jl029Y5o
RVeB8NDHuPkc8LDXoYLI4lx2/rngnTjtAaWl+4ubpjovyFhYJ/nWCctkpjBmdx8pWNAUVR5h3pp2
2qaf2qpjTP0F2Y2+B7wGWkFuPZ6sNE0W0BhEEHnpI0HSZDG7KnmAxmrnecEH5uGjOOaeLSY36HXN
HsCS5evhJdBqHslsdGlfaYVxvNQGDVcRaLb7p7iBgnHzpb/JsQAyAVkejHEg2ompcW3W/6G7zXzi
iGzhL+X7bT5zOruQEnh+lPY17Eqy1Cmktn8SZhKogCase3CB8rynTp7Q20wQxm16H6HgVdcM0Wwm
tE/9fzA7I74PYrIXnS1zJWgRq/yX+fRSh1l/5kTlHfo3xMcSDwIWf23eSRI2KICW3N38T8IQz5u3
FMQNR/pFufuTeX67ZVh/E+w0s+wgYT+bcAm72Ile9Lp2UTnM34FrtW0rD37CzCckpVXjQMRzAzLt
Y/ifb/WqjBS7QJSBm+v4RLjsIk1qRg37qFKGplcQXkAZPBKB246G8sXR2OgcRcFMhNBZ+/mvkhIk
0G0XxrOJnvj7onHEeGqN4e2ken1cn47ViQjaMXB1vLJDvG/uRVKz6iT0eReB4dS9c1kzsTHGIGsY
H6hdgz/G12l03ACdtgcghfsjWWwFjRNiaWugIlGenFDQe6zXyaC1NSD0SiJNo0XPp15Y2hry2Nf0
Elgms6Z+G20s5To9yln4dWmeKj7HGxcNM0YyemnjjoVPxgP+Q1Fx4boGZCQSW1OZu5A4v5G72N84
tHMqvQ4hX3xPkadpTZQeRTNpEFaJeWTI12evQ+neKIH99hNaq2fx2IRi9BJuGASkWFssttI6e1Sq
aX6JC1h+22YYcJnoNkZPHDIO/fmj3SxvUoy3BzjZegM2V+GuFvi+4pDAPOMJAuJtxkQI16BbpHOH
zhDXZA6WN75fdyg5g7IRWqNtydVUUipjbUaFmQZe9so0ssdKqj18tprr4QLIDbWY7xFY8ueAH9MM
T3lKIVgDFg9kzJIl4LCtZGORJ5VBYyjcC0vI9CsxVVS2GEWrP1GjYTZAioHmBqwDf7H8UR6gECRD
tL3X77CbiXDgvmL/i6qRZ8ShR7b/00uRHlAHsyxf3NeeBKRnCEd5qJriJjKWuB+QUzAc/kovvqPK
0qsLFZeOTNMSXczE1lj1JZ5H1x2cooyy3mI17qDavB56DbS+keWn19YQADV1uH5kBr2GZ0CkJYXi
2SY0t6wHcKg1KQMDeF7jk0Ag6f2t9AyZbzJa4PXeMWbYv3zT4FmgunDBaQNBUS++mWq5Y2KPj+64
dug6k1g7D0+15i+PDFGhVgeIGejSxhAyG9p1vdKs+9kJ/XZ1t3DbmTjR4Igs7JWX1Wt3vKjvaVQi
xtnCGGJZ6A2O+l0xxNK+ZaV29ueiFd0WnggjzhL+9oR1yU28+FVSrJlA40tlCb66bjry9Z1VsmOU
C0A/woXF7jlzF0TTIqHB/RVVT4tjsGKHj5eG8wquk16ucHmL9OVh9+nIgn+f69K8eKi1c2XkSdWm
WP4D5vNmPvUyg/QtAzHfi9fvcczq78Uf2TwGv9EkQjRglKfRYSJiPW4Cfp/v3zZGTbmGOFc0RFfv
Msw7/I6Xojn7P47dOkoGPmu05FcjHwraYtylEWmIBsk2h1WION6X6W98wWfz4+q+K2gXqVMEb2U9
NRq/dyCdNJ80GUHGq9i+Z2TYwYqLi0QBnWNg4RIDYhtSPawy8xYyYFv2NldeEfOvPBubNwQdB4KF
D8dWJw3v/n+m4ejgC0O1ACF8O+RGR6fpoDTNT/A5srFM8tgBFb+ssKGdhxqA9jug2V5QYsqcAv1q
0T/lwhUmeLnkEYUeiapfhwvR7xR++7olMIc8erBYWWjin/4HcxHb54Kr8BpNwR99ih4/zoCXUK/1
uvQKXJLRT7Q/lpW8s1v9qm0eCGKvaNV281hyp5omcxTx67QpvCO35XhFwRCvdGAmnKzURnEJC1Sj
qk5w+G7x4xfufv574sXnIJEEwV8BZgFBD5Cu+gkpiGUuRO0sFdccc6B1SMd1QKur7Pjeh/zYvbnj
fOgx6vVjyCZHnmhgty9i3OZ5MHCgaZ3xnUmj58v5NB0mtqAzAc8tvm8iKPFdi3hWUnjljxn7JvmF
KcZq8m25/s5BoUQkXVWNg1qM+mfw8cwqDbdwT5etQ1waJXNtJtpmvKWiKWoiLOdUAz1IbQUOu7iD
BLYff/2ZA+k6/YGy0V0FJUShQf4SMIIZUpUyIioaqr99lpEZdNvatUFyOPoKBrGlD0FP/fqrNxv6
N9es8ihsojExHBa2xKDmETs7rt0qf+gl0efEjDltkBAPqTPGmSUdaBZD2MlXOUJnWhMHJ5HJUoAZ
kr1PCJJlDaYQ+f6zHu/09rr4LAT8VZ/X+o70CyH0IiIm9bs3wDAL2PrThCa957BPTkJN9Rcv8AJa
5SgSss+CyKDDSrbFvxEQTGEgDmte15kPxHKR/ESDV6Yqa/SU//3jT2jxXsxSLnFZ1Demv2I21rBQ
NiaHAR6YfQdICe6jXKm3y8AqsLX/vaMfCvwS4iZJe+gpS7NjldXJ7mhJgjPSamr7JfeCF/2HbTe6
++fAXEF++aQN1FUr8ZKAOqeqqgO4MieShqul6i0A7riJJR4HUxDktDdT92Fqoa6aM6LUoopFW7Cq
AwxDBSEjmw30PR4kKPOQeRMR0qO5QPYC4tQbm1irOlY1wmO0XCPHgrlx1X2Z3VJeWTGlB5JYTOR9
9gIQH6IbyBYcnjBHs4G8tZwyuFEEsXgpvMBorXUYWo+nEikGNiIuAOJrWyEknBIwRoYo8hosTJio
v9D665nPwselwrWOcRuDozKNXkEB74S9vSRwYwF1ngHk0b2otTZJePtQ2b93IVhY4l5ux4orx1og
3WKTH3qKhZLfdzgXmIIgco1Ss09Gb6p+f/4p6R5dY+Td5vqcvRsV8GuHKZD/xYv+dcJVzJCVC2PH
SJG8X4wV20ksLfvQyjKoAYVbgNRgqJNYuvQRC9RU3G1eQMnCcKjdxdDPBsLMYO6Vmnf8TjWqE4Zy
X3QmOaqdjze/pU/xMFI5kvH8hhdgzVNdkdfZc8PbAc+mAoaAd7x0O/TBRmPihjgWYaE/ieBdrpXW
Rtu9TQlRTQ7/1DpCY5ZpYXZqtf9jl825OQPeyV55X7jJ7S//hSryD89nVUjHsvGTmYQcIPzvwR2r
+wulLiDGhYfcIfhj4o0RwWXxOfWcfXjWKjjq4kb/ppuN5pKWCNAV7s7H3t8iweF/SCR/BNr9XDfT
2EUDbEcYMhGA4baZmG6/x/qWJYhJqXyXTlKpbzs3SEOHPC1YT/RPrdDQjvjgeb+JBiKuacrOYdoK
fpNuicKplwadnGskl2JPFkzF9icD2JpHEHvzqxmCAI0bgiXes2F2YDnTeJQxQlLUnnM0QcJ2R8Ac
QtBzLfHKmNh6f72HTDjSLkYQhaUgYeDeIp9/CFtKBlnwYOKtoDANIiJ0NditTKfSNeffQUK2P4og
QAZUczEnPhieceya1XskeTvadf4eIYeQ9KwHHLqvt+pnr43wBBjp9f8nXlJbXqenLKRS9+MeNe1A
+vzZfXKVYjkDIm4gcXSmtCQFesHT+cHEpD7xSLKUHSuZL3Qj23f87F7UndV2vusbHVmr+tznS6TY
4qz6Rzr1StNxtN0LmMLYaUDb+R2M82fX9egEqByhotDaVE0JHjcpAidNnn1TRuVe/8jzrg4emCKC
hq4mberHguelZ8LtcZEoZmbAwK6TCy7hhPuXPPErDra7N5uIaS89ZeWFOEw/WmGmIOBxf4bvFmfe
UoGEIUdMfBu4aRNx8HNGPE8MMaDJaXpZePdMosy9S4cID2UxOm0CQ3mIc61CY/Ai8rMW/Vp8RC0p
TSz8qDDcvvsIofI94eo6gkP4KeqrZyVAS5d9bZHckJ8liUTBWJ6b5Jgsf4jKqxwjNynBFiG6hh9w
9rfz97IPVcbojSegcNri3xhtuQyMuY0nFUxphqkTLxM9nI6VOfhDbNW1AppxoSNzr0haKOaYLqxL
ppAFTUalMYih5Nz+FMa6SNJ7y6V2TU4YHj4sp0pnXJm/DH63uQTWueVy3e7f20thapdgDFKgBHlp
8973nWxqisGZpKDt9BdqzRwTxq8E3cr55jBz4DOW5rImAyf+hWT03WXzxCmq8hx9+biNIuQ7Z4ZZ
BuBFPWBtKw0R+t/Py88B47aiD0v2KND0gO2hJap9YMDrIgIEYDRSZx/VtoWcWwqf8cDgXGDiHxNf
+f6OWT6NE/AFUgpQ396t7GGZiBHDJE4Rn+312bq4vzZbdIzV8KQ3w+hBUUMbR3KwWixA8rxBHfHX
MEirmK8LYm7AnsOk5P0kom02BrK265u/rhoTBgKQSu4Va3MY7Yr/htNYdSQuPJ3wnZrvOj7h89UA
4Fh2rz20aueZ0nQLL18snVtt6GXaBtqkP/K69JNmxjU/kGmPuc60X6hfzCfE+7aNsDyQxJx8bfP+
yvRNFuDxbO9c7kmaGQcj2XjfpDFDHg75DcowAfzpIbR9f3Qj27C9Vw9Y9wSE4aYlWDbkh3QW2ETt
+V2P8iH6hyOq9toMNJ1JYopObjho8qFUyWF9AWiRSRNcSJzev6W4w+TPMi7pFrdXJy29Cwu6JZtp
6C5Q14rxuHvttUOnPVusRPzu+Fo5oZduFUwLs8XjVlDz+jugfhIrTSWJu+3HEne4wI69cS510PgX
+kN5q4ooTMYKUPNU1poiwxvuf18T0XrvA80Yy5739/kdaA7DomL8sxt8SToLk0oCvma6uq4le4r5
i3rO13ptAvNUbUo9TC1x8a7blS3650CWPwpTpeFUVfy/U536rnD4OLewz+wGVToyq1mY+AtgWTbL
+u4n1c7wt6kPn4jEnWLL1CIVFARmCrZB7WXTYUYXL1LwkoW32CzksY5QqubGq+NQiP+4rCcFscYf
M4XCxq1MfNmsJ5BfoUDE25w01uAYm87zYxJWVnlvbqo32SaknLxB8TJAAvNSrCWc2bonAT32ih+f
b9Tw+gFUNQrYJYnrTNZFseaWmpKrDzb1s8dMokDrIERmVqVIUiW+xgVduoPmplVJTmdVbA+Y+/7O
+DYbRJSVuA2trAu67UbRJYszw6VtxbRg+YRr464ur4K/Anxbpvo/06njpQ25HnAbFi1KLL46jxfU
8fqQcE2Bk4Wsu6Onbc03VgJcPThCMehp3dhrQgfr0yZX6IYSolxw6Sz5wyCbRkgfU8OGF9uk7f/8
buVdLCOSLfhQ7yh0dw2vDkn7sfSJYRWAh+a64hGE3Pvipaa1b+khls57+kKLex2npEVKvqYH/74o
KaorSVWLpTHuCTI2Wft1S3KL0JT+hTCe3zSmO35W6CjjaUz+TFPyn47rPmyOw2fIte/oB+/46AjN
zbu4Z5hIkbQ13FZItF7HPx1hhrWV850hKJvXeehKrpvcOu7+20mHgrAiEmkvQYITgBQoMpSkj1O5
QZU69tgfT2gV42dVnuAIwsX0HDd3snGQzr32WtOEYie0jBBcLW3xOhJbNWG+62wKSr5zcGvab1pN
RoX6AkGUj3V6rZCepr4Sy11x69ptH3E3MoX4G3swr3Ir2CIZzs+fq6p55mmYg/JkFrXdZVf8YXMF
FDgw8CmWAWchE57Tp61Ya2gxrJp/UlL9NkBVHsyqIgXbtfr44b/nj19/Kr9WhYiypRaENK9Nsi3I
uNa+F2rXPjo6P0wiczUJRVfIEpHtIx0aGIAQttVkDdfHfe1hhQhhYLJVg0asEQebhsqCUunCnQFS
wLXGJ2w3ZtEyA1ecdwM08Rqfk3ECF1H26J549+h9ZVuLckjH7eUimS8O/66udYd7t7VOYBGB7obK
qOyhfqgx/TtomTd65ifZVO+TpSOfUQvVM1eK0DnG7GgqyA17VtcBdxCS3FlJcIwMWJWIEeKjwJKd
f4iJT6mn7ysGgt2TvhOz/Uvx466aHRdSh0H+Re9d7Zc+wKAEqFY3qnJzCwWahNvAfFUhkHjK0CLP
sflmzy4j83pZb2ZB7aNlE3xPVOg4a+FDSgBPLD26wMGp0DMobd7sxXZ2lHnL/ybJNqk39MaBJnNZ
QzwwD6TuA4bN3OeblsfilCIlmjA1yMIJVQ6O3vR0cqTXpljMLFgI1Djaobs+ojZSuAhgryBNaQvr
YQCE2n48/AApUyVGll89AhxnHEyxiRPblNidCtDxxGKPEzX1wNJbLmaBo8e359j426iMNt89hcC2
spc4v1+bgTqVgNcbMY6XcVrjphu9YErnxguQPS1Onhf71y+YUjJLH7a3cH7tNyzohXrGcwyIdK+Z
Hh//K88cj5MaiX+bLdOzon8i1ORtcR9aIwaOrvd4f2BuEh0tSJ7VVCWSSWQ2CezqYuQwCHGIBg2p
Qt2UoTKmcyrDv0hekPKKuZQ9hpS7lMpvokcNadqEjU877lPtVOOKAlKJq00yux4Pc6OwQrpFw43m
84Px4WlSV2MnJ6zgSblOPvrTNsXkWGjSER3c9AhlAvtsQxZ6fqqVxC1NpptkIbtDvysHIs/qUTQM
KB5jA4P4qRaU0kLxgLNuXXnqhls22Ol2c5hTFAQRew1lDtMJ6ewDqhlxyCiFTaaFiUTzj/aEiOX2
BM3Xhb75YXe4jhaPffLslSFe5ERFdUYRYx9C3/nEh5u4U8RsdIfynkZdt0PNX41eiM+MTRjPCA5F
1Ffm0sCXg6W7gl9QF6/+1dTHh6oWOaoukfUfdC4JQE5ZkZlJs9QgtA2zCFgCOb8FO7PtKtrUwhFR
izeEt5jvX6DRM9wcmAl+CoV0VgaC5sY2wEtuhcVuLMm0GoQxDEZotka5zQye2kPLYB1OzjYzOLzY
CMjIKkhRYOv1CiQPMKmuxT3bvX0ZRV2wSi+m9AM9MVWpM5DjgJHVbbRddck8SgWEKVnMdi5aYzsQ
vlezj9n20DQ1iRaCWVEZpVBr4LiS0+Yh0Qsst5vd0ZpjktGNCTWx45Zedsy2p7LJ1gkKgfxPZL/x
A4HEU5c544fFCLjYOpSF5yayTAeMGp3oEaOU34rW9gbs1FPqWxwBbCYGyMBdEm+YqDhdKFxCiLCk
qPCx74FAel9O1+K0fCD0TDRPeHbyLMo+5J7zpMYk+WMQwx3zw5ovV3PUlXVKGrZPlLd4tNZCDV8a
V0mFY+OX6skpSfi7TI42RJLws6ZpQzdisRBc2iNOrOYK90PyPvE4JCfjSOnST4pcfxW5pA0UgN6E
raASL+aCbWhDej+nbTTnDXPJYaa3Mdi+HLWmTj4z+/DX6VNzaWyb52GSM5ilcosgSwmc2uOFfb8T
JKVVGjjEGwGCr5F74X57s9JZh5qz9fRCUIf60Se5sNTFQue/xF+MLRVFlkY4tP9bhEDa5k1HzvAu
0HmUWKdiqRo77vAHnqYqfSnqaKKB0RJVBSEswMCoU52Cx/y/iavHIEPftGV/j5bklijQhQar4Gwg
7u4Dg+Z1/jfm7XA9Dn6O8bYy1LfhgRAc3zePXghtdXj8sM8UgkJS8Wg2gplv0Wuq0R4B2MnUv55y
ykb+XmXuCVX2udlJQ/8lTDH0gBpht9L4F1VvAqIeidDKOgx5QJFpx9/E5TxPHfpIQOSQ6WsDBPSo
ea/iOtGlPa7Rr7tmNC4IzLbEnD00PUdpC34FOrFL6ddxjVqPslnGRF3XT98WSNCLE7i12yKE7Mce
8WA6PAVoxaABGjUgJYlUUoYMoRlmpBLkiSfujHe2xaum2RqsgU1Kifv2ca7p+BQF4qtAqQmgYyYu
480q+3ILsUuttD6XOHlRJD/+XbC9gd5UtueDnED3YhGMCfEt9mTu0Lzo1Tpyf8OKulpCw9KGOJGf
jmRInoyLs2uzvHpS1ps+8hgxxFAH0roKs7QznP5SxMFif08GjR2WGDGc4aGTvaQ5V7wOzAzXIpAi
SKiuexEK9RitzoicUF7kvf0YL6X86hyCnEiJiSCwwZO35dNcDNuV5kn745Do5GzZ5ngFs9aOtz6g
WRuEvB56Fb+R2oJigo79fVPHe+3CX2LzSRmdieq0JBNO5k/g3eg0d6MTlqmFTuVMz1HYpfDvGDAZ
v1/P6gGZJQ4KVb9XKsWQT74YIo17wYQMYYZQ+zBr0EXRwFP4Wd41IsR5/kj+ERsQPi4anllghX5p
V0ZGmeve+M0DHanrh/To/z2zSa2LjDICXIbWDBerHjj4keLRn/KNd+0HOzERX12t1UbFoUyVUd+I
q0ZgSnCg/SLC1cbmNmzyQy8+L5EA62GixvkkfbK8WbtU+NzmTO2SqK6hnhEuMECf1r2YRb1D6CnO
/4fM/ZH24S24ALLbjGfF/PQp+iqrwBWY7N9oCRYa13jPGJCrrT6UNNoCyy+q63qmIhTGoGOHICPr
cJO0BZUvyHx5CA45uure0Rvs2tMQ2p+Sb8/CblCISeB9sCv1gB88rCiS6imPfUs7/kbhHP+3gqKe
C/29X1wGFJvUwBwIljNVLfLkCHSfPgkkx8LRLPMm3fXFjTMdXn+aZwF2eyo8xjpb4puBmnZhIT1v
z9RYKOlpFTT/kH7sGxmi/G5mpAjKDSJEzvO7kLpMGFPSsVny7b7pnyfw9O/VI4Adcxbb8q8rN4OM
rMVFPRhb3tCvTcHUjONPJDETGrha1Yd5rfKhPSDmPl7bX/muXCG53KSsSstd1RdBhGkFN5uuxE16
+vw6e7caki/nWC2LwsBokvlK06s9CSDyHScIiPu+fjMvO42tZgulQTc1vHSd7/DjYmAhCvCcSWBU
VEEdSjkzDH6DkUlMsgiEMwcHjAoQEYdk4nusW7wCFI7+FBVaBiZ+N8Go2JdGk0VS41fUdygFKiep
EGX6p7vUJTqE8rcX0gmPbSNya5oriJoOXZVt9GwFYEvg2R4EtuW5cCbP1gJ8I4sT2RxgTlS4o+l4
93WIgZmG2atkGnlzlx/G6EoDbQZfvu1CQQrtBC0wbwSvab2uaXEUzqhbseptzf9LolipoGM/uaTG
YOK8wihfSFQMV4bBn/Ef3V1N/tdjTwdTpQv8thtPV3GaOGCZEGCQEgsD4Ix4rPEluB+uFbvYCHu4
2D/XYL7oINfjzBjVKmi0Vm4UerLOnZ/k2jYxsvj6dRaIuaNtQi7SFFTyvIjeXL8h1TZ/zm77LRKa
sB2E/StSl5R090n+NNbeW+94qj26tweopKJBjHy39r1P2PfMp1jlp2z4xoBFTpOpIN+0ilLJvhaJ
p9+vX6VBKoolvfNeSVCiPAkFlB+KzU+HbKNsKN6VKkpepvhyrsMsq0V+in7sdlpFgQeqhBF2pGEd
5mmP+35vnDqDZCs8yazSqqWmdSNgqMHubVhKvR5VJ6dEcFjzD/+uVjLzAu+zPfvW/rkPjUu5zUYJ
/9AAI+PoLViANmZIT/z2vdNOP/ynS2jwvyjLKA9Qn1Cvv8HwEkCpwDKXnpFJeO3HEadznaQRSsBJ
lw4u4Nc8WniNr6NP5O5LWUaGFtmlQiDNfQ0oGl8z7JkoNssLEC7r0HCDTugBgutrFmtJPAjew+T3
RM/A/bgc5No5Iw9S5CenuKR5F5HuLvBBqNYkyHyDcATwfLns8HG82WipyGtRBhNTkBLKgIWpS2s+
Cb5c3r5LzHPNgWlnFuE+quFUy3zU08z3rqrApc1oxFxJcq0A6vOUowVVK1JMWgntcI235n2fzFN1
tXHT/YWW9ICSA4WbPPcLeJoahaGRR8CabxlByqToQv75C+aHt7rEFtuYcuxAUKNi98D6v2+ZHtOW
Jrrd6jtwU7jreqBJ5NpXnLI+41DdiaWKiwu0d1ySRZWXB2UX+oRMiC8BKRbzsKy0eLrIWIKIiTzs
U5k1v0IKrHlWatgbU9EHIyKuL2LDUF5UdJl2hbtikwZ6jokzbOL0DzYseetpuLG7W3owjMpyVRV+
r3dX8XbiGchdpy8PWG/U0DSTiLfoqS6SeRa7daiV4qYUo3g+ranThIrig46dFOx9S/saJAhZIqOJ
Ya6BZLU6lv+icGzOVJTC/TotCsitseib/awZo61zTV/JhJElc08IsX2JvY0RRsDPKfk9kp7HcwQE
whIulNyPC5rQC+JnR9CN/DiL0h56bNNfJ45lYJFieuPtVnmztSrMNS4VMOGUy67JEzh95QZXhsZW
E4XWBeeERY2jboSrCsWCUupnlg9vUwIPn71DEVD0Hztjguol9Z8I1OjPjvV8JdU1qzRTFUBLMfOu
3G474+AwK+UI/qpJCXNdZWFIaEF2j5HjemvaCjr3wS/g5gjZ4lCSIqYyQDiwPuHVz8YEJSYx3z9v
O3NP5BDXPeVG7Le4nItQFopehwiA8DhHJ5nf6JFb2NhXqKWejCJIJSpUe2WYzC+0qa1IrEikN4IT
qJshsgoU2n5hnB78MeT/zTr6AyRxsGiQV2+cifQMFiCiVS99z89dsAeslnLhuwqfTHjNL+CCnizq
m0BO/bqRYTT0rUcUCrsFASS9isqiyeOzviqbLW/m3CtwYKRod/a3gRcqiBYfzpwfu4b0lEayJq4F
NNEQeVZsPnluzVVQ5rqs4MlHggNkD/au9/5/5piCOKSau590FIOakcZkumqJRnqkyaYU267qbPSW
ZCJq/UZCsglscl4GCihHla3Mtc+17NXuzLiUFDynehuBETSJVSPm/mNIoke/RV924ru6DyifkQf8
AXqt+zJ8eDpoecYeyiWYryWrf6f/HLu7njXYXROrXvlT9zDzqyMaOpLiX///BBt70iyRbzle1zWr
XWmUIYevW4UafkMwkmTaK6DG/hiCKmQiBLddmBr74T1IX9QTAHE9JuFG1Qw6HeU4lajvCDdggNtt
MBJLSGsjo3Fe8HytNkg+NYt18fWTGO8PlYTx0fEBhw75NdyqTz+BM84byZXurm9vTMsF7LwcczeF
SEn5leslaQPG3V0c6z5h/XYGmVkEUA+V3Q82ixVT7a/n2jIWr/Dk5/wE87ijUKrzUqikQsLPVIHd
XyagsFfrx8gymmVBV92UVfyTbZ7uPEYR3c13sidVEEV58PQWxYy8Y7QxgSA4MO7TzrNc8yQbhbTe
lWfFdI7mVy3GHHvCBIuvKut/U13KmvK9Y9KQm+TUylexbVUJh67RbSzDk0ituQ/vKrxnxa0lh98q
Fu7aTfxZGGmYvwSUYGCMw5nySdmhCdyXArwmY61XWu8BW+6HQE5NxRboJNTZvQwbmv33jJQoTXER
Eg2Q+u8C+dGf8vmrCYKDHglkoRXRrobV4duPcXyKNyZ+CEz1ttHap+REx+IXAY58BNECMuizhUzn
26TD2laGxCTIvVZhNSUVi+NYEsKgycuX8Fs9vIzqBoXwl0L9xdTYO5hKi5aMo3fAXcw7De2SPVmC
NIMIiFODbXg0MoetvcHb5UTkyEfvrqtE4wi18YavsmZ/rIplbgEDa5Pi24hB34SAhHWB3ncaLcQj
/zKWzScClndHCEWxWdnW998Hp891JhefzW4G/ahwIsXCzZbzx6DqIXzrabGh0KegkBSmw6HwqB3O
VtViBAhpMs/zFZcC2P738BwW0HlHJ1/DCsCRu73UadXr6u47pHWTkD59inpJn/f5icM2jgcsujeb
DIgAtCqCTVSzswP+25NvgftRcokNf29jflyN5WH+ybfujkJfGKFN/ZqToE5CZli7xbmEuAJ8FZxL
v8QmFPnSof7ib9U+a+wm+/5wr0ORQlK5XZSDzlLAY8Z0chobL1I4GNftNieUvqJTBwsnulJC24p8
EnIhhOM5UvlOXPIglFUtuhimpFGwWdBopoeb6QlLigZzh6W+T8uXQKmI3WeGdEJiX6riA6RXERLH
h8DIxGcMha0eMDJQ/yq4Jrd0MO2tfGDytJe2irriZmQh8+9n3yKtI/v59eY3lhkzulm4BGRM3Xra
Nm4p20CUTQdiDbKH4KKvEiXULWi5LEilVM0O61jev/4HBUy4WcOijVmtRLH7tGd7L1Od9hnS3v6E
Ld/0K2KIOjhHUGVL+H1emLQN6008rZiCv0e73+W/eONN8isZ6Xl+liz3U3tZJHCs5qeOYbu57eO9
M4LA7YNzZRO4aLVsagzOVfJjoPOuvEaBeK+4/TJuX4IJ09TnPN4MxS54GrkilAbzzDUgP4s3FEh5
2hcwrnP9FyQtbGe7yM+1tjsn7mmnb8+ubSogz2H57gd4DNXbT6opnJZjOucX+TE8qOuuzkFKOs6x
uzkDPv5+noeq6E0QI29eflAZnmaKjBqrUN/yqbvK0YwHuuwqoklkc6RgvZy9SLYCACiuKQzN0518
aPBRH7EkV/+1Z0V8qsfV+bCm2c8mOgCdNH9NVLUTton/qTpzMvTCYcvH89HfCFKq9IqfhnEaoAZd
xRy1Jv7zfV7iBOejqInUtxK1x8o9ixbcUYsEVKZiVrW6/2eCHL+uZN7w7Whhf5ziasAYFPPuUfAG
m0YY2oxFrDk7b+nRUGeuv2Mz8VAhJQsinR/rLtfSK7vcncw2Yrt3+221MxTsPbuW8TtyLwwGz8H3
Zy6yj6f3crGwMsVweW2bOGVOhDZ1BgUxrkjMoZhDATnWM97xrV/pHzTIfaZV2Aeg7aYAYyxCBqbH
CXtlqCeLttsQY7+3ODO6hLCcL7P4XFVpxL4fnS9rFOkvpHcIlyB3DzDJEieTYbOeBR9QHyYiEhcb
CMno0jChslBXpkFtkJ4Y7M4e5nG9IXa+QK86west+YpLiBJ5slzAj1hufVgTLSuTkvGyBqoPOxGv
IVoygETyZHsEOSBtjNX/o4sZ/PiLQVqUx/seT19/Q875O89FAxKFxQEXv1vQbgVR64LIt5YlFwvn
2QnpF0d/RfwrvIeGVTeX3vfpnxu6eui072SBrB5GCOdccd1TmrkeXAESkeOPC13JArjc44IBFPK8
2+WmL8+6t+VOIJNZY6veL7ffycnyfnfzhRwnQfc5DqnDdOhMmHxzSqcMtmqdTm9SmGsGCu0j0Zgx
iiJ9c/EYVpBV+oIRJMg85Bn3hXwTVe9cRVtx+FuCtjo0JNxIwpYCpaVpUVNq665GitJMa3ZXqxyL
wF3k2bC8fwW+denz1YjcQbtjB1AmKXY1eWX6VB6BSqKKBGiCZhMKQI2T051N40uQ9eY0LVszKxFw
uEjX3N6z8guTa69VvQjHnaUz9Hb45EJRN+LBroN4/UVCy1uEGKqiWBzl0/+VyBxcm6SaKB5MiJct
1aQXkqvo3uzcAxPzyHuqOS+7MTJy+WaoftANzbHn1kDMCId8hN+FM4PKqhZZNnS8l9i4wdUkG3VI
duTS9DaLGc7nqoKZt39HwEMPcGE5ZFQGXMmQW3NU7M7H06FdNlJqv6+tS6GjRtGis/vwPODNNnS4
XjLrc4fy7CZNNF/LJxJi5NmvWlA7+USe2c8TsUgsa4sY61qpEOIHpK81dcroD7k7/wP9Bdd8tjZa
Bv9qr78NfmJs/8rE8QqIN4ft1uvbdB1AZtiaL0MXXo11zm1X0KffArO4FFk91+PXVDTqWdO+zGE6
+IDJKWuYBWLLwrE+sD5DcvvaYXzwfnOJ70pSP/TPaMf4RhxMF8xemiRDc3+x9wosut3mJdGyTESe
CsUyvPHg6rhrAj1Kb3ZZmJ6/h1v6pxYbO4uGPTo/Tnoa0qAV1GYxr04vbe4eMm8EWUrOsh6E88IN
clM1EJ8Ream9rdHl6R/r9APqP0IqXhJf207Z+6pJsVflUZ3ohlv6PMZKKsnSpN5Qyib5MvkEAgM9
mnBLTfNS9N94EzcT7V5I9i8ejXgB/dzkk+HdS8XOIKytEISJcCiLZyydIR5zkrsho0sTYPUAQPGn
cjRrrQKj1z8s2uW5YAZyGHZRIqvQSv4dfy+cIrloAq/UN0ALgMzxz364qvVitEIgdWra9pMTjJvL
rKUxtddPu+SJ0znNwZvqFL/Qh9mLv/t5k8O4NDE/QymnMIb7NqAQdMnFhLk8VDyRW7PJbSzId10s
Qgp2QG1Q7ivKPcHQnUhz9Y6o/L2O7zGpPdCfENMvHsKl7at/+HH6YgwWGSE0Jfyz95r2USsKeziV
WGjik4f6UL7GBc8uv6JGddFez4tMjZHYHtSQzLwF30U96xfkzEysS2DslCYBCAJPB7ztVpOxB3R9
GQiXtQRajb7zEXu8fDVLdZwm0Lbb0rluhsfOLbgAWLTNxT4inXdViTK2+0PnmL4bx1rELyu9sJwN
ZQLC6NtfRMbwavaulInMnQomLiAzODkcV7V5hUX5yAc+Lcz500wdrTsD92Txrb2KEOM9pCsf/+OQ
cyblOiWhuJ+R4AV1R36Id1O1P9UQalA3K1pvNMw+kUv8HuD1zCqioOZGIl2bnxQYqM8qcMGG1q00
6uE9QcUInlzRyCX/Sa0J21x8weZtJhTLGoBvDz53XnNHawaFpCTjaUw0DOdocX937IKDsc2BAjVS
mcMbPZj+T2ou0q1pwWkC2j/yG7MNF8OQcHgWLQhaOdhaY6C6DB1qUwSp/pZcZ6aT9SewYgkROnu0
6uvNb5Ytp2JQjlkuyTEcQlSSPjYVoDkcL3rJkGoYLSKqbwvVXyeeDg+G6KvLWAMOmKvzCNGipGVe
TKl59rsACuUoGsFG/CU1AzFkKfl0X81cxdsLtkGib3biG8iZHYDBRrT/NLgpo0zL1UHTVRUGoyLM
h4Ijo7/maA81bq76dgeDFFZnhkUTOwThsiGpgUKY7xfV+7CEo9NSCghkYKnFemYJgXwRd0v0Kyj1
+HQcoMCavytYjs6SMOmLa3+Zqa5/hAmY27sh0TD+ZvezLA0e9cdzqkaKrCGQ1lbZzvvYfr3Xgnm3
OiarCOdjXWRf47Jp/xB++HCTIniV2w5XCPjzjF8wdsY8qyG2idhNGyoWwVAUbNopQheo1BCsAXHn
NxAluxM6ep3TLP43vszNz2K2QmV9B1Zzx5jo9o49zuH7f1Y3R//pb6QzsvHM9zTxBWdM3Ua3/uGR
wsjDu3kTlGgv6VP2EvCRCkexHE4gPr1YWZIdg1Kmgvrrnqbg40hrAgER7mamrEOH02ZFi0V2cNkl
HTMsQsdlIF7qLUM04pHpbMeMcZl2DU0HNZAwWjlKOKxQ2Occ6Jt9ob22mFsMFtkoaOcKigb0QDHN
Q8vj0sU80Zh9nYZfF22Mz4l+X4Nikggo/mcmq5s18UCh/dwGOkN//4byPjmRa+Tg51RS1Jbiv1mI
HiOkMZZEmw7BaehXWHWnIt4IJeR2LMs1LNZ2GnYjiHpGUPDJ0mhVQPp1pO2Ea4D8w+d+uQL9bqJN
Z43z4n+epS0d93gs9mjX17FGWwk4HAeL+HFtum4KMMoMasua4chydMPoN4X5Z2SC/TzRCxNAvVtO
n4Seud61kUqC4iHeQKFzCwG7f7CdpoAiljSTbxbGKXown4HYuB6zATVNQSkIxud5sLSqvroxPmFG
prZ9nZO7nBV03XrqKl9uyKFzH1SGSO2/9LPRB8W0uvNkoVd5bPjkkfEIWRfDK1/AcCAUp6Fej6r1
FsyEUMcHAWLmRkgy64U6cv9zwutE3sjdl3v9cqfutMUx07IWB5wFd76eE0ka2kJcGuSDTxweLORB
GVxcexOFx9QZs6EQgWhE1L6+JGXQIV5ffdVXL047EyjpVPlSVJsXwr0gksPwG91opSbsJrHyDGFX
wdULW1CsCAQqRNIVXF8YCJ4TvFgYWdvpMLeXDKKjr24TU4jYhA9kzJ32Ckr40KRO+FLFtubTD6wy
+X9XlnLJn3+0ZqG5vCTKWGqdwC+PNaJwmGTp9Rs42c863qQuIe7XzzfPRf7LfdeYsbH8nmJjgYnn
8GXCciQXjeYcykJ+Z+CwgS4P38xnCmFpnCWLfhd/BP7Zo1DmEdssAIaixjAG32K8V/QlfCzFt6pV
No0XETYV3A2PapE5aqXGAnEOcQHCXRVSpfSVaVn2c5UuMVpEa/Ub/xCcxw3cM3wGsRSWORwaL04W
zrpRLuoZNWnB2gkvzbn007VrTNWv3h8jeKl7Z/zk9SmyLpA9AhQAkcDjetk71ZMY2MF4ztI7UcgE
9WpbBDL8UKqEICWjq3nbe1hfgG56Woix7QydH/4rHFbdjAFTokOw3KFZ9exHuFzDPZ9NOr//EL1X
RIn798dQwaUdqOTl/RJEgLKU0xW0GOqdgX171uzsk32CDMHqdp3QtzZMeqhoMFFpCuBI3nEeCIPn
uPWZGnKdNcqyWNb3f8EIiPWMa5edfh+c+DFaWt1dSZwU4jNWitqX3gyGd0ekDvBr3xFHfUh0CNdv
FEMqlsm/794clok976bx3lm9cW0QVNpHrE6R56X8OitYtmbLov7Ug32EEC5HCydiw4RygIVsiN0T
3TBNf6WX69sv/2gUs3bzWtIuiKHJeMowjywCAofYbzGHJYu2JGiAYiYlOfY6yRApsoDe3yk+B8zy
lgq/lzy7quW/+DqZp9hn8CmiPbxAfE+bbdKM47gdPgq3C4UR8yqQxP+DJntuAvhim3YHm6WCBM2l
wU1F5wGEViseGkLLuFmbahuFlIVkelDvrKOUWLOatRqCJNJVvgwNGbHLYDWe54PlE66KFZW6Jvv3
DHC3rFE3JCP7qOR1AgRRlI+DCa+qo4J6dxwY5hBtjeuKsJUk9fpD3INktg7rwYEg8e/uV2Zf0R0L
bwml7MTCJq4L/xmg7YhlsJOLBgRZKKKKGDPfBp8lcAAicUc7Ds+qAiUXVlfQuDlU1epRWe3y0h5G
r9pziiAhW0L35xLYdEO3HbB8gCv97vEPD/0idDY2uFaKRnX8HFYB6EK55b6A6rxrQsRijMxZbXQu
t4Y+cIq7e5obyC5L552Nsr459B3q+5Pat0WKhrX+YRL8GzodlOEhd39+6+lP6XrudrLOdyyyUgZa
DYwY2j3mAQioUirtgRfPWjW+yWdyfXdVl9b2lDznTVc/BwcBQYtSpW8s1kTA0FvuwNg/9SGtDExN
+ZNXLfW5RdGifMqBo64tyrbt5jaRlJ33/n+HR9isTb2kKXZeB/3KwRInwS+in6ujrJj1hrzC+d3F
5nD61VfG5u/vNT5u5MXQM33SHR7YvzNXipKrCiY8blkC9XY/NogZEeMDdv2duOhmSKuFcYLS48Na
gjkQTuIjeubSSlKfQ4NgbzXPugaIZfmtTrRheXjcmvEwxnG+lo94gBhvLC/jR8c61Pkrl8UaKJEJ
/yBWHnrO+/63By3qSxWnJcfrVZJ45PJTp1PISXE97GFL6AacVSF/2SQwj73wejgHUqPLkEAWd+3T
F+r0dHlUoWNU5BwaU5qLK67PWD8rdr2GPzTXVIVHuqyq9UxG7gqevryT3G/FzOikP9ylkPgVinES
0T5nyKtEiS0tGBgvMwnQazc/kCWGs321ZUyIWQi/uQ4y3w5/1hopsowWK6orhvRBkBMbojvUKS+a
tvjwfPVs7R7qIfgnhcFv+/QbJ8GoDpXPL2DgTGAqqOES6bY8hXUuy7rtcidM3wjcWfSmnAMVO1Br
gVIuuO19hi/rOh6c/60Fd95I5VVnNYb0g2KrTF4zx/9yVxV5vUtGZ7Ws1SCByL1ZS8LMSUaBgJ5U
ETnXKAMjouHbTFVuNXVpC1YhvJIFk5GDRno6A2eQTPXq3uwCTnUbUAY1kVKrxhHI7+GowHUxwO3c
PkXD6Q9LLlYwnKaIr/bo1M7nUqOyRjEYnhecfB7iHqwUTrJsKDjtvpaxacf3YButh65mxkrp9+vb
3LdvFXQzqgokoPciIVSF9nOt2tjqzaQI+lGknOTAH5BzkL3HohmcRmzTvRvb9W+cP6iiZLDXRZfi
8j4uHqhK1DHXH9yQQAZhdfadtQWHlyu0tm69B35af1imNSwaU5vpPNglT5L+7IIyCBIWpshcYb+W
bdGar2w8JI1h1vdeSGuywjMoUYOmdFrzdo8Dv46SZfiaQbOajh+ASp9NvNehcgjngmb2b8+S6VUJ
1rCcFOhI1/fer/hJ56DEDcen/kcth8kd9WV6UfTesEgBjwxO6BR8zYNK7MnB/JdZYIU7b6HmYGGe
1sRXno4MdYdKPLvR/3qpEsOmFgMdrr5f8cIStOSJSMlbWTM512yMBpkYkc5ZFp1vof22pjudsFEp
BH6IjB5DndKYCYHbKjCpE4bXhVsh+v2aHlSPEtOw4bAS9GQ4jLLP5Wf5788JJT5suhoc8D+Cs9Sf
j62X1R9Qn6cSQd/+JTNNh6v5472uRAyks+XIiILKyXqmB/DGgaVsotnA+NV+fsV4wlBuZgz8I5fz
d/OfwHFECh3hoQdS3WbI9G9UhZJdArFfw7ll8NqIGZJA2CJp7ijSeiGqt6GVDIe0euh0C1PYexNk
HDiidZwT72BbNYQNopmuLaUvkjxkkxl6GJztWk6RQkXBSXszoZHL1Vpa7f9Aks1dA91t5PE5KJyx
NTm1FJWREEDRH6EVOuiPjDs5XQtiZp2Xe+fGndob9RMQ2NcukJU5SAihCh2EnjtnwFAruNAfxrQu
PlyWRze9RPqaS0agSPc2/mjXdUqsYj4u8S+jerLIXe2g/U1l6szz8GHyYMnHCUuW+EdQki2OsRmF
/hamZRl/OssX4QbAUpAUkN6tp7c8t6zg/Ogg0+y5jfL4EloKr1TX9LIKXQpX5QMY/EwOE2yFfPWB
EaWg8RFWJHxtFN/AUL78VUwO1OSewv+qYX8dlDcbyPDATzwTEUx1ke1uM4FMdg/B7XlZtEyC0srW
Q6xO+f07YPI7PiDxZetT3V3kTjJgluGRLJMXIeV2fSDiP5Jx22oUfF7a7Z1QLJlkcNZeMlvEkfOw
DzkdGLO8FpWQAnM4Gbi6xHUYv0mMkGW7GMHneQ6WbbnYP+bQGw3dV7w5oJcebdbCgsjkQcjAiF10
1FHnJsWkKC4Y1XF2UYBWxz2C6WnDgE4cFSr/736UVfs1fOCMUzzlbmDRqhTjCf4beafcDE8i5FJD
9RJsjiDmb2ih51VGdUfzfMr2W1wEWOAyPHRE3u27Kz7x81zTb5NrBaZn05vnixpDhjg8umE/Q2in
tXNuDKgSETdejvDCycViXQZYgObfNSisoVAl2P8cuKBph7giq8YVl6qc8Dp3TmwT5OAvxoBtMY/8
bJMVSjCbjsx4/hfnkkiJW1uDWhSsRwZbVqSJFt+dyDVa7w0pLRqgbkwuFhMoBYM3azOwZ1Ntz8nX
UAucolXxouuRXbq2iWCaNL6/UF+oN93/w0pJG3rHwDO4vEX42UNzhYfHbOlKQgYNVwpurwUxdJf9
/qsmWxa/ZsPtui4hBCKtvcH4lPyB8vE2y+Em5nE47578+cw57sfDdIpB5PBFlT6NTdEy6QfVSMsr
x6hQfiorXsBUblZYQKaLTKi0f6O+hT1FosmiEtbJhh9WRMKtqX27Ln0BVTpvO2LYbXMzxFawxRhc
Lab6ViDvQyjgxOeuCE8HH7QcGii3JTL2qzErrQjpemtl6cUPy/KmPfHlLVDqGHeneuJASGA4n99k
OqVWlXAeTAw27sA/TdGY1kZG6W5J0eSCQxBfNjvDvS3nvFUXHlQ5i1Rzo6q/p1sTfdlDskLvWQre
E5yhPTFBRmSkn61RVw29SYXMlYzdHYrEmC273osXcFlNsw7dZogocYFLH3Tep6nN7x80exOX5xnA
vmluS5A+yCfHCzRCp2vYgcSKCwbfsZK3ufHpK0uWn4gD4n7jDYK0WG3RCfA3xrpMPJfcnd7B4FUV
Rq6MTkVAbS/dtBLI+V+9soav/DR/oBKgxJlfNcyhcLZYvOA6HIaxuHYf5HoSuRTqt/kyO2fC1Zrn
qnK0F0n3YJOi9cJFsHWZhNMl4l3TT1qHUrRl45wMPmeqp8aUhUJagw+8DvrZP6ZEl40+gkfzA3/I
CIX/CWFq+dAGepXszT0uaT9/mfM657LHAy6KREsCkj/7w4lvmJikfn8nLGHso20A+m/afp5zhC+d
ydY4VwrL5u7McnAIXdMp/k53txBUwgo5GBdapkp5xFK2G7JExYvvY3+x8WrgXiKr/ojIcznfnZhZ
IZ5NbG48Q7cFIhArZMKZNusZvyABMJzNW7lVJXz6HUhal8OypMV0vq539jk1TLtsS5XHmmy11wSs
9Zq15ONw+ikfXf6+o5mqX+xRh0O2XsWWGaEusvUBxVhecqSTGj57jXk/2OmrONs4FcU1Y6FXl+lg
66X3EFwUYRFhsZHmeoLC+CK+CieuZL+bZpGVSShb6y6FKNfqn3o8XC832+X6b+wjTpqxOKIfKS9j
qaoMn319WIvXfBzBslo36pBndhQza14zYAPGdKSGRvbb0kHqDwNXg3v04i5zorP380SqpdW0iFJ7
aIcrACr3o+MgMRV9YxHnQ6HH9FilIpybhbHacQAVTk373gPVwCpLzoUewGivp275jXw1yIVViiey
BU8uS7BVQ0BvWWKAGQcyE5nSkgpS2k8yqrGm9UmBXP9++vFZZTCC5vpN2oQjA4Iugu74Vt1tLy3H
4W+B2KZPA713fuA2jqDBN++6VTyDBIrwu3SKntI47aI0ciXFfdXgmzjaeqMQpMwbW5rPJ2eIItDi
wgf5R/SW7W/8zRqAIEzAdNZ/K9+j0peUzCB4CDMWO0gRMC/yPa+jFcdhhsy+5dj7vBntCRImjOOX
zn5HY7e1KQwe9wdcNQaRqwhOFBiB82pqElGG57Rp3jRd4nzuOMItSf1AP0HgruFkNm518X5362Ny
jaBehbJwm+8hKDFiJd36i27WYX6cJcQ8rOma4VCR5Eg2ZTbQPwhImY0a1XryFm7KfNuQEdxepQ8N
eoFfgFlc6ObnZ0Kq7qxIixJfETWQERUUJJ9W2gSYJnL7CopjlMdlwmxjY4sufGA+sEd6BaGUxkXR
6gHW3ZtyU+FuEilAJeKWW70IvpE4zjZ+WZEn4hpdw1SUUG8qVBpyYhEzGm6VJUvLLsczro+SoGM6
/rJ9OF+JffBi83u8hiecJYpM0qNr93Mcimmx0IguXjjeNPUNuioW9maMcN9RAGRnIyty4aGAZXlf
px/uaDY3VKPOOxFGrVaduKv1Z2zPUuy7/lnNa4qKpnf3KxKrFkjY7QMNbrY2IzgPAk5Y/tXZxEVH
xh/kEU2K6ayTFpDXwyob2RksdN5zPWUvacjUxSdQB2jaoBpVO0z5p0S8dPgKmfeCu3DBw/ZAufMl
Uycb6FL6+x90aDP4ZkmikcmdR2oMpYBXpfqfso2S4FPEkXEovTgd383uNXmBJp/tIRu3NvKjzQdK
pXeuSNKPzFRusREBqx3/BTwMNZ9h+/mlQJJCKl6ima/EiQXdd2/4L2FkR+fqIHvF8jTzb2c+C6d5
3jpUIwHsMLi8unCB3yAPZatJUKrkS8h15UUnz7kYHtcVubpZRXRQt+tBqtFXL3auoIuFokcNzOim
YBp2osP1/gyCOjBf2sRg0gQ2tiNaTWfPXn19hwII0vpDT2HiS76z7ml8GnlWKjf0i3h4OTNQ/exP
EiMvbx5UGf9XpBEsmN5pWsphCgqJegX0CeDF23b9tg2W3cxduyFC0ddIxO5cEBo4ojNQ8yf2pKK6
/2/AHOUIShKrkYoix6k/PIbrocf/X1f6iUC99Sm4YzJaBj3zEs861Mr7ZLOr4DucSFxregCCbXYX
HY6AIP8sJMal4lgtTEoxDwPld1uPgXXKzEfct0QKxcpADTTT/GPoYuetMwfSobQ9URtClMqZfbNb
0ytLqrXVqQGIjbWo0SwPnp5hOSWSfMOf8GSqQGFI2t28iMcFSX2rPJlGCc3kY5qbCZQsOvVEIcxz
FQ14+8z50/oa/knJjCsgTe083HVslxa1bFSt5CzvRjc9MjO8YsvkjzXtuK4VUCTZJh3OjIx52rfl
4H+tl3zaX3diYOd7VCZXeNe0zsqABKQlVZj9gv3+SIRdVx/3dE0NEbz+EmRZlhQg3WLbLKhTQyyG
Cm6VRl9loRZe/0N/Upr6oOoFMxeTtl+V58dhiSTyHn4R7x6d+qDONeRG8SWBBC25mhTfndYE7bic
i2FdqpuECU7+BLbS9qfV/LlRvLX/WkLdRt7N0SyJSrV2AF4eS5QfKgURslfgYdNjiEEWHdhCzUJZ
9l82D04hRu1sL9i+ImY2B/5i7AsWydxisojZ2/TPfg1Gnh5rJB2gqgFbWR5Zep2WJq43lxA2yrH5
l0w8oo5zi+JkUoC/MN9R4mENS/168JiGqEk/F9/oEKsy6bi5UsGrbXgun+kEyRtGqF08dAaOhHjf
9OxGNE4KSJAYjncVbIQ1vtLXWAzK3IV9eCFl5osR+9/ZFIobReGlThrASAY2J56lf+8wM8Ymn55X
a/PLmjvQODZBGqMWlTkccE4nYpypNCGTshYDBjsl/Jzst7xtKc/WHZQRF0UjKXQ+PeJ5naeMLlv0
8jVTKI4E5VWRbiOCg4yJ8VbW72itDu1QNrfm3bIDjmucKNLX5bpaZSNuTkKydbzlGyq/25RWMLge
cY4ZTtmZorC3vY/9PQd1OE8AjWM4fxeCo9Bbclz+MV6Q4IJZyP+PBz1il2a+uaYjUzKXNwdja3B7
pgB5gq1bQwTcXOHZDNRiWOpS0JOQnZCPuKRMMT6bvULlcqzeeRZ562ccomL1xvic45RZlD6fsJaR
YhmPiyyGZsZRK49rA+vqGhOH3XcG2474ONJEHTbm5TrpCLpdaSxw7reprIYXVjfAAAVhIe+gsGrW
qVT8wxcZZ1tebPCnneQ1Meehi9FRhX+fEefarnGZkCZGQ4xL4hVr7tUPPSHsTZFI7zl/IukQnIsN
7xODHUIjqVsOWlgmmf8Wdn5W47+Idq4CSvuBL2hR5Ew3WLgnup72hfefarCNKTRedEcbNz9EngA7
TdYZ747vUorDIJRpcjD4//3RHVKCzDVdTTCjP99B0bqW4yNg6Sx18NPn+WBIidgJZK31vEG8Fq4N
3U2fp71Dv8xp3MgCuaQQ6ShtNxydq6q/Yr5MCZ0g5N1w622kpkgxiOYETDeeqyTuMAjrvX9srl7I
H6EI72WShm/LJyoh+kWC0QLf33rvSUDMn9evpLGMnpPurUvEUS3trsMZyePadulydDUMejfelx78
gWoYYmV4M3oC2I0SuvgAI57GsRrEMeC9ErudPYywKqge1OWF6FEDhs5nPI6dfA+p+9Dlk/c1vPs+
d2VCDABRTGrIB/V1tCa8rAXH9tKRahUR3qYU9TukkzVeyGY79+0xKJBx+WsMknMHZw+woYOW5oR1
6uKA+q4FZeNjUok2Hanbo3QG5ZubcA03OIygDaDlowBkvtY+9cgJFO4HITaFB4RQDkoiKtL5eRdK
4jF/Jo8gbrde45zdXB7ZfLW1mpH2L5361otfY3FI1Cr240Dw0L+C16dGRbh3goAJyr6hgCHX068X
K6qni+cfM2WkesL4jYSzsKq3K63IjSZnTv4BGYmASkMlnfZfgqmOuA7hvR8B+QB/HrI/8OF5J6Ft
n+Cx5nPlYBcPsKFh7hS57mRouNWHGamtu4N2DhCINM7FjnsdxjT2U4VbjCx7qcL/UrXTxBvNgYxw
m0RUFy+RP11PZZEUXnU2WwzSNPC0BiRj6itvmAJDkQ0ql8BkDMv7p6p72AFnGFEYH4H2iCcjc7Qd
9vC8DPvnMSBmc2DTgmZFX6dNcbj8JTIDpnKL+kXoitNQZU0q+LbfNrcW4OlsTwogTkXFNkZnxeHF
3/4BHcmiy8Z2ZHjkT4IN6XobYn2ciI6nLrA36dayp326Y+jqILS6FfI+i0frTrcSYC6eHqn2gkUa
8nMmY7pGyuHFtSXY+/uSu7JZvySZ3DEu5tSqKG0C5LV0c+tBiX5rHiHrHvbZStZK7FP8NbjXCkqv
n+4Diz/Whz75W/T5/3MDWxYM1RgKMfbhemUqUWi1srJbSg8bFgojO+NvIAmDXaBMvphCGQ3Y0BwX
0sz13LSso3asLvDDiGCEB1EUZAUNvuHDr81eXkIjFMiINoHGvkGZX6efqB9NfKaa8JC9WClUNbuU
63NTxujEU6C3HjFFULxjuSgMw1ekn5S9zg8/e+tSe2oj0SRsw585NVOIapSl/ErotjDxI4gURXVp
9xN8FgpLytiD7dhjEhvCeIuF+n67F6tA2SK8dwPb5DGuw+ytcwUVkcmi8TMvXLpXitt2RTIRN+Uv
4gjwlKiHDkPElNG9EdxdBiXstl/plEVfH/MnkDsJ7gchGacG2Ds3sGqfM6pNlOY6fcuveF21Jfl8
hIl3yy+DvJS12ZIC8xM0ZUCc698h0p3Vz03LJ3npldo1b7X0Mo3Uc4hFfMByNQuzuuiJBBuntNxu
gHx1pQHRcvNWsdojHBYcrjYiTN0sPdNgIB05skNo3HyC33NH5DxLqh/uNrqw6+C5SbYNmqFRv56u
SpIJIO+DBBvilvAEPfyLY6rU+/SwTKd3myDh51EkNUChMa2jUlyN4SXexUsuyFKhjpPtKypBaBHQ
B97TiagW7mAO1uTm5NEIzLZvOYTWzatmMZQLIaddNRu8Y50qKhGTZPPltkStqQ96khZjkyJxUF4q
Ema7F3JSknPF3s34jlybnSECYPd8ufNIc/QLJHSZvRAdMsYz9Fjz4bwLQWl+40LJtFEpTF00BEbV
6n9QzlecRjxXdU1Y1NeK0xsYSkRFEJttAje1ousEqXcJhNnI5h2bet8hny248pn7tIP+pV4xRzim
I4jTf0GJmRNCH+lY7KojTYFpMmH5SrHTmm6SoukhPHIyePWtxjdCr8uPq9q3nMO/LuFtk+rKgfBb
6q0ddufXx/+xRLCwEdDROC+JDgrNlBSjvniQfWZja4Ain7Lb+O4jV/OOoUh5nQ29we+FRxuRg78W
75lPbgBVM5yAlliWn3u5LDr7jChGer8qpNHvvPFRHyLI81hyJlOKbx2qIJYC2uArXbhaFGR/8Ps0
5m1L3rOlWSkR1IYOJKPCEvLmSJOvzIt0U7sY8bKpXtW2fh7Ary4dWqNPus4R3FHfyYuiQh+QlOj6
RUPeiLEJMDO7G4dTkU9K0NyyoQQ5KtNDoM1eyzslzxQu2YnvofvK75fmLxkTf1YojmwaxDa86NZR
LBbSdO4jENLWwlG/gdRAy/ieiOQ5BsM8Ne7YyE3YkrCTTSGVtUX+QQJqgYjwfq2ubUR6F1w34Q58
BWcv5sZZDJteY1XImwHoOSZXF1EEwgH0MSNG+Oy7HeX7MbLy+Ckm849bdE2ecNQ5KqSaRLODyUnS
Xiscx9+HauwHduGLu1O7+5Cye2Tz9BiiaOomd/ki7zojb4mAnDuuz+9+0eyi+nKNJJvOVctmvCBU
2UDgxZY4xfJM5oMQwalBhB63nbeXFE35nUz0/Ck2k9ENYuit4nP68zsPuS4MPSE7KeYT8XOEP/Dy
IBVi2VUqYi6EP489f9rsbv1gDI2Rx4VOkj26kPtUBvwoY5+HWtN3/95q2dyCisA4ZrBDxc07sxvQ
xI/Fi6qnSjhdNhOuTC8w2Byb5c+zk948lLqwbynEZUNWjAm4P2Jfie+bE6JjKC+MPwuG3pyxGIwC
bqmX63vF/8V7tarZQPOOVzt4jh4ZhFx9n5iTITxWUb0o/sdWRq+XA/Pv1nK7p6wTXk57q7s8hIp7
BkD9yicVyBjoe8QY42CwKcKq2njMaYsl1DlyXpO2S88FLyasP+1tNPfliKdoQn5CvX0kfIQTghL+
2O2HCQGRhQZHmB7ok2oYba9FPnM3Uqd8JoW0wZDFqFGkyWFzasPDT0i6pq2bmlOKqdRZ3Q3PaS6v
/5pt7rIVM3RE//jhAKYsFpgnOht6qCPVXUC44+h+ngdI3NJqCN+3m/W7XLMgZ0Q90AOKwZStzNYS
/rrO2aZvG05x/WiqdBAwPBODs0WxPn+AA091Dg/NgIV9qi5eXofx+oUQO26jwXYfY3K2/oXWm+Hv
jiUM8za6UZJ6JW6ca+W/1S4JqxdfuXazVTlWmJ7pA73ryPhg5eSzjN1rUZTsZw6H20f1seFBFrvT
ogyZ8Twr+kV4UC7QUb6VzrdvCpvSDls3C1kNoFvRZa4NA8T2nEoLH0jvWdnCUjJYXsyKye7TpZIF
tmgIByJPUd1ztL3k2abJO012BGgSlhgm1f7Kgm/7ZL0zP1amsCrdAPCF/a94GN6f29hEbmnyzBjY
t0FxkyjhtSiRHvWEs8YS/mXWcy+Khar6YW0Ah2aGx/+o8SjOnYuxAmXpLWTipiQHl1RyCQP6YfSr
27fM8OE6wvNQUpZyrGV3LJe0OL5E955c35Gig+2M2Q1lCs+v/SIkjQ21LymEcaSWFZbnSfhixM/g
i3dvZmoAcvfR2vxoYqkdLEdAFRWGTDHUMZn1zsr4X5p2KjVtlF+dAUeYwDu30PmuCIC7UeZshp96
XVmURdI3wYJsMcEHgsiMgMckXXY1iedOY9rAXhcVp/LVYsCl4Yv2SNblhTmqSGt5wM64uMTwbiQ6
0hq2IL4NNSgK2LQxiLMYjTtrTYymB122+o6cAsQHV7eH3Amr6v3vjdZGOMks3tm7YbN1uJIbT36+
pXeIo2Zq8YMkJP6dJI4ij9xJNMCX9nhYo7aOD3NdeOphTiRZtr85DzDyRMWR01DX6gxKGD4S7W75
siO7iNqtrBZIKBH0m4yA/RKJgM85qx/V4WvQsEDY7TXu+ztBspPAhQlNDutgoQJqBjA2inhCCrba
DEUBrcPRNZlWm75yMJTJFVzfFfepcStduKgGlfJZxzmmetPXWzzG+iyI6Baq2da5oMfuuVPGW050
cAI7w9Zoc/OE+BYxgXxRJlhU1gkKGwdXWUhOe7h9OhOAC3B7Sm2K+el3syepKp5Ys7pxcUFlw+MH
0e5PZe/pC9V9TbiJxLGRQ1k6X0/gM1xIUV/oQx3eDA+xpFqoJwzT74wIHMqgf31bIIHm97Jn3LVp
SvWLYmVX2ogJs7dgOO7lgF9t07mMKmpZUbFQCVEHi7/UEXj43ghJuSyfpJ2gXsT/cWleZW+gBgED
Yjgz0yAKOoUb4+4gwPBkOyO31B4ciZhwam3bq5JkhBaIXs77rpPfadNfvHP5oBDeiTzqjg0emCiL
aeLUCMeVYKInbmv1OklsEAcdVpv55kO05uIwZPTynmNdQpxTnEMyfDwLyUl0HaXzTiAuvHlUlf/k
HxtDtOTARH8gdDvUUtEwImdKtZ1PxLy+LZOvLIGrUyZV+nTOMZy6jukAf9YzuLbrAeOSeU57QGLR
wy/uDADWFuJXbyIL927sA3rTF47hmuRU5r3xuBi7SuOM+pJN0ALVVDhPVXZd0Q5qrcsO1jZv/CjO
l5xl2bSxj71vfLUakedgHUATsfsYFf4EX83UXIh8qB83VG8CFTA+ey40FDGP+Q9PiOPlzmgRmPMj
lziUqTp4xgQBXbs0HQPAj12gP3veQ8ZcwiNXEvhFjJpforpokZjK+T45gCCYOZw0ZMkTCoD98lJ5
TmcuCdYBArQgmEkDYyT3coM/sZs30vFmGt3ZjiU9Z+lvKCWFHC85ZQJbhWRLhyuSV0nnaOpvGJ8b
D0IZwmxMW6LIVLjHw3LQdPhLLtB63I+wtZLEfOQhC8DykozH/jf9KElUqHmpAqcuDNgaUUm5PuKM
/titBpv/sYjxqPIjB/zwD1ZZPjX6hRjjEmoti/7FtsYK76L5usaqw1qWi4CM7Ac1gWHwGMuNsPWK
1RD8zAsLVfOOyBtg2GG7gh4ouWlVOTUZfK1o2zJ4qyhSYGNJg0o9bDP0pS31NFJ/SguCanEZsjjy
Sz90mHrJbXVOYYwaiRUlyvpiuB2FtHtO055ug1dhqgL9ScFli3RVXk2Ldf2uzOv4bhYHer70hhat
wO+DPUSvY7cZvrlyeMYlCY3eTJWhtA6Fo6OsGKhguPktnOuwT2q+Qa57H7w0DGpDqDc3wieFAyNu
QgvKS+nktet+P+QIVeyWfSv1t79qrK8euuFgQrPVLFEvadzbUvq78IY36nf+oeyyvylOPO8czHz3
hdVZKR2ElxMoI3Ez/FVQotCSQcy+o+ThlOa6s5JbaFILSIMx2O9Wyl6++8YytKui6SgU0IIvvOlK
Od6JG9AhbPcXAHQMi6MXskqcuU4tCppI8gY1AeDTZ162UOpv4yUiOVh3jqA3uTYvMz80McXqiZ4b
R68DIvfz4y++P0idBQhg/zdqrJIjkhLLuKZvm5fanwZ0++gCinSG0pWnNynV5yg2S7XbOGXNzJG2
6gtwcsOwSX8FnW1dpPfeFp1CSs3dCC5a1NlBb1kwwSKcADWaXvVk+Kv9h+Uxe2cv9bXZZ3JMJ6nQ
2C0ZE1Eci6lW9TDpimA3kQS6L1F8B8wRqmQFOaW9wcyJleN2Z+lLSJ5KtW/7GTrM86/ZdKapljyR
zWExYhMZloBq8WoOsdEI0QldTYrODvxR3nvVd+TLdDGz/Wyngsg10HIj6O8zjLeF5VRQ/ws0cn5c
3LG7y4guwcggOku2y3EoSNflnfyi8P79vVbWojo3s1Bs4jy6TMy/WEZ6bS7bWUeKEHDRB7KKvq7p
Vs9j+eunLbM7eSqhgVtNhqzjoA+SGaWLHuf8W7/CyzHt3fDK3RS5NZuIn/FUG7+3/Zl5puKGmaRV
Bbm0ecjvM3qUiqZUtEj4gPLg/sxPl+ZlTC5gjBqNjIT+AsBMhQyYykwDdZRISkLuzXZ4M5oxTdTC
6TcWsYlv3M5p4b05JUoScyjcFwnDV/3pkzyAt7vBA61wNYczZhB4S4RRH59EBxEJJBdpnAXFphve
VY8kbz3Q5hDyzKpVdvo404CfyI/MOcVqrKyNBj8N05YUpzysxPrqdkITfSM6ur/1oT9tRol0IBdU
OFxebxrn9Fef8mCb0ONi9D511LQrPB91i6zxI/J/9x+zyoPBBulC/xyyM52Csaxg8WzOrwBi/Pvn
ivAe5nq/o7TBA2+uiPTHiN9rXsHcP2QmA5xyVZQhL4io27SXkF4pphTOgZk5nc6wB2ow2j/G6qZu
WKKmTVmsntR/SuNGvk5twWTRXDneLFz2MU4RikzmvMvv/oTxJyoXH2xfjEWc39BYOaMFBIFsZ2OH
wsyrB6JRonf1MOW0CZmfnDExBwwCd7hoOhH8nP00Tn5tLvK1POeqsebmS84Jg6O+vgLvIK1Sfu1x
4ymT3ZQj8vHxegSHWMpaC8hfZNLWgCr1YEMtzG3bPwEs8Ps6rgxwITZng4m/ARayItRocdDBb8ZM
zUsQ63/iGcZ59Uucqw3AWQ9Gji0Nf2B29+byAnKTxQ0uoHMH/9i2t4ob0ETlsoIPcnWHR7FZdMXf
XO/86xXMBDTvVeq5heST8SNhgsa5eVWtPyHAZJaF/THHDQ+/gC1GPMbKSbAMWVeDUFLKLyAxFLbC
W3bhWgZARkpbLXh+C1cr9LMzDXqd3IQmCJ/mH45FYCxiDZ1v/HYUG3ME2mvticbsDi+nmMpTYjgZ
8COg6gynZNYZGmGN9tymRGk9aVEch9Ntl7skGmIeAiCdOabjM2Dte4D37+S4bYY4BtSU18Te0of0
xLnZ+lBiRWUl2k8Yt3e8YpL007zy1Mvf/cMYCySBnbpf2EvG+cEvrCw9mmixp7yvC+QdfAm1QHJR
bbh8k0T6zZY2A+WJjJn5iDZG/L2+g6792qXbT2dpcpuMeI6gRuoH2nWSYsVDc/EVOjOzT/mXcEz2
EQ6hsLXB1xqPKNJYl4v+avcJOmD9OfhGvLaYJ1RVGhUxmDLgklwRA1dnigrmJD2qtQyP7sJBV+wM
X+oJsqYPdEWfAjl2V7yTcZtqxBZ+/DwgDUAmanpWfU8P9+90ENb0t2xhUf3xIKeQNtkZ5hn+rfCQ
SSHcFFgGFIOeL/Ona3k0F9dI9DVpBfPpwA5lMYoyy5URi+Zze1qysYNpsBp/7wK9/+3MoDFeugUy
pIjLTQpa40wL1kVIigyRz1F7Bl4Wr/rq4Kz/Ak9EMXXk61aGNiR33s/MRn6iuB9zKPmp475FGKp9
ngJ5SARsvaiXNGuxH9qzimWUitcCfbIA2KfP0ajC2PTgIVlHfAxPM+BPWciXzF+e5cvg/DwR3Y+c
bKs63BqencP7R53RkV/vxT04268Xf9wlZHNatTqsv0t+w6HIX0Sa/3VhzUnZIna8IuF9e04EBxuN
zHnDTE6GlnoEPai+ixan9N/9HE7eY27TqjAkXDmcJTuM9wFOmp+UCC/ssFgg2C7sxUB31aLNtwhy
BOOZHNlr2Laa9pqVz+3ycLDOMAgugopFNAIl02xHS4pyFl5RW9fSMBlE62U8nAOQqRm8CTIQVsAs
Vn4Vqo100qLF4PoOgagMCY7Wf/+vh8FGbi/ZCKPwPlvP64GGO8gBpaktJ36iQfeGXVaUq/xl1Njd
AEo12p7ErEksgSnuPtmYpjh5GMdqFZ0jRWgO0x3h4tSEKx1SSEEZzNRz2YQVvM2FLCHdmN3BFNyR
vm/Svk1KC+ba0ICzdjH7uo4kX4sc8kkYoyBW23arNGr391fK+IdD/Uyep3dLjc6vto8PqLIKYjeL
k0fUAR14/2fl+tQhfdaP2BLtboIhdJCnw+gjB15WyKvO7dL+ZCEqKr2cKXNfEPPNSdXiL6VS70js
bGMFx2M3YNg+cHE9Ba3lkODmcQfEiWrB8nzOXdpMVeY/lMAizDcbxqwBrGzRkTG4MTlysjAZk0L4
wJhdYhqqnYx/lURjUOXebpZyAbrH7h1QXz+4x57y37jF54oB3hS7Xr04E98ziBRtCk5MWd4T7xY5
gen0ZryQlW85YK+oVENXS9aorkcc5AoQd92yfBK05Vu+G73Su5XCO72mzyCHOG84QWFXDAMGDiHY
dFMvY9BTzroOfeKdtP7RDryljHckb+St9a5YY3mI7L0oD//HC5srzgI7miiwBXi1CSn3tVMkCvc8
hBdKW0Ya/NCJSCBaBAoTQZJEwwQcv8TgUU8MwhVr2sS34uhh8XsZYRrF7xIhgxZa0cGQlIQKvtaP
6SOgoGfbR4yxSDViI/U/kJj7bAjrnFDlESJTkcAsNSIYIc8DPM24kdDpOjZoxseqTYBh94qzTX4M
RXUap8EbeFqC8R1IL85OqhHZ00DWnJpPRcRQy44Mc5JSOKdWBtn/RgyITf+zGl5xwbIpQ0CgpW5s
yC/HbqTy5e+j8uHu3zvsmsuYHRh7e+Ncd9dEUkYmJwWMIc1RTlLDJBpRFG2rwAY7cchFHxUVhftV
zOSh2Tdvo/EGchhxFLCt+IJB5p3TUko1hHF7HokYOtFlGJ14bY/9vYEkK2q5dAW6zFuSOh1027OO
DE759MQP8Vsyql83ZCtolKANkuxf+ovMscoaLdaxUSsPBK395xVghNvmyKAzkixKiXv20b+eDIgD
knOxdQXjX62IZuctHa0q0iKPN8dvlhPHpxBM9R5/ERkh2DvvHph4b4im6RdWUOTLYYZCf51yDJTt
XcnUrCPXzP7QSvipMr5p3ew5BNkrSFRA/iAOiiPzyYj4WIIb0qUQ2oWCZz7TVkKqXa99vRnCFQlr
nhnqmp9UkbXw0wbWb+KJu1KYtkQ/pgB3T+bTEyaD+0SH2TrTVRHNAgyM2SaneQNP7HFdlcobCVCN
r/D1EkGyE6gQ/k7QhJfOYzvl1Z7KTNz2v6mHxas81IWIyvOPIygvDV7bjNvmeQC0f3pcxrJMZ+2m
DX1hjcJhlqDf12V2IMaxkYxszWcAWLiKm1vncvxaGj05H6UqcvT4/YSqfBWxwlB384E3R9J+LThV
zAjCg7tXgiboqIBTOtzqJ+S+LPIlc6sijLLnVvwSuoEXiXIFhMlbfXkBdNUJ0qHxz35vCM1mYKsz
uKIj0klESx5d6ov/09574tOiIH3muU/FysSoKUZeR31ohBlYIdUgbZ/1h54oC+w2BHf4qFnnYyUc
nRtXL69ZaFIjvHDQD7CZymmo3kQU4UVUIb605CykxCDBBIFITQenWapmCJg4SHJTtBGENiTZ+3xB
1wzW43eCct40F7yIBN1cOzahjbx79S3cKMHCoflHCmndbg41F52BwP2bEkRhU0o0FYN+zPlx/Bh0
0m0dR+4Ttu1ccXeBZTHlD9Hz/PL3jRHTsgp3PaC4GRQ1yF99HKZjRReDLebR0Tc05kDlVmMage6b
jY1rms2FU5U6+lFACNbAUuTLZKrSJ1+Oqe1OwUrT2moUTY21yQJwHgvRoQp/KTYaLWNHcmRr7auw
VEPz8PUotszsjAwo9OTYXh2SVUy6y8CB5F7C9sw1fM0ftfh3xt+vmjg4SYq0CIq2nMhP09qR6LqO
0TrCUjOsiQvyyj8/VYnFGhF8HkLiwl81dl+z0BQxWauN8Y7KXrXGq2fpVa7lwajU7GxIp6ZM4Pux
f1sqt2EPfkeZOZjPA4VHXS9TD4bJUEcGc+BbB0YM5uZ1yJKVQ+cvTHvsYe4c1j3nLIdwgc1ev/n+
wNUS/x6bZ3BZ/lteJAQIy3QAXTpAeT+JsPp5wtoONv7mTBIH5gyxP3IZsE4nJA9i0MQ6aTp4b3RM
yUh7Se4PtypAX49+zACDciqrgqsJvP8vwoMnkC3jr1Y/zDzeqyDTGLFtSL16N3Bx4dxT0QKeVtlV
KzneEqGJThWrU15AzMS3Hz910cqK8gQNJkpLhGkBna0WaoTUqAf7/wu1nH+gLYGtDECeYfjPA8cM
uTpp1UvoidBwVpSTqOZY3hkrYhH0YBFomPIEqGQgUbG4xi4PLs/vOCLUncXYx2yYfHpBO+zvKmUA
TAq3YlIv3PLdmWw/vm2pDBiXZgKujCwLEWSMBWZ2qBu6mW6vbp5IFFx6pJcwJMOtQ0t2tOtJSCV2
dyYStNG45ToEWvIy7Wi0qofnnNEtPZem8ZHxavGQ3BIzYRngFI4S1uNcIeLfW7SQK8yHXDrKmKYU
ujVZ5FXE1RSXFchPIBCmhU8/w+XkVxC9SgIt8gSnzYQ9A4121UvO2z8ZtCNma93bI1+Iq8ZG+rsS
QgllnVX4R1eXE0LTYQuUg8mw0Rk9/1NAgjdZpvyeBbzwvIwAEE8aw6gmkdkSFRJho5BAG2MKnvI7
VP4/fLettQMdiDIbdPB+besLaSINy9/Qu6v4l6KhdLpDvpkv2z6sb4QFjEBsH9afQS27MIakCeKO
WErR0fNh9TC5ForCvA/rMHL3UIUCtn4JcVAdVpIGGb8N2D0wg7VlGaaLw0zIbOEWCzbFPwbbvsj6
PlqCML3GfS770FYYaRkZOIk9iA97z46vzxCdUHBwGvGVB1+5JhngJsZgEQbJ+ap7M4zEgB0BXi3/
PPRnPPe5R5HzEpdB3KgykFCRmR7NQoPrHBeZSgxQ0UPfmYyE6csW9Qgcrq4oZ7Wk9iziVPN7xhin
zj2llFVV2wI5eMWrmhFAkaHk4bVxfJpOYWvMhRE98R5Yiv5quu/uC07dWjRRRNZrXvC5OovaeXa2
vYylv8JLJPQdckChu9lVScu2GIJ4sePgZbqOsc7Mv36SCfEoamJ7n1RYv76Y6hwBi3MnaEtoJsOO
dUTjzxGCjZESkzL824i0wFoxlGhfU1OqlJMU7RUXlIFOC1c8oEM0SmAe5YJc50u5SlgK1p83Sx7W
DBS2vv4/UYqOg0YLzN+kgeKDn3a/8UsSETZ8TCEdJiGrnOAX+OiNlISnYWzMqjMvXpORQNreJDXi
jOtQHYghxcPuz1oBtB0UD9gIN5X9AtNDPZekuplUGE0hsqKGAOQq1ugsJYnEl+BQZGIe1mkto4CR
1pwJBhcOIWPsYRt4hTNpH5ECBZZB60RPT+hRBo/q8bC80SR71xJpjaqUVfrlTFal5HEbvrcabSMT
Rr0sgN1YB6zgrpRqi5lPywXvNzfpN48LOMk3t6SIVwviI/tQ4jnbB9hpFaNv05RWiJia8qv2dfws
+u/AeeOHt78MjAYIglz5n2/ebi4L2lwOBKj6x9jBRzNJ/yb5B20/5FXXBSGUcuViuRyjI4N4NDCQ
EE+IzfQ5saw6DNhHfwfLAUKoZxatLETuCHQyX/+zLFFoee0nLXPcPO0S1V1hAxDMEcGvOYblrw+b
PxHeTRb0fILgS41jHUkB38surPx+dBJVXsazFqPYatxvR9/+ZVnPmZun7wDZFlD5qnrpTqyxTHwx
8pfb2IJp5PFEIxXjznrJW/vlISxfuZW/T9Qdi1i5AejwM1QuSw6CS5H4cipkr8PNJmUd9sSRIVKX
bzukNMrdg37ybOIFaXZ4LcqeJrmbKrogSv6Ocu6RUElWT0a7loBO4M65EQhZLlIHlq83qrswQMkw
hA5b5Ww2nm87c/uZN7JIvvtEjrL6nRbYfwSptGlhBpklDsfJMqvT3WHi5nP8zYVBle9qSQzNrMDr
ZltGTl3WhsXk6FqdNVGg+Lw6MzCpns12DPNJH6ZzICAnk50ibXeoCOFmgNTJmjyLA536B7Lhi29w
HK608feB1IsgduPHhhv4UTo6sajVFQVwUyHfUX2z7ipeQhrgFS0yOzQvRUzY7hxPtJYmvyDcpIRr
z6fksf/sNTcrwT+DdfPHB0ZgSJvW3U0jBuRar5P5eaqaibWHWV6X9YDJn80Fv5rNUfoHDoa/gSaA
GRoVXJ99fu/UhKytfsgJymJ3FJNNRFGJJF3hJb/vgGBtuOBJqv3Ftok/ZJ3k8OQFCqzzrO5JyWd8
7m2AiJIQcvFdNYifiFMOPM52saF/F3oZ/GipfvZKY7wsbnizd3P+2ukVylPTq9J0GKKKB/8EhyfA
4yNzWyB5UfGZIdFad08KyvSrNOi2yxnzWiZeJ6w85ZTAEjEoLisKggiUgZM2B8nSzi9e7HsAbcmA
FuX1ZB5QJ0Ftx9OocGDL4IrE+q57FwP6T3a5tBEpiFVWfUTkVTBKyFGjH+AiBbXZ6fNlyp+MGV2j
xxg1E8Uy7o5NwoHa3PfwB6/1VIlJxnkqXEaWsw0R1gwbX3Xqz76Ug3SaSkYMLy5AQLyGyCC16pWR
dpLohGCG1QKk+GHLCIqKXQktpsx8TJixRBvF1dg4WqY45bDUQyr2DJSXEh3HUZbOz4Z63ZeR9wih
CwCTPppj4GYZCgdUhjyQqZleooe7Nlhq49iDoYyB378/zw20e6JV9iTEAVDtPIshaAviS2gSrfJM
4ppo/sDd3kj6Z1KTlrgkfEv+hs8a3TeRxr//FU5BnJjx4JARkkzCsORvfPfG9ewERMq6faCAYQve
XKzufaO3gWPpDWcwwOlHU5Nyz4TdYKgT8ORTGQ4+CttKxehUgLILhPpy9gwiiGPYVi28+UmXTgjt
+tiMJb4RM1KAQS2WmGP2474nFaEg222NciPgIGGE6aR3ag9JmGBgcMZYLPPBxz40CNhqlQmcXBpy
dyPs1A1MhXdBb2POrLt3GSdcK1Rbpye3lD7pnfNE1M6ZOBO3CCGIr7veFnukLCGlS054bKAmMfNW
TZEadRp1fhjofySX3oxCyXq1m3spcTwJ1P2jxKxehyTbuoQMmU6n+Z8dhfBXqYK6g7jtr335N8t9
PPbRmSsl46yyrTOBSMmI1OOxtWPXvGTLiiCR3/LDXyv1z2lSIkqEqn580fieP7e5FHgvtaYJHCPW
pFVFD7jTThL1txwNK32ubVc+kyNbPMsiiZgXlm/baOoJMjdNMRIOWQVkmsgg43lqV2PD4vzEdbBB
IJR9/bt0xsZTP9065++5Cyn2SW/yeXZzNgmHRgo/4lLYJHw7uNPHIkTOw4MJbDY4hL+262avwVSp
Jd8TROG7KdvcTS3v/YLGII4aynChsL7I0t9+57XagtadT33Op9B+xWdrCR4sA90Eli3cuCfA2ji7
OmiGv07OEyWUSoBow+6dW6UT+t9x0LX6nVGESgpWshbBFDdpm4lsLUSKvriC6jvoVXx8funGbq74
n6GA4XSjeYmN7pM/vZvcaFxJ7fQcfOE3K+UhX2qveUATt++YLUDE0k5AYDMcd1e/M9qkvSxMz9/G
ToW+8LDu8KNp6VIARMh3W6UCVWY5IcYxwvffh16RanAiIuoZaZD3mA5RfgGlv8OTKaZtB8LF49+H
T8YbAPqtoTDnXirueXxWZXS2HznUOb9MRRGARMJUPZs5D03BOD9a+rvEg+o23TPW0ob/F9ZmgRAO
MI9fkbgC6RE50sGpW4gpTQnT6e7eP5Iv5ZZpbTcuS4KgNidJDL3qXlv94A4Bf/NcTDYpXpEoXyCb
hNAhj87iO8bNCVxGq4rl3GgimL5A6lrXvPMHm92TuJO7cdU9IStI5c+K8d2Xlo2W+b6So5XskvU+
yYS1+aFotsYkCCMA6bqMKmGDnusDxFML0mvetx3qgx4DfshK/3dL8OlyWGYFEkU7nIJUGt1bdoLY
9lnEDvmtzgPyW6VgGqTuoUqGCU3wIbx3SJ9NYUPse9BodCIsPyGrRt//7W9g2JP/LCvyCebGakBP
p+yKQeEEF8S5+ljvQb6qtFPm7zl0+zlYfJyEZ+uP37iavfMI5sAuJuXd1/viOX4s9Id1iQCbBDgz
aAkcz9ph0gNkyU7Gcbbb+MBUMG6SVy4V8mYbV90Rdvh67yIp4rWQ+5FnX6j0PHHI6mMuw2IhgSQ2
Uu15KkKJaUxwE3tPNkG85T5SAKZaiYFEkke3Ph8w73NGsBc3iojAI6yEwaP7mZc8HiF4yg96wgZh
U/Qok94MY/Y5B9oA6X8zwbtqOisOCkUkNlJp4Gprx8Wab1de89i8XoJoE4L516hpVWmNDt+drFB7
y64aGFPejnw7uK1+aiFzG5T7/WdR4FJ/tdS/37wBRnuq6gqTCQYyfV5/hb3Zenre9emY8XC6JZ5u
q9mlquo6PT0Y6mz6vO4gs3mUILS8TWJRFWOGUNL2ADRYHGAoM2NL9jAEn7WtlTaWLERwJ/2UYWsE
ZXDBl1xv0wjclrPM5vpFjK+9Cc4/9PtY3eYvuy7NJaB/n5OlqIiivP8yJ+ev3Hpm/+eiHjNwGI7H
ztcMbPOqnzgk1tuqsmiE3xwIo/ylueF3oyXbchMnwUgdMBKtOWivqaMghXR9hcxSPTQRZLiLfG7v
Ot03/DORBMyxxqHqbKkJSMsYGv1A4Z9YNrUfKhOAvKEWoMrQelqH6RPB83qari9ecnzKRa6ffMJe
kxyFXWm0jD+ZtqWbMjXxeC9Vp3C0Qm44wSCKqpTpNbwzfbfMr2yv683h4oG2TFlUSelD7Wlda9Ly
ys4YMAwf3oDfDmSOtibMBn9E2mMJs6fowsPtwWZQ0YgUJZxAZ2Ljo0aOGhBSWY5WBdyFD5w/tmkP
PdlGcxhZFUBvJ6FVTWY78FTFFQ1ctfw8m337KoaYCQVrjCjmslxfzjLV46gemevASPk6ludtX9Cb
7jxoCwTSxKssWA/Pk1/j29ViUlIG0TCiTr/KRBCuNXHJ17eDMZNA+qZQQBjMXzwHFb/o+PTW7Ljd
a62851IuPp9vdyZ0T3sJRqzjm9QVMD4pRHgLm+IW9hgho49g91xZWKIbo26C3KvkU/ar+xT6h1CV
w6uhf5ko305cZA9D0mpyPOVOKRyomYcIF9S+XNgaG4SvXM6COqiodiWNekbJ+LRj/6azrZ6DYxe+
/Lie3quEJA4qCoA0huRYpPFBaSClfgEGV115Qsc+QZb6a5oXo6UEXAbvz8LJkGCRyEpsVfs5OSz3
0qru6Tf8XK1EdAUArlw8aaxEwctuA/vbhw6mx5lNg7IQZnrQW+8x7TP6vjSgqs7dAKoKD+/CWbvc
0G3xBR8MRYOeL04SYBUkfuV9U/0GY2PidOD4WD7LvEy5oSPskRp6jRl/qRAEpMrq/5UCyL3H6U50
aSXgbKNvmHkJEWpgiJLwB/RS181zZ/khrxGmYCLZECTZCC+/zRGFUba53P7Sj9Zfft9Xg+DZ73b7
MHBzi1HgPqKTRFpuxVoeSRZkqqLSOHK8UMfTf9AlENRg+TXUUMnCDiNxA0p//xIYAW77xLpaVyYv
sHPteVbXxwktJH9tdaJy8CpEHKI5M7o9KcCjfZOlhv1TeYPMf7WzdUSZ4ctpMkNEEGKfOfSOgchD
lowknLpdESi+EvqPN3aQU6SlKEAivhWkuU5dN0RUh07bbz4sSz3HuRQr4tIR73OPEgyRd5zhjFRk
pBl6sAsLw26W5g5TwJa1CP+9NrDqtMJNhlS7rpUijIz3mSNhg8NZqLtPH7XkP1j2DID3YjRUFytU
ZckkLLYeW4Vethj4++AOmIPO1N/vo9e6Z04bazIfw2RGse1SHyJTtdFSiwnB5pVs3/eIqYZi83RA
H8H8+YdSCpzkZYvzRhCBbFLGkVycICswFJFT/sBk1Ejygnz8pbsjX/0onS5wCwn1FiitJAJUqTRg
EmWxzPVYZ45OMzqlGLrStE//yuOgAocX0RDretp0bwVw/5NdqX8KJQMEkQfztOm8GXLqPbya62DY
OUv67CDuHmGl2LR5/oZrlHGohIP9HYlrHnk2v4PWWBUkQLRewtHW0gAgscahHPdVkMPTSTdJUst+
Pd4YYvxoo7/YCgyLGG2PAwHD8ainmC4xTXveIqx2zMHkQijFQmcyuBgmvS1uTL8uzmUdL44qp5tJ
EVmOU5LDQOtr/lHQd73Orlb8Qj+uXnRE9TfN/SrcyAjXO+ucu5kUvgMy9HsJzg6ICVFH1U1EyE1w
pNlZtDMgoVB/GFoyPyWJ/v+UArbJJdGbf1aC/ZrrT6PzVL5t6ghxuzctZDd6/glMlpw5qnIBabHI
FDYGeh9QcGZ/wqqWpd8iOHlrnaTQ7DFcsDFqUY5Xqe6OaBjalmv65Mqg2Cw77Od1qZ2b7RKyKzrE
7aleDMEy7BEXAYFi3o6L2lgoemK3lm7VTJk0Q1xi/n/5kzBQm3fezQW/mTFVSb9H8nMVPUaW9yZ/
wmdQq5VjQVPIypz3gTgbYm1M5NCouHhySFxmMtp0BPZ1MKmsCV+ymSyrZGPBaGLtBEzaqaOpkJo8
C4FcEkdzO4bW13r4i/SHBb7oeGw6gItOQQsaovpZO4sipOX6JTT7JzHJL8Vm8yt3k8bacniNwDkK
PKi4cRRmDbEzorZJ9yOqguIDJqiy3R+2L4ebWVcidb/y+TaEx5bAccnZnDuI4FLvB4+Tmu1A0y8f
J6HXxAkehnbPreA3AiihzLh/e48Ojyf0y7TOjL9Ebr0+q8FRhDzp5jXBloQ6XJr5/7P8o6dF1dDL
W+LbbWtPFhSRyqBx9nFoXaK1tCGElbqxQo9qYap3pb05zIz3i5IHobb6FwouU5o4YBclzCmJC5aF
u6s3/SvcnKrfBzTkDEWiW9TlNo313iesahbl+ycQnpWJqM9YpetyfaRlM2XF/r94Tc5QYNQgm5ug
zLKDWZY9SbogwakC568QGwGE/u1kj6DJQlIBGpj8ZQYJIKLwb4zBK219zlw/w3DhExwV0XelragE
Nunbr6VkVMt5N8iMlhwWa20sj54sproWk2s6Y/ADTieHlagFTamEtrahaRFtiZcJ/nZMCSqPbhs3
fMTL7SajBibcDo8C6Y7UjrI3Gf0gTATRwrtzgrtDJpemznJvTa9pln15CKSrqukVrvDvwKaVro6w
mHPN0ajMiPrXn0XsZJXk8WSKlfzajiVXAxJVi7j80LXCPCF58T4QaoCSlvhM9tjpcXsMNruM9szi
JZJiiCamB1hmT12kcnr0e74+DjK18TH9Cz3x98oUGDRewUONzHXJpuxLZNtU5cuIYP/CCd3xsPsM
yvAymMlHb9lgH+6xqaCJnfj5HORvXXdvHDKrt6IosZU2Hp2lo5/1kPc/656w06K62iSeMgHb6HXt
ZMpqene+mEwKjcaK0JfnP4Kl4sd0V2t5BicJC8k6QT1sn+Y3o8yZG249X0UvI4UFT+6QeJS3ynH5
CJOUiwjAtxtMGzO/4hMwxhiRh0M1jq/13qdRJEEo1xkir0Tk8wIy1RmvdPKRfyjpYuSvzb5Nrqmh
Aqs5wEv14u5NcJ/mwiuzmEZgV1yyxMKXhwanXvzjv9ExZxQASuLLTVNZUg2WgwqKPt+Anw39IWS/
eVgij+vQMX1wG8wj9Yn/L5dG0QZJ1n0Ld9uZPNsmNOEucHUvcMVUNLR+XIZPi7zuD9LgXeY5Q7Id
yaCP9+zvtcv4NpMkVwk4ym1S6kcI7au3s6Y+TZpRIIPhW/fcVywOKbSSdMe2VC2pE8ETq7xc2Y8g
g+2RO9JOPawQVlogE2pP4TPnw4HE2KhGlV+F5uZ4Td3j3Nmko5QFM9T9bA4aRGF5tZQRHSiw4u8g
oSqVLX0Tic61EMpd4rog5ayWYz3mDxdj+IyiGj0lyMKOYHaldQK5NsRAe3lfkk3IeYyGBBtbfaCl
/QSuUeUzkhVn0w9uhbkgkjb2TGGxLwnhkmKGmrDdr/1+56KJfVabmz8e4hhtMT7XMqn3f+cxCIty
6ASOnIvRAd3BpWu2d/picMAC9eyjC3D5GrGiK5PY+ZEbfKLiC/mogHRJmh4tcm/uhWAcCaNxS/Gz
xvlkFhiraAnVLMgFfE2MXgMJ3O7nAO3qANwMWTxU0Yhw+c7L4ooZsbKswPevfzr0RXZ9/fm7YScZ
czBmVY/rxY6iOZQ6y0O69qlPivVe17F/MRbxTWqQ16IfOO13Xe6rDgpHRm8NA5//nTiLLvHlroBa
sMVHbQcH1dmbhxSv085eKgvae/lp4FOT6FDxZDUAJAgl48L9kuwJAuzFdWGrG4L+L85gyFI7SHzJ
UOVaYFWMAINgBG8Y4p4yFQ12XOO8Qm6SyfFBaK4CkhcEHt9+NMxLbPjaF1kCJ0vcbOoBf/564qbn
II+XCK4D3rrEMNQDWIFN4ecDU6FU+slvZwKHOss8cRJLhCMle27r8+IVwmojrH+vLFIP+USn0TQ7
fUDtuzEJB2Sr/ydbxToLjWN2AZFSPlQzRRXO6qPIDj0dZJPLvC9hen2XlqwkMAu8fInI7Tl9nSfr
pnDf+GO6XhNq9LmJcSHif6vRPgAYzRMMvujWwfrFWlvWSSmvJ4tm61+S5DUh0uOwrgWLbvfFEg2f
kHAJWHcsuSCm1RDFq5RDf+0/uA5VYY6Y3z5Zsf3AWovMvnqgh0djaeA1unMcIIYdhtvezfJemuBp
0m0dSgvLUlQF08125sMJjN+MGdgsLZoG8alRbPS/WGBtzH9L+Qt6Y7oTZ4oLEwijEDpMWlq03Tzn
V5WGkFVcahLotFwPhkFH7TbXT+I8ZZqz5xYQkW3Ah2Swg+sIbI/nirZFsvSJu/OS807cIiF2ipzX
t/Pe/hYq2XL1Ia+mpuGv5wuSNjrbdsE+oQ4KD0dVFbY3o4PKrTcStYOs3M4BFRQdH8C4Ve+oWTQk
/BbOBPZfVSUajdJALF1VdDFR8n8DlTeEHkADkbv1A+HJDAyoJ4PQqHk8KpOmhvdnDoMBHP9pN6HO
vuIh0sTwA+ExUAND6c2kT5AoN6DNRSMw+v/acXzX06OCIw1dPAeC/vW2TjX8gIHPQk2x16+l73hh
MGKE0F3ChPyhbYGs0LfVk+lFVSOdKnAI/WYRpbffWAc7myRyP7H9e+2rn+Sk4DK5qouxFeJFhhyo
rapAn3ZvJbAubl9SBxIorPVdaLLtyZxITgAPoBEhkV6C5JrMdkMiIp77hii5zxwpQZPVUDuFpd6Q
jKivdc+jThXX273uloQk9VMbTi546eElrmWjuKzDD4UMl+uwD2zJaQIsrWafFZUS9gFfD0TppgWv
oBoSGMGFKnAXGlo9Ajmu2OIfsXrtVjKRg41CcxMmOZSu11NhAk6ngCHHNIVmlC1aOrFXN4o9QWE6
LDYjXNoe0aB+iBMIJGsh1/g/PC5EfpS9T7XJ5kiDZXEvvB4+tdpI/3rPJxn7aufiumZatgdD/+Ef
e+Ilkh23Nd/k4qyEtyGN60d/CsWYISVj80rKBQBqaG7K1XlP8xVS9QrGNOlDYvaMbYbfkGz1wRjk
mHaLdfJqGSMId1OmKJ2GW2BxngGR2vrWSehLBXBKo5dVhe8hi85qPE3i95FKIRCVGGruEnS/I1av
OrmXJ2ucf1aDuWQI4nELijrMwrVJ6/lfcDLZY/uVD8PT1qG7P2AoUWphVi+3GoMc7jK2rqc7x/l1
oJvUvKHWGyKx4y8wP93Ag3D7PMbLqRjl14ebERytmfwN2TQe+WvCIleXO1aN45ehoLUBIl822UUM
bW0OV2mL6PdDRgns8Dr7qVDXZRaeKWwmZV/HAEs/DgKv0YHA4K3nD8z73lEkQ9L8Qo/dU1F5eHX2
/MzrMyygK971GUKAaElQ793r6IJMNsG4GeMpndfm+/0O++maSkyr86zlivNvYpO0zGD4aA7643+a
pB/zwdh/Np3cE0p9YTMbzlw+pYx/If7+CHo886klRp2LRHrvFapJhuRRhcufwvOw1iNe2P/yPwA4
3Hr2AV1NbCRhLEhiXVewuQKvSq0a+qeBPb/xHj4eTt3DWqgc21oT/0hha7oZ6WrFLqvQg6B3eVhB
F+ImIA1sqkU9g36ZZ/INA2D7wSfsdMZJ7jTTTtVfi+MUYTXgFZIWXUS0s4Kz5Mw+VOFCK2frcCQ0
kxOQFmQV/JEV8qej9wv0QeMx6A11vU47Ndr1RpnXHl9JI6oJpMOk+Lr5U5Qa8TzwQEPqGsD82KSH
dnK4vyvgWvNzWBFxxsq6wgr85t2jfK+wxq6fYX+D8Mgpd9pT6M+LVhUaSvdFz6OUGdxvmoewaJO5
elLNUoJoicH7a1ZSLEytE2asKI8pIyqFi1+ITARMJindqyI/7BmEBYD8EKZrJClyJsFuZ4zTh3C0
UhzediBMZ2DbJ8cGKSWbzCLq9c4UWs24pQUuM7+CvLXEugV6og3mM9Pee3sn0P1A0wmTzeY6dmUN
mAS/FuXrJ5zs9HbtjV5JbDFy9s/Sc1/zxXrh4WMvQHbFusoijAV7OIJGWbq6j3Aq50zFqZoBzGGP
b55mApKR5RVxNViVTLHLRT40Pjyhs+WPSf9ZhHJlnV6MIK6SpWu20fCh7sm2CHSDSZicbyNK5MaJ
pW1ySWOICCJ1A1fdNLbJgKglP649xNLumz8ctpyAUdQsZgcX21eCKURJa1jCUy40AlfiE1/G6L8v
xwUIOiIlCcPzYY0uxR+uOGz+bNV1JjnJD4+FXlVBLZ9HDg4mP0vpV9CrVgbsBeO/DOreFZmgAheP
ENA9XJn4uKmKaKhMx8gtj0e/xice/V4NUvhBhWF3wZTXVXVSZmcIJvDI57LOcWvoKfgR35FeBr4I
pDInEud3I/oVS8vsW3JrZwdyAdRdziJAAArqvKvqFC6b3n76QiDMHdVk0qPPmeZC+EN65gmtsHfr
+/5mEwK93pILTPBLggEFRTYN5H1XVaxT0ZGsMH2oOEsQeoCvOuF5bd/0HGUTbagbo5/LONwbHw3c
YQ76VN2cvE1HV7auL4G30u9PYvYCv/5dMD0wfDVUJduTU0Mgtu5UfzxynICHao0WgsDx08hABPWj
jh05dhUaAM43Q/702tW/CADBHI7iTGbGhJkFvZrrisa0H3RD2blFs6livA1WfXAlKHk1MovjpOF4
gZP58QnDj+1FKuWrJnVMshuBnwqIIyGmNU9QExpYujreKH010E+a5S4+y5w15EQwPBF8NqH8JGKC
uj0XyKcei0QSQ0lu4pHePUBa/4E5qMBa4vz2MAth+vgmSYmgxTyOX/YyEwKqNqrrcvhMFmBP12Bg
Xf++8bp9j5qXLPDpSEG/G/XmFmVJ+74/AXYKzoWpauvnH3Tb5+1UQWPb3d85zCblKnZw+PXiDZ2Z
SqS9AsZxaz1LRkxXbcgMaoUKr9jWoqj5PzszSW8FltAziYy2G9Fam5uQynAa3Gn3Bvle0zxN/bEE
hEbyrZmrzifhnhn+MOk1KkNP8UHmQldekMech1CWjZmilrCRdpd1PAyfQ68eCO282pCm70jtOmnD
UmOOj8i2JxBvkKPsGDTGxT0rUeP9/Z0CqWzp7x6Kfp/GRRclrxuIo4sNTxVjXaj7GHYkGwUdHONf
4Tf88RcQCL1t6m6kymUeyZgecYDeP2Rq+5On7Vi4zh/2enBNiINFCe7zIb3Y2YUELELRNA3z+3gJ
MXKnTIQUuIxrX2vownIWqnATqT1PqzVSuMZ3zsneh7UMakh0qhJHD6OQxdC/GzI5AIUfFKW49nm+
tEu9qzZXCNqeJlIDU/5f8STl7Cu7bikANICE7tTwMCVp+w7nNPGBrSmLZiUqPWvttwSMLL6/JTIg
b2/l3yQeU9cR63cbUq849xOdYuH0qpYYM5XmA7//QQp2t/+Hk8FljOXe8pDSPRCIChiQF+qxRsGQ
D8sMQSA5rERF4W/a2TJD2Ca+x8hSwV4XghF6n9I8cJ2/upmZF0aY0yclsXeVH2lcKjc0cg+nzu1X
Qv6pW4kiFKKMQdf7OjszFnTzEMQBPr8b1Ho0m2u3vGyPThsi8qou4ElQzE15iPLudnIEQLX8Lx1O
qI27DS036fOk5Hgm3gOJiRSnLTgsDl6Qv/wtuDUsu/kNRdpc5045+hM+LgIlVMvGFmp4PaXIlTNU
4NqicOSy6Sx+uYlAALO87ciuVGa0XWczP43Y5fq2X6an+ktFzioHF/vUiE1p0jmO8COOp/c3PZch
a1bC9fJ+2DN4tU/YjFfLvs0M23nChRmHjqGCdF705aErkbXIpoOHHoCjK9klN6kEzKNrMkAw1Ky1
0+qI759ouOM4VP4O6w1xkAf7H+ZSyR54dVo+czOg28HVpROIRJGM6VyZVGUrysLRvJ51xZQdmmYa
EP64MTi17QwxAr428BibjEJjjo+QmJqHBaCOdH2vve6J9Uu1g7F0R74hRNsthlXoaidtqQ8oqEhd
/mlmwEWdHXwe7MMrWF+Vluqkxvq0D9JJIdyVh10jl8TvkZryzwMeW3+Fpdj1Mda5L8qOrSatLDx2
2kD72dIB+YMO/caMCPje8fNSr7G5KiyZdyzBZD1gJQAe+eCeLhOEL8AfhT1ufVnGIreUcjnQh9Mu
AzOaykod0s+aAj7wjsia0UZaxSMOukvWQrgNqlfI5i0R9zp+smaPcQQCrCnebFb1RyIY0yvz3pnh
vzSTy9VxMCi8nVN9OHohmG/9Yj07PZUvk5UBborU59He220uV81dalpQYku25UZRRE4gBZZmM5Dn
Gmq8uWLKgue7XdnI1k71GEirLjRAUEtUHwDBVF6oQR0AljUWt8OESEkp8CTukkup/pVBkiUcFdvc
8IdSiEjZokJVaeyMgQym+HEwIRSYTLE+h9ZW91sQDtDIuBuqeMszPE86flYvsfDuTgCAlMTuSPfB
lSdtRG8g/OiOeqODrla0GC1wGpbQ9PAhE9aziuHDQswJRx+9A92KYC1DGMYqHCHgpzHwj1DWQU1T
3M811NFb1uwtNcPWRfV9nr6SROXa4zay+O7hoB8svzef6GBm70MHmHz07Gy6XcLrmlxERkmT3te/
5cnJYfJDKBghlFc8myEA6zTAd5GzGyYuUBsZCrSwvjBMwSI+wxcaTDAY83rRjPqFjhRA9GPLvh9w
7Z+yi6+nfKG+q2AHPLFSHlLHuhioBvECKpOVBub7wiG8xpx0iT2FJgs8ii01SGXtMpIdrr18pmy9
979DWj3DF1lMP2CKOWOYYi4D1LzJwR2ry+R1IjpTfYWJS3dj8WGXI+HfN1kABJeLnYcxq1N5B2pY
ghANYhomsMl9jFx2p8QyfiVrUIMMiEMXutXq1mV2UcAU+1so2a2Uct1Jci7H0WeTBOQetX39exz+
/6LpP8HNkpZClV7lA9J4LLm8gKqYfX+S5crBQYMk2l2DlNU2DEjOZui8jhtt6WJBuyc2StzA1u9P
Svy1+ybkZsmTjnZM6y7hCGu2NLFH5bqCr+qxfSY251lxXUAAvuyW2+R9xulegZHJDmenvZANhclG
0KrbaEET2Hbjkqiv8mkkdBAUHhd3xpLE+Zede4MJAyJAobThequNg48eWKV2J/Oxkj5uklOmjS78
g7/XKFeTyStPKrQtfMUt310PWRj3h7YcmP0sHtkbL1uX67s2Um9Mh0TUKufg35z3oCA17S8rIbwA
zSe7Rvm1ganJ5HvJrbxSYRqIgS29U+i3Kt+mAGoOQUhMSx8ZGeP4L6UUpETJ89sfn+rXgaIXa2V3
98xswQfA2+DQ3w33eG3noC+JHD8IeJR/avjr9rPJuwWRcA9LXCeMaVWLngJJhkbOeSEs9omNQOJt
8jyCltmEo+Qlj/cqQ2P9kfTxOv65c1IPPBprWMYiukNLf6OR9ve7bv++tsdQtAG3sLSp2mEgt4+J
m/m9XjiG0e/8du91mr6eKYyWca/MBmm14ooNHq2NCd285V5w5OwgUlexNr0J1x+8VyMJsUYemXAO
yb7gFdasG8aWfT58vVBPPWb3UWJB4Sq3saDhoOJaDu3EesetjlojJT0p9Rgf0y2rS4PIX7R7z118
vdYMpoyCcu+fMiD8RYRZhQp2pwLMZaUVATEUBGKuxNz9+UmikNnF62wlmm61TsyyYT5q5OscQyKn
aWXjKxblw0uaA0zSNLiKF44sq+/RsW6Kg6UlzjxFSrcv7ey/dc+H7WQoROPrZCXdTPcZi7vuwqLA
P87VQSJc9vVpIH6MNxo4BpaViDpMMtTMDWxVQgS/j7LiuNqVCYseqysBse6Bie1MsT60UBOdoFLs
xMqJxtFC7+6W0r+iRB69izj7S4BnqRP7m5CRNvky+P2Y2yYvLigxiTYhLGx1aqdqV4ZUuzh8AEyt
hkDaSKCsEdNf1goUGFZ7TLFU3ECGT7DIqSwjeO7MYtstkd612MnO2dvlsI0NidKOLG/CB8uU1Pez
xulPTWrdYxOyCWq5ZGD1qpj98kFe173fHS2UpfYaV/+sjKhnkMGhq70bH6EM599YY8ziokWe1v5f
/atSfx+JOalQAyxYhfJwwH+fW/+q24XHnT94LWtdfOa8XH1xlRrykSMJihubYqkBkbtYTohM8So2
JXv4E4xjC2TCblU3XIQ/DjHn3D1Ix3rkuzlBEDKamYoT02FvGFzwSjZIOVkwP+ZgvbnPZYIGlOFo
Q53e2a3Y+0dbdRkMch+4sanb+B9Cb6nzY8WahDBWBOzarX49ilL2L9gp243AMgqQ2q7fwlMyiC5u
rgdrHx8Avp/sPRru3/EXSMfDd8KeSfEvu0jfbTQLWvvzk89OCAbKXtOWtYt4DQzyb7b95aZDIB8x
t9XPGaYf3Bcl/yrw986b9dUEy2CsO5vyw7u68wE6T0KjN+HGhwcHqGym960Jwp2CYFeDbSH/Xfl3
Eil0ldubQzeIPMgyNODmB2ce2mUeSpLsy3Jagoysn6j74XQsyWraPndoXXhtOLhJt8NKEiIsvykk
Wgb+UltjazP2z+gaqZXdclGhpPu2O8h7dnhn4qh++pigFsZODhBnXT8G02QUeqjqj5dx0sYPIFER
+g0e363B2uHBeNFGR6sqXsIBjAzC1M2MgVKLknWVKe8mGGXIIT3V5wFc1PGf2Bky791keoDTzP3T
OpDLPvcbcmbF7d44IuSuLjyyddRXzsQD1bQQbuOgq+/M+PW8Zf77ow1w50Ami0MlW0fFr2z+S/JK
WMsV6EacvAwkY4W2hlhfHxl0lSe66RFJSfQG8lh94F+uhbQN4+eYuqbNznHEyMyNKPjdn9waa+M/
CSOHwkG0ZKemXSlTxqfc+xmBv7DLtpyOrY9i0UD1p+qt6UB8xQGjkZoc1LVB9elw5aO+SLYyRFFg
Kt8MW9X71bfjhCl8/UAH7+oxNxeB4h6iR/KvWfiZeO4yk/ZtR/IaOBXixZcj5MrtEw1/OdzoM9R/
DhCo4IyHlSVU/DXQnNSOj2KmhbIiaIdgzjI9n2zMQCwTYg2LrC8qF6tGyHSXJE86qsvr7B7dO9sT
5bl1kAxwbtA0iP9cQ4Uvg/VDKWO1u5fU2Ue4KLer+YsNs7YcVX1XraPkbHc7zgPijToRMGvs5cp+
xtqY7Ri8CCeclwMovGwQwYQ3KoPqHwo6Wr+AIUUfUJsrQ8E/cAamHzwssvI12i32NKi29E/6V6GD
LyO7hQGNkSGW4NEaEWbtLoqC7EQcJTNhTxTw346ZJj5y/LX5aMioM+w9orUaXjTQILrz+vHIMzqT
91ZG16nntXS2GqFQCDQt5aqlGNV+mwLPoXzpuh+6mtensj5u6nWFEQYhLVF1MBGydWSAKz3kfRS7
6lognb3XmLILYWWKgyDbQcsaeGBA56wFi3z1NKqivPLZ1sYQ4Sk9S+2IMBuafD16Ov7sdTsp5073
GRppj0gn9IsS1C0SHJkR6enSj0YZoTtFiaDwSwycu2lHz1euMpELZIgkpd0QSr8doZSmkY/sKpqV
MtO3Vmo5xTNkPqvkKS8GBAOAuGW/cbpzFNl+sXordGQyAMqOQsKESPqt+2zgLcGrjUKblHrV/uAf
q4sErrRZIvYcu7AKCS31ggXL6v1ewYvVL/AAJ49imUT9WHRxowGU0FIZOxDKm/Y69vJQiHUWeO2n
1sWU5xx4hJInDSybIrtuqsmor8H54J7HJXMlGQ1liqTvd6BBoHYbH+N9dIcjcbXn1HxbJbh0w9l4
deHM4X3T7NJTyBguj7gxBCIYhot3XwzZF3uTLppHAit54hnSkalevoxcop8n494SDl6ITuwfNIZf
uS7DpQIRe8iNXreBMcxZS9VzVq1dha87yKXt7QYeynFXY/WRbRAr4NneUzkT0RoKuR7FwebFjDQh
I1RQbjQrsrxRfwlJCTW8HWvaSuxuOvOSAxG+alHfftVZQg9Z2LYdgmz8741E7jNvt7f9PpTEXLtV
cC2cgBYnyBEdn/uuSuQAsnVUQja6lvsY8d1BXUwmr+V0ox3sYRbilVfJ535mrF/uCMxj+2v+ZwrL
UrIo13QE9ZAhjPFnYabCarxDg79E1l4KSXPJhvp3Or0guxRXZ5dsePB7qw2W/tXO7al8g/t049y7
tGLe3k00OFulz8v2nUTyzPKc8dGfT8PwyIo6hnbBKmnpeCQflnHc6sHz08aRd0cP3HDDtNHnQV+k
d0CxS7RIWegr2/oyG7hb7Yc/7oqGC6whEsx7IbnDcAeKQ0X+tAaLnLha56NLRgksIg0iQ3kSTfK0
8xVhKzDsjefmSArGK05+voeN+Spf4w3+U5OPDm01y0l+faInjMH+TbyQBDO9gYWwm0Nbe5ZlYxVA
WlGdHBwXG8pB3CNOG1k0NA3ktyiDSeq2XpLVuafk0UvKQdNWHa84v2UGxLJg2t4zyeP//Jl4E7Rr
vpZ38pg0Wx8THi7ojKJ336ygmKTKbQBIuUCXtz4CFgfENaxa42aTRAWTXXo34idMlmb1qmmIwgzy
rOsS/dC9Fpn+YVf/vtdHWIFxDymNb1vXYiLfJL6Iq2XxOMxms2Xi8QZ/YkV70QPwZM2CTNc169p4
WY3wj70kDV/fvso0ojyaHx3bo2YVuo4lxbpCdJh9QC2bNBmb1mW7iFXgxAQ1XdJ4LOg0Tlyw2d4P
2xM7xGXoHcEwjoXXwDx29WMUr4uOepiD4f92NtLJFmX59/K21uTXtjUAjCeN0xCeY13SFZeagSWG
kao/jUSsaBB+tKiSDJHiJLrU9QVQ+1uFhAuJFUafx9cHvBLv4yRScOUBIAvKSt1y4b3dkDkoGHPi
FRbubxuJdZ6BFHgJw7F0elhmTLJk7VE4cpFlEsdYuh1Y39xEcY7ObosVfjddSop0hot31ValODFK
jHJIARSsvf3ue7lbAOgTalcU7c6/ksVR6vGgq+OTY6e7+2VT5yNKWK4/OYGHtvg7R2MXbvgaZFRP
VFUrJZZVyxeN/qy+RUu8XpgJwkWLM9GrDzmbm2EseAs7aAvJctL+UelHtZFyvZmMrFHrXFogCLjp
vrMsmGDDYced4lxykdCQCKinNvcMd2bDKjFkMptmGEDTCbs/HJm+bSPbU6XvPPffKwN5hBRgQF8+
OoKHQqAIfQsLVpZ48yKg0UVXYOLke93zfJX8b1doVP34HqXoQIvMYkVvhnQDp+xolnZHF/qzMKN2
cHRhqm5j4yczbNkeCvZqRXQ0OlyJ5SyjK3aKjhvUqMn+hmwaihEh7S2vtrxLvHc4sPJvPCYTIoIl
7J51ed/wtUkqTYaXgSD0TJA24nXrCxvT7ydX2G69D+aYWdjDjD41wo2r2GBhEfGd4KNijr7dFgaT
OyHe9f8dzTXm23UWev+qMrg3MBjGkTakmiBHgiy6u4CEbkuBEzzixklXzZlVBqFbcBYyCdFTeu1E
Ra8KOhOiVu5F12BCM1LsotFgN4xsC5jZVmikjZgmJIM+KGAaNHaAPscLcjHBtJxRV//9chBOVJa1
qorbe+j1aHjssciy2rLYf+fAJtv9e+U0BArbdzf+/SHC9vsR+ZiQ557iZ5rUzheYAJAQnv0oYRAy
ynBMx3u4BLPTOIqkJ9jZHQhPsM2gr7tmm4RdGphDlF2bkZBf0+F9CiYj6BxA4utWwzo+vieGIPjF
5ChFXPRgFEh+JQEIyVLO28BvvmZHFaDnMO+452wY3uQW4gkc7V3Zi+hISKo2Pk1h3j+31aer4oio
+4CgahcKrgAyFJe68ppuV9QAzz8SPiXLlVAxwlByJ7VhSmlO4l+J+VBUlFLt2tfChPAIXx7P8eIB
7gBHsJzCibHI3UbAhT3++K/zRxdylgegYskVPlgeMT/hB3FnABjwIXpMdOyVnG3pXQIcdGs3G0s0
sUS5vhsI+Bv2/1Jhh+K+26U74Z6xXMYjzVB/u7oJcX9ROmQ18I/F8LWb1XLsur0ke9bPZooQErbG
d6OJTHGovlJi49/LIIaUfF4Lz44mwQt+EfZDKg6/0CEmuXKObgJzg2ovvOg/yIZ/PEvgmJixAxXa
zMorUVR+h2tlbQXKCg2bSwqEH7fU07RZb/WT6KVt4xtnmjumK+uxSFclzAyqwWekh+Fh+RWuKhHs
SNGKSBS99V1gv7RYGf/yBtu7cgLRFHH9yDYeIvWbA5Gv9IoJ9dsQ0lZtLQA+bddW+2k9QHYo/ZZ7
OWrgcAtngtLOGTkBfLljEQfT6vNklpci3nNdXsTBQh1GrBJYK4Uo/tLYwGogOnfwFsGkal+ZV7k1
rXwSSw/5SBeAf6YE0/IVGuAwtqFQt8zwHu1bnayAQwBDk1vrKB2MrYWLOLvGQu9JSDz4IhyxHTWl
peoDwxNUyyY1DhVIC/PZgarF7/pzVtLI8rCSV9jpWshmq2Czzl027gdIzBBsTTG4j53PxPAPjXu6
elNCDFvOnkVny1LtgGxEPVIQViaHmPTuNG5wnJKFkmDqIb08CTNwWHfzXW9qsIgHdY5BZfLFhcG1
fQ9pfP2lB14nAvbMGrckX9xsEAxbWETtQ3ANpTu/W3Mf4tLbXCW5VVUi9JjaJLzNQz3OXC1yOSIw
bnkqhaUG3dyoGn0utsUYn3BXOvAIPALvt08nS3O7LyXRfligmW+jayRxeXCsjfMIeidP6lcMbzJI
qJg+M8K6DvK3j1ndmHO7kk92qTvHDB2khQmcWnm5NQtbnwWyVdA1p1IG0Q+UMjmzFpLbL2OO1ibm
/x6+HcFKRp2BRvpfNrwIaoh5BaiMXWzFg2AMSkrDqhcjUyR7SqUhhNHMBnfmNT9qp8CCspjw6vwX
Ji4NhMyXsNC3KAQ2DNTshupXOowg0JP0wUtRwN13W1fCYQK3GctNtLp9SlCsGvOWYkjwqx2pKzDx
4M+H5VjeXcpgYrKYA843uf4ooWNyaEA34hJPK/h83s2wGyHlKGJKLWtGCb3/l9cB1ubWF3FUYD3l
JohELxJ0AYbPnKMRptSw9ALnqlKv6ClrtLZ3nBNMLv57P40p+hbKQCrpCk5URR64uIfM1oeQgOGx
CVUnwBGS4pkb/Uewqpq24YboLJkcShtb6/v9ost8X3kf0OSYlRRIlnIICZ0J8jO0UbunBaKj6VPw
4Bizlk//4XXRgx7mbDrGCqpR8qFPymc/EPVEPBdGb5z19Js18IlgDVFO12c/vOjFZnBMoGyYc1sZ
/MQXivIpv3L4VS4b5H1W4XcY3YLQnrkrgNEBUsHknlLN0ZR+gG+wSiSlGDs3GWtkkw7YEmGKNUjV
zWuA33jbMAREwgzLIcIwuGSdvv3eKQNc4xH0ZkX6uvn6GKlcV1xl09Vr2//hQaVx3K24Wk4byApm
36gRbPAjy44Wgnusio0+L4CuRmWaI3gein14zxqHwqwGkXLnPkQ80b7y954cvFkWECmq/SUHy2m/
+t6jzmIojM08pYzxXzcGKet8z1sHbry7M6rAe2p2GjeI/ZSvJEwuM6Yc4FEn03VrohJSJYabugdG
BBd0DLzJnSxOykrtxxeteDwzo5eKOYOfq6RWBNlBLjkqb/JroZakd6EyM3Q/yiGrSfjvEZP+uVm9
YpKj5UEpZg9oo2njKSqP0NO61Cf9rcpiY4MddKpz7O1J2xWYnESOpB9ohtzZA21STeEMCsun52cY
Gl9LhGA+yGUdF+81zpmFgZoJnNFsh3tNZj73b40jgMFOeRtXw/q8XNA6yVA8aMujk1CUkrBZ3rUJ
NWQ9DJ8G/jXDVAyvcVyp0TgM+YmsD/+WO9sTkWvfh7IGcQ04l9yJg7J1ERja/yb5QM+Rlg0MLlVj
D6Cg9p7XDVYRIo4J2DvEDgl6P4xgspi/0f6jlIhjOHcrADxe78Le22xzAtgAysh7BNj+L0dWJ4eR
6URW/EgfaHbXdTo4DXEOCOpjyTYAqRrGw9Ludq8AOkXr/9futZJfweuwpZlVlC9DJ0jyo8SH4Lrf
WrVjpD4C57rZuBIunCr2TcW23Tlz/KFKe0zAgOkDV7tadHCRP5g9NXUoYk+sC2a1edlDeyRnqskT
cV6Ow3o+R2ldZhH55NoZdSiOtB7M6+Kq9gSW1rqf/p/sxTIx3wAdWPmyi6DJG+UfJG8cgI1OvtjM
xjhZ0CXbGpW7mV2elbFTxNETU88JT+iTB6ezvzk5kX+/tZn6tjFyzA/JdLyY51Yvxxhuq/AqaQrC
v4PxQvX6cU6kVLvmnLt+3WORfwIpGkjsEg5gFytGYH+Eb4Gmrw2+ByF+crOtc+Rr0hykVIa+DOhr
2P93m13SDbnhjW5v2qS7It14C4dd2p+FF2GPqpZSqKd1dh5S0aKlY8zOXE/7LqZJVibE09pj5UMf
vJFnJYUni1FdfnQlnwXUZyq2PObHqSJBIQBTRAKXUxTTURW7L77uBqWcdO3MufdG3RAO50cCDPaB
+dP7OFTXa/gHbDzA9l06GClh0XcZiUD97eYcuyXCri5x3RPXoR89lpTrDz7Jo1CCFtCfa9jiNLwa
Tw15+TIyVO4BvmEgd6XVEAt4G8wG4W6WSu0RV7KkuiEbqtbF930K1uMh/ZZ9LKmXjGWwZSSomTDP
bsWW7bU36dueiFAOX0syGC88jUJfm/CSGcKEUsqD10ul530939b3BYyAn4tcMlBjjakD0lCKbMCv
b6h4mRE9x65zDOCUvN5nRc6L8IfF7CboWqo+nUdnZm0m+pQbC9YcqTeLVk8+7GacfiNTPbtO5CjD
eDuqAX3gBw8mmMzXhTXwkXa6vdCSPxfrq9LnCs9NiaVHcsXiqvZhesWBQOPTEvXWdRot1oSxGB8c
7Qh91Vinr0t1Fk17WcvLUqaRTUQ5bgjw6U/qLWVKc5GpE7FtuPfRJItfcj049NwMJm9muEocoIaY
SUSvIgM+W5lZAOZ69PkeJzat0mELqcDp2NuqTCPHX1YkR+m0xFmulSEn1wWqIP2+cIPc8EyuW+7d
peI1XNtXGlsE/6kqHgNH4gcIbrb4pil/6kjww/mZMp1ininRcFA0kHFRehLqIPHBmaw/meEt/+Zi
W+g6ZddIUFfp/fat9UZWLrtJtr9NLtKe+h/jEIrjknVU8kSn7oTONrGeOXNjw8OCe8f4cQm8zYDm
i11TIMQc5Qu33uN6bfC4yHMLb+D7KoF6xMRgArOQzqQxEskVxo6VBvksAGfH/4sCwWBQCQKcSxke
4czfIm3LbtCO3/4u2rztHu8rJptbMqnGt1pejWuYR8O40ZF96ZDe97hVsXr42eKUNtVimJuJsF3k
+j2tNGEGQRlhO9bbS49pjEkkg3i3o+vT8yeQLadFm9aiU7uUZEHosBA/zPkV2m69boA0jO2ZxPAZ
UiY+Ont7HjHB6WpgW90814R9oSkPS5KcqL71keaUXsbk8VoQDdauM6L3jMGobjgKtMilhQcMW5rO
tz6ZhToUSM5iHscwJ3tbcYx6kveQbMuUwWacq+QFwzjzgebqwWu40Kjx7AUuQW9JYNnt2xPXpAdj
0vbLJLCpwG2tMAnxvUeUhFhr37odOQ5L0V01vObd0FgkMLVY94g5kz1UwsKCMcT6EtW+lywwq+jn
0by4vNlRvA1ER7ygnTqfClRdqHrBp2w8JnduMjHQumJVdaaI0+WchLFUdpE8cYaLV2HwO1t+77eP
kfbWsvrwXJulp9SGSqTmn70RUv6W7FgN2YBst7mphWoWJnseTWBYPiFGeYlUYf+vXF/4bgsl9vPa
ee7AGLLAXys0HdDDbB8cBAPpQhamL+2OQ8Sn0+y2+aR0zwIqkKkXn8IB/ajdx1JAvnXyk0LgSwhD
gmETpumYGHw32dN3rsksmjpqCVuIgN6gAkMwKj4NXL4juQB2V0+U9IhOS6jH/pxfvOoNMpKxthLh
hsfy5DLx4zTbubnfs+r2kx8oAn/LdvcvsC/mByqcdNC48ONAAs8FKQVCo5yezwBgVSckXucqPcub
U6VfOdkB5Fo9lXrq4GRxqk1tLMsjWZALxeZP/3X3VQ3sZvhCWaG3/ykMJTZd6JPj2PtFie2N6lYe
nVfVDRLdxaLThqSKpeBMu5yaYrksBBXDljknDVjaRA/Ut1dnYdUELGAGb6ecszwIGw0Kfoh7v3TZ
FnVrtH+ng5m+lM4iIjlZkbVeQTI8qYhypZB7VoK+H93OegDPsQc+QnBKrJ0dFygyh0tDVBfEKp1q
tRRn0ZJWz/j3zHWAZ8d0xjTs9XfothZubKLIi14gGqjWlt4xdZunGaaC6rbVS6u+yJyOePSqwNjE
PJAiQdCVRqSTdRHv71orpoEKPL+JfU11aoqVdGpQeHsvYUnlrfiu/P9+eFMVJBplyPqWQ6tDjJVT
bx3rLMagkUcTZF6mtZZjd5OheNxKHTQGAAbA3/C900HUAtYNjRtoIEiXJS4QHhTP5cZkr32RPFri
r97fNPkwTCOQbVic+j9ZScNJvmobtkjXoEn/dY067Bzk5zI+axIJMb4cGil5uk72ws4w7U41EdcH
+hbU9nyoVsYHUVtyS8Yv4Ehvs3vbtzj3nUoyF6GGZMQZCeiKkxjJef549cZKXSDyw+Hqg/32tFtC
S8sVstUIRrh2IzB5lHfOm4wlr7DdW0Mr7S7Uac3gwpwbQ5mB1t26j/ujLaYLNBkEwHruIoxC9EdE
HLIUKaBZ12ZtTF3IiUTUoREson4Wy0qBrF4X5PcJx1UNFEsyQoLVsAa/MaiVgNejM9P/59HFMQ/6
jTQtbe9St8xok4qrc5IlrWER+EaVNlGwrJWCTirH35tJYxGKFyrf89RIwsB2KTkyfHtXID3wuoba
mZxMgCneMDVN4ZoergjD1aE8Ss01W+IIc6fMOiCxwnuINIctipAxx0JmwaQF6f4uZs07t4NipyDO
5/ynzVFpZYH2kmoEjStp2zA62XecE6hhZPM+TChJ6qvoIbmNkxu/NO1Xlq+ys+kJCOl/jsqswaFG
EHeGAi/ETEMMrfmQh4QJPpDpGEQYzww8NyK8nCCYGXpaM8z/fYnm2LYAuEpuEYdJwpq4r1iARfsi
0cI2db9Mecp4vKc3r34M8BVt0yrH6ojjNvJhZJax+ICHh2UzfJXcOn/GjXtn7RLIjbYue4YrWLKB
rsrDa2iwIzaTZYnhI54yUcs+xmFISCuptBksCGLmpkx09W3GB/ClYx/JzKWI+LtVmnlPtzyUO2Mr
4sZ3dgwA18du9ZaCFXvJOydZ8R8AtGE75l0JyOuw2qVKwd1X9gxrcTkSaA6PnlxsPN+VnuJ2iU9E
I2cNrLXXXExySeg4soGywY9abr49xR6xw3Z51xG5bFqhDLj9vsjqjMnDX7XmNcPrnLNt8kmPcIDR
9W0C5pYKCV5i2KVTHELgTWY30oAhqdDDNYG5zOFd0CGMIWX4vWaqPNfFRhUVtT6Aa/Tc2r9KgsH0
lBOCh0TvvdZ2DrIlWwnSMERITNAcPcPMSu7GF8Z+0MRngLBRnTKePTcSFLIfpik0XXuv797VzAKM
vh2brqpLDi+D8fkmp4wCQbsq/nkqgooBJHfrQ3ywsC+TyIMjwvs3d9uboXJY+B6wOcxSwfHxS1Pi
iLfRf9KZdaxK4EPMS8vnAYBlZau8DhCT+5gdSVxVNwF3OYht8EfHwV7excSWFQBxaLHXtQ2ahCBp
ShI82ueq8q3v5boHPwqNPyYRpVNTroPojYYDuO58zJgrFQ0FhbAZCttpOlsShpTfa08tjwJ7rIFR
uOOORtJf1fR2A7IcjBDsXDf+hU8wmG/HJgtEmTcAZisze8mzYRHvsHljme5OflubQ9k1hGWz6dID
wzaUk4WYV+UngmmtYuUjgnejVnuAGX81o2JxHjTZNmYI1Sdq26ZCnefHGOfwgHUg3qlafS1jxoMM
ZZH4ycMf7ol6QiZwHKJIJpqemDRWWBk105BuqOWf24iuLzwPm3XhULWqtTPsN1yx+2ed8XVPK0bw
dsML9WbmFa1nF/ECYVdl8wiR5I0wpHgFqxCUHVra1Na3+UpbI/F8DcB28YWjolAvP8pTcYcoy7vm
snxzctMM/o0XCGbWemLxmjhHUPWDkne1+n+YWNW/oPL03VriM0EP+yGcQSGJu0uCciFXtUfPojH9
6dBzqmdtaHNKdsMzzGU2rAG6lu+TUuSNzd1REjV0Vk4blS2jAJXxbbB3ToQ8i3Kabc4iZEwIxU9l
yfm3/cgrJ2iiCMclQir3+aqjlYs27M4VS2XV2hRMH/7Xlrli6nZ8daOUpI5QCM9l0E6HnMjvSsE8
o2QIbqdJ5ReOsa7N8spBrY0OspIAKNUz1Q7StCD4yxnTPzg2BSergmYIBbqNE1umUgAq13xt8q4T
DuACp2LwxmJ8WNiWZm7y4G/n7Wb3wu8GZ164c/56nA5/VR50lQQuuVm+1RlL9Dwxj6k4sS2rX0Ep
NlvoBFOtU0CvbCvrw6MXAPefxy0zibJGyO/xm+R9rn0wNs1g723lUNCTTroUYfkKFbc8jaE5Kjju
jsd55+quaLRMwxjXReAeB3v8uyzw7j0WORabm+lAIe+UV+8D0ZDbEVz6XA3d0gyyjQChIoui2066
ZY9NF8yOB4BI07jt65bFvM+qkv6ohxtMggeGzUMFPbXbBDVvNTvxgzSsl6dDf2O9MUbI5H4pKRGz
CIm/eOmiSRSUTlqlcN48FsHANT3Q1ZLZi/KB3qmSAKqnDuHgu04atE4qcmf+2Duel5iPsz09zawQ
VUni3Mb2q2l4K+18zm3XbxEpmndpkXq7AXIBKE64Odf9IQOR3bCQnVAkpcjNBagq+8CZJSOHfOes
SXvCyN/+WTGCYbxtHN2zkAmVmS/x1/AECcuRojFTShax2Cw2KZ6QmtBZEpEKv5dr5OxquTJSZC4U
3eKcpAFKfY2THOHhWdZduc1uaXX4MvNP5rkDU79ExN2CNWx9YsdLmYBXp7HMczW9ZwfiDt3XtMnu
I+sBdm9cI0IlQLRs0tNFPZzQhPCwT8xGTpq0LrK2ClW8MNkTk2qq/DsZoJtl4HPwYUKaOAwz4p2b
A1WwejPw5efK7RhN1UaJFZlbXOwMgGUBDEPym2bIbc91ODtCk44yp339TS8sC12WePCbm/ZDpt/S
tN+IhsiFICzSQt6Q0yrqGYZlPm5vtdA9Y0/S9tuTqDXSM2OGcsK5zvvPbv+bDa8PL7J7foTjLNMA
G1zBFFTNOv8bcyJQ4J11VuSeumaVbu6bIYrjXLd/xKWjoJ1yCQUgnnOTd9EKeSkiSJTv7rMo7xoh
0vjgPzZwIlyoANWY/BLZ1gxBGdXpWxtDHBXkgY5b3/JNQv5JQBW2X7EI782jwjgsmwy4Whn09Zcf
M0KWzZqmaczuTXPWfu8aZGyK0XASQM2EkW6LRcCrC1WagQGJWXURw3vxw41n4mkFqIKCewr8OU3U
ileSxRzURb0kuT9ssOcPxqXqwxikv+eY0/lkfpnCBr1PNjcH7R67FPSXVJZgtm9s9SIYoy6ZKH1k
9RAGwYChOJkloUPeZtX7G6kvf4pG0INShrGqCNhYQmA48IJb8CJtYn8veRLSFYnVnydVJ1jZLWEe
TEGgf1rY8vuaYe8gRrrGddpikAfQkxWKhQ5lvVuzKh0dUN2LhYNa4IthWGMkUOFoNLvH9sqcZmze
rmH+xhZ7VbKlf8GayBdtpKKRy3tKttDWlQ9uPJSd7L8SeacYCU9bChu7qa8ZjQbDww/1ifdIi7nd
puJLmglwGwSgeJLKrbLnZi+xo8HwFno6McFoYJxHAmsT1Ztf/KAb5ekktAqC93wX3NnSFhhPKtE9
lcIyZLewWaG/VvEj+ACByCWE6wpArii2nGG83vSbhBXBF7jHLk0vJA0C/1l4PLRrI3cmWOInBgF4
oJVwxqrb3izxkzap5oqyr8Xuz2MoX5q1SjIJNBlI7OQcvuQfet5h/1WODrRPKQIVCLgxAjr4gujf
9vGT/baK3UnnJEg5hHEFHhc+v/BXso2NNmESFbKn3dbJKkZchMVvN7JnTgoN3d0PgN9kvSnZW9qe
ZG5HkjPfdbv0SG2NDOXz4huMc4TsTeQJVYAs292xpdeyyCQGiV/aRKqm5/sJoN7ulhP0VP2Ho5dj
Lvpd7lrd0lVoogfCos5Qv+wXe+WWX/xZfZ3/ztfGzfBxDhP5xo7E3AVvoUW5UyNzcJdCw0FW1iJ2
AyxTd63YJFoeZHKlOutj5ph8X7azK2BA/RHH6nby+zU7ParwQR+7bqbrOkNsIWJ+htldAPZxoaZF
2QTIXwkBIInQr2D1QYa8IWZLvikg1QbJsEFRaI1topoF8erA8NTa6jPH5iHn8MR4xwhhhab5Ttqy
udlEXls+70V9F2rMXOdBZegthBJeeqqXllz3GUR0geHF6S2Gg05QM/nUxlLCXANfwpKGhg7Dg8T0
E9HIFbZVOliNM884C/BsbzbZinWBV+eXQqcGtnQrKHYA0FU/K8InPPa8PYXJtaisJHBdW8t2kEIm
3E8zKERVrV9KLh576RkxQcdtQwe5s47q+6e2+ZxqwprtTu8/hVJ7JP8s+2uyNcLAFZhXmEGJ+8jX
CfzeYbYMnUmtZ/cydcXoIqLVFLvSt6zoDrCou+SKNg6IOC3UHgKAcn5dTYIfcdqznP0PtBMc5Qgw
JFzzMBPsxtx/D1KdnClZB+UUuYME2vk88nK7JMJkRjoUYgjrMz+HZfBxcbuN8NI9f5MUJR1IAX9/
1IiGdc/QQePQlKk+qZl9VymiMWwuL2f/Fh3hTvaWhKiLZJmrbV9RUrU4TAl/GxW7+yzViJBgLXMs
+54GYN+sS1XZrOHgoi5VF48ex8u8rQVeXctfn9ZLdEf3H4/IvEY/MSRUt/IcR8U6HH3m06jDOjg6
1mL6iaq4rmEvNTUo9dnApV+z60YitBMMNAiCG4pyBrzoFD+osZCBLVgGr3oOw3dPjZ5crH8EVAUA
4EwqceCUAl455gfIA3Pm7GPQys2CTrsKswxqIm8Wqi8xq9uMjUjShZ/4YqLoQuS+Zt/cusn7D1GO
m9/TuYKH0ZaiyZsm5kAz9bKwj0iv9AEzHzRJ40E0PmjQ59+dFF/kmmfdEkzoXNA6e7nNii0NEexn
zRETacQ0P4O3CTW4rG4fwxVzyk5+hv6j88ArsjipSHq5twlZlLNSEPosBgshg1FlRqqxVG0d8+rT
QlX/karoq/BVKqekHlLE9HOlNkAC6g8ynkhBxA3GLrIMDZjKcLn+DDpNdSXzycZ3Km0b8l8bJLMl
uHobeqiWSF/XVuozXuY7P9GZozUg4BcqqFo06wr5mAM0SbttJnu77fgl8IZKt5Izf5iUPWjvBLwa
TR/kuO3cYjA7TtfRYt9TobRQN4vz9aoyrHZS2mZHYWqPWfwka7Wqv2f7mDAFqhMPdc80VD0ahM95
I0pF0TFBYZTfpj3DNqWrPytsYTziJ+UgPBN8tJ67MXysMg5KSMvLPJIUykvQzuW0ZI1xxCZ19wk3
4cDFh1IV5DaxOFRD/zc3bTeneEjCHjokeTd7xUgUVbpguKC3cET0TD7b7RnWdDLX/JUGmm8i4kf8
omeztqp4W7mYJYMroODOK/C4labU0TOVp3HBapNysawNmPuB/E6/NtWpXji2v4earqAFksO66rEp
tRYLnSs5k07obIRfu52U0HXmO65SONBqqqaSTZsnXnCI3d3Wj3kTrnsWsnx1eIj+BonkZUxaXhC7
Sr+Syw7vOWy4rptnXMit2UVSrLvMzF8+NoSSpph5hZ22/CIr8NdsToB0w8AWfyc031NtLkr1XVyu
u5HzaHX78HRs842e8319imfdeh86TOQGkfud2zrl9uDtWrLfq2g71okbMHff2vLpplfpHHT9agPq
TwEYeyQUcAp1VZYLIGMudiAKexElLieCycHYdtsqoflp/rlZQutoF6ef3WN3A4TlwNiBq8mh9Mvq
A+Hc3TZ6gH32tk6lLOEOieHx6D6D6sJEzWrslln2WjmRn+84EK0Og83fI1+OR3dqrQt40qNyDRRB
9qxvdaemXRCxbc9KMDK3JKo6hHKDu3nbKqVYGCz3lm/LTWOc5XmZVqdTDRtRzMaNSmlrJqbhDR0r
ReSQxYk96i2Kpkp/bQumkpPy1EsyfjHECV27lcGpKILqIdXQTYgOuzDNfI6A9HxjV8eLf/dwrdAo
gSDTG6a0zJkuJ5PdMcoSdBJasm6pVIGV1Dns+tUIsg8BQSaXUXmdgzRxSZwWkjkZn+rvsjEg0s5L
nereAn2wg2bE6y5iEDiWTkibX7YU+tlkgTu8YiVbgrR4ssjrc1PQdRFBqa1L1uAiT7IS4Aojt54V
7AFuGVL/LM8WR7O9aay8S+ds8f3hSbL17QFouwWXgHo/JK4Yq/WMIIB32bLE7eKJ1hDACfn6zd9S
JXPcvfeCcvZri5tu0aMKHUIo8M+5ANTE0kMJATtFcMma/ReSSFKBjvsKoP1CsrDwsFU7hrsaoHtt
jW60rD03kBObHT+GKAOmteYOEWJMDDn879QyzfqhwUwGECVUoujNVigCg9YtwcSzdfWXqNccsQzf
HBHeK7ot8Vo1sHZpz4yRTXx9gT8Q+u5QN/8pbS3m3/hf8BCNkRAG3cx337z3jm3QU2nWR//LVfpK
luJl04+U+Fq3or7/ssIPDv+BFAA1TpP1mdfReX0FQZ+7cOCeEW/MIFvz49sscL9BjvNBLLDprcI9
Z2SP55U1N5tl5SB6MaUDbGrYKxVgvzGa2Y5NPOHQgubMesJybWGEKwyWJbwyNJxpbz3Nc+on8Akb
o8ezOSu81OoeSQAEP7zBvUq1mkgNpjtPoSJsXmzBwkslF4LYTgxqFZZp0SqleirqDSd/KbyS9iAK
YOL3ORtDVsjV3hyK91watMhqqoTaK4HQZ5dQn76ObA44UnlBJj6X/RmxfoNGVh+IIrMPjQq8TtxH
S5PQDD4JEqUEMWd4Q11hc+4QG9j5D69Zmwo3SETZgrAY3S4qNr5eEePIDOGD6KcdwBk7JgEmXXmA
7S6NlsumoQgVn2baROklZwtu7CtauOqsfmZ6TsPm0mScGBuMZ0LEhCxHRuG/YKCXAbYA+Yvh6/VD
LR8M7SkRCFymKda9g/YNOGXeiSlvHifjJnRBrg8pxd3oMOl9SPbUE+S8Yvipb8VmKVTElCOc/26l
bpp06gdZwuKXd23OyxBp7MYQ/TiUb9jsEPXqgI/G62UIVQmRxOjyrcmPSfaWI7x9rVemv2HmjzxU
p7G3ZLNyA/kLo2ftEtVlkCbUHL+sntBcXg0hbxHbG3Wo2gDvBRKDYzZ9+kn/8v9SrxbdHKw3uA+p
d/4H6PObVeEmlwHvnY32CbzFi543hGxUr9qNS5GzsIrOlVCNd/avj/78XBZBfL7/ggR2AOQoqMNH
n99+ojBIzR9fdBn3EyHYyNfEf3I386MwWe/UbkLEd+f/3zmgM70k00Fu7hsRnEWv+bZNGfKTQ9Ao
WXnRmJ46fbjyVBsJYecArDWkHbPL0/zO5ZaLXq5DsLJzzTXZuI/AraYBy4wH0hzPI7aMPLiergy2
gCr+SQ/iPX70bV6Ta9ekTfkt1ck85HXv1mFXxDLu5siJfjjHDWCbDRBz1AvhLzBElg2/brtNrmRg
8lo73yY1VCzQ47aEnbkL5efXKl7yj+bZmw3KAWHw4xgekI3sz7Ybtqa09PKBD9VkWiCQZ9TPS7uO
OmWjhH/bfE73co/WRjXL53AWuh1Z69t3FbVFwcXVzxD1N59JuluFjjA3RnAE9zH9Cv1+21rHOcs2
6h1RRukCVb2ZMDh8UjqhxdU7LA9fOSKmRWlj6USfS+9nah/hrg7eptoRsnh3oFApugYa5nGEUf00
vDa8QxxDmvhRDxrmm5vsJNm/OFXVufdUgHl1KxkXzj/6trlWg0W2gk3BKc5FxSiZ1raPwGFHDfNm
IIvkSSR9iudrKBmpuRZPXKNXygX6hiFoizb0qmh/zJGDDTPJofhVy61eACeaAgklB/6pj7id2Z1W
m5CPdPAreR41ewEYRNP3gsPsGMJ/mQx3NBb4Pu0hu/MVfjzOMBOAtYT3fh+y1sFfm6in2KIhFsTc
vD30VDr6xm8W12iVc7jYREgxM2dKB3Fx4IxNNfgPYatdOtyCsWMNzpWqW0ovch8AG3A9sqie/P7c
W2P0WkgUOV6nGnqDxFZir+P2p02bDqeJIse/sv8/F4jWUwyHuFDRIa7t6SwXUw8v9MX70WLOWwfk
BC0Uxe/57sHM2UvSlOR0cmoYdx56CcPMio6S1TZPA8syzhz90qsSbAQ4lNEf34JXFl89GpbDSb9v
JLfOGFlAchuAiZZlRo6xxUHmENoWW3aALBHBIK84U2NwfpxZxp3wTwE1+iu5KeOIAMT6zewb5+iU
xl3Dc+FpSFOQq9LMpPP0uwnE4QWluzVhukEAlrRr0heJoEbAQuDIRNmixBXO1sNv7dQhgdU/bTZC
25BC7/ftH+IAZjTaVUuOBtMJ3jTzds9zwEFiG/shHeDPfz4TLRFPQbm1+562OqFimjYg/8OK/eq/
47beDo2JGD1Y8NmFndejGEwh/wBTKp1/g1jYa4OEjNedeQgQpbFKEGFH9MMWrLIH29dVSIS2NG9y
sMyNvoSnPgrSqV/dkI2MKdFFQzJa7EwQob9BOHeIn8E9xrL0xr4p2VyZduNQW3Dk1AfbCvUHvjxD
4Mv0YJmN0WXwVI2OscxyekFm7dtd0/8lXu7JP3Uya04xeCY7hqFX24usrdDkMTD7ntJhxX8qp8JH
sca4LRaCTqftoFovA+qSnXxBf8nDnJxfI0k7YIHqw3zclmSVHyiBmbfQ1yoqOtNxaFUqTn+0YIDT
pehk+2/r6w5PC4d14GU10QZ6WeZnD8gqPrJZUeXa20xx+xDb+tj707uiagG6uZ4AVqlVx8Qei/Q6
q8raEpvQzjiCKb+3i9ij15wJ33tXjojLkrwynRYoLA2q35HYYi4aKNLaQ6WwTLdxyfgO/SbX0n7N
7DvuZ+JXvyiuJWqSWYdIxvYFHMbK0IDp36YCJh+Z+AIUJr4yotL5DOXhlAbU/UwDMDzZl+hQmih8
x/eUeTkD0g5iwj1gCa/tRb8zJ1qxf7VgHWkxjhhGKn3YE8PVHLU0oxY7l+mxm62WCvmznnzMGalS
NJzOUiT9nkjfziLaZf5+GQU3RXrTKHkU5ZllWCeG0CXQtXWaEoQSNyTYsgZpwvYVctsuIor5uSe9
4l9Hbyzvav9U3lWsND75kcyBvXWhYSP7KqdsRZwiJX/ZPtcsnbYZGAydzKSQSJ39A1xVJEQHuxYo
CjXumiMmcFjCrHpGkwZpCZpN/vyqE9HIAn21NB7WfLWGHKsQZa/a7RvBef1efPJWMGix78WE45ne
jZcXiDfsjhAaYKBIgNxMu77ROgXYsZbxWHMEnM9kUbxveqShS6Uj2gAVzDC6Gv/uN2+LwbO+xpda
vLAwAlyWLdDlkaPpVBgmQaofxDDInHKflqKi+h5FxvQBJWN9btuGeZS+Qj0LUwyyiwOygx5L17kZ
hWdRF/Gq9NLuRq9iiEJ6ALxLfOSV4mS5BTT0fvFWESpSOuW+XaWCNfYXj+JkFfDCtuookZN/Xcaz
cWoaEzACe0ZbNtNY2rxrEiqbUfXJOW2Xfl+NYRnh9BoW5GRxMsQrsxJdHbspLRl2/tIEr+Uy9GiC
3dxPEv7iIxEt530EPwilN9NNFQBtQ1ozwC7zcP3UxLK1vu8R8AN3/itLZAwjjK/ZrneuXUJ6pVc3
nrTVIDW3LCx2PwYFhHVKLeaS3fL7mR8I0tLYGvTHaXIZUk015cCq9zIWwxozN5jaW7DaZ4TCrxj3
BbNyRoWMmIonZKEOE5NKZcp8KTvNIyuqwT4S1uoKAycWmmC8dUrE1xlelIPRxLvt7vVnBypyu1Mj
uIRsQg/e2h2cXrVmEW1WW0RGtHaBqGw779oc1zOK/A6U6y0j7Z5qVlWmVnIoDh4IGIEGDyHXm3eN
18Er4z8ZhzaHiihfcILaaTorJZR5XrVY1hOOVNMFrdK6+zhcK8qkGrTTpY6zmcsxM4QKMgFnNN4v
BatgJyhkt0XHhm0djd1wakVneCeSqbAyVCbAwDQc0S8RzPVbA+VTv8hrYPlWGMip+vAaFr7hd572
wHb9XVxCDx5dRFmeT5drOcKz1PRyWAaIkLo+mAG0C87f5lA4EeT1nTEy4mHLpie/PF8WSyhw/ndz
Z1CB5CBFRrNJk3M9fJuDZ1D3peLZfqlg5DnlpC+U7G18MSpcUcgDrZiRgxobI1BwslaidDbt0Dae
NkT17RzO3M4EcQfyjEwQa8h4cnFPcy0ZR7ErsBEI7H029aPVzTWWmbOvkXVX2FrUrdTr0je3ssyG
qmSlT8oYauidz04+YKPEoRtgA5yKO/k0/ZirkLMpwDibuC4KODrEE7VyLBZG9RKfsjbHz53N+fHa
ozHJ1WvWxw76O3MaDAfvfL4l6pK5N3BrTeFkWCFNRK2+R2/K0wXAXDDHWhLC6Wvx8gQ+3LeMsI8Z
ML4LHiSQLTjFPyqUgdk7FvJXr+BVGqaX4yPTmaqRBXTQpLykweJ/AGNPUfn7EEwR8XsLBIjd1il0
rj53ky9MXcaoRyb4ZNxlmGdCYLElRQVtCVMEBdIkTuUGk0gUJEgI8CfKw6cE8aGm3zOOGU8fpicU
V+idVCNJ0PyHBJW5LBoY/YJZGHMWdfdtJWZorNAjMHSHx4ZSqNddckUAUyP+Cu6qhYLcOJLqTx3S
XdUyz0m/GYn9DwFGUs/FuGgBzCoVHqBYyjYCgptnkGObsXnDF325Q8NQEVC1SEMTNO30XGp3QNhO
Fa8BvlAkE5dqv4inNP4cn436MXF0zHZInc3Z0LTMu3U0hnQmuU247r2K0/DKsjrNJPEs9Jl/prLW
UZKUARXTNLAbIQd6VrjMZ5bigXJfoCOVVyOBCJ7zxI5qunwWbUPWnIZcPYm78E4MN7MaMQqnVFyD
3xEunEZwLUaUYOD30kLzy1UbEh0UMQ+Ur4/MjtY2Fxa0qGjERL7soUHftBW/mnGd1S3igad0Uw29
fuuLuS/POHXVA3j8ua3L1kJFNb5VEQy+T7kkOzJxw1V1U1k2+UyHAhETDPtfZSPTuR7iTkx7rrFg
if4K+QLCv/Of+QP3ju4ECgSL9J41NuvqwTtfviRQeV2Hx9qmbKVMZBAmh1LpnNO7/+bfs5BrZb4P
YnYVd4Ar52o1kBu3W51xfKoOAvkMfcItOw36c5PlAPOwoQHtYJYDFCTsVe2TFAGUQNmj7+jiosiS
+atd1NoK+3iUN989GvGJDrjxzI6/P5W+LI/2migmB/63QgC2ZUej1fAKCWjm5BKX2DhvY6Aj1HJl
t/Hm0ebzwEsdweqs7gFvktpoEOD/BkcAPBStqppOmJdRFkFrbHAR9tlLYwFtW5rrnU4zM2DLPu1j
lIbeJOE672wIxH3/NVls4KmAJ8UseTeWhaK1EzepU8AWiLA3PZQqVpNM5y+D4MOD1bW812GUZIF5
rqCJdZaDq/9uVijCpZ6bHzrlrrr0A1Ddm11T/4lN5/0rXw5xK0gNM02mMpEGbsc9rB0o3nEOfhUg
dfWyc3Yra709njwJLKmKC2ObuV/nEqDRAw10Zmz1+Twc+iqz5ZMYg/vNrRZx6xjwEjYxhk0JrauJ
hcdL0FdWRj3bdJAEURZAN2YuchT4dbRcol+1hZf1GlhJdUDZqv72pxkziRZAugDHEDzW93ZtHsH7
65rGK0KdTsqpJsM+vz0vpO5/LNpoT04Q7ExcrIjzfyzGlILZT29CZckS/VGEinDiyU0HMO0bYWJB
KdPTNNVUC2j2bePkHEamZ1h0kwyCG0c7cMB+/Xa1/4Icwl45bvc3R53pCBgzvIwy1PQ4oK6H4DWE
QQYMb/ZHj/lEwXhaEeIboMPBV7TmL/VxC9om+mv750EhCYZZIqq/kEiXZ7s1hJKNWpOrPPRuoX/M
NbVgOJkhXaYSDJdGlohSHvSvu2MqedDYDFu0reWYAj6swj45Dp2qvX69exbMlPEGe5IyhG3A+mAr
vuMRN94xSPMy+xqOCI/Wp7QiLmQQO4REC/NwQfV872TBmg1a+qpQs2M5PDhR9OkifbCkRQxvQMn3
qDLRnZsJEnNq3+TBbwM41om2BhwnvQKWaCw5GPTgxmNdRruLJ6lL3jA4byt2tjj+aHxZLDopvQ+1
DxN7UDWAQ69xpsDJ4GDIU8dD4gQ816ejtmWGrxBbss+XuGibTFDMeGjicYZdGDYR8YUZhnrzH7hv
aBcKOej50z7XbCFkbYUyUsDTpjj0xTuCZTWVsPUN7a7m2LoObdgijX4Oo8XUKT9/njxHFt2xXaCY
uE/ItOb1bFHWahTQbMRsbhltELEHzZwVoGqYQnyxp4uRNrBdML7qVqcPP43t0qcq74Jo7l7Lr+1/
RT9a4u0Gy/8SWspVSQMZhji/1UNrC6DCkqMzd0y2avaIqrogFa9o+yrQ7Gqr6S1lG1AhDiVQAhXm
LN4gMYMgM/o8VuOg04PYNQWuMVeblOgUK2UjLfnoYhSCCKG3FuTd/U/CRa5pi4Pn2CrC+DPwnC5U
xYf8DCbc3k+1eBI7vWxLTasErE+mMf9sJ261DDliT9ML47cD0jcDnYpzHGiQK5XiAsK74mg7stb5
zDKG5Ma27M1O/T0PK2jUHUuVIW+CQdE4RLKnZKdWJDuSRd8x+W+N70LVvvns8GDtd6t+HyxMBm1u
Y75iNW5YPMf2/ODbe3RKsNBaX16MxTap4ga3vWDfvrN5GFnAy0I51tG1Yi0/S83HFjxeVVJJUdCm
2KjWQnwOt5Bo4x1Nkcdr9tUBeF5GDJblRVoLFwTEdp5sfNhOjdO+ntA7sFYfbjZXyj3AqaC8zjsM
G86Wque3k0twH1id+dzs+980UtCiCe1pwhbo2pBszluR4uc5SFxzJ1H6pplTXHhcxd7VriOdvGzI
WAJOmlj1b+BM8wavBjw1PBMCKFwm2I8elunFkTNpQqkXZTqxCIwJgPhvYnv4HFl9t7rDbx4FVkgW
+BCgl39QKLAaMbiGoAVdnBMYpMcBirngnQNl7O6mSdPIxJ6H+teFwBPE5809sfS7bb1V6L6HJ+4u
kOW4BKOhKZIG1S9qub7207sV8YHkSp4eMba9YkFj9b1xsuzQhi2IqwVjWhiHlaZZFPIQiaGezBN9
BS2T1nT17Vvia3KWB4zp3eQJplpjSsfXdRd/9grSF6NoOUCbjY2/rCIbGOndj8qhZIZfPBpb+fGN
Dq6hUHHGGU4DXzxD0YyShr2xu8T11VuBQI7+5d44IsuMZiuEXkmetSVVqiEWw7wWtYJr+4Brcog9
WfNqxLk8M7rEJLNZ8NzdJokx5VTFeMrcX9VOV9AoCX7VhZSx89maAH66RywrJ2Vqqe+mi8eqkp/5
HvcAv6oncZnELpNAwFosrT9mq19/dPZscG+v3QotjDjitUJbFJ2OeIEkwRQyfLPEmIhSj5i59HZU
yJiJgbigZ0dOrcPH8qGlbsyBezONUhwtJOS7m+Mg1ZD2XnXPhaxTzVu2rX+SxwnTzmSrgtLZEa+A
DAcLEFYVWAfEv7+CzzkR4K9HIwJI9T4EFSqPqlbl3moFA5Metc/vKs83yQF4etZQ1Jtbrfv+6nNY
sRneL86lV8LOIISx/bPdHs74Ub/UuZgE0bI0KMqDPEeUbsjKgZP9lSD7NLsblF2M70ScdcX3Pv9U
jkW/q/Van/g43W5oa3vSfK5VaQ9R81fpT8FZgrVbCuI4in+PQL0j5veBLvXERTyFwS2rIjBYDAfW
6hxuGPKGwrIbO3RCVW/VPUlM/LCPqf3eJU5O7hmnrySncmovuCuhX68gMtJ2h2PUD/gNwch5aVCz
KVO/FEAFnDm1t7sc+jCOB4qfV2mYtuTDyERMfGjky6R0z/3IAVyVcFCgIUItyKdTasq7hbVENjx4
gnEPT/vihOkcc+Z/1jfyYkBls7QdnesWZJqYabzqLzA6z8uGVgswQmHZ4MdaDaMC7B2lB+ai7T6j
Y46LsoX5jQkFcIvrv4Gg/yIcAlcecDb9hPNTTjx6UUiDH1VeDmTxXtYadR9PJkoBk6XzH+hlEN15
J9RokJP4yjzNtQMw8dHs8rBZM4yyr4o/Ma425cy2/x3jLeoBKzHG8tcQXuz4RV+KsHbw1t9P4Xj1
mlSpXi0XLtkt51MZfYAZUOKaz471rPFyMM5KhSRRu/NbzTIJ/tNsvsEwJ0KiCJpQVOj4IWmj1v1X
1gA3w9qT6pzRVsJZpUl5+43TDIJb6pKTTT96vXD4V78tofdEmUS2cQuXX68gkt9KAOpo5ZRtpT7M
uHmzz4spwfKVCNCbZXqDBUskbZVqAAotlI1Dwl9s4/XJ7Hx3KdrWpbvcgt+8PsNYTa2Nv6zlifle
ndiTTsnClGQs+EpFyLVQYmMx4/0hfccBaJjBLTkzCgnkx+BOjeM8bfwvANi5/ZONyQ1ID9V0iZzX
qkt5j4q8X6lW/lhQNagUrjbd0qVkfZLmgpDuD/4+AtMYnu82buf8M38iWsWmjzPU4JsNXgYO/R+E
m7aS/7oT+sE2Xc9B8Z5PsFTUCayOKUPWsW4xdcn8yva7YyMFo52u5wyIY5jjBRiBndWlWfLTpNzg
g1lAuJeGOS+ffUT8DNrY+VdPn77dsiUGhrKT7n88CODpSzPAbENA9edHxOFpVS1fi4Z987lZ32a1
9s7p+3ufBQ4gZkehTrhoa09pgQofWIMjLrDdBLsVjRrpF7qjfAm1i5EiBS024aih6aZmUTXPJn2C
HggPgJeJRQm0q37ALDvYHAbP7BjY36AeKIcTYDq16YqoCeQUGZ70PGUNmYnqzap639ATaW2dHUId
aDzDyj34Sdun2vOrSoq6/PTii90lENG37Ht44EEh2KzLH0PaZgCXeVhuhytcsIZ11hRVCECBRES1
nlu/3vc7jx7t0shVFwRR7sHd5JLqIV0RD1QxLXl95edRi0qurrNUhnOwZx8gT8a1sI7BhNRz8Zf3
JcRr4hkMzp8L5dJJGCrUZvfI7gi/ehFGXrTX4ZbZbWoj17VrkZr/YCroWO8/HkYuVK34gCObMVUO
OWQO3Mzzj9m9F7Aj2pn+GaAit9zm6zEXCaT2YPCZcvM/zeEht9Y7Td0980UuDbCOu6q1oy+/g7Pz
f0i1JCGSQf/TDNscpacPKPxLUga6RqKUAGRxbf7T+jB567kQJ8a+vhQamuY3UI8izxYOzkiADH3U
n2aYEAuJr+N5z0vNRCuTnvFT06Xl7R9ng34qOrVhl8h9nLOkbszM74dgw/KniwGv1R8vAXNuskzh
Ehmv3MlU7JjRKriZ8gUVoMn3iUah8nxx7BggR2P9nDOceda41fPUxEAYzpF3uxr8gOjw/TtgCniQ
FsdWgTdUVp06Iv1b/5NYAPUkNiaMCkRTtF+4ykuuMxKjnpUl6pqU4BsCPhVYWlMaLgdfv91vq9VJ
94P1nShazv0DLuP8KCpSEykNTLmLQiCLYBrEn3rskcDRoxNG25ulRAUtl4FRCX/0jq7mIGM6gcyk
TNXiES8VrVldKNFBDBZDAnQGKxo2oitnImnWoVn6JsO6d/E+F1OISZNkeHZXsVJ0LzJ5aik85U6X
8AUpy3NvNZzzTEGAn2pVL9YdSlWP6dvmhvU2pil7tq5wxR7lfRIoJ2BLKqyb29S5kLX5qNy0V3NB
IvAbdj45sWkCfIrTeR49s1pP4+stQLYYeld/dKfuKT0MuUlp9VUsKrBGJHG8pvFtPuvvP/jAvX9D
te9jegyWHHjoi8j0Fu8alXjV5YPLXt6sJAt0yPZK3zux+u6jTWhWaGNzY3BQChN5Eed+78x6dVfU
RGPK45/wOaEuY8+iqvyAOfpF3CeoK1DPrUBj3iiedx2ICvlcCwKk81obSMpc9dVNxRkASDcJhWm6
xyzi7RlVCXwIg/3ucumHsb1Z4p7qx8WK3wH7zs3HXHCFJPhnhoST+j0LychSQiH+t3htXFYQd40d
bFIw1W6unSydReWGetrydWvQcjjs3/KzdOdlPEHfo9u6UfJGTIJvBc76T3MlK3cne0cmtwbC+NJ/
TGAMSI8iiCzExD4XCZ8oq41BqgH8BhgsUXwbdVOBMZOzPVF8bpFD72BOWtInY5Ei5PUm4NImWlhO
GeK+kuDNcq6LJFXJ6Bd5W+ovSiqZtc2e0UKtgkw18Pi23sGv+bCjgVod6dCelLfyK8Jw8EZrNcPF
izeyjgYNC5CaXW1nmV4KzoduRU4mKpitC91tjQnokhr1J7gDneifpng6xo9BktuUHYYv5l4qE0Ws
d0x9Nk+cSFFzFj6uScL9djmHD3jksWuIuaRUP9OJ1rTEyVKgB/VbzL01oTpVuQhgYEFCSCbTAK8F
mFXIKQ272oO/pv9Tn80I1rxX0RNqFp7pzwBchYto/kR+5Lo9xq/Ep8JeCuiyMwcuAL9rxpkj5FYi
P1ZPrXMnFFHe1FlW6g8fOtFUH2xG6oe+r+a1H+UNG0K/8oqq6vuKh+O6nh91SLk8q23UbQi4V6X7
uQAQlqqvM4E3wlVhatMSscjjqAHN8klPEqPfPlLMYgjE6VZ0tEUvnJ1y+dQm8J9xrALK7FqQnz+w
pcjOc19zzjVf2ZNgBG5HCR6qkqIqZMfVWxt8CtjanXGC9IHdCtobvqDFPTmMkhHJsBk61E8q7HFa
48fQxn+903UoKHVfKWpfHFhiSruuA6pasOZ06+gMNwE/cbE/KYsfuE0gKfzetwCwzouroKQYDo9N
PD2TcwFQ8JH9xRzuCX4Y73sLgRnvvU7733V0k3kaf655OuqasKwl2WyqOduM7qn4EjitYDZ3W2tB
iThJgczw99kGk7IGU/RfFbSnsTmMNTnSUqqluT84HuLeTFEYHuVwIeynju5lf2n9SjbthYH7mIFu
3iCQ/YqrGbc/aNNvRDreERiQbu5GYSlbfAsUPvYvuJP9tMVRMfWoO1VG9MJO59/AfEnT51exiV+Y
rX3OpCNs9RDVIl9g34veNGUo+Hk+u7XB6FN0XWXnmwy5inOz8Eb4XXErSuEIlBUB1+lsX2CpIcE9
0z5mgp5Oc1mbuKtxoPqEO+S4pVwY8pnHgcmE+GfgohfFUfiLoYx9HPy4wDaMu5fQzRYglZsHVQzs
FKrrolGNvaBD5WtyGuZ74O28D5NKx8qQ/7Fgu5qteuIhQvx2loQ71zM350/IICCJayHiBaCzMXGu
xQceVS2r6oHuKUvDJc6rpUM1lsy/Akg03An7hwsmgNd7aMfUEnqG9t7DCfAU4uzCIfUYlcRMp4uh
6qTngeiQhA0uXZ4ssz6zWQc6Ql6RhHIVLrcd4hVSCunoOxOfe3EAoaiNdR3tZ87ts+L7yuh7/LN3
5Md/Ko7/tlJlOjUlsHSINbd6BFpDCd/OtLsyFvZh9VKm4YW28X96vKPUrpQRjUA/gtMRcXOlnhFh
IiFEhhSKEWWKMXoCko+kAhhNIPfeFW5GoiK+QPx5Vkg2fWB2rgsiwHcCSccXmUga3DXN0GlS3f5Q
PwWQvm++alUwbShWfYYp3jmdWzOlMNgnm8tV1mi3AocaAYZLJ5hzX2KtpGVOstUrLd2UGpGPNE0C
RDxxpYjLL3ZLAyOtFv5LuLFOWFWoAHRhFAKXSTch+L8uMldY9SpdODoPi1F1cntKARfrQe0o+vk1
afEeIFSF1wqPHKtQT77rN6XjtpxWxX8guXSzo57lgm614N24j03MbO7FaGqVQ/5zVIic9LcwJaS+
it+3yW3dYXbciLMOcPDAg6pPbUyt3Zx5ul8265d476ScPh/OYD/1B+focYRW+QoMDO0LvRYYIMIT
FiLLYm+nGC4wan9sEIz2tRBvkinhFANwcG4hd2pKz3QtFtIwkQroxYcEjthd3EeNVZaBNuDYM/gt
CeEU4LOR3uBAUF0d2jMB5jHrKpbSXg8JP3CmvscuPvosVG26rXe0ZT7wTGVMftdyDGCtMoxLkPuj
IGNrFuI5BuUq2/5MUofYZwVnoija+3wU6tOREFll+ARlp9FNqt9frwrTwUUueeEQjQa59rId3bRq
UtvBa3elqhOHt4qAZkVproCXOL/grEDtGAs7boJFW1wIKQSkI3i2TOZ7iFqNK8Kqz0h24LaE4PVk
tRJDBDd2cuGQQ4a5jSFtN9Aj7ke3bQCVjx8ENQbk6pG9QTGKGNi4IwLMvgKevbFs57O7lM6UOqfk
xvb56jCxC0dmmcBEvnIHuq8mYxhwuE/jn2oC0oO1RlwMJKxilp0uhMF51i68DZ4em0szCBpk9eM0
qTvMOYfCsP7j9UOmCYSfcMnpj5BMylSfCqNGcm4jjyFpQjd9et+ME2I50PE0KiUSpZlbnY7sxPsU
E3wriviz2hABjutBWE/qeiMqKGD0rQWVRMZXEP/+fFifOwWerpMfuk3bMvx3Du4i/aPlk0VOaT4p
6MtjrsLTJ0IO4yYk6KrGeY9LUjjfH/mv0JRwquHNaKtz/b2MbQMLsPEuLuLWEah6Eh/z3SmG3jec
xVr5eESYdjIHNfHqjtfs6oBdr2Ff2jvNSiujugvL9n7N+8mk2hIbj5V/L4PRdj8XEvpraWjVvla8
G45ODeDymUnaQIkw0Cv60EZhU1hvJV8HBkSPt9jTiVtleYO1nnjzDnJrs9u2Z5uaSrYS2m5h6diX
g4KnRuInFtH2DXIKb8N0gl3iCOwLhbCOivSRmvpeNq8lKB3+XaRLHhAvQidPfh/7lNhOiZUknTbz
VTLDps+pyFVeAwLCmB5w7crGfKJYc7V98TMSELiO8QAUQOEZTAFMVHwgq7dNFt1y6f4re7MK+cRG
d7/4Gar8SJl7Ep5meWTDhNgsplKha7lxzbR8UPWOE7kJZJAu5UuSmvnIuWli9GOiCmSFLEADO8jw
2LSgcTMdPnv5Q8pRq9ivgW2Mh0uWm4yQGV7XaRLgOq3Yb4CvuwzZM985bMlD5PTj3nH1z4SVe7JY
xbL/BHuEoLkQ3xtyhEV9yC1XN1XAxi0aGBeejWtV542AjdKBG1YfXZ84y4rDrFsS983wTA75eSou
p0ycqcpy7dlBGr3PkYprxBGr5jL+2zT1zQYkjuZnhb9Y4uNU5l1WH8GtUqWu59KNVDWSHpcrKuvq
6S1J0akx12bUNC2R+b0zS9vUk+779/7/Q6HE38wbl31rCgR5wEkoSnYlab6+D2+RFuadOjuRto2V
HB4c93y0ONS5jC3k1P5AnyKjhK1j6dSKXZ/rBa8lisnOSvu/Xsx1zLrxPBPOcrtWZYyEUu5H9Ivd
WXIjxYP6KYZfzjMEq5exu8C6LALw0AhwoMcvu3GUpZp3tAurf7a2uanCEYu/z6JbPyUmYB3Rz2X5
YljnKYC3whkf7LNnaBBRh+kvQ4tE/6uAhEbsbgborvX528i45VP8DXVzP1PbLxWRjnhfjEx8fNLK
axtFGJmr/imQYjxND1TovJ1+qCgyy7xrbMmJxMWwUHEw5oxtmAXVdxkbcTlBYm8/JJR3OHvfnjDo
tHsfamiHBKYFeG4pxACrwl2j4/+6uHnhh9/iCRKOPQsaWcXztmxJskpm74k2AgLp+y20fXLj6W3B
bsFZvdV/7D2zTlw/BvaKbDg/Qp9IPl4tXqLvGVELlQ3YbYJEyO1ykHtyCpuoo6/XObUWGly1ASz7
I2g8aPaUBqS6PenyAoYsWx8JsZ2twWN5/O7asGmDPHAfU3XYl30S3DmKxERNQJAfOuB8rKQ/366g
4XENpQHffjgXPDp7cuLsLpogHGYfDiQwbqQ74XMIIsO3uZjF5W6bpKY9PzPQKDNhfVc7uzvkt5A8
jbQrcjKGEMrClRFgL5IIKuY953epGN69j+dWFLPVw6YugFjJrw0i03WkxoBCjmlCiTjF7nMEHFmy
p5ClOcVmK9JINKfa2ir9KyY6CnsECte7JzK/HIhOj8bum3GU/TV63LfC70+o/s0jfw6xWZcSmnbO
JMTfAnuyNWM/uzPj+mXF7y7dtniymg96zjvpa9DGsGL9fTcWmq0cZ4cGKrdZMiFiQamBzpLMO444
mjnp6v44RyzfTvI75bEJvOsFSQ6y60FBG4FB41k9KB2MsEQqolnj34B086uZ2yCbLEakaJuITT7C
U5lm53YA0ivAkeso0bPrsdct1b5NHv1OpWwwkiMqJGhZD15KisADwXaCkArAlOAh6OjVqH9gCvQ/
zUQZV0GGAyuJO781mW7LXDWpnBl9lKYCfEkMMOkPbnExu4LxyZP7Da1Z016EmraHENczaoJOaGDf
/D+cjWa1ej6TOGKL8oCEzuhYembIHmZdW6PSgv8HZtXurSyslI4hEDnjSwiKE0IkGvYB+1Onf4zR
wXhplT1PiYSx5/8/AcJ0tqnpa1Wcc0llp79HqSa0oMMjUNsuzKgZGOHd19nlX+rnAsqBnkUt25Ay
osMFa6QY/0euRSnLRjDT8UUzUQGR+cSZ0YXDx4gXSuiFw9K+kwRt/GBT1sC5bYALI5AutYqWr50J
+ouYoLn5waqNNADaWdFM7+xqStVt8MgwRiAxaSIpp8wVv8KGz0MqHGVJhxsBkQxnFASGSSGh3Y4L
TtiMKoZ0MPlTg7m0SPt1kYIz2bMJG8iRD4NKtQjRX9wNIv+1r4/9ZnBY5DuMkuu5UkaoT04dUc30
Ymzz5apGytvLKcnghu1VgL/51UJOICUpZM+cs2ypGqdXhph6aKgWIPqy+Or6IJiEEHhSgNmXaeh6
FlmAMp5vuvhh9y+odh+HfN20cmRmvMXUnLBP0RWfgPkmScDFcn6+KgF+FeFeekAW0MN1QDUq+Nlk
9fqKd1uYlX7dqF6t1SLpQefGDXcepHUzgnI9nGstQ7qiyPzCb5d7JjWtD9I/onAy7jsdLCrgdpbg
NxkP3aNkKlr8kFAxheVpXJqu1o8aNbdGBOhGlve8sop61cm1UJrJuQdLuUsXJdWPpcBzWe0WWz/p
U7LeumEi2TTpN0hu5N8ZOeyTfpYe18cCHU6+n/yA+BDAPIUPJj9HK17qL+iguvpg7fWFDq7RqnvU
22N//Kc74ZRltugfYMbyp4MkUSleLulTtDiuottLJekJqDEzRoKqYX0yXnunmaiU1TIjvXPZyfav
CXpUcz6pUVFzgCTvF3R3eWUUPbgcoqB4kjujR/3Of28z8m83x1nrgq9YCFBZ3T+6gi17SFiM8b7S
3YmKuTavWsMR8OwN6eMEg4zzjojdjlD9DbKSsCIYpTcMksAngZb0OSGxg08Jhgwcj1+OhVMHkAPR
+72Ad0YakJEBLlC9r4bbS3n7d/rCbu2OrwJLJqggyUoxVuzv94XuORWUWHyTRhkbDfgYlKJTUPc9
mpl2/NlnkYFuRCRSw9gntPpmfduNv0jPtBozY5vfa3SB9SO/NUwVP+gELpHW7/nPEwTW40Ttxinq
BhROUMkxb8A2oyU9Gi+0QXWgXb/0pt/fNqE8hFb8zF5GPrzGCQWVRuh30WLhHS6FVfcyZy045qjA
ZB6/ZED4IqzywmsWSCrukZ+jr4w6JwVyaLPYQaGrx2hoOFt12eDZP9+GSiruvtERmBEubkMI6/tS
lK+kwDxAN+YHBc2RFIYS5rEh6L7I5IbNl0KF7LtUCaVE6XNc0WNbCzS2fQu7G2hcZT/nE1LWEHe0
2ShJND5N5Cia4eza9vvasIEboiXEA1pEUjl3aZckHyfHweMm31O0Qtcp8LXz8RESmAMN9/J1WNXM
DbdLPnHaZYsNS2rv/nwWrApP9OfAKv+VNPn07QbGRVKNUMdPNWW/PwwlGFq3/L7ot+eWEJ7Hj4Jd
sp2pgU1TMJkuTpi3ES0Hnzk2S3/c23q4iuSFUMqgxLnGs8rsS+EPIgKslVQy799DcCD14HXjWY/s
qW/iie95DTf9zsGzlKOX751birXHZg+ITx4X/R2fDSkzr7hDTsNBV4GJOba6ZieIfvAo4X/X7KWV
CMnV9Pmc4L96XJKTVo4oU12bJ0ZRNUNtPt7EmM/2JOPTNuZj0Mp/KDi6lrIur5QNysFVIkacQ3fv
1A3LjxRw4fBwmA+FCUQex7zt4QnktSqeAn9QETP1fccmYeJ+sA/lEJ4aLZHK6XhV7g22aVV51093
PjfZ8oExSPhYlJuUT94a9wrcLRxaydvOJ0+qAQufvRmU+pZBXSC1KZSsFiB8hq85sPGGu7hz+/xr
vQQps9gw8wzPe9Danr1B344xW4fltcR6kKunBy2Cqv7d2eRk2jMiQB4tP+hXenHDrmOoJO044TSQ
RHHnyscA+//zpj9r6x7GZJL3OtljesLrruXy6eJmFhI4h7CcKM0WJa67HRvrsBYbKOrl6Zb1oz7v
mADcab13qHm6Z4ViI6cOssW+3KvLnSu54nE5ycySvAqEEyU2gkA8rf0d1m/2zpZRLOhJ4KtNV5qb
zI9o8lfr+zQ05ts82bkJB+yYYLV0z6pdlock8yO+vGrFj89pOjQTbOlx8tYBcvkI3paM6EI/rT88
AOiDnHnVx5l7HKpqpa3qU9nNchdnlHnoXNiKOBZN3uOxTiX35oA8gM0lpgqtYUQlS8ZKnJVXFuAU
hBjMMOEtYtIu7/ZV0psu1+lI6QJr3sxxuzNNC0/3L0+q6yDTub9GPpmG3SD/RVAHV55PXJz6ARhp
2GmargEa/z4lxFTlTXDxm580ZJBtx80y8qoC97V6KKxlvSlWOirR4Im7aNrKIv/1xPdiDLNaIRF4
uRxSxPyTF8XtZ9TvjcQI8RhGR1wWrfQtrcM6V28fkWEkwfIMRAZ2iqLfmuQ2kqn1feO65WvX9fIl
bCgfKrSrDafZzynmKyEQcvyNYxskwAXrmumFjjK83KwVeLvF4ok9kcmMpchg1o/Ddy82oVP1R3Lr
U7uK3UhucxYPY/DRoDPQbGkv7om4Jbv7H83UM1cglEU6d+yjlyE3QQhWQ0dOZ7hd6RAV7GV7HtYJ
w9hKdPkaHM+bEh4zTgW52hPJsxHK/f3THWv5zEHH+0JEsQ8gJ3tY7HsGGT3VsJ+mTZlHid0NuHI+
VvkXtSWrLd5Gvy4f5bDpEo0i6a3cKCOTxe+v6wzFgRpSqs9WgxRSCqBi6DczjYFRB+nhM7ULXHAS
I2Ec+D39T9168mXWNlOlBubaoc6X7pUOjB0E7yhT99NYXSiDDQub6ThuTY+mLJTCwX/IHuO37vie
vjxQ/8RXpfKof+IfESutSt1QZDRqoZad9ZDlQGQVutHeXQVdCeTwS7y1IoOnKB7vK4awLs6zIx1R
1EGtnte3/zyawstzwKza2uUWoqd2/1cCixNMTQS6UtHJ2RRRAYB6KuRvwCgrKtqq0oVn/InvtrG+
KpZMfeG4WBaOZthJ9HlSOu4KBkygzOJKoj6SK2Sy6aCVrITUIZe6MwtIY0ojTDyVkZx1NgCvGFoH
fVWBP1rIhgP5XTX7A6OTSSED63gP2SaihHj193eLEsMbTYRndnGLLbNNRPbRMxqqNipOfsdQhyr0
weGKxeYyS9mvebCOGi2/f3d4XHaLPxSlry5R1SsmvQc3Ud8vWGNIs+Xjo/xioEEH9KdQYbVVoWqE
dtjk2N9ehLjooPlRDD0qUPhd+CBwC9HaRpSROoa80slzN3GoAZ3JEpD2Ra4BCSPyLJaV/6pdUSU+
UvMJhfsTuWQpRM3MeMKaBH523mE1pMwRvMa0QId7cqEX9L9EVuT2FchzPSWBcV9oIphdtXe4Dsq8
hTWY0LztcV+9omrNEoveEoW5jhVHG+iiTy/QGp6ftEdWOG4xR0dMqrjm3l8ywoZtVvkyAcQH8nrV
I+FRgdS5LDnAqBX9W060wghdJUBvobLFFvV81X1ZtUpg/FhGGtIxHcz+IE6VpBB7XwnZn18zzZey
Uy1tJB+TKRTaeC0keG/2DMlAFz/MwyAkljYJ1n6EyDDm7PPTD0kxBB1oCqZXxIE5rq/wnoC+8bHH
/jt6NO/HHAqwvC6cYqFN66p+sppV2bez77Uu2MJ9GFQsGca3PL3WF272+xeERHRUIHcgh35KRQFN
+qKP+6lzS7BFsjeTSvDyjFXxJZGje3GFvL2NZXLqoov07ZevsTP0/qSuElL5jqCko//BQNAnx9hn
hTMUlvf8C1f+j+9OJ1r/1qsy9pjzho7k6ra4y8ozZdVPJtYVz3NyXM12yaLks3XEFxiV5bnlWnew
V9/Q6j1X4wCM41PW4oTjTXGKAnMjD5NlJK1z86IcHI5v3+9zH3OXjrLeU0UqcnknTzHq2OhWEEi1
04fdOPhdEZ8jya/1lK3o/zxCC2CTW9r39EtHY3D2ctqS/bRSmcJeS/0MbgTM+3VVQMkvX+nIFqTb
kcYZQwxNoFvW2YuwNACPo376s9Khv7OXZfIZSlFPWO1s49V6GXHYgtFGN/R3O94Ya8BXnv5Kz9Zf
wLlrfARazhT43B5j2Yrjl/e6SsSZsqkUW8CM9nZ9k+myysFkrsZjIkNkBryrNQXOb7NvzCVop6XM
tDKAG8dAHkiOJGBYA1deL+ALOXw3op5DLuYzvfl49Ej/XrYUqjF+wUt/aVawTc4lAQNvpYCfr2Lr
T4Jr2FQ1PcEaqOZZ3uXfc7Q+ZqP0pIORItB6hmw6iUdRptt0R9hokpq5qekG+qSQwkFBHt5/XrYC
N03fZlbep5bgcg5RZMLq3IxWA2jDAAJUwzyaZct1iJr4AOPr7n5ibVaQp4CSUFnnuNe2jbwzmj2x
TluBzrzsZBUsE8hfENdHJV9R3qlbl9V7dMEneYCwPKhDyW5Fo8EZQNCvlpirnglsWJmot/63kK6b
St41sQeXVlJ69KQJZl4gzN83DJ1CSw4rvSDcT42nMyhtI4o6i7WNcwOaORnKrXA7jkF8ApXTbPYA
KOG58jYJjmWU5rtalCLALplEBSTZPfk5LIClWP+MG2/Zipv2txMPEYoDyYIOkdzG/4e+Ggyq4SVg
u5p2FAHZ4XYT6KY5qe2N3wHF3hkGi+uJ42RxkVg7NjPputMx3WavaZBgNOYF43Zwiqx4YESV2B8I
JwbtqBMEuYA3eV8txKIqCmb1qyDkZIO4XgiMBdJe34qtPGKoaGVIW6om+rXuFd+ySFqSXiXrTgMR
S4UaCkdyLZY3yOpSuy6SZewpECu0YXeZZDIS9wFjtcGNyakMxdovT3U5ESZVRc+gALgYDYB2WL3R
z+B6lCA8NVtCyQ7gsJML7nT3lk1F30lkRNzznX410YD4Ezeyvdqw7IyI4aK5gw+mpTa+KltC3PNP
8zvdGla01Ou+T2jQa6mCyfvHd/Tvz2iXlHehjr0qpg0tehN3qaivk4j3Ywt0ApAWrrlSwLlZZ6qu
y5PXmCa+iLs1JJKk1p6pjsB8bK+xo/E8QfUcO+JU5r8oE6uF7MTC+m52fahJcN+jonnEvHcyV1LE
1eTY6XtAHS2LNZQ2EhpYEjkTygpedlxhwdATk3rCNKTZgZNtL+5BGzspQvHGTueD7YTuUw6bEufV
fifKZCNSLbaVpxdziPuwoQ+w0r/3EmXDQneoNVoTi6HDXXUWgoaUdSG3W/C60om2Op9NNCrzMVa5
i60m1BX2m4dBMx5+WBI5I8vSMZoO05yDF6kXIiA44fkktwCT/BLA/3xt+lHXcYF1ppNWcRfg1SdM
kmg3xAkvS0UDNE2uuGC9i3MGsjZfNt5KtkpccKhvw42YnxJmw2jlyELZeDNQQpW0jic1UKXZQV+x
8YyUxVwrytij4WAZ3+C6XKH0BQL3FlVBL2rjrio77Y8/NO7rwbrfStKC8H4DaiIUgdLY6T+f77IZ
6WvJ90vRWeLiL/qabgv0neEE43lT2dCtLa4CHTPLSLGEFVn8JP1IaF7dZnijIoE/mNdevyg/OJvx
ieIHzw0/JD+852zVZ7dHR2KEpttFSaWA9RcgyNdBUoMgcoksko1FEvkLNdN3U9iHrMI7LLUUEQso
kWQp6DXPbEy7vrs+ODv01npYlrEXM8Cptv/3e3z1q0Xs+KuSY8T2omUBercCdx41SiSlm+4fgh/3
JtRmtN3XgLwc2ap+MymMHCshG2t6d46mZ5le60yF5JlakY0GFT1TSV6tHuvLVRqFQJ4LZ1QLmYoi
U9F5o0UYWVVpXykTljmSxjRbjchVrXl1CNCteiorfQJTz2bYRcfHiDvmyKEcJBobfubqW5Q97USM
DCEQ0pgNOYYg3CB90cj8Il5wB6bcSQ4S7UGDTM1dc46OQu2axEgx6Z6FYrsh3HwmtUSum/k6WLFH
Ufs7wZ2kADNX5lGkbjro8ajdJqkZSYwprMI/KiIGo1WK27Bf14mq3KdKIta03PBSw5n0mW8HGvNF
Kjshin4HpevAyA8uyS1FCmyo5A4BXDEfAxeiuZc1VKs/oYEbVZNymDR889hjjMgWZhn5uPvknQ7k
LgaBCh1rr1tyqDpgm71GPx2JoMFwr7Sg1Jp7PpXpO2NX1pBIPLkxqyseo1Ae2h/ClwkvkfixC984
s+R3x/QNorCby9EZz2aURMETsD97jABxzjr+n5PL7IJl7E49s8rKfRDVhSPlywB2rrZXHmCXvluP
E44PLl2D5nw2uHnCR/k3R6tzr3eZgwCAzBmWhcJzdHbb/2F00GuEgTzUGgNFzzwPjS+PDH/IxyjW
XeeHsonjxZh+LciIC1mdMQOWmg7VxmDN6yru50OSx3DMGen83f7zWuKuh5ns5xhbJK28QuV3FyLr
ZHIZOorBYQIBxmvdzSX1Qc8+bfWNqDzty7NrltZAn7Opaep9FqpheMR/8i/m7ZxXMDiHH+uuTfdP
ucLkc89+3V8utwbjK96o5xZBnFRhziQi0lIeBNoXo39QYcqXhjAWFexMLlyv9XQKV7AIMi0ShThT
JAiPWNp/AngseDJ4qt0T6LKtl0Wxq1OfVeAtFNZB4Hql5IGJvyrSEQIXJnpJsf3otg8JwQV3d4H+
oB25bjL1vhNwCAGSjtNvQQLylsq2u6gvPCFgF/S1iLUz/gV4dlrhZr2ESid04fJbn080/tURdiwm
WdBmuRtIixGnkjHc2IcpYRi5J5v599D9U0+esaCYMIpz2k7QkVJKXugAL+E4Hlnfms2lwP0cthJM
/KmjjxhOH0/TgfPBfly9mxgXFTEhtY8QHl0hKmvZKKUfuE9MO4viPwq8popMwH9B/FjvjsY7ifBs
HfQ6H/2GUoe31W53RMszluIT2zkx+OkeO+LhP7KTwA1Z2lWgP/6QtA/1By9QyFM3Ru0vg4BmFg02
tTx+1gFZO+T6ZXoYSgBxnXgNUBGMdz2TPz3TaO4UriZrP9YJZLOCfNpQst3GGXltXSuPL2e8z5sQ
o0CjUMeVsO6Lc7+kgGowvoH9mXAE+/yTnCoBvPc0lbosL1cTSzEiYVDMZZ6y5wq+tfszATMvs4c7
taFuiqDZWB7+ZA183Ap0GwaQGdv1l8UHvJxJ2Lc0psP7IcvV//1ij7InaifrozUBm1e1z7bSRMWN
lFShiI1DNDS1chyOtwhXfRuRLMK1Lg1KBpyD0oSeyeQEVD9uzafi5WNcfYe8sUDEyxx3LkHvvYwZ
wY8El6J+iR8w9WSD9b7zHs2DTe7y+4yXX3JPITNkEccE13U6umok3+gUGURpwOgoF8S892RlGCCU
IFtbtCJfSpaB7+ksVRi0pI9qS3AvO859LfbSeIxE9MMGjys9A6vIm+OPbZiX4vJRGVEon/9smCvj
Cut2v6GY8D966pweJBNpSJzvGsxaXncnmi+BcGIDCUH8qePty96F9QQUHSvuiKRyVg3lTOskHgsr
FDB9g7K89WmKeE33z11otz6lobC640uL4WRPhRijUlJCB0TYJWeYCzA/s6YbmUIygA3bO5X4ckKU
suceRcdSXsi/O7Q/WC0vgKlNO19RHcVMDSpWmucNNfZmpFP6ZhwyqaGU5jd0JbRqYgjDcfgGWYVK
9z+EJJcSuwlov16e86bIFsbh0hbXaNEHu+/xCGH+ApN3fNsZEmnJkiXI1OdkM2CDAy5z4Jt/pP2q
MDfqJ2FvSW8GBVzv34DZDa5Evlu3nfPyMFWkz9tQioGBRVjUByTz0cmUdpkU8bETKcHnyTWw12Dp
cHJS6Ub8M9xiPxnqUf2TMlS0dOrog4ZVLekAnipz/Uafy8Fsppl/DYZLT2GL2Pa+NuX1md3i3+hN
AFqzQc5gaSpPRTVPrw7LOCTYU6N+geyhdFw0eCa9fE83aR/WWoOfznOK/m169viamX8rwuRFiQGe
JKV7R89ijR7uif0BmjvcsqRIXJcDyyVNj0O7Y8iSErpPu+p7CnxYUtv5UCuXwu4K5PvmhDfbYu+w
ech6k6JoDcUQaGnnj1u9IcCM9PGLZ27kLqz0++HXHm+Hi9XcE7V2E9jxZmFVRsD41YC5f42cJrjP
SVvQDwHPt3P0TAB5jBOSWTS8557wsyg8UhdZG5xWsz9Yrn8mauP6nava8P88Kf9yM3tX1jGDqatp
HJfhyB00t3QzjaUYI6mxmFtSApA7WP9wxV9mKT2SxTHrS+kwDmA3ERgqziD05XRW+0AaGn6vd98i
PyU8ghMR2TBgf6CGWFz6KA06SdCI7+WCDMo3pOMfJmHGcE7CcDu02D+mE5w2DeGeETUowAXPCfVP
eUTTWpdNQUHghTA4aHlDqFg+eCO4xfytj8cpwTy5sJ2uzl50wCnqZVM+h+Fe8m/UZhW7hTosap60
sfxSbNW1Qsvs62jLrHMjqAJFYCcppGrU09PtICBvVph3lZrm7KiY84x73nkbh0b1ycCNZELTovwG
Hf+W5QQs9TD5tmDf3IgpSo+PNpqC1GueeUAqvEQpXcq4FrP2X9+XVXAwbHbtIJy8rbUHA9BmlZU4
b+cigOs7Z700O73DkYT0fCSQ6aYrf90qhlI4dIAmztV31h51/CBVSYm9hbR/fcMTBOB7oxOM3h/c
j7Uf+Sh7tDAY6vYaiTHZo/6dzVWhrjFdmXtL8CuGVWxY75T75cY/JeAds2mBNrqay3ykXcV7me+g
t1WpJ1RX6Cc6VAAyf+zj4ldb5qdbwZ5ExDNimp1fsv+kCDvtGEUWjVOx9fOTZjUB7oMbe9IVQxUx
vEh+bC5u9MHvJRLtrD+W/D+hvJmqEHR60nBGlspeOGTKSoZiD+PFUFEPqweFH24tnye/SM65pOJN
Asn+aIFltYepX4VeFBRaBD436L0JYRYo91QNFmBYC04hjmcvLg7nLL/ztzhSvT7+EAV27hRr0rmw
Ebn6h9ImDPYfF+iJzQSyjvyti4LVrCE2OhlUf5sC263UaaEEwGClx+6+AHhwv/+a9lBtpiRwGrm5
CuctIBQCt0mZ1odYA/t83aYAt/qchpFBX0KcG4KiSgidCfTbwJjTjlo4QXtaPBkNJs37AMqfAmIW
xJ6lQl5+iBRhHFwlVXHcODd2Ol0As2cUrUVZdUnPKLvg/Ks0U9Xuw5yTVcmVTgma8fe/6T+0hao1
aAi/Yqz/1/erO2C9zv/TMeUnGzfQh+Zib97e7luTcsVjvhMcsaKfTDyLBtsSY0duedUwQSLHYaD5
OjVyYSzTKz/yhtNhTDc696zok/UQloK5FpSp4LPwxYMTuULIdV/gbEWhnFL+4wHOKs2pKBvjHg6z
cYuxOe9vHHL2oS75iNE5ZzG1YH/YBHpuTXIhd2cZJdRjzrLD9Qbwd77ruMU7RrxQeo7wMBrIyQZW
cwGrpfYx4lVQ1zbiYSnsDIuBzGAW92BrMJuAfO+gzS8Q1rYygUTEfVGiHF2k3cQ5WeKz4KSnOe27
kIJSqpV6MCwwlv8r56QnYoSsAVwK1saDrTWylI7hxT63I5kd+pIrNVql/vQ9EpeJZ/z9F0wPoLT9
Py3hIu8GsUp/Bu+/FstPjck3+L9Zvl5lXsA4LmTjeQ/m/DebJbKJSo/YSdEFM8keZxBbUTZYqKbF
uI5zb4xfnyyJXwL4vuxPGHMLsLoPIyotb7SuWad2hCRZoLlyzbTl13Ug88saSNO0DcZNliP/XSXX
Ol8kJSaDJr6qXn2SUo2xF1rmYg8F3hxGs1gIZHv0OvjZCQtpdOH4ki0T7OQF09rpolb4hLtYV2Gv
Vh1eIXcPoA2agEzYRMFoDBxlrhHlshYJtNObp/poHLnm3ScsxWIDx/+Nf8pF6DEYgPa4/lvEgXWe
wikUIup20v4svN9RRL1NUVwNPtekspoPj2LQS3wpB9JDnawCoblcdaOeCl6dviKh5NNFL9jU5efY
LlH3G20WKRojJI215u/DXuZ8JfPNmel+teYsB5KWud8m/wKpBPjvt94Y88FvnLIKtYf5z13VONgL
sbbFraOq/RigD99eSqOXyqFSqPbb0npwmcMi9oAUQIROpccvkQOVXxXvs0HWgXGqql88WuZpGZHQ
HU1AQYcydEikTv8DzKzLDrKkQ2QcLOKcMpX4AYUBRlqSaBOAFQI+2uu21TdbyKs6JBTh9hac7lzs
90tMOnD72J2akxP51AwW8kGqZGCV940aYeckUiOidZ9DrhVTwWpQKnQfRzeFYqaUf3aU2sWJF3nA
UHjMKbDgGVwz31Uc6zgS+DuIZxPmSywIf0atK8kEX5wrIvoDvbOBAmdBPurLl7kMyib0572v2Tm/
R/RD6suveQcBHNNf0yDNlGd6YCnaW6LrqJir4RCHMaiHNzKevnIuQ9BrYuVFhfg1iFL+16uGaPN0
+1ON+6qVdy4yMS3ie0YTsHXGco0xWGhSdo8m19XWS4IenNKHHCP/RnZt/2jDLeku4UXvBoWZS+OZ
TtlQnNW6Dp40HE/ioKw4FYL6rQCVO9HS1uNpfz7Nmla3Gw0gJzOrHsgk5ogbXujRfwHqOM78U/7O
JZJmbja71Xy/lg9GRcQ+PemyTLD7wY3ho8nL8GqPp52/6y6tL6eGdQhTgArzqvQaLnTeRVS0S05I
4oDgfvbBAJdQxDKWGdaJEB2POZwOG6xBlq/1YNPmP1B2/7Xs4Pq3U5YCQuzCRxmamWRvnsY0v/TE
1rnVyj0Z86rbvg+n23dUeTruiTh3hTULM0rxUQ8Lq5P434J3Fle7ns8IIwK6OC1AqZkBLnKwCgCW
YeQ1X7Dq7deWfL0oeylWsAWDM6OT6uSuzZk/yShfg8DIgHOrYZgCw0EMre7lArJ9xQyAbASsxGvl
3ZOs6BlB7ozQFFUzK3T7PveaoyDX0QCFu1D2sb/Zm9VYctlSfCd4oVaGAFDbbUVnBlHvazU+8pb/
/FD0III1avYgwTdK/83X+CNPztZ1ByIThvE89I+npJ4+f/e1SXeslpAcy9nWN4zn+GZsB5Kf31tc
5FyMorX7UW5IQs+w1O3aFZ4Ofxb8UfngIhUtjRSvkH4h+lUyEIlX/lqfTFib050565rIog9+EBXh
8NgcfVxRNJYDPHg28Cu8ybU6ih66H3VK+h+b1VDjgnvtkybP50pr0X5dWKLvrY1zRzH9/xaT+/US
dGCO422cFzTtUkmZ6Kvn7801ZBECxoopxGW+fmva7YipelUpnf0hCld0uKwpPmQ/KQJHG3SalDkQ
8FqSqJzkf7SL1kK+aJiqSU9Qs1ObZbhBP3a68ud5S8V02Y1S7cQ4AeLlR40wU/qq8MNuZBLNEFiV
nFCTd04PRcwvZpGaxhwied/6tqhcXqTHbkDu2/jxTua/pkkq01ukepfmEzGquy8FrQtpFxlUpAE0
Isdn5+hRCzqCYIXzAZOLtFy5YKeQQxepBgmk8tXzMPQtldJq2r4C9hBMNNTgsLgxnT/f41hJoNsg
wJLMFJjMRRlroPXybTNEE7K3y4dDvJj7cAIb23OxHHic/Hka/TCBFLb7kX4Q+4GoMHWOaL/ywbqi
sMxGWwWmVaZzihI0upUdO+SWJ75zPLkukZLS4JKy96qRY1h/+Ctz5gLwu1iZ2KBuGu0woLqX2PgE
QDTdg/YPsD+932/uL/JExD2Rnt8OZfPs2qFvSCe9p1AE+mTmMf/te0wFtscX5rqEy/oo3940wuLj
C9NX3qOxACzhtG1mPFJEHIzSjXHb/GWVW5fzRtmQVUwFvhTjIde1QT9sbTrFM8z6SV1g7sNRWV00
0Wvx0Y1Aue/1Uk7p8+2BB34tNVdokUh398i514yV0WtMcdXxz3FJc5USMfUxG6w4SfSgDalU2RR+
oiGiWrFV0661Ob1MVk4Y0loALpr7MHgZViCjAs3fzYdtXimyqC6ApghtHp37LSCNvgjG7lhBTNQL
VYZvWREmZYkVgPCpfnCIdkmLC7x1e0XY/lqSrXz45D+J3rIFA0TSMwROW7HGc2ivAVKrn+qgCZic
ZQbERABO+AeGBRSVDEm6t/5iRAO8+zSeMhh6PocvWq3C7yogJ62DmLvNG4XVpv3fEstwlGmZDcb3
gXp7NLvuAb/KfWy6+FHKYpp/fVKeY3A7OMJAdGBbc94LL3VfuxRcgVcK9FLFvQ+WZHkVvQFpFGZ2
guBDjQ2Bai55dWqRyZ3wfC9ctBUdseJaE4R9cGNUrXMnbjg9KhUYZNLjWr/MmWz28TiIBex2EreI
/6SnEQMZH5lrRUN4p21qyG2fAQVeYgvQ/MpA9uRLDlc0oy039MfjmyvFB4ZH0Aa6VolhneesPsrq
DywQ9b0hZNHU/epDrlmA7wx119Kssu1IHW4W/ko24yX/owloa7TZE8mb4PgsVuNERO2EV3NEZI7I
sFlbh5U/eDN+6gQIB273Q+jhKqt2Yyu4e3VrPuKOtoqr7yMOexWPiFgb9SuUTh8xEu3Ev/2vv8f9
YeHEYG1N/JPuinkr1BooMH2eo3F+VkpTa2fE1mLef8oohTR2+nBd5Snp7aDTdbYWDH+UZnUG4cvm
cMvRPaw0I9aQF4u95Q85mZWiDwgj2POQ5+mAwAlmGJqxGru/X5ID5KQw6zNtw9t3+neFC9DlCWMO
TuWthMDfIx22apT0eEAZRbXeSRf2EK3ULA2ruAi7mELhVI/xX2WGr1bV9YDZ8vYm8PRfNe07i+7M
KEb8tnTUG4VvmXNAThjDcb0NfamN51gefcpM1H/MR5zCAetYP53KKCW6q/s4tGCyJgW6oUvUWUy+
SJawePZWyREYr0Vskj5RCj3pi2XfT8oJNNk3Id5HTd7awHlpFfP3x+ZslA/Z5F+ke2h8za42TG6W
ibt4O8uvILva1zS+s0SqWnPL2BEh6cqc6GAc33adJJepEn8ZDegD9xG8RzypzYN0UsVbUMxFb7NU
GwnYRyCa0r1x/81Ccyx41Nx7v8ez/1XqSZPa3RJ9CKwmT06T7bhzGvZn4M1zrlgsAmIoVdp6JsRr
WztOkLFk0VCakYa20ythh4vbaYjFm8QzCilxwXimbUsdBhLjVrfGCenObbOBWRijTJ0SzuxetgX1
+f6lXCoAkyUnSR2nEwyit2/ftCQUh84QsyrdGy6IoxlOUrE2HsLPCgHOK+LhvOg9feUKaBgjeAJH
mV8/D1JxkRtqYcUlbS4uRA0JmDEaqhBJ2H0f/EQG9LY0xBoIJQESPskLZglDfmb3/tLA962FPWsO
ywr3wf+ys6NZ5rcp7L3peaMfHgIPLkAgy3GqDQFPXT6ws2+M/1YnPtNaVbNMxgPQva+UkhqoE64v
eS0OZx72/R4sP6VpplrPISNsmkHnL90gNz0R7daZj3O7h6gqRouLMb3SeZowvGElVHfPb0jpTFPw
cSqC3iXmWu+D9JcmiooBn2AaQCrybj/8jY9OIsHuAgLRkqIFJLh9p8DlPclG/9JfDlJ4XYd4TGjg
6N8coyTa6dDcEsHVqhEBLv083lkk6qF9be9+lwzYuJLdnmeC7nGbl43ndNNLo2X3xoY8QTppCaxd
chWt34qYKNe7SMw3tRaP/qwAXqCwGVFO8glipvLGK6U4gbkFdd53Xv4Bzv3v4OzszSXIOHdQ4Lma
jy+n3DWBsw93gsMfFoKgDlp12jNbO9xFnUgohRM1V9pIweQzi1LgezyoAeH1elJvHzEWjVB3Yks1
tse+9iUSZGj2OLAmv0MKNT5hqzV52z448PevBxMAGRh2dmBXiVn9gRnVOh6TYPnUqNd5LLxnU7EU
mrwuXVzxH7ClvLRgMA28glBmd9bnrrHKpVi7xPXCEhkFyXvbrIkuTREKLsBG+zAaW2V3Lpj7pMAT
cPeKPAwXGWECioLjDwBU0Yw1wkEPdYmMq1KpJM0n96MQZwTk5UdticVlk0TX6zvpOdLIcqLqqUjQ
YIqQQegX3DI/tiMVuzrNVjuJ/ukOkeCG1BbOIw7L6VVf1vaTwuz2TMPI4sumFWurHASH+AGHtPc7
zS4jGegYUre4RzwxcPQXsSYqbtEbSMz/Dd1cf+gFsKVZPYPa7qGkgj8kT+klv4uVgvD6J0ro97Jm
AJJ+MfOfT55gJYVAf9KkTovdjP9QGeEpP9lPjyhPu9AeqYWkOj9aHnIrEDNDkctylUBOdxbq7Ef0
UK3IZBkPwccuYorQnN5ZDVGODfcJenQrFAnuhmtF/oj6G3Ey4sQf3v8lPMJnnNn5dJA83So6dSAm
VCPKRbC6y4qMrcu+UxKKy74rdivnZivUjlQve0g303PPQbXLAjegHVyPa3nZ9/cyKyhUa+yI+Q3N
GdhIvZqQIr7sPqvx2F1/yIXFSKEEy9dsE8MXsP4rV4fEnBdOZ5I0P/wFkhKhbmZ1kNgDmyzvD84Y
cEiKndIhg8mp3NzLHVdHkqoFwtLG4dwlogk014v6wfp7aRpq4pFW9rRsomFnoMcXww766jl0xVGc
itwZF3iVmQ7lfzdVVP60Wti4Hw2EPFAkyL5a12mES74BD8DujYvg1xl5/ylr2CcT9Nah8+qEcVmR
61d45BOlUVqjunFmjOmRymM46xm4yXq3qTY8Ha2Kg2u5+0ZlHEQsBLvrMwmVnZjVjGq+2V8zPHsk
P/lk4bpDgVd3QmIsScpPBbB6GqhG2+Oirk6dz8RSD7xTCA+k7iAy+e0xbzyvo7nO7o2XDlmy8RJi
HXkvdMjraUv7WWiiNCtUzMwgmcFVIf4Aoc9P5dD8BWp/9gJ9JLUjCpu9ByjPJtQmjXCe9vT9NIq7
Av4mHn/YguDNXvRQDkbKc63rn1cHQNcmOMyOo0JY0EQ/YpiKBrCb4pBGzv6AfVZK/yVA5S/xMnsr
8ij10Zma5TeTlNLxCqXFSqmkOwJTQLsKDTHGQSKkj9oxGuU9J4hJo9uwTiOd/p3wwHx6o7uG8YvD
JS0/opzSa00hSuG6JxA5yBtEtc9+xEooEUE7/6LXFjgxFZtJ4/Uv4Hr4FtYiWZRZCy6P8lJvTI9C
2pjcg3l4V5JUqkROflBqNSpQq2j3Tlu+2XYUA4EIkvxd6W7oVsHbAD/uLfLnkCHjXGmjenxNMJMv
y24WN2Cfnc9LIpAWT0XInB5REKxlM0SG6lPngIoRJxtmtJH4EY7KOXw+tW8MdBeptAwcAx4qS7MJ
6GVT9k9tE17rTGZ8xrq75n79KP+LNZQxJxgUNgKbwYGzYbxJ6MS+Fz1+hNvHk4UDWxM7NSh3y095
g4b1bfH19LYAL1Fl/khp7JzKKQh9+vBav4qRUanctRCAYjHK9LiHJJxAxb8wz9GOmSpUGNhuqP0L
93VU2mQcMQ73ssUrN72yC/y0t60xkNR5A7LfhLMjst9RywA9MFtADeAcPQXeVIsEaK/xGShAI1/X
X5SeGZitMNNtyVoY2tDA120hwaAfIvIelyQTRzxXeF3Sv0UqqjJNaZYGGsJUjb2K77iKtr7GQDFG
hZvVxbxuDMh7SkFI7MOtot+yQB5zQYKpyJ8P4JYlV7mwV4geebb62OV/iuU5YJkas2yYU5i3Cdgs
UzJe1Sx5no3N6GuMFjypN/Hr3ru1ALTVhEfdTe2tfQnjpPkFq3kIY4mWnJe6bfAGuKbuz++P3Rvq
8ghFrQcIst3MgPcAkDb7g3ficZjU7ZHryGinbM0JNtECmPBxnbk5h75reWix1NfjIx4KbUuixpop
t1K98UdyB2vqM5EHKaUQvKrZsFQ1tjMdzPUnC6KHL8VCLQZnI5+SUevWMiARuT6JPy0g544tTOGa
nBnXmAXfVV8I0DH43Frmrvbh7GUpYDb/QD7nQ6UhF4tFZGWGpatJrmyFVmrrttIPfTxCsprlvqJ1
E9hS2YEihIr+eYOXqYP3dC+a5rERyZ5MZHkDYrn2yjuieRMQw2xZ7bcldEDfu2pSYEBPgq47lar0
Z1uzL53mtQd5Sh52CgZIgrb/CreI3phA4Zn2NxTacLyQzeRm4HFzHVlLqmEB8jwM+aSc4/QDPrL2
Yq4bwEVQcKe6wXPbUqTzhchsCFuDcBO8rRhZ5kjmIF6nkfqzJMzJpg13B/VZmTqnheCMspg1xM9P
rh8SUjxj+AiZ42gS27WBk+3fxHofUOgYrlAW+wWPmtFMumtjLRpyYk8PL1l+RtmFPvi7rFB53XUF
0/11PzUIA2VfHajiDAdfSGqiLBz26Fuveca5CM4X6OWMMJowAm0tbLbpq1OlRFUzfrSZ00RUbWdk
yqijEQ1x1KCQD3urYWTorGnTR6z8srzaVw7eGKO4TcASeFghJzD+0TpGgqpu6lvxmvu1XW27Iacg
pd6H20VZLDAYw+II6jHVdNYDm5W9LWX/v8YBBavLN6vTbCD+o1ylIfL7LycmrCBKWKIJpEg9Fm32
vh6R40Rzk3srr1SDYIr4a8aSI1V93HAYrgOWl5nKEpESG2i9PxsmQxEjYIqJnwVSjJGX3qAOPrHW
5+2K89HNVLHh/lx7Rrqr4FVTFfbID4iBm0nih/5E4SOSgl8idg88ojKrV6uzmFNVw45CpmisWLS4
HBR/A9uxNftN1AimKzN3xwNbpa1oEDGWK2m8SxhbD21uxtOP9lNAVVo/eC++0ltfbm3pTU+KP22/
BLnSRRiTE+E/OwED/CDrZ+yssuxXJEgG46mZSimhX2ni6ZfX2w+uIsAsh/xZBOrGiQI1z8OJ7vEG
03zV3Qr9uKMeEvbHYRs7xwB5zmXKQDXenecubKRkFlHHK0act5FYbK7OPJc4Z+fyZprR4La950Ho
L6QfY8mt/nNG9/CLzj0UR8I+K5i/YxsopkniJoFP9l0KhHF1QAWsAl8oNy3kk8CxnbzT2DJbyXMH
R1sdkmbavR4bj/fe5RfQZzz3CID8/0W/nus83zmkMfwExfNVC2SafoWE/mlypWvnCMkbP5qPrfYo
0nbUSohC8mnbu+9mmj3zfDMjv6FAyMsJ0EhQ+FxA5mc6CRogVuUXUGEvWcwW1Vw8Om2M8/MraLDz
kVXk+FGSYAnZGAXqoLfn38EtEx8JOYprdrKQAp6LGubhIpR6477vLjvcI2TmqAEynj6LkasUSm+3
svuqOZCt4ljldna2VQAboiQw7uQ2ob6KL9Dlzj3A578jlAzQ6u1kv0LSLdbWWLmUSJwp/NsJNkHg
avQhDdDDqXSPORpouVanzXEokIZ4UTNAKNsnaK9EybMdGRJFWcnT3H6iRi6BTAG6SMS/yYGtX56X
r52R2b8IK6HgyIpReSEv4Liz5nVz1Ye4ds7dzbIV/Vt0jgVHMZbTliI2MSvadoDvjGXfT+tUxGH7
SbsYlysV3diC0j+ArZm4j9oyI//O0TTb1wSjnF/4oJmI7OPfioI/YtjuGrSKNqN2OlZCX2w8dxgz
Sg9sFhJgqLSgQh8wV4rWXFrJWSnnyGik79pvZLHX5kN3Ufa7GazYuqk/AZgeplVAgDkjyXKphfBx
Noy/zqXFeOwe99S1FteoYFi1roKy8c8KjacU4vP0O/Y0+vXJzOjy0zXKYM91xwfEfKPeFG9+UOG7
dxBH0B0GquNyjBXc/EaHnnj9Afd35ei828UX0vBYbU+Nq/apnp6u9NcTQtWfvZ6axeIlos77rAYZ
NBDakNFKM6rJrae9Q7MxBgvkmFKTZVONCDvsTh4tV4gknUliYHOTNWtl14oO9F/jmhDquIPqXeSV
aBWqZ0PhJunTHjTuDKWT7DKC9f6kw6BMTRCepGwuKL7Dno7UBHTW2Vb/VpIOQfmV3Nl7Rg+70F2M
ig89ok7zjJfqFphQ7fiB8JqEYJZicuQ76ppgtUNMsSU0CKKgCLDWbnjjiCX8hd9a7YnFkYhKoYwW
zuOgJmmtxluQd8whVJA+q/3R8iuZxaGJpbWrnBt1B8q1cbvB4adryDvgkuVb0VsXgjd1a5R1iMH2
ei469L7L5+YAE1UKw3S4yW5XAKbVEu5SofN4C8W8QqIC9A+o8gvAzLzr3/SOdXrv3ef+z/0TfdGv
f1qfJVt1rZk1LnQ5bu/SI9pWClh2N6GW0r+xF0ltqtGclegr1Y8X6npQC8dSZPFxHFO/ANTU8rdO
YX3puPk5t756upRTDlOLT11MjtHfkSXvXTWcUYEuzkMskHA4hFf1gAuStKSvi8p8wv9LXCP+7/Pd
ZwiAuLSIBNFpkuf++8jhlixQvtx3L7djyCqZylWIK8sCtOWTB35DBcc5ZCBNkpzF8OcIo9aPUJ+p
8+EUo78iVWvFZqnW1rP7yLPb55n/VtlrcdUTD7oa6ePBUi+8iD8uDDpTZmS7Fc5/jYbcr42ETKVy
eRJ5E348gxJGuUKDhiFwTmgI0Up7hXJNnZGKd3yCkEueSY06BgU8whk496yKxeBzTqh4U+vmOPYL
iEfTyqS2librBu0zx7Nf8OMXkwMTlrj+YBkuWewVq1wcYFBAET0rbCa4e/unAgSLK67fNtmC4OuX
1Ykz0i30Dv35wyUqoEeHo09rP1ffaUugWbFG23utPJDXtBoXZZHFTnTqyePN0BGi615MvtodRO8e
cYmOOjMDSnf4F8h5zRmhZICwYU/YHmh4PZizf9SY5GSIbRI9U49A4ykKGUGQKpaN0CcKbeLm1Dcd
2t3q3Bsm3d2GtbojKD9mVeeL0pXd4WD6F79SoQrSm45PDtLjyHAgzyDjXMG5cns1sl4+OvOuCr90
PIP4//BETOMc07/WUoOkohGdDWHFhxPonD00nttDefdMzIqOq5Oh29WbHBuck8IaFyrs6f4QFobw
/S3MKsugjcFJLh3gTxxB1GpbXuLgvebmA5r/q/4HIPFw6k1MeOfzuXRDB3aXAH6MtFXfF6Jue9l0
Q2A3Pm3x18OP2enGbQiVpSUkyxQaQRXGIoed0E08TzJmH9UlRRcKPbXD6sxDcIxdGzdnkjt4aM7k
Yt84rHWkLGr4iEgmI5PkgmEzkVZ3m6Tw1djvTSJQIWthKDD0jdK2rD9bA6UC6cpWRN9e87ke/j1F
RZPRJl3IyPVlFkZnI7JesZEHBtfoDX+m4HtqOqWru7j2o3OoN8INFQRvO+FxSMWQsHZUxZeU8Sfb
UJfYvYdEvwm3I+un+dvLb2/2kXU+3VTr22tHYiqgLOmSnCVchpFuCznaB4BVVpj0eALCHz5Jhnam
SKn0wPnyn2A4ukG5vPjXCOvIUJUVgf/hnNLpws78YtliNpmNrqwGE8LmTltdMT9ec+fnLFYffUc3
K6/ufM3E0hOnHA6dFCllL7JmtiiEAjMwZIlddYv9TEuexnmSRsP7eLC5vXM/epvr9Wl8dMgNt1W9
8QRRjGFWlWLHgU3wow7owWQAJHecvlHH7yX7XtlCj15D38Pi8cJ1mKq4JGdyiHBYP1Fw9D4zDsj8
OfmJulmNfgiBxTgkFzlpm4/gEfdi8TKr4krEoVKtiy6mNwsU2RSJ63QM22jTnXvmYGrsp5i9QOLI
/2QGUQyltM/f+Z/44I9hgQ26lnYuZb8mLNj2U48N6Rd/G4SY5d+ufOFqdf3y2npthEvrRkoc4Rik
zHlfo6qB5zdJe9b9Ped3xKXc8eRbfDKPfzvtDLyB0xaoC2WQgoG0YXFG8jYiTJnVaNp9oaTihUub
lWGrWhmbqteHjRFzmAIQau7KSPH84u2HKqPorCP6gW4GVIY5ELleNQjlgrzB1YrnAa1S6Zzojcub
5OX7/rlgzFmBRKmV12gNBPcLT8jJOxqcPVxUucfsN03tP02mbAsmazGtUOQ92pVJTwuG3ZRbwVtH
sx4WVb2iZSdu+mHfKaxsHzqfFvzSFu4EcBiJ1/JdWK75TChz4J/lyCI6k0Ntm9NIPLmfGnK+Y/fc
aIK4/bfd1si6Q5aOulKrb4iGpVl2DWjGYDDa18JoKTyMXLbdJpJBJiJbuqKRZI7u1bvKkTD5ZhF0
FJFGp5YSihneWh0nLCi86ygN+aiznCdjUj6+0dlieVZaasSwKf9Gp4zhyVA3wEP2IkLCMAUQqTIA
eQCFCOImd4gIrvCtpFQVnR6SuPdH9VgGVB6st2yaDhaKKXaw7gLeRZbHrESPohJzTENct045F/RR
TV/KOYDTECMmuhKJ9m9xX/fAmsbL7nSuHBPpGdBwhaxzRsE4RcCFGjLtKX127XhDWs9hwE347SMQ
I5Z1/YiEaHLIhNNzwrvbrAadUdsdgRt2b7XugEpK8Ivyqiq9/9AeLkSoKqDHoZVnOhia61erB9ug
HX6PKtxQwmPtwTQHZAWtdHn8/VKRc5f9F4m4AFWXC0y3ZDGTpVUdqFUcOLfY0Co+xkqcb55+iDVW
Qc8ngueLMfF39uf4jzzBKWb7dZTv1ZqU54aZn8C3VXIWgZUfXaFtsmoHbG9vz/JJq5uZzcG/45mh
xAzMGPxMKmmkeXthrgaRZ1X6UmmxGfQrOTn3diRIHcCDyW6sn8INmYFY0a7TR5mTVURoWZBi7TlS
F40MECZCOwArO7RBtrNaQrD/O2jP2FE5NlagghCv/+Fw3NZw9mVghltpV0sj45wBrULJ8RiOwItI
Q+1AH8HWkOug5letd/MWLJ6zqbeFY6LVbZTE4aJt/uPBxEbiY9KSbpqxtXIEnmrKbH9T74R7HTme
FViEswc05BovRqaMT/uZT/6NEdyPSRhIVMHagW0aJxzCabKs7aRChx1tTu6FH/kE6a79ProdYazU
KOhgytHbkFh2fiKALqmGr+/dcCaVdZ//ZbUD0ie7KH0EK4O0s9V0LgklJOvMELNLo0McffjzMYC5
8gqLqoHom2B7bztTf0mBDu/Zhi5dDC50E9UaHH50cK7cbg8W4sjHtE0HzwxSwDNQHLMWkJWVeo5l
l7an5mWbLMtrSb7WxzdCE3UZL1Hqsvxcek3nNcFsMCWfuXo9i3D3r3HsZitwYfoK8sCNgtIoUU/0
stTpWFG0RhhV8EGiw0iA5MKJQRMHR3OnZefualwMVOWZT2Lv8q3WvNE5Swa/kQMhfegydd+SJV/G
RSOoJLpbAc0fHI4jJWVnNihl1j1ZGfA+3uoPIHFYWTpaJeEBHJP9YEI6T487pghV2dHhGWfwQzKT
KSyTzFMAXWSiMAh4FDaYINv93benXtU9/OwjhcHxCLkcdNaNzyv23ucDJHrgcslJdWknfDwItNkJ
JT2xTnmzSQWs9XQUBqJN2PpaXOyqVtwAp75THxxuYURDQnGW1H7xHxcLaoiJMy3zLVre2iwb6J6P
8ro2R9kL8ldSCwiNXg14TRBQnYoWt8TiTSG0RSWP7tAj05iXWtuuP4ahqgFwKeHE+MOX1O9gY1M6
3poPO/YbkBUSKIp+HK40c7droJA+dzX388p82SMjCfBh4NECcc1O2UiW+YqCgn0CZ9jLHweRRSOi
hvZdRtoZaLq4B1a1c+gdWsQVeEl9AaxuxdNdcN76iMzQxknfHj8Iq+ybhEOEfBqruE16DYqrhNun
koYFS71npIL8GNp6cYbuD6fo5P6jemSUj8/PkAkFF7WlWhr6pnQfJBU5gI5rG2WlLMogl7eCeKnC
gkLOcVkQSIcT2gX4aSNyzfNgCurYVjgEGk263N4PuKIPh1tVEsRD1McvLI2+4V+qAJFpBvUPhWbO
Pe5lbGho1zCT5QHwTOv3hlXlZfU8drtpVomtkRyluCdzIVM2tPY9CEIp3UKLGCnA39qaBRFSenVo
1AXtyG6HF/aVbcvS34hdmEEKmbMmvQuB/OTObLbFKgfnURyeAQv+lBzsP5jG4rmVuIW9MI31Jdus
GPqWUYPLXmCkP41lVTwn0lJxVmKe69YWd6CnHjL4BJkIOYtUtbHnZWXtakwJfxC3joxszZqowBts
FdT0sbNAgh3v9YRTa4acrB2QGWT1XKtkOslIcY64mDtoyfSvVMqqmVmh7yG/CsxuDNBf/GbwB5AW
B/+jxjF/UD+1iqlsAmvQFJNc1aG/aanVYamvUkojgxahA7OJdInxXYflA2oEr1IlMVT/aBZ4Hg31
e1vLiC5n9f64Eyh1YpFyKnjCVH2k8bfjCow5e1A8SqhTBelVwEHsZYVOuueZZanEsmxjT1TtsrZe
aDYDsNqrVYjF8spLxS/GJ2BJwbhjmXbteMFLliU/CxxJ4V2tUFxQ0fXELQO6SUNyHm9e46M/K0Y3
NAJBn7PV5/8vsA7JsqfZzYwMRbgYDLc8UmfB8xd2gge/TSK6uC3F/S+B/H8yuHLDEdBXy36qctz4
eUcq6GsFHefSndpHifJiryVi/xZLpOCAJt4PP13piv1Nh6u96f+yDi+GDF0NFT7qvzEYnhxAxTY3
rVSeL03QXPiCrneZ6GSJhpU4hERklW01ehwO8TZ/DmcS689qfMF8O4On2L5kR8AQvgA+wHybPss4
s5Z0TAlnCWiF5XlQejDSJ31jnvAxiGrfgE08NqsuG852PUurc6qFpEXE21uSdPUdRCYZJAet0ykE
zCTGnxFfyssXvJi24Xt6jmw8W9NtAXh1dCLFjPH0EVCIdlbR0BkhynycfzDqxLEVNLfL3EZpurqc
QmhQZOSmmxJOWKluW3nxLxfgKbeX4rKEDlatmuIG265fLTRSISv7X6k+K6Ws1qjatQyS5q0MjRhJ
POdoqkaNKpAY5NksH2GnALeBHlAfgNI+Fofl4iEm/hXQ0UF0dSfxwDaa/ExzyjC43O8u/GmDEUQ4
tMtXIBKMZXiRzFOoSf59RYEt+59boNkr8EkDz/7ukp1yvlmVscTn1a5SBhM5ZdfsOvIH2p3ounsu
OJTbcnLGbvkOTBX+FO9Eoxpo4QxiPwEkN9ofpviPclD/Nn3IdDESIHwja6RItxtg8UhGPkID6tSp
F82SRW2h6LhAJnWhbnTopuP8cbv6kgLQ/VYr3b5vAt0VrOgZNebHGhWPR64H852m9Ngx/KPMrL2t
ccNQDS2PQUtxloF0F+olnbh+Kh1sFmloVD9dBxNozFBnj1p1UY+VbBKuyp/jtiChrs6idaaBo9ee
uKuAnhCxF7gbjYJwK7cFcpOikGYeYQSG66P37kKR1FvZrt2cjEWqQQWmei56DpcsGABG3AOFW3QU
y3+9OMeLNO+pv282oDZ/0I1ivWbqoxVDb7D4q3d/aR/wTLqs18MvkuxxF7ruM4D3mrrza9g32Un9
Q6Q29ub2Nx6SyQN3TwpxB+a2a/ucioiQLbDIoxXIh+4gUBG8FBRoEuKzLPG2vrGJJ/O7CE67oKaj
zUjbcQTyAlaeK0aTd65CPil4+tOzhR5gEUMXmfmViQTKSpWlCGPSK5a76LoFGGXbIr8PBrgLMMrl
3vYdM9VcMmIsfPySTHKGz91ax20PaglKiGznrZdoMxiHZoXQWdCC2Ka0QzZcrrSV/UUEncJXWfrQ
PWMGJzT3NxzjOyYPoz1TZmVgqija8gXi5yQeVoCAplu4+xQeRlukE+B5QP8BxFwTlx0ZOdb3NGmr
A8SA/SRjl5GI2JtCwgLfDdtrrGEmVsYs18ETd1IpUHCUW4iaInlEWDVz1PnsnO+6CpwkYPGNYosa
2wyFQ5606tQmv3HsHKZV06C+Il/L3d4PLS7TpvWGe3oqf22/jxREA1j2wxoR44SuUy4qAnopWkhe
5EoIaCLoe5HhX1QKPTY1HklUb/xyRhEGScefIdFLB7urAOTgIAkSN+uPjR0358T8Puauux8mUAkq
CdQp9x6lPqtXy93SRPhBp/C9E3QkRLN4q/dsVPy8XpOtpsJ+bkMlNVe3JV60huclx5nZzamqeAGC
hvLgqs1B1SPloxwVtC87eGwv/rTUYMF1aLOTzlpRJ09fLZyAKdoE3c9JkbmM3KGxCShAua/73RKd
ngZ7Shuuo1p8UUCqz3g5FtYbDywLlxJdFDzxaSNOOs+4vtdH9+KNJB5D2DPYDoHPiJcua9wvwAiw
7lxLkrQBcEoW08bc2v07UZP8jnLER3FKUOBrrycmiugDCa+RVaUd68+k5QxcG3c+rNZphzkP5KlP
Yk7hKrxXMnk63dWzzfAZjh1GuKIGWvecAFd1tcfen22smSBhAjjPaufZOjNQxQAYypHsPpR/bSe1
Tc7vs2M9dyw/LMD4sxsPsY1tYpnREkgUMs8PAbiKkpfTjD/I6Wuw2N2QeqJIP4IzgupBrXKPr5nK
LykQM773iGhbOR4qAv4Lk5okqNlCXCt8vS+L7zd20Sv/TdWG38/a4aF2l/WE5vp2Q2r1pXW1VLIx
U+1Pmc7RKAcGVakxMDYmbosHM7gPI+dGPaAxnvc+x5O5oTj4t/z+9xTK66BFM00bvr5DDjSOWW7t
dW6UYr96/Ce2FtFJpkMukPd//gVocS4QRy4wBQc/EDRcCHBitBPJtaqGvT9toN6NiB9GczJYdi3x
4QVi6nYbV7Nz/qPIhocWRYn/Y52DqW+btAGncAEhakNGLyQzj+lrtQfuwNfY8fSy8Ykspz3WupPj
S//pqCMlGzSPtkZqXv1OG4TQfaGNLvg9ascOMGLbLBXLxJvRKp8NRqx9IaDRQW+GZ8Fd7LM9plz0
5TX7V0t2xNvuaOkBB7dycco6uoNN4fc7n62lk/lE5EQGXExzi/GdVX6U1I95ZlBNvTJ6Fg7Gixmr
9hG/FHA5Dn4Pe+HoMJcTYJLZ9kSYYDZ0hcUYYcyGCjjgdsbNWGcF4aCIrnFZ6RLNUGJwbh2FyKcQ
No7Jj8oBZ3yshO9CfTy2DzJ042L6U1eZOmjHp58lkZEbTQybcdiXnplmZUn/wYdF+Jsd+WjyRj9m
EhjgfCq7BEA5xOvdwP3NuO6RUAS+eBfhFI47rZiL7KITqUa/hFLi7rQmPR9Yp2jqWdLEcAvavj61
NFrJaSLVdUs1QUfAMnJ/2qX8MYy6C6sfzkHE7fNmqO6QGoSF/uHgVeglBNkcsv249FXt/hQG0LKY
pA803F2KXufhT2D8CiDRPMxKwB0awpIsFscnnbCVC8SM4AtohOT81+k0vAeYeDSMD7hHxLA4nn4d
UATlSsCHFxbl3Wn9BR7i0PYk4O5nQcLOHNaSxU8eHYPCvVAMy+siAdUV1V5mbsoaiR8euwYxxlRf
2kKMFWlC3+Ow1EId4BXK1WIHlm4jyehS4l3tIhidiivlMTUytYY1rU8w7RKDR9vaJVbgl6HoITlj
JQbASidR9RiQ/m89u5kku/2Mt06ChEpSth5ufEZNxu9DVUFF4Tb8wXhbi99C1Xg5XDCTtCxAUgcR
w97qQdE7wO2afYoLLYQvAzQyzBYEgu3ZpKcgiNfKI1QQeycccdu0zeZT5ruJCQCc0LC77ubTHMW1
Qrx7UYYP/C2P88LaqeZmxUAaqxkjkbOWIQ5vkQXJd84ZpexqYIh8bDahG2sseIck/dSTeD0Syii3
QmIoNuI3PsHM6F+lIQridlZoU9aXFTchDSjg0GgVfCuY3p1taqUpeQ1OrwX91oxgh4NbyyXRUWf0
gDpbUkOnYqgPqgdyHmiSxpczGfyj760CME511u1s49MqxlQ5yIgSQ+N8cS3FNQvkWy2lLYRXZHDE
ZPBir8tL5klEPYFBLCekbtpLQBoZtQN99399mvP8n8JlFt64vlTwJcXqxaPUuLF52sz6KBdPTxLb
jeoReIstGQLKXHbiBwVxOlb7xjTEW0dJQZl6rUmAFEJVkzpDW3X3vFo/mAD3ow/BsOiA6s2przMv
x9rCyONNZDspgzP+Qe4TEyJAxrOOL2d2PhsovYc88/ZYKatHm6ljzTo7BRaZFHxIKCO8CfHkx8NY
mZEbmZGbKKRX7k681YD4IbsWOo0N2EtQWuWnqY1GxENCOuVWpqjHojhTIQge2QCuFmQW/YDjSZgP
j/CPZCAuOEFsGZAoEb0Zb7wdCIyG1v7E7wDU7qmWLiO5bXnM/I9i8FVPTnJY1IVgzc5I+a7UmW3Z
5snu6s9Vg0TZfEwJzwM5tRz9QULILwAV7riBDxmBPwJkX8K7pb9KjAHcJ3aHFZ4WjPJCKRmVXo6E
4Y05OgJLmiwy4HvKbKmvJ6ZX0TRulwIdagtcIefFt2vNTNcX5KUjXSQlb+afSqOS9rjo/fd6bMrY
+KyG5hguKR7gXPz+/1G4XJnFQ9XE2bqLJpTSY9bCY43qCOC9FDU5up7hVfwGu4Hbhz4nlSMgSvd6
ceH3ZK8hoQBLNFdbkm/1dfki3+G8HYyNa7/AjCIVmshf6fPiepYkPZ24pWqio9dF8zCTWLDDJzYc
Wo77tmhdQA566bKSysdTl51mTJcDslPQQzV7tf7at2O9DPCUvHWs/UteWJkj2g/Ok6St8jaS9Z1f
ViHgdR4nlTs2J7GpB32V4nQUHaO6KjYHuWklwCF57PrTDE1cYDMk5KTzZ2APJUM/V+PGyjWopjgU
zd1wGt+kntKxwJwxFX+CIPIihXYL55B4n8l2P9Z+zQzslhQgz0WsCHgiTqPBuIUpD8hymK6cXcuV
sHFQHBvWYrwOuokZxZucGpjC4GGCBeIc2qv9KMAaPrkOYI9j4c+QNCsenx91PYfPgIYxBxpbVLpE
b5nZ3nknm1YVf3LTBTZ1fF1U24FYmnPlPKYVrFtAJD3SZcdjFm5yqzw0sCsl39zhKoL4vCcG+QcI
YxhtjIw3fj6vKNPDcGuoPnmwd6lpj+oc3tEqH7Aqb17vpYF6z9uFPpbbUm/xKKqO/s3ErUG1YC6o
NTc1K3aULpZMRRZLplUPoAkvl+4wxyf1IrfKgshuPlEAcudy3eJ0wTwQPedXUUGPnz1NX0YQY/8I
SXW2kpVhrEY8dEKR6IskXYihoDjCGCh8xTs2aYYP9aj3/NVvOnWwGdqmW6zZ/x80fEqp75hzleaJ
CRqR7AiL6ym4jSsO1gBFkmA9LZgVJ25vQgEljWaI7IFukLDwDIow7f9OAKINSXDqAcQmUl4B+O95
pRKMFsAVeuWZ11cvLMq3V/JrIBrMH/NChySjkAGWimEeOCON/ghq2JhkXmSmLxtUxim8Ou5a2juF
hrPS+eBUJGP385Za02CMTO63E+eldl9cqomUY1EhEz7pc8zIvbq6LlBo/fSE+52imFQz3uBZFlHd
4eGXodytYFFAgFgig1e1xAdv3efSz1i1mBJnLGYE9VkYVp5Uimy9JZRvAJ9I9PK/WoFYMl0FcnI1
RRMJ1fkuUyQyVMvT/uJyzf/p73n7VL8iaszuePfB76LifQ02Fs6AY6T1gC2SSsSWqrzvHQhvcd4n
xA+F61ywjC4I7oKJ2mAMHRae5A2QP5uXt/gE3Y9JD3s+lQxne9Hxb/zS1XN/uLLr5MIinlpsJz5e
56HwzycWuJWe2W35PatlpMtzOa1LV/Ra4QfQTbrSS5sbdV/nAMieiIIxLv6XWI65YCsPOCqPw9aC
lxVy7O6b8wEGinvzK2UW7VyLs2t3SZWLqm5A22N2ETgOfBHDt0o+tlqidtoGjbjJL7E9oYXmMdoE
r5QZVAZrnSDFc2qhEzgnbL9+wV80+W1r8YqlUT/GGEKndSZCEZYEiLLpW1HEI2KSZJr9uDmj727T
Ofj3XR6/nes6Lz3IlHo2sP1CQjz02uBTHlIYxrdthr3Wx24g382IEl0YoqBgFn/nvklWgukdl3TF
kE+oCPHVIBr43Hri8JgXQbdIgbeAp14UXJchQTHXX9J60EMyn0NZ3cH3zFDHRgZT3oKstJQIb4nO
/xLEC86EFbiFlzU8UTr1MU5yzEgHaC7v8wTyb2riLHzG61SkJakpiKniIPtfhd9f74/ErWGm/TxU
9I8V8DX6MUG/y8PqqtldxSpUpZKWvTVy+QcBS6nKByfAwAJsp6qX/h4jryaQ6kgrrzwZpE+P27Wa
FJsmGfbMfkEFf5418Z1th0inWBQTG6JNM/8cjRdu5GpHmOH2BVf/gPJvmlbsxQ82Bnu1ma2iFgkK
Z4/QCt3i4FdNOJpoWkk3u1bnZzDSTV8w3GIZzcDW3JaIKbZLVPmCqXV7HqLR2EXj8SqCeyLY/BiA
3dSiBjB764erqlO7Aeg2/nGTgQQmlq54f6WX69NDuuLVuYZOVpo1BzDkRI5ZnUNIswJK69T5ijio
5JDHBEZSyMsYPDIivj8VTIRgKuJCVSsUp0CWrOkGOd5zJmjrvg392SwleqRxUDwDMIJiWgTYwXyn
Kv5uLm7YulgNb2Q+4OHWILNa7nASqBzO3sQ3VHT259F7ViIKtfRFc+QwI59I78XfbM7JzkamjVWG
n5Rgg+T96LQZ+n8zB1ozLsAuk4bx1YbgzOWKtorRgVRspVPXrjBRJO1T1hVnrtIGntvUzGNeZKbN
O1F8gHPVTBS25FDlFTakPU0Zuu7XwByKOrT/5ikHwiQL29F57OGm1hWwK0w7LLIBRouW/c+mvddJ
rj9QSKLveDcx58JdrcM0oKR61rqigirMn1dSmcc3xFtIMNmlEIahGFNMtXaHqBp+IEimKSJdrZev
JbbUmupGEmnkOcq+2Bfe4WDqTCL8xq814wQkTHCxrudxenjs6PKVc9fseuUrr/DG6vRVG5w3HlXA
AoDinwgeArO8A2PKC4K7zgHO7B3Rrlh6rOJae1H+ZG7llY7AwWwjKh4Ki/WajaluPAyxCMKMQR7C
EZHZ70tyMsbNvxnFso1rYDSOsgggNBI6vGtaOiRXEdkXmZwcGyH65xhjMGVt2EE9CHAdS+aMcSFS
uxSkJlaGZqOFjimcFnFiXaHLVP8EpQITT6+dPKkwUvMufQG7T5bdi4jdelMpuDj3RWdAW9C8722A
sx2/UN+LQK/p78pvOyp8e8f/Z/nABmwHMCI8YDd8FLzyxvh3ToWH1CV5nAZokWDNVcpcSsto6Xcl
1y2I8hXs5ykWO0j3kZoWBDpnRqOr3L1X+26AuD0belHqdlrMkm5WxqKWMwrMih8zKN8TM6djFvB/
hyiMD2viq5XSZq87Ztl9ZjZ08OzwRvpD40CnFbbACVzdyWttk98d0TTwEJrEwHJikAIYApJCdOzt
2GoKjFxT/LGeXpISsr51KRU+zwGYjqLYHUXPtJzgh4gezJb7hL5M8lWbWMPhedyNxBQLcwc/EUS1
1xQsELQU6PXbhgGCjHePQnDmZx4TSP3fb7zwhpcVRewk2LMsI/cAJx+IodG4FOVMp+5XS9w5qfFo
vZ/PvvM3TIrG4W2WsX2ZcdD6dg+Un+tDDiUxf5YD94Laf7JTQbEexptBG4l/fC+AStJ6gPwbzFqL
4TjlLkjGsnA1Urm2YfthBFmzJbfKpPjWZsSTDShXP1vJABspNudMfGmWbnhr0q7aIYE5PAJgLO1l
miaE1/Maxdbcsc/hhDBSa3rO7jN/meQVc7m7ymKZvk24Q3TVvAGxlZ2jQUQe7YLQieQyZmAz9U81
teoGfHE5cdMCLhuhtYP/ZRkaOW8W4jSgjQzcmlrg69w5RNUOaaQK27mKpBub/eMOiHY8iw4oz9Ur
L3hjZc2SNRe2DDDBpdgqnEDA5uDyHsW/oW3+1A2FO8pHgOBFW+B3X7blEawkYOj8qOtVcXB4kMJ2
D/wxy25XtMFYaKzo+kIzyFHZw7JIacUEyvIOEgEuu6lm6IJqxRHQh4cExuf4r4yTj+vPWWbntK2F
eW1p6EiJQRljjCVFdbiKHTzzoEvrjqChrIvjEnNcQGysWK1lciTaXU8jLkCPld32cIuY1/Vnn46p
16BwwCKjfU04+5pJL3sTUywbJnmfEysJbGEvekeiH3BbqJAJ46c6tDKXzRO0MPZyZFCT9uYeKxkV
A14smuNMf72/3odHBrL12MlajgZYylRnwUORVOBLNf/vavPwhRxbe5XbLtQs9shJiXL8Ljwa6pUe
p0oqLlXPsFk9Si+nU3UWNiW2q62s7aUmwjocqF1q8JYjC34BDSEcXv7rl6A9cXGk9lPlDr3QW5iD
MWj0jl5c4RWgRCHwSieXmZnm1ySGV+UdNaAatpvcVRJcKU+xmfJy+RiixOCYRyXuBQhbKIe+vyaJ
eo+tZ6pjFo0dn8GU9g4SGoyycD6TC/ZtH8yqVCeCxzmBWRnSH5l0CFB4yL5YP9n90r+SQDz/v8Na
pqvtW3nIi2EKgYXxNHJNdo0HcoJQjUmWa+tFR8jU8YyivuKNOtqpBxhScUH/lihGSdkso4SP9+uM
gKpWGtQBr63ISvhuJH/pUsz9xpmHOOugUg7tePbB470h05P4JCtQQ7kw/FeEYukbcSDyNOcQ5Ryo
8YO+gzlGIS9d1ZcCoeBWDfqhNMcSpczB9akPZjwlQ9XoHiU8Fw+IjJdGfz2F2ncKdwKKSA9DZpz4
7vlsv1PIbsjlEyb02J4x9jXPCwclpVnQcdidamkx1FVwvDHbMez46IrxrDzb2uzXpss9+0uSccuq
Aksy5vhH4sMofupbgDE8J/o/Xr0XmvClIAre0by6UFgBmf9Sud39NRBn7WE05eyF6rRcBgJ/O6HM
+mmghhORCMhk8RlnhSOrdx8nEr9ZDNCcEY5w8Xj6unQRegViOMcUUYiOsVUv194jINOzyZFeHR5g
KYx0KEa2XUEiamJLKUzNjKH9TWJ2BrJl6/ltuy3fvXJnjaVm1vMDEdo2/d+VEBB2mn/ih1LlOxub
xIDDm9BCJQJ7fZ0zLjj6/2q4NV0G8kDQ7t8Es3yZZW0UzRyFaiAiSvaCJlT9YRz3KsKmkrr8ONol
W9Gu494yRrkEu9ysbGg8ZDe+pwACMdnpgOkIDUgQ7e6t12V3n33ulwU84YUO6J7VJf1N/2SyEq01
AefcE5FOwtKTtUHbH2Ua8kBnJagC7PELKc4tA51ttLG7SY+EyyMEwvBtjA1pjHQb3RdPvPhFvvk4
aVWGmpUhazVhMO8q79X3fcolwjME2emOaa8PJoyUqppPQIKuMYCejKMSVhpLRugGiidIbDJZWBcP
wgYGximgI2BZx6t2JgJMJ/QhGSScDcifpak/54fdVGZNYFgvR31XWVik9wsfp4jkRCOMjrWQnP72
tJdwlq3a2VoUgUyB4QiXWIzpRCmT1QyLExn3OUtmSMqvG5Cm9qBSI794ql9Xx/KlNvv/HpVUHryA
793qt6/S1MpxhnLRESpFgNGECUnbHVR5xoILtn0ED9V8ZKDWaXbzoRzpEIqt3glXG1ju1Kc3Mr3d
sDLvH9B/WG+nXoBrP8cibz5xbSkCR01ck4ZiGBmpWGcjJosyVudB9km1itUxt5nIw1RR7mO5+qGt
NRBwdcvw/ADC4W9oIE1z/wJnJAavje3RhQXgqXJlORpbmhfniXVmFR2g1ofc1z5E8VdNlBP4ng5x
j4jmpRkbEGDOe2X41rnedS9A5m3KLhiqBJJenQeitFJ7G3rPikeqAXHTUdEFsK9UyShByfSS+C9d
FRhMbyf6iTgVqQZ2xFZE+pFurvdKI+b7iRxXVoEMasxXGsFg1wh6iwWj0CSyjh/mjpMVfltq5ULn
lLMVRD/dVxB3WQtS6DXQzVPpwU6rz/SKKDYVHfRRn9aKbTKSr5dekRKeP+/v+hDfEd06ZcXMGJGq
l3hXcuhYIEZsRwuN0157zdey5ueAUwNGZC46OFq+XrsFsDyL0d0rZq7ALCy6gx8SW7RTWMhLnXgE
0HMjvefkob7O9l8eKj3uFU7v3Iwhc9yA5IppOxyUbK9EAt9M4ZbRrqK5HOj4G1FZ0qnclTuQEBn7
jLWUxlMhDMyp5FEX88pM1IzkTpOVAp6m2KytW0E/kkrg+CY6nSTApFIklge2yU4vz5OW7KjRX/V3
bi2bP24AwyH8l8F9i1QO16yjigV0jkwH9HU3AIUU7vIQKD3VpF2PSSR/M3FiU82JLMpUbKgK5Nz9
FTH/4GDHa8+VLb9RMPqwRwayEUXwdaqWd98BbI/k47JOK2zADiWFi4kNeqCPIHX0yHz1cASgTjrr
avhnCflS9iU5+30uoEdOD/fTchDLSj4JR7h2JxZQbmJAw+MyClpn/SJg1bfbL8p5LxJ8YTJgQj7N
MZTDUFVTBrMX2aoyYV0IUYKF3iqlRtBnm5vZiUzCNwGO2jKp5bJcxvzeUuBAqWmEsVCP8g/MnwNy
b5pBeyhMtBwl8xnQoGwFP+3COyaRt1bpaR/P8QIr8W56H6CoL+7fmD3kkYSzQrX5dZRnOPqhXPnO
qaDr22TNgDBYDNi5i4HccnKYPgQSr7cOS4ScLGANa5AfCL4ZbZpvvuf30Y+45DIrH8PEB0XXxuCv
30nmna3Mj0pxdIpnLToaGfYSZItHjE11ihsf7kqhpgcYbWjz1G31XzQUyxKT0hRDYGWePEi1wHt+
k3Pi6QgdelQwU8r6A6slZT+kC7qgMJCTd7QZLvEYfMUyXffooE3tQtjGdCY6wXsXDF2oEaeJ8W9Q
G79SgHCAECBu4gXCx6motJ1FU2/BEX2zsEI6jAfwOH7GNyebdwwBRBB+eVX+g4iHBaysNjFdalW6
d2KsmgqVi2Qa6xfZw4QuDo7zJDG+feC+r7RPbLx0MoGHaiaO1kYXAslF9r9uc7z4K9u05c61xj0s
n2AG4yW1c0SxwiyM6Bs5mJXTwvwgqQJdyDb8+R6r75sYjYXr+WImQZj0/UZACzHTysHxCnJ8kCz7
zr1dst7vijTbwUppYvieeTjZRJp+7AXD9r7qZw2HZH+p+i81XXBpxwPF63hKDSCZ/Leua1AqM/5C
xuUQQTH+4oUTk34G2dFrB6cReLHMBZIj47eOHn4Pt7bg3ULmKCxmaxXB25v3jP5tcgHPIx4mTFan
4BCWRYT9v8J/OigxXVMEH6clCPVQeiKn1YB6DqP4yuMYySTsl3MBO4paaePTySkoy7R4PS6JQjvc
OPfotNhQwB/7Q7kW5vEpGGbPcXdyGpXSFktlhQje5RyMfsW9H7Oegp3106CLNjW/r9LFPmcPm1K3
pw7HIC3EDFi07hn418HeCSxp8F94hTVF0F3CA5d2Tt3VBze6qi/cT45bvLXOoe3b3yIUtBYhyzIc
eZSRbhFD5n1QdPxqyMUM6+GpanFfBEUgtJkzbmxBlA0RjM3lsE0PRd374v7QXXN97AUMVHoBqF4W
E4SEoAAPo0LqSeiZdqptygQVKqdj/9zhQXBdya/mMaP4327uwN1lbnRh7SPUhipRDXTyMits/eY3
dmffNtrTl/1ycAwrDNK3ET2/aS22/ER4XGBIKwGf6ep45RtSjzpkrRs+oR94GRWR8pDJlpG/hmKx
oS57jV0TooQ95ujr022JtgBk+E+S7QFh1WK5L1tNMCSaOAzRioymgBUD8DTGej1lT2bokgrvARNy
NfbNhfLrAxdqEJJe6iQKIMZp2RqfX4Dtjw5qd2wJmoqYh4MVSIbrCmoWG5rIFzZvcpx6sHNX3e/R
F8xDxYb7s46A7elmbyU/G+rQL6tsFCRMhfPhQYaLIl6VQqMKYaze5XT7kv26CD4R4Uo5l4MVYiel
SV1Q2A9hSSu8NMH1HLQ7f9DRYQmU2R+gbdFM5+jWZzKU8OIe8SWv9Jc4ZtZRPWgCO2Je7PTVWb+V
s+wDtqX+xpuwCOj1tOTP3g33fHC3CSTTjFk1lPlTs39rotVitO+YzxvNZjk7899zExeKlvMed1Yk
zdM8PZSPZCQX3X0JXo+B/5u/4TCPdrfkOGt1GkKk/VXeno+QHmjbcHFDe0z9QcA68o5EmZccSTBS
vwu36gAfW00yE6VCnG1kcn5g6qcz/d9Rxi9kjqB+MiJvaOldOBYoNlUN5XKlNeJvbxxO2O9nj+Zo
m/P3I7DXm+wwgnZXO2DQME3QXG6L+MoZqB49KB1Trn5/XL0cRc37QInjVY/CIKiZsx1gjtnx8tIx
2j2Jwo9RihlvmvwaO39VtWEElWExItBvtJky0SUrOt9zX7hb+s5Wrz4ihcL/VlIVdc7z3sNBV2KT
UKIb3Gi4Ycj1EfrYMS4L5hVe30rnD6JX7qkohpdbVWWkOmakj8sTSgvh0dqnNlQH3E6VjHQUVbSq
XLpmgIDjziGwB6Alx4onPTPddjkOXqf+s2aHOQnlIDzkvuBnJDLtNSONTSjU5Djs6rgIMMX4H5sQ
YJrC2/2e24l9pKnwGvHtZSU5kwOUPX3xsXBKzf89Whs2Pk8c7UW5cK2m39eglsBb+3+HD1pczQTJ
vnE9wl9JTwRoBmMTHK0EETcNB0ZfRyPsfEI7zWvVeiXQC80EkU52e76aNZABlBHhZG1TOKmGovFC
HvN6g15/Nql6Hdsx9wVak5dgD0z6CgpDKNCz9b9gmG+fgUzqNefIY9vPX9UxMGHwh2fsp89uTKee
4orEWb5JpF2GbR9OyKJMhax3nhqdgp4xlucVIuobNimGQ3J3INMyzPK7DsKNj7BjzRbOzE6Z2Os8
e5P+xRL8uIdVM9EeL3d0s98leYHOGUHQ1FMYjXtT+PLIHfkfliK68c4slmh+53+oKreoQ17tddRI
CpMer26978qIBgSWS3rTvbyY5KIgYitza23QM77Fde/u0GGvcervIIsQe24l6gRFYny7VuyorFka
W+UH/KWb4ybxXSOfMScteUjqyp+1f+TQfQr1uE1sregNGcco18XcDt3fuPQHA7v7ifZJM9Mtg3SN
U/duNmUcnUpxw3RSjM5kIXfQDE4KHKTR/a0hMpfk2vBz7eA6FZJTECc/8jDhpxFhuDo02jf+2LM+
6TmpTmDQtQzLo75MO8kleACjxPsDbapA3f8UmaFiZ3ElmTmlVqYI8wGwgeDLpfp9UiF48MhhwgNo
8s8nXarYcJ48dN82wkYnSQdx9rAstok3D5cW1pBllaAwpkza5U4C32xPNSdjxJV7CktfZfWDEbM6
lCN72UDnMk0wpACzu/ZDUoG52KJxSaoFaefv3dk1kQqYSILJCZZj8n9jTQEXCF3ktWoiNmk7DXhK
WR/SS++6awRkgcL4E36M2aGPgye2MnmrDKYjpUiSy34DsW1wl2h8egZ4wZkFAmRISgAuh4TaOcYC
5vocWbDhf+ojIRmMKYMP4DTDpZO1/8RAI7TrMSTX+dgMYvtUh7jz7htkX/qqCT0T1yVrkeRpioWJ
b79dnx8Zyowx9MPxuw3LmjqK4sGtjyoP+twq3Cr4+ipD609PlHGyS/7ZvXn6lhB+xcES3GfUzKca
g6gpF65q9xMMehiAge+/5xwsZg4CVhvBLCFRRsO1GSv2uY44GeSaiSEVa+2YL/fHfuZ2WB2xjKP0
edBq5Cj4E6Q70+5dpgtXsCH6lZdFF24Rp866XO/9MkHvfkmOBb6QexEb748ZjFJGkmqcsu75czVc
6HLuaWmtjKlKAXHqjOkKgatx+1h5paloBU+Sr9eWZo83c21Eypl6SRC8p3P4hOy85H3DcVMDMU5n
xMGFqFQNMyw29s5ZODJYJGKOTQwY5d5+6UwCHExYeQ5aTbeIv2ryNjZUbzDqRtdovDne6YUactRm
LRSCu9VaTbPlzPIUK3l2zhO425bpkIbt9OSIFVtuSY/cNKlWBFxp2aO13lEDRfGMhmmmEUauDrjW
nIXrumcfqlB/WdepajKdGI8wMBBtizkgN9cVnhnUT+Q6b1Z0MCGzhnT1/C0lm411CFU4b8mmoItI
7XZGPVmM617079ByyQ3K+ysJkN0f3dWwT+XwVnx3F+7gsbi6BMdvOGLz/aRLK73KgqFPn3UnEMf+
uRnwts1V0hVvEuhEnbTO9VF43HHDZ4CYyQUhl5fgu2HQ5gcErXN0u4lGvRHf9HRY1lvk2HHsVfCJ
13K020WfKc3m+zYVvuvy8c50JzlfwiUmfZI6Ni0SE+eMAT/TIupCuO34GoSXWy3GmkbqphxwsXjg
bbdBvFqIiHwW+2G2G4rxj3bZSufb3fatwFbPgNX8dANq0uEuj0n3L4R4t4DdrVAq4dYiqrRu9ZTi
t2CiiTj1FgviOY2gLqs4qo6i9BSEDbHaRqWrWzNO3cUk0/cDgvvGrd8AkCeyeFkGX2Gtx+bQzTj3
c2TW5y4an7k8uTcC/f5YZrw3+Q7WcZPpdYyX263oWtAynST08bPvWZmyJNZonJQfNoFbWP6HwQlE
mFzaaEwyG5v6JYy+Prm82xVzk+JK2ZskAx0BDAOwxyd6U1Q2WiDlHeY6LUNFs3i101+u2QzRH+bi
dcAA1veWzpkP9Og2aTzejj8ZUop+oN+3zuwqrRzKtAdXOhSFMelE0mcNpe2WWGZhgZAsZJODoCm8
oohYzo8lNgLGR5rY0aOz4kNCpRbHlA16kcF34Jzqop5aUyskETclBVGdhXMhW5H75T3Ds/YlIHx+
nt9m/c+S/UkaZdgtJhfKVY6htoIbuOGBxFVOWGvTfx2FiP6crFGLGxD4onTFkbgGtAyyMb9krlqJ
2oM3FoPUWs/t2UhRut9CkheEX7r4ieDgfyy6q3Z7bgSIYqEvkR/2gRvvxbcMXKbWAcnnaI2Ufl0G
BKKEhwWMe9u0f8D2VjK6w6k7sBMmAXIstg12asXHQ2Do4hpoidBY3ARHpYDjDHRwCCMe1x82PuZH
BZh4ZRB95UWeQM2GR5FapF4upRBNWJfl83dYrHBK0NUm6H+ydQVBUfuGRvzBwocepnhCUYaTbB8g
P27SLA0TE19NIkub6sra3oaPVXbg/TbiOvyq6dkCRjNT5pUuqqbmg3VExB99ecNrPHX+aiiDxuw1
U6h9KKr2pjSOTQ9UpZNUaGa8QwhE78JeshUkr574BO99npiBmckleOKqMF01Yks/5KAklkt90JUK
AXK5muneQSK9rEueho+AH1iQk9EWsS3S3hXxeYKxFVGgBY7iY+8Wxid1FUcwkntP829yo6eFwfI9
yS05E74A6hH9INMijfJqMumGKo3GzpoSvy2/vj/bai9szU/qWs4KknvkVBjT9jBumGx1f1ECcv1L
BHP7PO+NwZxJ0ho4wT5PqDzvA8BwOybA0uTRJf/8hzTUtFOU040vDKJOTptJRQDocLJAUK+oSdIB
1smbrzmJZ56NyA4A8f0UdrPYHgzbHNmrdjlZX9UAo6bTJRCpIP7AIaEDXYXJd1jPJsmHG1zTo32M
cDch+sWg4q/EbjVTSGQ5QnNnp1/ctm0AM6dHeplajGYgab1K3VssoNxaQAEVOvCQRNwsT3NcybpJ
u0cRKPvgUQ6J4Q1riyWyd9ZuCvPtZdPrCx2J4wuuwx3gJf1STBRuS3776yKBuc8k7qNm55pbBPGb
qQsWb8zt/LNG4XvFSwAtEEakFsJtjViXBVrwblG1gXKBL9tdY6tjKgAG8RBZo8loSfy8HTMWcPuz
ojQpBRtcwLiaOVqSOd3UxzRpCbXiSf2q99Uy6tGIdIQI0Ls8EEDLNi43/CoJ2+OORdWgN5Nbw8BB
0IHNhcXF8A07PEbCOnOP8aNjSNajIkralwmIvMiSiDjI+8xwohHuNtB+HF8x4tcdmut1XrG5BanS
BrA5LRBHYGILm899sKe/MyXjUeXj8bkDQm5i1aviPCGXmm9BiY7cF2xETvdtA82gdfwNiDUIWeOF
eG85zGQdFI2nAOJjF6o8xGjGXMRDHeWbtUToJhN2nA680PwwZaNCnpM2N3bF6FnCgaGWqXCsXenj
pnFL4TAV0S1wF+tzeARdQ/ud5d3+lkvZIfGZaoUadCaeqWV4/oHfwJDUjaiB3CdQSn+RNv1/5/+g
YnfGPXGcitU87DpTOQLCJ6j3IroQwjobLAPilwpdlgsQUofPPrKwysj+C0UsRAlpFnd2l84pcWyf
VQjd3pL8aWsveKwk6cOCswo1YPWrp/3Ckbv0Aq/iyqI95uaLGJYYqmtsjEkaowO5mYTC34uJ6Aes
MGb8sFJ9U16N8pQRTkepSy/XXIsMLdz71e6ZgKHPjzFx5GDY3OHCjffhOTSi2400IeDLYi1cdt0B
D+OYo60HFhTxGYhixa3JeloEcDCxG7fXf5aZ+1ZVE0tKCrWPOIwqFWOvxCNjyXNMLzKz0Ej1LtgS
zoPvzcOiKRWeNIAR0l0Me5lrx1iS4mxeA43iDHeD+lV8YexJUnPDgLP8zpUjl5lh1nUlOZQltSy6
ATl2b6IULZ+qvPGMkrzM39dDpRpUJgJZxU1VOornjpojaZ/pmp9PS+WJi+WUKp99aR8tk9URzL/v
pHYczITL28seTA7w864/l0XBgSD280JW/P/7SC6QLL8BvG6ItiBEvZpeim2zyxCFwX+Ucx1NXs+c
MducacpY1yULtu9D0IOQPRP4miadM1/nm1+Di4fR+50suiMX09LpOeJVdwiEO4aqec0nBbdyXP6I
Gs3UoJdX18iwEYSEtUZvBnZXUiAoFl6yWlRrhWKprkl3o1ySjoPy892FJO9FyRF+VUw6vbS56r9c
DZS87ndrBwhno7K70TfBMMoJU5PaCqM2kesWsLkYWrFG72UJE8s26qRJLMotlwbwJp8XCIJrvye3
iJq+gfc02R4o3hdSNQUF+AuuFNY1vAt8xETL+6uKLqfLQ4OaLaClFSvWcSGh3UB9GDdui7LZUoAn
rMRH+sPlNbl0KHatvY94j59uzZMZe7UT3Qgh4I+EqIHJXeOtpn4w5JVEURg5d92KxDisU9RCSk6b
gNgXwY93yFESOXWU3tk46qKAJyM70sxIXfGFR+meVwxtt48q4BEU73pQYkLDbg3UaFuQqkiV4WxN
sD/yW3O0s9ix5pNEtE39jxJG7ZToQiq+XoGn3IWEJCfBPcLdEHW3z/F1PFh+OLkgDuA3zW7NuNOJ
2c+gXuHjSDUZv1U89m6DSp0EG73E+uARAeyKqW5VnQmmtcOLd1JZjGANh6nf6FFLS/kvptF3tgr2
QK77nob5/KcKCUqSs5xB9q90m20ESmyXhWLiRn4ee33neC1eU0t+MLaAHsoZ1iNQqzz0JCraXq9k
nPqaHCygjGhpiwzYfWL4l0ucmY9hwr+uZMbKv11X5UG4JDp/9IbGTG8ZPLHuqXw5KMqmhhfgLAod
RsNbO6P/fnE5j6WswSfn8b9ya7wf/759GjzrQUT77V3J1hrO1JpduOMWp7vG2Rnib+qh+CD2xT0v
Xkv9++UJkWaJVSizEGpRTvV7L59QAn7+9cVV9xaBQYR5mWYytCpy+435PTK4PocgqA9IiRoayQAg
4lbb2Rj+bgB81QnUFpmtl0c+2FfBn3WQHb0Ha1AVl8NvppOZv81+xYllBVVtRnBo8xqBTDADxxBZ
43z/BNzmbrnFeTCyQUBI+RO0KJu53a8RBP17lWb3oJSJE00XPzhcOjBjSCC9eW2yRxyklDJPqJWb
3HagXBNpB3LCUhy/9qVTA1eY2KnAUXYMRkkeJtFGnRworYyk9uyLedqZSQrRD1V4O3Uf7IwiGo8W
10CXv4XfmQ9zr5fo5TOSy6tlL2AY+/QYxoZP11ymxbM84oy2L7LsHBFZOU7YTcGncTlQoYN6Y1LG
hrekF9jmCgAmbAu+tJNJroftt1NHy/AjulkSQZQ386ihYFDJWQv8cgX7fzUqmo2C1QcwObb5rRfs
fywLtLgapQhRhoJNXzpmP2XR9w5RrwxmJVqu9UMndWNCDcW8WlMHSdKQtlMl5RA9Sg7P8Fx19ReV
vM2GQLhLREvJ5FY20tRkDTEYMfKrIVqBrTrVjeq21yfPNzX5tzZHyenZEw+Lr/uSE6kV4/Ac76y9
Eu+9DkhESG4AL8W+1g1zmLrGuGoAYI66NVeG+EC1ZkgO0HyFHSbDwvZ02PDcdNAqNMlxnMOH7Lyy
gbzqdLg3GEB/oqYrQvMi9CDVfYsXxYFArELcnD27+bi4CepNR/+xDlQXGQYDT6aUTJ3D5leOj4RI
Z7dHFw6IOxlpFNztwL0yXfuM/wNWNykoSiL6WxHzxzxJiT11j+lbwYrLD8GQ2rYJTnsIhS9A0l7p
NbuRbsooTpNLcg5BoLNkvdUzSkIyPSQkQdne/3foNEnYyFHXiBgznUXS/m7QZnDdlxouqOQ4SuK4
Y+g2BVby9oirgUnHOeTHP6Reh4+jGl8Rpfn7FZPgkz2bbIpKvZxLiKuUuRDVJDCj/bNfymNvm3r5
AZSaKxwjqylLSLYtGix9HWTMuyReYwW9/0glWTmrFM46thqDPnJc4yHs/N3eFATDG4immNkQLiV9
PyjwCuqGAJoo3h8h9KSml9OAV8PfJZiOQczU8j4K0u+zJkw6PJAQEUUfzil5jLstWpWDievtSdZd
6R1N8fbfRAgbLHfP+S533cWb3zl2D4RCuTpnxzh+KY2mceErmrRmMiYecdj61Bh1uWdZYfidrQ+5
ydY61wJamYO7AIol/jNGE8FodqMhbiTeYIcf6UNWM69ciROqRvwu2rAA9fwvoIn97hgS+JBU8ygr
RwsD6vgMfylU6VP71+mBvygxV2vTxJhkzdH4n5fQk/pl7ilkZtDDonr1agetvZI0gFJrwV4Pm7sF
dSZ/YLiYTfk01Eq6ALexxeJbLdpbvwwqEbcHMQNTF3iO4dX9BLd5hK66nynCKYMSlKSDmDYUbhk0
+8yLE2OVzVNG4q9Zqr/PTMj/7yyZN2TReEndDBYjjY2Hk75bYHsvU1O/h+r9NoxF6QP8TFvfSI11
YZDZrSc7TL6IBMk2kOJdHVezb1pH2ONBSqAxoME4MkH5agspp29mX/5dwX4WYBT5uT0UTisCC8Q9
4FbykdjDNDRLzmXEtE0fD7sSb1UKmxLRFGluBwiaxCrnz/BK5UrSiLdHd89gmuIeKvBR9grH7Mod
KtpUOdLGBuJvwt3Vcc5yQ8+KujYkmZdGMmPlAs0dr2YY5LySaMywniSeaTHoaHI4BPDi24zTgsoA
duS44oIFaNoQuyDOygqDUgw0phrHNzh8YZFmWH+kLMXAchvzl20ACDmSEOKB/s+lr9iqawZcsoQo
mqqRnD+Y1SiUaUe0MCMqLpl1mFbfGtbonhXkaomjHzup17ZopumDvdpLvgTSrsOc3ACdh9r6UP4b
6ElfCKncWTsXy8cSPHNERtUk9euvvUyYVCI/byZ47qvkHFj0OlygM1+3rgIC4bw4ThfKwq73L5Qb
S4Xbp3UiW0ABXNGO6c21loqjE51eVpUur3WlB55ZMEyau6eRIBfQDNPq2cmja7wkdHWpfxP3uAxd
ul8q4xNUIWyhtdey51W3845Mur3hOn1641RQj7KrlXSwxJHfj1aITaI/mD63QnnpFJFwUQltxd0D
/3ISZysXZfv6Y7lzb/72x2n6H2gr+gepm+o/AX6ZFU1znrWc9f4bhtGQJpeMmj/gRbs+pKvfsL4O
00ykJL27njMw+TV6SCWirRBK7eOpZyjwoFXK3uy5vARwXfqj6TQIUCFmRsUttkC8lF8I3XcbNCMp
JxxeJd0P6akzqR2u3GRcHHMqi5X2CNwTtABZrgyfswEPwvl7NAYH2g0YHh0swnOqnmOI6kp+LCeX
BgN4HhBHzg0OmBvZk7WBNAw2Qyw887HgwVsb0xYI0FY8dDdjgybJGzbL3LEpMFEHyr/ja8Hrixda
4O99fhvoo0wb0weY03bQkYnBkmPcqwjIosuxIMi424/3J7IK0hDAcyJe4aBk+L0qbAxlGgnEaTFL
8oroSSPNNSBYKCMQ72j9glfFW98a2qK7aT5ki9udgkT4GHAvjFiPFHTmVcuz0tg70fVPsBW9qzT1
ywvhmleK7UsiyLy5QYdh91zT+EYu7twFPaaqc3OGPpLJUqr5cvBUfjB/h7IMdB3m8VtVLRZDL6rn
ZFNP4zpSQRWQplVOU7ZsAlcxkfAOcsYCjjP8sDj1BQ8BSWCfQaDj/79zAD1PphELrlJ4PXPRz6q2
EN60S7aqdkD9rOBuewn7E2wv3TlH2K4Cy2PVVovV2y8yT2rk/RBP1xW9GgJbl3u23J5vsBMH7NSd
Cw3R4F2u4RlFA2ynJPttEb2ZKAngOnTzF9FmIuDAuP+Tk+I9qKlioQv9VYUcpTe8LqvtztNj2t4V
nH/Rvpl7ZDF2vvZ41PhNKqh3TgfY3vX4CTH6fZ9JDfMi7Ia6HEGK5jNSCsxNGMUzHSlsxhSsJwdL
K98TXONNXMdhxgXOJW+3mVFOsSZ64/gKyQkqVKrZCaC8xbvB96g8+QC5KHrH2nvyio3XIREEp1i9
+UJeoKNwrAiMsbAYt27pSVVwUsqoUr8NQ+XOGvMa0fu7QEfoRNeFNlFO+1ZEG2vP8er8U14H91xX
l+jHCuSR+NugnRs6zRjUBHZX3x2Eqfa2N17oiLQrwWCdpxCPBxorPSUEwf7CbKoBMI6bnCNLU82c
ZL9hFLxqlepAgjJMtHFLXTcdqgo5k2flTqb5DyaPt+zCuWa/FaHfefkBnLxtLM9QqHbMfCPv5yjA
sOSPc3Tr/OghxwGFScza8KmyiN+EebnmYgrluzeEjnOrXc0Abvju7no/vxBpEiWZRVGQwf6oMkaY
vH0XdVPWgnYk4zZioI9lCOiCEKpc24pbzINqmJpkSLYgk/uVp4tqppItKju7O8tjosy//GaEeaMN
vHG9AAYNdRHbpa1b6WArzS15tAT1M4DW+wSqmnxjG/HF0q25QC0kdNglx/fHUCsnGQqMHvj/CHCh
cFGQVmmukfVpTm45OJN+bIoao626crmcFpxhMf17h9wZO2O9uJQx83luXo6DWO/Vp+pWflQs7lWq
G3l93QsTEfI1vT6itoUMQ+sNsK7ZEgs0JIN/GvkTrH3YwlpOo41u9plerQHXVPu0W6SktF9Isi9i
zTEctdnyT91Gbmc0aP24dPjUTGtQOXjqpM9fhqlXj0Tm2woQp61g2jAxiMvWOuPhofqNFNwMB3Rm
Bxa/yBHqsvSjWcWfAlQ7426VxnJlqGTfFAHzBxFidt7R93PEJXvf5F5ClTBu2bI3yJzENC0mefYQ
wNyihtrCWRhJ0qqY2WyqSboMucYQey/udEBSAL7QltVlSwPl04MD1xWjrO1Kc5e0dSzVFcU3nYB/
wTIz3hHv4fVJNEfqqzYMf4CgkcR+3p7l07h6WTPbcOvnEqwXNnDNo2V0y9Cgii3h+Ed8fCrVzne5
cNAk3299SNxDF2kUEZnLgT0wHzPoYdq/QVV4XO7iYMy/3WzRKZfBQiZzYXeSGQlzPI3jzEdkt8i7
GGZSCBRNILe6a3C+GxOIllm6DWVAufvhDHa3P440kWoq2iYyiQYENUHP4gdjgbVfPbCXO8E2Dxg7
ALj+XSE9pSk6sm2qDL9SmQjGX36cqH1000gkkTaQiLVcCUM4OOSdmA8ytax8bqu5xt6+squV1gCn
OhqHoPRto1jGgTgmQ86Wy8vKZoNYpIeC3XUnzlGuTaFL0oasDlV6JUCxTouRnPNO6kvOkRebTKa8
ZTtQHQm2v1HqRD4LeNevMhqQWfJ3sP2wY0u2uXCHAn19Idn8BICfTlSb9C/OwVS3j5Av4rtpz1FV
zZ/SAKwUrobLXpPIazr0zrFTJwIN5NSfJpepQmvXYDjJo6RF8eIEjTfzERTKm1fAeDMpUKaqjv3H
8wRed+Y3f2kpVg6rLQpdlvKiiZ4cDfRqgRFr++MnmMM9J5nyFL1dfg/6Gfq116/RKCDZe5Qr6lj0
YTd0x1cAJjCvi5S7mr0JkOrwgBPlLOLILYWAnKUzKR6oEE9MtLQ0BWMKFR8Qbwcc/yHLT15CxGC5
tv9xb/a7vaA6ATXb3Tzur6EcMl2pw7I4mjioiof7BYjI69Q9LkT/x9PlsVDm11r0ZNObrBi19B+f
KAvcjUvy1y0jyH8dU3YIAc+Koo7YHPFqKHIFXtteNPVVLoFv7CvBeoIaHs/4dpsvJDwJwHxdLzub
8BQ9oy+UnTDe5dLZKEPltyoQZ3qhdXKlLkEhzMtFAKsdkkqWou6jpp77PxEHpVcgr8MPe//voJvE
/ky8kvWiqsPGGVf3PB/UoSvzV8XpTLuc6tQcaA32zbRU1aN118CYM95Ewj3BctNgXfvskWVj7zsC
0ZN8T/dqFj629Glb3AAKWn/3p+MIROMTWpOA2ej75r7FIyiZI6V5nviIXA34tPDHO67B85/vFUpN
WYxPaRb0P2r+jagj0qlMsiOomt1xcmpAy8GXqQYiwpIad373SjgK6VtuHeA0lqyQ++vZ1m3R29No
x/SPWjYjsdwJJvEdTnSjnQ5XfuYhP+LeZy8PZnNGxVQRtumUlbdYo4zAaNSSvKMe3bVPKnEquJSx
cByRA+gm7CYstnbaHur5oDNzL1f2WgqDUNNqNZ+Iw0GzQzL53DjT0YPmigy9T8PgA3cpFxR03/D+
aIznanb62JWEjPtndcOayh9N1+JlCAaK/pmJxpkF15+jJyipFzGMwhsQB6QtB+cmFV3EilKyV1Bz
cvl0Oq/EZC3pqrOGnSBXYZcDI7ahWbov/9YCdlhuw+tyxlqfWzrpwZOObhalkg8ZJPyRxVLDQkPk
TVPbYosCwc9hdLBOvXikMW47BwaglX2D3WgW00coGlPZVcML/gYHGDvgIxxH9VnvyQ1evP67xIUI
5XZD7Oo2N8ipmAcQSn1PS6XSJLXCR03JwNYMGmP1Lvye+4gKMGIKi3ubH1zsBs6fsxgHJ7shRMFw
5cMGDPqTaxMjJJIMQZstxheBLigBApIgwQFtsoaJW93w3hDzQtw78zVgduKU3Fqs+sDqrUGrg2rl
kXOfSOJhJvPcmE2VV7PoOtN8k10X7YY4chnuecJvic5oB5ZcfjGU8VNWMvnYzMIA6HGPF8lZmv6A
xEKKjuk1xQWpalECfnefjvBolNbeZa+ymoKyeXr7cCArIA43E8UMToPPpxiEtwjKRpuEBKhYZXu1
Omk/rNxD0eYswdAYbYKVNUOeHF10SzArfLFj7lq9l9R201n2I10l4cubGrFTbs71f7hXYxErOUD9
j+IFAjGrfF1SOmgIVY89ji4GZn8oBmGnQcYw4pn95Z0z734MyJndtzmWZB7ghEQsm4Z6Mwn5lxX0
WmNFWQXmPlWjZJ8D9tCG+PyuOS2rrhnW4IR1TM+oupser6X2tYakqJbcxinMwV3gRiwK6wsu0KXd
A3kgQMsxxqjPeyxKCHDyc2r0WaoRkDtvZrK2O1f0a/VbiPg4/OIIZFWZ1Kawc1yOv0gp3sxzLJI1
Lob9huIOlY1QZawV0wuMLIoqqF4kQnRSOUg8tM1PLisEtjh7AkkwTCTG5ePvq2cS1pvYw+nxE7mD
WprjrCM+B4jfYCveiESxRGtDVAYG2Lo3/NmYqh0nzbw2bV46HS65o621Vm1Y5n5sz9Dav97WEP/Q
inpSo2nuO8QU5Dn3Q5DoOh2o+eiaFQRQXxBSxo7r37o1u67JQuBUUfZkMTMD5HdWFsqqN2Uo9KII
WfcRUNb6ZqEcA+tFDznJE+Bpw8RyobBlj7dTpvjgKv5pxPqR7y2QSRipuzWSUcbFP7YvW3ReTNL6
IyaYUldsxSSN1ngwa8l67rzUb3gnpXx8OM/1Tvf9kdlPABZ1kMfcZ+omtnXH0GwhKsYnjLCxAZRN
81c4/SfZNR4GNfMgiMXV8+3HGdj49UU4fDWpOaAwpsa9FaXclrp5lOV+jOlTuvFb4vp8gu6CKLQa
5ZCCipbMCCJEmVMwOjhl9fQwgfqgbFk6jnSKBbjpR4aqS9l/OwKldz3JTaS+mfv01vW+2vyfIk7B
NaFxTL0Z1xdMOMdtzymfW9cmuFDblF3Zh37txs49plUC2ooGKYMiY6o5/JPhR3FYzXduq8cb6xGu
CHK7TrEyV8T+0btCmJxtT4in5t6pMegyq7sq1ZD+aAMC9XVunCfBW/Y9keHC2DZRcTRRANZh+gI2
FFnm9/CxdQnTImRBMq9+jwqwjLJFcQAC/cWuDyhxQOaNBla4I5XyIS1QKirWfSfILDf1w/UL7ztE
yBnd/eQp4RuGezdiHvl3RFIq14nRlJonH1TkPQJpf9FjhhX9Ha9TTRt7vdtnhO1BpdH3yhcIVHIa
dax0BW2FZvS2/OKdItXgO+LbnsU05c9l2//In8YY9qS065/ZAc+2i41brid8QfZDuWAkJTm+KCCG
BL2Z84rQ/S5E3USWmhViqMclvmxnzVlPZses1SjNLAOUVPU5tKO1UeCQBYfvOJZehOSBJSU4+GzM
P62LnRXS/Muft0Y/pEKvz6gQ8e1orTGTa/08h0AD3cDNVJSLXEhFtFF+FrlJhtwd3tVNsjNuTDrj
wWYj8rOVm/obfoG8qlkCrAzUMHKAvzxz831XjC9eC06s1OgLYNWZEYJ6AVOyM0KqQdxXFXEb5ZkE
bsmlSmTSIaDCV4uows28ObALjng1s9mz+KBa8HJtSYpWwBB3wP2VARg0ForGlwkHGRsg396qnIsK
BuPrnJNwy4LkneRF0p2UpjfHjS7mmWbicn8oYh8n8mS/maH+CFPPiHsE3ZGrdAxMO0Y0H2A+vj4v
gvahdqyfNKp/GIFEPh8rVPDJDdOlF/P6cO5nEDVrvQHWvrrIyLixnpGVE9DSTl0uuDZEwWZUy4Xc
CbTANkoryTPtJdRV9cOTRno8kyysE9pQjDfcpZP8rageTg/9DKYCcyCU8vljrm35/vVV4ebhwjJB
IQW1GBEdtCsGCYjvNcJPT2E+a75ShPPd9dcC3KN4ecqJ1KpsDFncYZixeIvNz9JR/c0HphthD8Nz
1PdONluY10qadRRMrKLL1hZB57ZBNniX2RB9YKmOb6O9FRvfP6Sl5pJGDZXB3z3gPPPHH+WTB7Xr
ZKqznOCZFIeVT9kTvzyuf3G1CujkHE3WMIuCHqllso65jWgh88fn8WDlzC3BtKTcH28kUnhVJZEf
encpJSD9Bk737CyaZiDz7E1bqwO2O1IvXAaozmRotXCZ8/+RJQvR/GxPbNYOAVoBNpW9qVb0d2+u
JVWnsy+zmDDUMSp/Pkt0nyNFzEkzUIknr+Blf61rIaCWbkJr7qHNZMqrK9uxjVgpfnzABPd8oT6x
wiG7wQdDrz5HMLO7KA8WhWgPBnev+jVMqqHAKRVypf0c3tiAj9Z8WWFqmh/7v3T9sjeFfd6i+Phn
Ce0h068avzDm0MRtoHutCB/FiOdhTaMTrQWlnX7AyiGc6Rq4GvwoiINLPS6BFLhEJoVMjA0HqF/c
uQYf+KK/YUPSVOB15WNjwLXDtUTNueLqlHT8ttcfVYoHV+5rCNvvKcCtd6R5KepUIU0Rzksv2kFA
q4nMFbITpMd40ObM3gLd+DWAJvRQAc8dITegRQ+ABoB7GLu4eQvEz1YAdihaQekMSxmF2aMfyAKU
Q9ZbU9dW4I/bw2DCPrL25F+JOva3AxzucQliK53L+M+8Q3KCFR2BaxV2OGO3pPn8A2TcCGZzi5m1
mqP57MWhgdWbFPgBgW334nvYpOuMUjwISmfXZo2F7JmKDKLFW9/vw+0yH+ArjZ7XkdC5zW10eFRR
84adXEoABhewftkalE9JQV10h4/C+A8t3liQkkwTsaf7S5TBTRuL7mhMY7lLzmCSwdsAqw843RF0
1+zpZlfoGIYH4UUzkMir7qSfiWVB2ADGmOdQTHT+cspEgUQYorjc1ZbEZnlMW+m04ndx5ymCNisD
0QK6EM+4VtpmdeKG2EC+QQmMlg12oR8ZXMKX7Rb+oqGEK1wV5RdyDxXNOf+nY2dJvSjQhEbaTbdp
nTV2+ahFVk/R2mUiq71h22lrTIE2ZkxF+VXHiVbQRC3cvS4A9pbGRcv7gNrFuJ3L9wBZOfim/vxA
6GbRKjsBUWgcdVV6dW6+EkuEtTfXzNjNcGjFfuvTuihP7h1omlqpBb1WL6wov0MqTLxRxh1shruD
LDtnrX0Rq8I1ZIkIgkrT2RRcwQdjs+OYfzdajCmcLYk64OdJLcqJtuvmEuD8E6tgbZs5zvg8flV7
ljwlmbUN7TH3fPuP+hGshIlob4dfKEz1gXB/GZbFtGwwnr0B8xApE56yHSNvmW9zIibkFrVmQDto
95AF1saMJSt1IsJabnFsxHLY21R3IJFZEHyUDcZMDcDn8Kq5gJaRuOHm+gKoliV0N0Mykuf54hCB
zlhgUFqqf5cPIhwq0ewr+VoyLbO3ZHvCPq6Zo9Xzg/AliPKyj52h8AzMT5nlkUwxrNu+syiahXXj
e/KdkTQALXYZjWs9hnGTelXZX3TC2Oel2Hhl4ax8rAGRwV2/nxuz2wfqX1P63aI8me22XpabXHVl
GKbHT3mgB/qF3Ij3RQwRf4+0xUtDyPUKdAr3Ij38onTcs007AEsJF91IEH2QNHXg/zJPAJnAu0E4
W3r4R/72ycMpaG5mnjlCzBv4hZzJM8EiMZ5DW/qkHu/D/991sf6U2XTgBkys68J0amd7KbCZL59p
p8fv+YO+tKU4JE5SWpsYejE8snda0jwo6KkGHDk+CRN5Ehak0ZTEbQX1lwcawtL4g81JFPOnhw9U
EPR5oTZR78etww2O6m4VldcwYlkjjG+xipE4LQOfBx0hdJAXsbdMgakeelUJGfU1D9NbiScIVFzF
DzAhVmBk49ppc4533D2XNco0e6FYwGCqRsZtyYVPlJ0NRD21OrEuBJr30k3TbYXWVRM/QZI/9v7N
12XqjKTxipdA/5cToxY3svpy0+KnvSnmKVb3/ven41i6+yjUvIzqPhpEtbcQxDAcFQNna/Bow9oh
7DJtsEf0UmiAbq97JMcQBH2X8fGE81ec3dmDHovyoXWIXCG44kHnKSZ8et12GafeOEFM5h6WeZDC
BBJF/Y2GoiM8Siy1SHDH3agQQegDOkbl0yu0Ig/fTv/hDY7CyLGWjqZgZ5kg+8wdCOhDzhPhotRw
eqRMoIPvxMF9zfZ8dM2YfCfUOBXMD2OigBdhK4nhxskMBo5BrH3XXE3UulldNFfJVCqTOzPl2r17
Z/Up0UzxsT5oHbXBcY67X3wtP6gsw/lhjJB9K/U5kDekeFIsqVRhs7zfhabUkGw8mvgpY06DgFkB
nSVjH6nUip0Tax4/fSICBWcRE+1PVxYZcJWF11dVsaX4DhD3/K115Ax1+PpRSbVGsl8MMlRc27g+
OI4KFHp6uNAGZn6QD/rJnpOA7f1aUVNJccYRd+LedcyeUs8KM+gN68gc6S5/Iasu4oaNAnknBxY9
j5nQgZ8RmNdRiZTAcZBtJLJ7/lqD0b3f2ihM5huJwv+NDACB4WDd3E+485HhG8j1sZrXz7RkL/HK
IsNC63ZfQO0ez00EV/42nXg3xTgVlwMN3+rujeglBJe+lX9RPN5Zz+S7PRHWapuhay1TekVXALHl
yCDJaVUhPV3664YFKChHZ25j3LJXgqZX6YfxrZsu3fdk3okP+VmJf/v0J15KhZbqEbkrm/F1PAsq
cUXSsvAmYbp85k97Lq3mkVa/+IahOIPjzlf0QK5/oEhhgGtn1WmPkADl1sg+4XkoAw41NWTHXE/C
eSS4ThjmBCTwBPSWHaWjdwl9llE17x0JXwmitHXAyCWNlGShMhZzA57ko4G+sv7/ehMX74HyAjlI
G7OskJHTJdgJqP3o3hTfv4mVc19/p1VxeZdva0YyRBSQ/mAaXnRZU62dOe6s8AFB+aimHfhoF6lQ
2s+vzlfVp+ukGsRzrnbzG12Q0jc2NBjaEz60iadtmR7kGAjurBsrX4rKy2za9MMEp6qAlTmguu1F
78PHFpHhYtWfuFs1y8tUv6lJMOMzkyG1KclmmRQvGoIAi2fyE+zGpfwOEFsjQiDGKSTiV9Agoep/
apDVC6f5gLhRPjdMcx3FoMny7bsobELldc4UQ90s9VSWtqduHXwveBE1yvJ54w1psHLbRLf7qmbK
Jv3A80AlJshKrZXUWBMKORU/xhfTAO4DXpdf+lxN9C5t0WTQLq/Gm3NXnQae87BSR8+dbYvXKbtG
q/0la1K/zIR+SbZmI1dsbLTKiVCADoyYU+Pf14xvgwbRUph1yI8H8SxUHsIPxN/bn8r5oYPjh2tA
HtI001BmvIodBHO+pXD5RpCc0QB/m6+fdUetKr5qooQqzLun0oelzq4tmnH/nMsLQ1tH2fglHavm
DgML+fZaqJW5kj8S535eIVCsIdyev33i6tnJIYqm9BSc23GzSLeqa4mDjZOPpr6qKIoAyp2opgp5
dk7y4I0i2g63BWweBoNPa8XMjFwTAGlg0KKNd9FUzDXSbS1wzb6069lQHDSuYEWTBVGPuu81lEcN
46Bp0kX1QKvNSGwP9zBe7cEmiCXxBa0+0mAUyDaJoFK8/6u6nd2mLjCAP0P3LzZObaxS2SBSUVxF
d6vt9wReFqzy3CSoF+CErSplMowYZqRyHfs2TV4jK+Icd9bDWdsN2x/KoBut4AvYSyQk3nDsxuFt
DmHKKEQdX8dxKQ+1FxkU2aJy7GCC3QBYe3CTMkDtx1STsfxsF6LH7F+piB01L88Zg7yG4fhTOYMJ
U+cuAmVlenFlZ2qgt5d/q8J6W01WENeiE58KalceGcUB9CPhVQ21vW1YIa5TxsXBX0k3zjj7MNBL
T8GdN0M1YP4chSpC+jiC0+5vezKfZwHFvhro5c8ZNAwHujnMJBa9EPAnhsgb176P5QZSzp12ApgA
MzI4wc687P2qGsK/SpGLiJp025J4RgtmR3tMxc6AJx9HAw3NpjQOVb/oHap1CyoSZGfSYHjBXk5h
DATmTyJRPEYzt5mKLkeypPnBbNM7qbBYTvbPE7TSk6w8ct4NgLQlE0LHG+PxnQDX45eGCNrN7UYk
ofjUDx/h4QD5nZjR77FfAzS7d2p5LpVBVhe0hUbglCNdMiRPZrBejqvhIauxiyCVfFSA1peSUABG
75/t9Sfa0QcsnT0M9KBF2FxZIIaccxaaZ6x6/2hTJmQ7YdmsvEAsjg4/JTqKuIM6QB6h9s1UriRA
xHEwcvWj3z8IhzH2orwOo2gBngwbMaCAFBBsMdFKHyRWTvSmDkML4rzjPmc03QFxLr8rll7Ai0NV
2rbueqJb7XhEeRBAcA88lSSg0wGJgVTvG8ELYqrxkkLGGJj0mnKA/I5DVzSEgmZM3sPEtsYpc0AZ
6ugPNT92dNzPeI6oGvG83K8Rdk2sWHjgKKGk4CWrWLBC5grsOQtvkTw2kUMQYf45x8Wj6dnOCDmc
u7bZJ3qJnHm0CwzP9DcQL7o+uIPgI1YWfhr8XGMqvnskAu2C0kRI2g+YteUxqxppFd/upoT/Zmnp
0EsxKwmKOhh+m/pFcGYIUj+WQ4jK2vXeWo4pnW6YAalLW1GIbiQpts630A4Qv1TfS+yJhCtpfxjC
oKHGujNBTOD19Oep1mYMwAH8+OtWGLn3i0vcjKiCPeD4B6O5q8Jy6K+5P8IjSehrLE88upPU61gB
zEy1JSH7W4Tci5uwhwtwRhqrAzAdNJ5dLEo8/IJcx4xjPbbHlwkx1R+ur6JzKuTuMtI1vBfnntFD
O1ZFJXna+HLw2YWtv+2bg3YJabq58qBcfMva94DLkUpzo5TwMmEj3tXfYutmCIdjNbJScab7DgAN
cu3bC+mlC2M7c/JkUcH7gslyxM+v9lglVkI/zwsSxccsyvpPxMdonCBTw2d2LFZkNsoQUshUxJ+a
sur94gvfwjkqq3Bo73CJCDnNxija/uYaJDQr319SE+JjHZCsCT/ArLaI86yaukeTfIzhL0WEOAwh
mah6wL5ft2Juz/4mQtmj4AnNmU4Gp0gyshp+FpeP8TOUsIasdVAkZGNkECRZJ3VqlGvSjrOIHfzb
uKreKErFY8kchIGrInspHHaS3Evh5B9yyTZ/euFkVzn67ILWieTnRU3pF6XS3UGTodCXfONeM4rZ
PdftX8sexW57fHiPlcrdfGKlgTWXpyX66notQ3EgmNm5OSGPJI4h2HVLIsNlqDKEGAMfgPa28SWY
ThVEETY5tvd7l08UKyNjwQD3y3MdOdG/zDHcNeJNbsEAEKgE1FgqWwEt7CFWuk5K5tx1okgbG/24
P2c9CxvBGZiyq43JWLXQ6vhPAmPFq9naFQO4RWSAx8Dv5PbrYaQ8BRbnUxLbld0Y6Rwt9fGuYiMt
YZBuShYNhOO8WvS+m35vhlFa0Y1Lu60ngXL0fExTdbX1/++XGC7Smmfw4S3iXgcXl2+uV1tWR2ll
eHkLLtmESy3kvrV3ywubSz2VsYIJIfD3NvVlM5crx7vCqBYXpPHys96mW9xgYlEmSHayv96FgjoQ
/lKRTX4JbwFoDDKAxn0fB3zitvCHMy9ETWKJfX7Mb9cWTFEO7caKmyHcYMu+tyKQrmvwhCGftDZ/
PXTl+hZs34Rn5CvDpxPbFieFzHU8HEFublgjAr2UODSZr6GQ7jrssVAUlBMatGGgB3k9H/+JQLk6
o7Cn/sDiR5Zug48yc8MSqVJm/iN2qECxbvcesWxuAHG1Bnh3ayw3KBzIsPFRibWbBrXvcK2rCki2
JhqLIBqhJP4XvNzdafGF81jlBbWwg8bUbpH9WWH7sY47e92IiVzT7tfKHKptMGL2LZ8yXT/J9gL+
T2YrPUSq9e/eDzJTegosN86f8xfTJoJNY0CksgQfE8Efn3DMn0hm0nGd2aNDApTitRYXetgT6NeG
CIIUQcB82lJ0NtrXhRlblGlZ3scmgBss2VbWaCDJBapOhXi9a/QfWZqp2YpcDufBPcPdXnOO8oBQ
2FL0cJ5Q4YmlM3bJ8kde2cpaW7ik0Efb/7+dDGt89zPaGgInhz1UKtnuMvEmUsPlDGMrrr4Zhpfc
DDT1ejO+jzaqAzocOVZWJMtw5D7vOasSX5bRiM+5G2Ij3LCVjCrDXspbdmV7HZroBrclr3gOiNb9
Uihs5s941JBQd+cBIo2wj3uKHc0hqL/tolHxEpOTpqB1ae+us10xy4Z7IRxPMVcNlB4UZ8Ro3RnB
9SCffGR5gRsZLR4VVhy176qwm6Q750VHJDCednYRKHjUHLe0tZflyZzR0sSmkqeYLi4/gzRCPBbK
PuphwfNMJUw8F9T4eHvNOT0UC8IxU9zNQ06K0aXMYgF8FaXxktfxvR9w5PgfXmqhuia9BIHH4eBh
QHbKHME3sjABXE2UmNg31ysqfLgLq98VG3Xs81t8a8u0MtugNTUB1+gEZX86p66/4juTtEMIVxEf
RXIPOL0YIZBWOdXAu3gAVNVd0ZkwP2dfxn+AkmuNFGQNWC+e6H7i7ClmGpotzwZ6vL9zLKvWF217
SDYvq0ObdLf0khakypu7e5vq0Lkfdq9cCpfr6mLx8u2DCLqRHDWuwiU6HABTBfUL1Zk2OfVerg1Q
iWnRvJ+2xA+K8el5bbYRDbI/XuPjOgW1VNyvWaf5lKude0sC/9jGeqSCEgrKMkaK2NEfITDm+aoS
WFSJ/m4hgBCLv882xw5bmrd3nGaJ4tpNXsj00ky5Eh0srBHxZNvu/xcFxGANyy90GOJRy2UwtWln
XD0Ie4UK4MUAnuVqIgpL2/vJk+7u79ZIZFz0xUMB9yu3D6KJajAXZ7JnWMEQXgh6neDxGNcLREyj
0EvJ15RCiKQPW4GujPdyK742yq9nURr20zILzgW9HSX6iOd/qZQiF68tgfNuwPzwmcxFwAXJ6U9y
UYdIhSxOlbO2256Y8KdmROVugsrtyqzYiQP/gLCsAVOa6RHKa6dG0hZUFlNSliEfjcoGEnCoVbJ9
KYjr2DmWpsz+OHafP0CpFhVCuTJe0IZiDB1HTytY6MJuCzZ6kK2bYDygj2wiHoGr/BqEJtvOr2z4
hvAFU79yMga/1NNklBgNe8MAa8u/gj/I2w7jgytB3zWYzBLWk36zyXCwEbs/YxzBxS92I+h5ocnW
fU3IObyC7UdEzVHUMQok0HFR7aWi/0Cbu5QqEPm7f6QSWzcXwR50jtw8rFsiDZsPwTkE53hh+kZ6
MIepcwzuflTzTlIHFv5HikTsECNZLV6HS++2zLRxhhpGmUecc5sc3HaGg0EwifOR2Wc2KIS2TO7R
GKCbXzEV2NBN13qCLd4BdjhvHt0VuLS8me1/VBhXNZ5XK+HA/6uP6LcfwpVFhKWYOehrP9cO2nUA
us0i0nzj7vDMASxDVHMIwe+ko76zMMHhL4jAFwAAoBEzfss+VHIAsZFNZdm5FLa3d+8nFybdCMFJ
kQ4CJvaRQGUNTqS8FIk2TXQrxYiSIKulutuNN9SKyaSvdY3vfTdUyiCum7wIoc1F3iUOwuEXcxhq
6GxjQNaft8EUyUPEYu7wz1iHyTTnAMoiK/tgMRmMrxCBCFx+vIhn53OwDr/36Ar6tZdRpXFkacja
4jKfLF1j5WhbP7OKGOWFYhD8mrSUxIMBEU+Lgw3ux3Hgg8gN/selVS+NXQTxf0Ms7J8k4tvEd4/D
by0DfuKBnMfxI0n6ucIt8k6q4DjJuahO2McMVObhb3zYWJvyfSHj+EPV6mxm/0I6hoYOUCrO4Glb
fL7jkuPMkFQ+z7vh9q4qTK0usd3UyNfu/VTXI3jbt1PQwiQWTRiYdk0RoFFGzm0M3JDpnak1hiE7
Sy4uhET3nFFK+EA+0wQ1upTSj94yeQaURPQVRFhdRXIVnASp0AiM+taslWKNpPbRcWzpNTi8krxo
7lQnmQQAGPDcexAr2fo+QM0jj1NKC2MpyENqZAU2F6wwfa+3zSGQY4floC1cDfVfR+orJU9XHZIS
kCefAjQrMWg7fygWMLV7lVqfOo0mLu3fgONUjK/eGlc0Buo82T7H/PV7ZGGuqbJMLjjLCt4PvDrr
x6XIYtGeCr055z/HfiJPbkME+Gd4R+cqyHsfu0N2WIJ3D+NUpM9zRFfWlQFk8sLBdV6qN/AgB9dx
5uSkjmkKio0oAIzbFzQDV5t3CKyu0HOhAFEmDNu3hZbZ0kao7LQOPaCaM+63Kpi4u0vR6BuvDqOa
C2EwG3TVm5bGEqsPbdj4LqMz+SGj0RQiAd1YBhF0gHKPaGzVLxrq+Yy83+OG4ZEU/sW6cAC9xRN6
nXmQl5wpvoCo/LaJfpXfvVZn8gnXrUwAJ3F73V8gX6GkYcC7hNgZhFXnKdTgxEQl4z2CesyxkJc7
VRiHz3jFyxH9TJ9vruhhl5zePbgIlj22JhK5d3RaXSFSYP9bUtd2xa0u/2k34HvvHOI3A1d9KLZK
PANg0VE8MeApU7T72NqNanknb1SEi73hBwR9IDpDvj11ljQf1zeOZJhYGPctV/kTom4nEoVZNydt
7+Lnnhk9FOWVjol6ATE8mGoqorfWuNKR1WrOJStVwDEHdq6j+l6ShQU3Yd/xRSC/KP2MK9hzHfyu
i+EkYvHTySCfxdMBwBg2pOhdilRdmPB4tyK5dqktQc5l4HSUQEx/mMk8PH3wGgRAANOfgH5lUh3a
rT2VMUAv4x7qtPDmPFIkqiB67zSLYemm+gU+mwwpmimD9m98Lj6y7ScLMFK4hSDLPai9UtJB5hwv
cjeP5GoS0mYaCockhGpXjTuxUdOjag6baES8zhfhx0y91OlGRcL6Nv5zxwzrgSmOW3dSMAestahR
ialO7t1wUiMiIDWmSjU4y/bYbdOWsJKjHF3640oexRln1Xbn8NU3KiYdGga/3nee1CHIl0tpkhYy
N/MQBtO1rzCjdvMSWT0WKkPH99YDWsQWeiMY3Crtttlfdn1nWqTbz4ipDNRdkCBCo21ZK4nbRYcp
KwlRW9RaphrxtJ0FBrYnz01LLjYkfgZNqdrYhSNKBjY37eKximm2egj3TW8rOf7UkRwLnTjZ4/PN
ITCFP+7JKrBO5bUvswdSD2ncM3U7a1fHVM18IjrVdH/gux7C1Dz4vHRcv85OcRHtWmvIghiCpFvE
13UZyuqmABuUQ1AvBqFh0kCJAfndE0r174vTA74bRlFoxos4gsUXklzg5wMHrHrhEs2YED8OxGtl
mjoovaV1PvNp4Kcd+C1zRmZ9MSCbXsDgOUyt4Gibzl+Tc/lvI2cV5gvAvM5lIp6wCSJVQBUAGNQ7
YUxrxU0W+4S24nL8teRXfKd9iMQdVJPSLgxDG7QV/dgV9Om2Ln28Co37ANVcIMzn41CYT1+/HEhM
hky/Q3rCo1hoy0tEYPBYwfsEmjIr4kBVCx7ClJf0YYJ/tP1PhVyu7k8MjfZUC3x7Z6BJkt5KkB+0
Ix4fOje46y94idsiLSJBgZKIQqOCeBtGk3KZZ0yG8lOK3rK8txsk3/W1lanXirFB+zCHk32lRICR
3gC0qzIvMVBWwB9C/NKOzlAClo1yKKCzYZdUn9pWsANYZ1Y/MuaIvFmN3HTldB7GMtt2IL4yxJYw
+YpOInW879keYvFUMOcrhPf5uuyoozJwjW36g30JUisRMiWlRHO73TIjdrqgm+3FyH5l0jlZi+Vi
gbFKbPkmxCxgQAx5F9HcQb1pV4M/r2X2fr3+oadgtYCJDiwSUdnHeSLx2c3uePm3We4R6byUmOAE
yebMt/0GhsUu3AAC0GSzZSvqYT7cnW60j82p4LRV3FIA8P8zpMktm+g52jBl5X5yzhYkcFvRp4ig
7y2WWxRuDBJwsPxMEGDWcJMhxkm+j5OqAEvD4ys1bOqC77dzYGspfA8HalbXDE1OssGaY4dDe+Xl
YG7nueOMyxUbbSVXcEidJEQoF0WpeRCx1rI+qYXuzmWnyTftI1tuAt1W4T1v3wCX51ICx3uOsZOm
kQrytOraEll1t026ac0T4VYTbM9UcDckkrkEbPt/29rsi6evFZBUTbsMd2FBQ3l9ixB5vgMqBjmI
5MZnzgR14W8TBYKlDJcnoEMoxwo80Jke6NQBMSH2cE7n33gScII6ylQtmvYgrxoa0CC5EvzZJirU
y0fBZN/tw0C5Ilnw/AZTyiTLKbszZ2evn3Sr1v8db4n0c2A611Og+T7eScWShJG3FTul86+iXOf6
1R6sRfkxNN5KJvtCTqppqn4obY7YcuQYgQOttp6I7X3MAAUTrI/JBW/o1uTw+J9REF9em62D62iC
k3Y8svSm6ZwhjnbURbpgaFov7OLolkRc2HhuvArG4ZaQOfMfalaQMkueByRevlwjH1qVRwseJj0A
Vb/Pyh3ULxZhUwJfI0GBqskjY6hHKBX1mLVvz0dLVZumnNGFAkkyQB7Sga0AYgR12+xSsRQjStZF
8T3zFynd2rt5aVKyRuoEm2CsEdyqiAwIIbnAidszYO8JkhB1VMK4ysL0PpHPmSzCDB85PtK8Htpx
iMcRmOCoD5bo7gSg2m7s0D/QdVK/9Xq/7mGKztMYfD+yr7pJ9kaedPNlLkBfYyeMkhMFiXxDqGph
V8giD4CqCsmPqzYXeK7CSoJXkhJUQ1uv3Ru0ltOZX3ykUvZaXEo5q6lr2eBGO5nQcOGAFjPZaaTt
hBq9er6K+KUW1Y1r8Lv5/mnWNmdNecShIWX0/dyujT4CaBkcdHf46MTLsHLO3GxfwMCUwjq+RhC7
+yDOThqqaMa6pSTcREOvfijhHZsMes2Q6mUMtS5Hr9EIbawU39XYwkh6IBU2/KnCj3sQdQA8wc2q
OUTUohU/8u66Y4foxxm1GUfj4bN+m31pdoG74nDKWKZdzi19t6sW0bIzB65Ppw8ijwDcyTuh0CTA
G8TaPHxoFG5ZZdM1XvgJbsA7btM9iR+fCMsUb3x7IuRUSytXo1eoN4D8a3MTNgAzvUnV2Ls0TV3L
bkSANe0Um1BD2u12nk09/sdS1K0D0hA/UpIe7YSkPdLxguyHY2lC++EwomnsL+39RhregiNGFuwu
eqG26emGyCF9CaTq5p5BbDRc+TI6K2X5lUenpnuP/RPTagSjYdhTsYq2plexvyH5iVBDckbvnQi5
xd4Wv3+cdFGYet+OCVLx5lUXY2h95uSTH9tylEcXhl+ZC5Z4HXs/uupnhaqILeOQFg42d9110Iqf
tOybg/YUfIdpUlZ5S8nOU0CpXWBfcye/T7YRDVxAz8gjSvQFAErLT8i/FeSuf6SS0Jb43P4wGJlU
nvFsUxEx4HjmPbzNaJXKpQOSJ5K1qtEUbWtCZQzy0slRzzr/Fot3PhksLTziJQ7XItt/+e/IEAlF
WWBUndPqcyXiUDRRnxLUFdycHJofVTB0dQJ2B9XcRilRrujIBGgK1mHg4xVtFd0L/pPo/eZJFXPr
lMUpyWdUovsyHq5qGmc3qwp7bNw5KGSX607/gzKG52CSSNIUD3CR4JtfnicLnNsqLY/869WP4eY+
OsQIiKf86FJCJg20axGOzDeN17+//EhKvSPYRsPr1ppye0fy6NGgzIF+n2g8Bmq4E4PIAU7qyn5K
nGepb7e+XQH1xTCq6HoniKwc/ApmPhkW5vVoV0l1ydrjIrJ63Rjhl7zGIEJLD/+BXSDbiwhkQB5I
XaG2xGeGMO4OEoGnOpcMoZOLN/NMexUMPTREuUaqvG7B8IZwAJ7nO2j3ZcoYw9dzHuVW0JvmAKve
m/rc+Op0BYF2p/qn0oX4nm6a5GwDZzYed6mifX/t9Ob3ofAoBOIFJjcnM+h1OkLzeTTuolMVNrI1
SUhDTVTeuR9UxL/5cySQPgKYy1HBJbrvyrF73f6O0D2/aDLgWfbOrvQd+VBs0EBPvKOAiuQnK2zP
oIeNoI6ndYa4qcAd8Bh+dnedZa8YocyUKJM+SdE5LvMwzgCpR7YDhlnfkZbg1Pvw/W5umgsT0sR1
kPBo+t7OczedNNv6236UkbZsVa1OYj72x7Y3H9b6xgegxlhY3/ZKfNF+elvUI4GUUKin197LKf4c
c7TzGQmpbYtVR5dR4eZGd/7KA46gWl+W7ck8yS6mavOErQJeNMSAPnXQgdcebF+R5NybNRcRMW2Y
sGIHnN8dESJmkBp1eK3JO9jzcSR3H74JHmfKM4ApwY8gB88UDXmdGsuzpwF3eIRgPhNZ6o6iSM8R
BQ2x0gYjiJIGyAHNBtv75InGHh3uLEzidlKuDs4fsS4d4HZOXx+ustEFoQUhtcOnO8gS5HBxbmpc
GtAf8oaPxDb28f3IMr9SeiacDjvasXZBmOCorPkKqSUkJg7Qihtvz0b1fQtoVBQKZZtf6M4rshGb
D9qvDdCT9YR6QHUImJjm+1RvqsrbZ/Ce9dnSjRObzYuxkO0hiPlMKRippeJjeeD68tj5kOEroNKI
ItzM8ztmR2f5bgLDLc4uZpBP3ggE956n2Mmizvw3GBU34l5tl7ZtdVxEZjfqoiymmuG26u285xQ9
OJ+jCBDcuAL2WSqyUXw3Fcw3jgU/9/4T5N0cYSFW0eKnnE8MlWi73Fpn+D9ZLyUuV2EOh7cPXDzI
ncIlKlyXbNtHX69LdhnMJXjY3HbBXyelXQ48x21+M4fdnS1O30mWAkoWaKgrhnpxGzCHATvANAwy
aJSaDJGE6Sv0M6keQGmQiKODnOHL+E+Q1p1SzzNqizJfMYA/1SDuWFTgGf2WBegkNQt+WQrDcr0J
EJMHnWRkqEPqGBAHvrZydOu9zBrezyctyurse56gJwSTZZc6smRo5zaRyGpl3MvYgCYtXX+RvM/0
ytXH++FN3C1NEA7BtoOdvI2YUacgiVDmUWCwfFnQCZz+Gzm2bbQCjhX5xwRGrEJ2/9K7WH3K/mj9
hjDH47l6Z2smf+7DoVjzBxa4QcVxjyK7cXR+uXDS7jkuG7LfnoW1y0Ng0UfEyxgxStFnWklzUpwm
u7/ef3/0yFfUyTdRy+VbfaGFTAZRhUiXAX/EO94kWBPh8hIt0rK8dtuZ2N8RhPziYA6heBEemlJ3
jvA7rUGY87y8DigiaxPmM6t2MN31LMJGLUxw8OCvPRxdGnnDnO4vxxa2S2q7Yk8mbWahLOVnT2YN
qCEJdhDb6QUQ7QvTkR3snr6LlzqGmX/Dn+537oAuRkD174kDYOb1f/P7qqFSZJ6ZAjUtRavbx5k/
IUPRcuJLVu35mwwUhS/5HeUaebH3LRKdMivoJNnRMk0Wa0k8a5PWJfn4XOt7x9UPhnuiOdUrHI10
fwzTaTM5b4gtbkcXJMmh1ALZHKVjAhYpzRoPS87WMyfREGjO15Bs24nXLoMXK/tjD+leoCzG0ar+
43sALO6+IJsZ3UG3YzAhgHeK35QHKKwA2SKmCPhjGWCUyq7kE3jdKMP2Oqxi15daGzaHx93O0RPw
EkD2rjU/b419cOmcj2fSDz1oeSoGMnM+cJGamfK3LxPESdE8uB/XDu5frx5ptDZBgOPzixtTuS8N
6HigUZTD/4akEdmrQfgjBtqfYHHfpTmPK/W70mTXa7eMUiXUufnIlntdFdKUZC3sg48gntRZxgk+
sIgBXRnxHYN0uLgaK0G17s1IuSftFGsJKCF1xchPTYS2xo+Kd0U08cCiM2kp5rhPKV165ZfA5+V0
Ah7H//dA62rKfIaphhyXBYyYwjbs42OrInhjxwU7RNMtfXl1deGYPNXBr7DGtqfKMQ87U3dgW+1h
2gBYPuu5hJS6BNQbFiwRCWv+FHtK8B0HR2twwhL55zrFkUTJI59ZUgOjIqlqJswWPurgjv2iQF/R
0zXv/uRWnyUrSQZ6Qo8ajX/rEkGVnmVUulQJ4Wl5YzmhtF4Ouzz5YvGZ6cVnArQeM3hSm2LaODlb
yEH3R+ySLRcqsGgFxta2U/GXMk3rlFTZxKdS7axDJFmsR1JP/UVt0os3HzHJmaEQzEC3oZKDJYhW
U+pjdTxt8oT4EMcqjEJEPASMR2K/cz3Q+Onvtnt7cBRJI6N195CmIDWm6yIpL7zS1PwzWo9o9+o9
WbJy+R5qfm7v5ep8n0ejkbhiXnh+t4eGI08/MQBHFiRZ11gE7tijYsb3PwVp8lvtCjMFtKo+Tvjs
xdB5NemHdTVL+OR35SBo91+oKZZkkM3UIY/ocqXW3RQ3vFlXCp50C997l7DmmWpO5/fT5Z+e5ops
Mt6DTWdLt1uQeJwJTceZ76lakcObULGdmfs1qv+fWuEsWVTgF2w4GLClO4A6Hh6/X0r+xLnvdKgy
FXMaePmryg8n/sDmE00bvl+VU8XkPXz1B2J34bhRxPAjwPob8/T4RMN3BoDfj1PU+XHjKpxHdb7u
sxVvv5Zf1xe4T/0InH/LOlwzn2EEBHVAxEhoHxN1Mt1wwERTrCk+hwRCHnvKryOrXncFoAxvh7L+
9/G7hD19ufZ72JMP/YSl+atimb3nnR95lb/XTl+EE2qWdHkgkmaBA3lCLeu/FPQkXK1cNfbpLElY
gKStacSLzGGFRewq69FE4ZZCH4fohXwNZF/Vc1+zw59yVoU5cVByMkLClRzx0ynl8XgnCMKiGaih
4RBx8f7gZ6Pqvlmb75HIBXKMuQ6giFKm42KaDoDKDdsFUwhq70B6qkgKeikQThe+TKANH26iSFta
EDovFcsA09cfIwREnoC9S8yLk6M1MGmKdUiglCPRXz8C/s0eqYMhb6Ud+l7Gr2Gv1D80yHN222cs
eiCioFGZuschNMqM/E4qD5Sti2FjQi3+lZlKAT564gxYP65o84xsKB+dY3HNiXOK5/zPBQuxUo2m
MQEz7yXSLp079fuh3OUunEQoCM9bB+ygOsNdyMMAUPr4gTtb6ZJk2bstqYRI1n73jidQVmiP/u3C
MCYvJd8tol+NaCEhV6U/38alqwAERZoVJzX/H6IFUc9otC4yG1R+9H7rNK8c/HhSk+L3I57CX8wf
UwtmJ/80RIk+YFrZJ7zzNawflFs9tQN23SGaIKCIyK40cRoO3YzNzOf/Y6xC3Gsibro5q0HNDo5p
l+DYEg1N115kBe+WsTuYhXV9sWtV3BZtwZC6lfrdhcR/d/V4NGzKqSBdOBuj66pZ3SFt+MhK0hhA
+p5tr6R1wBpIyahNZCJkUK43PLf0D1fYBcL//MmbPisXmvbvPDS1u19XkTOBVl7gbhAmfNn2gpOR
qKGjTBNKs51D655fvJqRxoCTSMjJ+DyyTqrvNuj+mONoSV89JXHyH1Y0u5sXUHUdCYpU9V/7lK+F
uTc6XPdVMOkI8PHvm/oQiVqimvw+gOUHQ2YvujPOQaT20m7C7pNXIb/ggZphkCbap/IQElHOMfoq
gzQrPUnJQuMO6Rg9vQ9b8Zmu9GkYrXXIP52q0UMhpAYAoQerTBrcPeCjPZFU/Nc6NrloxQoUH1VB
H85yqA7GuBfha0FpwdWuv20sQlVvfuXguFuvRUE/Mf2nHsUktCYf/ACBe8wdgM9RRGvzCR3TPNg5
KCZLVQo4D83fj0T0OoK5MMYDfUykx9YcLGJNFXauGCU6wow1xCQek/iWHcO+jPmeMU2dOTrrD9CZ
8LBHEOQB0E8ELfRjGE83Nt1L/FrgeftWMY2kmvrW9VfevwtUv8megzBuFUCFx6hq0CS4FC49ICOz
8za32FD46DrzVjRl6Yv5ytOke8TaWUG/k7lsinvvCqIHDVCbG6rS8c62q2IdjuTjIDWw3h3Vv7rt
uuh2vg0UDf6TJTeRIyFYXBjvllhfuGcVFfj76pzj2qpQxIx1qmRqvwBZNpruxPKnX7yySSUT2LqS
/0A3gDJh5ZLmRpCxDW6kVWXm40XIvHEqQbdW2+AlU1H4TuKuc63tJfjryTZYJBFIcZO/pwSl0Hjn
Vt17i5TVRGpsQ/rcyuKc0hSM/aNQfRjb5fpTT9Ruvxecq0N8tVMfw3RDUOHeqTCgc1yzdY2FiGwq
RTOL6+HXvHxip0ixA7ckILto7sZ8PB7RhZmPaTvnATI5Of8usS0QQkJcdSc0idQQj8oZDg5mGZxS
n+YP37XRsLKahj2a/az9sMvSPb4DDI66USc+1zY7r+Y85q0fNwQPNzkfKw0Ft8Vgm9GVkEDrPmVo
Lt5YvquF5P2XaKFA8MqqhF6+XxJq1buQ1J7jMC0gXAXSkJ4/qa1fku8fQpz1GJuQoXN4Ir+gd/TG
7vC1P/OIeEO90ERcNvIvvubzK4pfTsDCNL3mVcVuNHDGE/T+MttHdff4GWPl2rcdD6Rum3E/p1lR
GFyZgkVQ57PMepBokVWl7yPGXEGIPj37X//5I7rODH84GfrRh2kYqBwNMaRwBugGRKodmzILQ6j6
rRFl11ZSqrxLXSjgNqVBvhOBzw9dTx4vKq+v0xpicqPAe6p6yNDp4hwLmm1zpP8UdjsnGGSFRfKd
HKmP2feOveHydNRvqptPa/837gIfAKGwID6Eg9S/uUnwzUOnL3BRkUO/SJd4Pi15zGkzGdFBZlIl
pu5pcYRvxJhV/rX7zPQ2qhcVQ/o3qqjK5nNQmk0EvctIvFTsjXIPpoVR7xY3y5hdE0jg64Ic7/Q5
yfm0xG0huydiwYzZgGQvdIWXe9c/t20wOaWk3vzoprED7hhdDczPUKUbrXJo9Q/Jc/auuUsCNaLe
4uPJdUVUNzpQIWCT/yRxr+23Hp+vutWL2tHyKquds4NeYJAhkjiFzEUMGYOgGr3s+gCGUUsVFRDX
DDoUHvCDxeZX6SL+PFxRRDQtb65i/0nQg91JrZ3iytFOSKDXPRrCROW7yo3mSg5W6qN3XrGO879Q
MsCKLliRXrld60IYe0446MSg+lnEf9t+UTjZJ/fOGlauBm/+Ys3gPcYEuoXzkOIrr/oRmc6TmhEG
OX5oirlOMwWz5tGLDz16k6akEb83xSMlWjeCdzK6kEY+mBawE1cBJlTr/jIxMSyr4PwivCjPiV5q
jM73H8ORm4srxq6Eh2G25l1ZoCX2iXBNoa1D+B9DI2lcXYp0EJfWiRKQoP5Y5eJgAJCBKbldZhaL
cdHTmWbgh2x+rTaizObf+UT2CMhM4yFOwp94HhS5FWFn+m9NHZrYiTDJlTuMUCyrugh6K5Gs+Yrw
2ZbhFEI8+OgiQgMz+OX8V0kCvQgRGhi58GcHv8pc+tKeQO4Z0eecvMgHqSBeKJPNL6wU5Y5Ji1oK
OUjrw6/Piwf0mrz5iD9lNbdyAcyA5lYPz9/RPAbTWlwx0lHA082VME58yVdg+Op22PFggZ3bmAuN
Hijq8KlTaJjtAUx55bR5zPT25HXz9qpqMpMMVSsDlxW8aDdqZOBrfvKxVYrYf708HGe7aOPvVXqG
M0XfgzEAgCpDkD4by+yoIu5Z29942V00gVoAzhDOCf6aEVehkp8GqYH+zomlWlP9pkgkqmviVGgB
fE62dx0tsfK4DQ9kkS+aqZmGBGmA19lk3hzuSel6VsyaJFC1YtZHhvK8SjMAVWBJLyXKxOHzqdq8
Xb4fFF8ob2sYMKlRE/dE0cXW1uRtyd4OqxBkROeU+dDwWYEz1sDHWwxhlg9KNR6+Kjte6f7/8uAy
dKDC0+40u4pKR9Q9x6EfQrYRO6/RLb7VYaDcsa9LDXGNBHG7FRM04jDqEjadpYttsLkk/heVyAcw
zdgPIvAr/39wd2xbNnqGvjSKOJB5c4ZHt69M8nTsmobYMqe3ecvo6iDvqnWJneQBHNC47U/6L3W6
bOliya7z7/U0ftLB4bNydX2cx7enHrM9VlKzN00A3+3OYfPXDu7bz4B+r7N//LRCvh1CDYOj6xl3
UMJk4wwlomRUBJmIZGPMdlzi6qZM3pwhVJFtEdMRWSGC68l21luQQRMJEZyIhTnho94HD5nO2HlC
3m9fL9I6bV8u2qGbnNqAIhLEdKakif09ZceH7KizPaQJ1YLlkXyfjfsQDsPqGyMCpzzM0cFpv884
va14PCVTx3mx9NLyVt0COuVMkBhBXM+qRYXJFy3IkfJYVyo0M3ZMWO/lwGbbKzKBs1V755Kxc/dz
p8Tps7o1FF+2MzrTOK3CNjFv7nf/aYFbjB26FwhSRfoDW9qtnSTARxtkS6ge1ei3jLvvHmtCVnDo
7oCcHO8e8nj7iVa4mEZHtivK8SpphNAjxwbSPsdgRlmDm0NUFAyMelYKNW0EFPNsHBGR8WRDll+4
qjqEp5Ny7Li36bNM1pVCoNCWMTH5wzRraNvWRpUzfkgt3WKyd3yXqHiVOXeZZzJ/A8msKAn11FuI
B8VAM/cnBRIzkyr9NPnXSL2xeyqnexUWsbTSgrNQr2UFOQerx9B7U6237wiUXExdr3NMyyPeJHsQ
2wQ2XsWkHAFvumoO9Az0EiUgM5MZfI5oxr8e6kG+JyCgL4VAp/pRi6TA46AqaQG3eWIG3VuG1DRP
FJcSDcc2DI+7oX74U9Iav/NGMLRkLwfzO8sVTnQGBEZx1L6WhqnV6ODnrwlsyi4lAcpeJK+e0juQ
lJSgrBgd6/mz931/FWZiQGZcsdg4y34pNtAs7Fcx4Cpc4X1MlIoQm7eUYAmsghztfI7L1dvLPlUr
0MQ53mHL2FtfK2XInXHOZs/7nSLAFlIDlxFuQ/NKrVqUXXa0ZwZ1+GXW61U2+sq7wrB7nw1LfQ0g
DC5lvtCbMM4HEO+IDf4CCbe0n21pJ0e10XaL5nDwUH1CYN7P7sZllCfA31KoIiA9aLJWjBCaDafG
9ozda1jKjrmEwldz+8DzmqvYdupqxjRViDZ+t/JIFs2vlbwdKj5W3ZMjeGCG1iE6+uJ5+HgRlgYM
uzvvs9+wehZx3nrk+kybG85vvxtynE2CG8ZYQ0DXR7ZxArfyT196EEWRei/bZxYmgY1JSRH5cQWu
o2bRQOJOfwW7tFDdBMMgCWKlN1JPkYqA56ksLZKWLgQ+qJwSr+wrbh/UxtaImLKPswwdwNxLWarT
n7mPD/wxplzgT20R0FFyHfxEEiFn2PLrvlJ5VATUtKd9tA45710by22QThEDX8LHSWwFAZVE51Dd
kU3rKqAqxbZ8eNEZC6lJ0DAWkwaKhhFW25mcWCMxHUdR60d34hAznq0DHPX0JFiuzfPmH9/4uH7h
euP7jBK6121dOAJqYDySP6jBwack/AEX76O5D4jlsII9OwJzumiOdimzaRriVtsBgr83pUwkGsd1
0RGejW3PVe7sNq96yIpMlS09OGkCBKGmNm1TPe/UDrFDE/8GaYNMBui48MMNKVaDbcTw1kxa5KXT
JSMyz1heFolKdLTZIoDazs+Y9Bd1RE97LvxPby5VhUaZR++ohOfcOYleDRdO+dkRcm2d/PU4JMv8
36nW9ThRZkep5Jy9AIdPS0xWzTFzYZDQMrYPZ9IVmbgzOMAnR0afM4y5dU2uJrz5gXEX+d9+mBHE
qb21FF24zYnVjQMMfH/cSEXrGEUncB+y+GHjfKwaOp6QqB62DaHIgRwx3HiT0uluUU7iZLzSbrKV
CgLgNiO5z70mFbm6iKvTNd8LOWTuMnEyQuzMRs5ejfGLgsz7pFSfN/0bAGarWI9uOX5qNqBys0mm
jGrV2t5UJ9TGka2CYvLPBQDKbPU8dcK5GKPHvXMnktqMBB/ZGywqMySPp1HiSqu2AKEIjTeqmZ8M
WyzDCS9U6ePcEeuspITlxSRTqHn9AcRIwqgBzgx+QdpliqfjnCValxsb5UEUAxHKNnPeciRMFX9T
2jiTBTtlgmLmlRy4Nfj2DYnSMgPPZcFvAk7c//FANMC3/Y5WOJabkqnUDHvj0/xlp0Fb+iWBe9EB
++E2i6n5OAU0tLrBjwtVWbrdoHzIF9QXByKIrtb93Z5vnr0Ji6c1KuTedOPOlqhZ3FEqUnOWwxrn
1hTb9hsoobjk36pf5YAyjs6hXZB0WGqF96u6W5yD+MZ97OT1v2wmUJAfhgAX29MCO9gpMq9soKxq
lavyLywrXYN42DX9FJ23lWU4wLHzYQut7MyWyD4QkT2H1xKvo1SEWnBFZIRfhkRcygsVqU9LFYq7
XNEgOhjzClPfPqJx1CX7lwewxAJFLbPDhE3I0G3Hic4oEEQXPlBD5RBfjD6FOXBRiIR8qQMFprDI
GTZTLTFmFUTBdsFecOMfleytX0zWN9IqnKaiYS40WfcXKdsJJhyswqbq8RedMkZe5ycau60sljxp
VXPL+w+1wrHcd50D0eVUqgHw2LkwoyC2KQKnmfSMJHkSNgg/BPtt6an2XOP78CwzRqErYPmsYu9S
DHjjBwqSw5GicvDhsraOSE4I8FIQgyLtoVzW80Owu3+TDoMvDkdl0+QQyvE/jMtdEs77nVarY8FB
dB8V7qI1LkdWbzgkJGHnHeHWzgOl8M+WlGbVUxGNbbNVLSoojSN+XJlYaQCMLNjzdf0/RC0dOhTX
zYZiGk35KloY92y4YaQ0DSMUK733R512ITs9N5FRABWzJVRHkrPEdI6rEx2O8MfRWIK3JD74ebY/
vXlnBEj+n1SESlXwJtqZLeVzA2KLoBHkmAEMqQVw60paourdnC/gm9aLnJf7T+NLcINbk6qH8K0L
e3jasFRDVxc+Jp283ZAyO2frbgaQ0RDKsrgM6xRNhrkCrdAjkAAQmgeBTRTOHPUqDzbfiKQVup9i
gUOqW2uQ4X/Tg/dujUU+Qd73p/hSsIY1lv5k8RspRwZSOE+MCySQi/wZuQFjLZDR+QTaWUjmftQE
KJvIDHXZBksynEhvEiqNicbzW3dZ6Ilv9AIcAkXBz3TXfwugBSfGBcXYVXXUvt1GFqdmOd9axpN5
+atsPmN4N16izM+XhFl+/I9xFwfzZgabJjIielnUUBt0upQGIlTpu5LxEbXjc9peYyAbG8FUJqJc
cTdBCD2IJd3Mh0ARS8FfUmQg3DqlGKXsDVNUp3cY/Wk/JrKdsUKx7jfU1u6HVg2PCZbQ13AArkwM
BsDkqaWgWWnYmjegM2Y3OHs4XxxCv7pxcZfx1m3c9+oKIofwcj5fneHrWrrCUWRXofqh7MqbFWfu
JgcIEdaTNywhuFvMtcg9sb5BhzCD0pQTabUeJQQxiWrefY0GnlqvCw6Y40b+A1yxfBMis0AxHalH
WV7xXo1H4QSWRtFwPu43bUH2SrfVH3Ina5fc9kV4mdYEncWUk4052IymvW3kEUgnLYTUw4/+/T68
YwKD67T5XnFd1hQKc0iM1lQVuD3be609ccoGoNBDjPFLJeKkfMSFNNii2Sb8+/thLajF5e7V6iXo
EVewmHwbw2hrj8DDzr4tZYaVCau26iHB2lYQmv/meOdTGij+bjUeFI9F3YjjjDvJFGmDZHDHiaew
yqYTpfb7Fm2Rh3Hm1t//GeD9kpstN/4U1u5/CzxRvTH1WWVznqrMYIprU/CprW/RP2vJjsd5nY4M
f4RCqZaCNP1nOWG4symr28TjFfJv/pNo24DvCPO2DfNDlq1jxAV9S7hanGhThIlxvu1gMIveDynS
eIGL48SeXgPxMfnEiaFfYzO9l/7Ff4IK6w1GIjOIjr6+ZjWEPIY+qFK1UezgZsmz6Ykb1kucbwAt
0E9a3IXe70ex0tOheZuZIigp1/WW1oZwpcPF7WjwH5X5igeGOvYepjc5zm2w8Hb29SoJ3uEq0syG
Y2ddyk3TskQpMtUtoZd6Oa/VUjbLRLyeOvpLeuwCdUYjqGBpwSn8h10Dy83nvV7AHwXyrSPf0KWZ
EGA4lnajkqfI3YYiySIjgTsONKfVPN1zvt19we3uQdpw7yIm+opu0GAR7w+lVRkUoVfo7ZZkcxc+
XjpL4pxBvE/owLJ/Iem2oMcMI9ZVSrKEcOQnLLGQozyF1Zd1+Ep9KMKMAZCvT+ThYbjP66GW79T5
FguE8oNsYyLkNeSaqTlA6lXwQOfbW6j6f/DMepfLh3c6BCwfFKCbEMIln8ZixLRPqmdnivK+sM10
zTctRUuSkmKqJnNkNmLaLaNDUFzK9NWy3Oa2Zg7j0Lm7AmSma+V17WpvLS6lD4KHqcFKomBQDfx2
foQ3tskOfxbu6nPJYfK1VZi3oAvB+VbynHj1oJ8QrI+Fyvznloe1jJlmdu1/NMWfP+yioDaul0bN
9ydfPpPhMbLmaq9g5faBNtAI/kRkkRuQVwxeyoDCySeT18GOrHbsg5ygA1Q3OB0jLD4uidR/7uVU
CyGabI5tMdz5b47MUIbI17F9vuKcBAO9C3nd5VQVft/7ero+yfNrMyDrKHGgBgMgD74amontDpaA
ylycoZ+UPyJm5kiu3UuJlTOIuum+wQsv/QkYOJmZip1z8Mt+JyAeyJkUZmD7V06iy0z0Xuw19EjH
qEdjmIkGIBzRrUlci9/2OWO3JNF2LbrpfXdKfbq0wnRuGPpPLDy89ZkS40jsypJYykBHbkFSDOnk
DvIMjwIHHhXO73yVKYwfxn47c72pkR/edO3CXuKNjya+PDfJfD+AGmAFiH/0RXZVUr0uZbZQvnXw
vnKx4ujgeZEoZB57YEG98/DMKgmLRvJj2my1M/miUZp2m8M9NsWciX+YctmXJAGqi5SdzoU2GPA/
QTuLgbF3TdUzhi0MfNbQvY5qDyrukxtKSwz1WdJVEa1SnIwgGmNczlUew84RaZo/iJIK6FSse/ug
gUrKUm4wt21ehzJIe1wmJ9uLUl97XriYyh+gUx7lbz5NeWntq8Vx/+rjCBK5eUhWudMpIZ2jUlco
+3JOwq7gyNlkIWfovPTKMUt/KTaxhTxyRqDG9tf4jnrXdoyJ/XrRjRBcGrDAUUfG/O4WOuF9afpI
ztEJBJadPJ3SqgXf+0wotqob9ezncrs5tOebk9iryor+JKeY70fczligBbUgI1Khgcpy0AJHmhuw
yIspreae+xLU0xxSFwqOGQGGRgxJO83TP6BrjdENnOfh1V8opupvQjmLNf2R4+uEeMvrGhrWWEiL
mdhi3H5LpPC2iPiLqcrfjKrxc75NA6b9m4wVW7CibFDf/vmU6fdhde8l5C5OH6ZecVhEcFcbVQi7
L5UrX87oXl6ILO1Y/fB3H72EpyqKjPFOtc3js+VwmhL1wc+xrz9SG4o0Jb9MAqhdwaOojitItiLS
8CmdnVV6yX7JogPHHjegP1yMd7qgPCLpOxp/0qOVp42eFBtW28du5WQ391w9UMjcp6Gc7EVzRdWU
wxXeqrwPV/HOmFaJxRb1/gbqKjdl0uMEzJPqygYi+VxUtglq26226Rdyv0hvGo0dRhe+Z22VZA0Z
rrxmotkh6GebBUcj9tDxHLdCKjfhQmKZE1vQJodp+AOL41D8m/PaSiEyaeAIxAJIyukLV/Zxg+gw
V0nCxNv/aVzLPC95JxCJyyQMUv5EUWmgZKWecdVybIPWq4FpSu7RqNUAJObsvlHOLhCcvAOFy136
Ddf3o59SJ/WPfSkPwoSsDdJr7p4UyZYdKtOoAqTPmjoYQvp6QcYOUFpwbVGub2qOZt74YPtZFBRS
iCr6ZsSqw29M3ZPX1h+7Fxqns7ZpqAnPYKHYIE0SjwqU9yizGl9e9abw8N+AM/rZmdo2IO0uk6a3
LIWwPCA6WNFwzZVl36bbNzZSJUpfdkHS8GTuXIoCPvlLXG7GFXCST/eT5QsAcAl/99vxkJ6YQNAt
6WEte+EbadKaemGuEE8CaLSiOhkmb/Cptm7t2or8miYYlvTI9vCv9WoHywCHv3EceH9uSl8exKH1
R2tOerDre2++NAw6vlYPdwMEVClEr7bdVDArQTPVD/rIXR6nQqNDME0tmD/+QuH1MnrpyKVzhWQb
41hYor7x8HAXu8S+NnHKTqFrau3JVK7N6MSt4v3JopvCpVa2XIuUPqJ097A5+EXu7JhKYIENv8mc
fqf/K0NBZaB52/L7Y4BT9EvvpmSaW1MY4COLAkNOzUe93fr5raEFGD692D65mWCnazmlPwXXe7Ja
W5j8vOargcD8yANSf0BkbTU+bdjv8vbWqB+wp3BpvFjtoMk5kAdMqXafa36xUIOfTuhYEv3Cg9tQ
yfRanumLKxwkQyt0l3I3xU4ZeG+B6beCsgctdje4hfdR4gFH514P4WsDBUIKN9s6DYdGg+3pgEch
8NAIdzlb1z6na9VCBwb7c/EXJN7GydSozKesl2IaVF+QURSek81sBlo287+Z3vjdPiCp7boC997i
ZpmDPlyc8Ml6DxQpXLEcnP1dk6ck5aytCd7ExkiVT6lX87zi/Rbke8HKfOS6uQzLNapz5XqOz/8d
8sNQSy4AatohGPfmW+pN2VV75VdKQdFFt+pJuJ01lGVbRfuBp0PQuQTv6jsZURFDZioDgMmUiWXT
TNC5VsWGBpztHNel15l2uGuuUZrLibfR+fS7pz2CI40Yxtm++8YhwNsM2/KtGzszSU+bvfDcb7rS
1ACBt54HSBL9bCNds8IqaAu1bd51I9mlsHsS8dU5rlpDQ3zNhtLPHzIhUQVKU//Z5ggXLxUpAFoF
/J4+iosP2vjuFMJtDpGrNAg29GtLdLvSsK06gJVlvYIG8EWbbfLf4AyG3xY52CCy/q1VWzs5j8qz
O9qM5KuTIzFiP+e5FC9exJ6csZuktP5nRN8MF3BSToEBZAItriz+A5WoriGRDUwbnU8afoj+geXn
N8/55/2YDrekaSTSCB6w5+wXuYUXaGuT6rCI7NHae+qEFHc9yvOYUuKYOOZfDAGtOZ+J4Z66qea2
Zabi6wLwNK9von4/GeVZQYXnN6vVogEFHpjmLKctWCYYNlwvvLgWnhOxoy9qbiT9XKe5DUr62tbM
9wX7npEDT3wxlX1fgv2kDjEUFmlSiyRRBHZfaLWpvH0KRd4P8qZ/zxH5lzjVGAp4Cnj2LDmR6YvQ
jMLc8yZO63h+LhRfGPskpyoDISU4n1+L1VJIkbOVwt/fXBxgF8YsQuHXcCEKI0mTs8qSallfrYbc
cgGHUmO2lz77XYJCrSsPEA2b3HNW0H9m2IPaebUURItpnVcJ3Svp7YIW34pqOtFS8Um2ik1d86FC
LnFSiWsOjPlaO6JYcxdbDO5yIvxnEHq7pfe+GnbTRL2H3caXbeUaFSRRRIBrb4cK40ylwPm5HSyq
Zo/d/DLnLS11dM3B7W0CZVtBXs1eOcbb60L3UrPwmHV8zTmgS9+jpdhMEZaBI7JqTAH5HuVtNxxZ
8AIyEnUDZduvI/tckkcGsq/iDWbdBIUkkroLiMArKujchEbNSiabMiaETC/PfNFLXs2cBKx1uDTO
HxBba/7WufCDI4ue7jLSc7YI2qOpGYhPYbudWrzAMMHF6FCvOFc3Xnp+EkZm7aVNVHUJRVTBdEaA
GfdMPxgqsMxAYhEClWNKJC3QUR46yjw1gui77W3vJ5EknzzixNSs5yqGO7TMYEya8JAjrVbtilnN
XQB8SJg9o8s6+dhQGMLOU2N+Unf5Tr0gJeItPhKq855diUySKnO363hSLS2cr2lDgOCqh6SbIFDc
r6wPjOnJW/fGMqNZan74z+dlb+MQjO7DHk+J2X1E32fHLGnhgn/LJwtEnLekIVwitysxwIlChegX
He0t7bCyirJBTdxLh4PVE5lZJSnFolzEegsw2DdiHQsVllv4CEnqZvbo7V09/qQKUCRFmqAHNajW
ABZKjsrwSsicjl8Ucn506CIpuJL4n+reQQVzdDOKIKLZdb8dlmSeTQF1l0hMg0KIpxkDTUOuUWft
ywfu+UdSc+cGnmnDVjjk/SujDRe0hqRxOgOSqpb6pv+66DMlJ+jfYkgUMpQkPJuarJxmtt8gqJu+
FsOefHW+p9io2ctKuGoaHJ1mOqdUJOtkwO09o+XqED9UweE/PV4HlwPqVP0FrvUcbmlzjsvSmXb1
tu/KDAAQlVz6RbKOLLkqAH/yixM5dJhHsXsHxADACwt+LaromOqXSh52ecsNECar4fA4bD7YoVcG
sP7qRe2OuQHB00LhOdX8SgVCDgcV5jNfLHZrJilRGLfDXz4qF6vzgrNR/mnFi5EmL0rtLZ04Ivl3
ntW8nf9lzxKY6Y3qZeLtI6h3AwKASRZSc8Aey9smqZwyn43HkbPf2tbT6jpQDNT7Qev1pXMODRcU
A6WqONVj/Isap3HbcSH2uDBqHAECjUFYHwFY/EHwgnw0sCcRBkwAMuQg/WYGYGoDgBXXJVFc+9IH
6E7qqDKOyEdIMxmSm++GeZ9EiA6m8klaaCsX+cxUyk9IKTEk/k9UN1RH/87YhlBo6YYEJTZoUhBg
kCRnyha3L3HVuPqIYD8gwNwT8Pi541FCPG2y6qSSw28HeUCzRaMeYVAQ78qGL3UMWcNEtxFqbSl3
gaMRqJYkt0oTB16+FEDakkuKgkoDDNhf5DupTtcgIWe1Bi+nVQcyQJt1tX4cvPh/Qs4KZHFooK/k
XxQXhosbEIn1Ks0RVoBPQ0vO7FQuU4Oofbix4wJm3Ah4nOF82hdroylQ9zc3xVKdkkMr0WeyeAn0
LDLLl3sj/aR8KsW0TD9v1hh56XTFiQUqo1PVUZSmGFnPiRXXQiXpH91ODd3zOtatC4Kii+zHWmBV
IiaMCSjRLAxPkUOkMml6uIqnHIvvV4oDDQ4c04aVBij4Ml7QRonZQVlRRqopcncyZKZHrfEkRQqF
o07oT11wH/wlzAMuOjSprkcTtpBYKE4mn5QAB78Ab2AAiJbZKk1eHd2RPYh8fLbgFmBBNcEh7CKa
hEfiX/zxGqXtvCidgECzqjSaQyIlF2ojihqIsnHlg1FhlTsYK41Df7mMeOpnnSXSe1s2yaBCdJpa
sPTNxT3PiT1lutlFsLIxg5pP067nKzAgGUQ/Q5Bu+rv2QD858657QK9heqQ0Byp3GZ1nWoRsYTTB
0JgPYfEeX+6Axj7ojY7axtLfQfjN8ppNM7BJayEqgMdY2ZYgqxZN/n2gdTDDMH7Q4cmtWUAaMXRE
VVRz/yEwbUVEapGFgxa8a1KbEDIp6jgcAc+77AB+ds79zK9qV/2jDT/0N2t8rh6U0MIbY/jIns8p
KTb8Ps4DZZKEhR7R1sffEJK1YGv1Nwk/s1ElRdaZ0PX+hzu8/aWP5sbz+I/j3RBVJ6fkPEetPlYf
qSt0q8jEc4Kwf0dMJH0joKeofwBoC869g89YbTWSN+DU+rRDz+VlRgT7l2/+KQ4V9wURQtv6R6kj
8SW59yJGLo3emAxgQCakP8I12qWtnW/nCp1dZnvnPqsU+AyFBSiUBr6PW3C4FSrDlGbUJ+klIgIH
83qKaUhtyA0Rt3LQAI8uq+fD31F6oSJNn9ltAfyqkFYRt0EHeEebj89If2T7P3Kg/48cve3rPSoC
D00GNRT6A5TdWzNbrYpSOvW9kJAR/8jrqWn/vHwurHJqpPFbw5s/mZLPHxUG5/us1AI4e4y+UdGy
WLLbJa2DSt6d2+Kz2SnbqErkmlBaRCuPmIShiBd6jNJH/0BqXX9FeV4ckXqkTnD47zWIukauK+kt
YkSfsV4FQoyRb6XuVPM/8j3E8YBEmTumeMJ04iHO1AqwpqHHibjfwojaKbA2kIj5gY0AsQy7sg2+
t+v7viCRqVwEPZDl5WzRA2biHfC7xZMDAvG+ufEvFjXuheqyLc/PXTu6nPjm7c184UpNYZv3bL4i
0gx4YxKuUk0AQy7o7x6xwrYXszP+ccMiVGaiWVOrQyW/NzyMyabRrqcHaNv9ozQmSD7+eRRxxdj/
DMPTwcSywoCgSYKRe3NZXlWfKK4+wBdq+Up1UKkULodqgzbZ6rOXjupt4/nhGonkhKZCDkjtSI8i
UXWoDIH8id1zxePU14uTyHle0GHa/AP8mpPkdV8cRYAdsBeiTCQ/kepv1vnlmR51uy0aSTvZTLKY
stIvitpQeXYuVahs5h3z5TdDpvwFjbKebo275jVJpV4Ak7wFwoamax8ETB7M5IKPYYvzay7ChRah
+rS5hy1+cfwenOSPCLO9tj0MamP8w5xDCmRxTpMyGb2Vv6kFuG64ttWglMvaLataZkLN/rS6SMic
hGlR1Mf6ccmsN9dbvQkXUjOs8z6V57bclInVrVnV6SLJwEjSC4jhuB/DRm3hD3+2ccNp0WP41aQv
bGvpTnJT3jFft4Vlk3czYTPALInikG6dMYJvH9ujwluYeFQNwTUYDNtvzNcMCgc33n46RR+mdJad
fmgpBbuvXp5BABsJQvtliCGIO3rXQhn9zufPuUdgUJJcGVM6rYH+DbMqc9CRQemxaILxalXbNkJO
pwhydQVt6RxAkR37NGkFTy6/6PC83IjnDY4Cfrsnxawcg1sk9KYYU3pKXyHxBVU652ZKPdzo7Fzc
r1R2aUtODX3iQNc/PaxOFGBTAKW4hLVXG6HN5zAfGxkJSWG1BwS7QUqVeKgyqYqNZCse0tWo35xv
jlRDck7x/ct+b6Ft6blJZwyuOECQLCRm5YtoQNY2qRmkZ8iBNMTsh9xzIdhexiOWIINYLcZ1s4av
AaFsl9DJW2QSX3Et8zymIJjLFnE7ZT+5G6j5w9OxSlnslzvO8trC8GHXYNcBv2WLscj6UUq3I2Vq
RhAvoeMKJi1A9+iX6L2C2T8tc+PYflqYz/y7mhXj1Dw+PjVehoAzoCHbW24xxmNRcy4Rso0Ce+Li
rCVji2vbl1wmD1MZ+brHnzRDxinEzv6d+yJQk2RSsJ162tfCWTv4II3V4DY7YW5RJe73TL9Fjnq8
qYDlYOLXMaWRCNQQqz2HyRBgeiCU4Nuxc6rcuNReUXaGe+W699DVaFgpf+N0xlCYSNV7g3A6sAWb
cSzUSbbinPDTWJ3lejkZQ5bbxLN+J7bMaH7QwWwj9fNrebvEtjAOlNO8h6eijFnHlYguXU4pQxZA
GgoEET6xg0SzRxr9okqje6EHDIdAGnXtS5dxMVvaseXFbAicWEj4/6+rj6Is+40KD8TCxIjKBw2Z
UTGMm0BT0d3qqvJzvCHiEZ6Dha+64+tCkVLGKJsHuQN+WqEdDL1y93VZT1mdkvr3kcCM/iuSpCpx
KWL8cdlglCFxIWQLGvP4LcaLp6T60/LGUtZE6q2rH0n89PDbv72q2MK7mXFIGS3X7+EuKZHnwTxk
mUfH0fjnjoFKc8bfKdhsCvY/bIb40mQFxgEYEDYAlgJhTqfSFVhCNIqBX73nXKpMhDH0epcRRhH1
bp7dKi+LK4YKeYuDw5tWKn8eiyNxirNEGfvoawNQmxVkc2LZMSkKf7KNRrOyrCgfDdZFFWWJ51FY
h1jTKDCgYZMUXlJUfEI5sYv7YnqviTSe8RtOFndRkihiP5i+XBzjm8OTpl9SYzlBT+Sgil8rMPKm
TAiElzfIWQ6Q3GDHxGmvpwkhb8pntr17tKdcMQiwVZ4wOGarqIhmY3CKwY71PueSWSHeT2cJG+iT
QJRFoqydkvHMoL/eb8vPVQv9cz0m9ZMHY++pRfDjnzalk5SdiAMVwIwsPjQa6UwpeUrrUYAO+BBm
Fxryptc9ETsPjn6urVNnm3+XycrKryZHSJ5hhKyBnwm0Q5cX8QIoQ78zM5ZIGdS6oj9TKEopIhEC
5/uq3HfEVMty7duOuED/svtf5Hjl+6BgU1dqiBJ0yQTU0vxxdYO3AMXaU+XKbTeKSRiaKnONicuw
xB+YB1Y5AlStdpf5qGmcpBmuReiRv6RXh1BytV6YbG93uhdc54TbusKma7fj+vydmkDCpeonOO4d
aCv0XZjGPilO3i5cgixhTiZxAjM7QgXUKzidiQdCjlo9T8urGNGOyPtIamkhYporH1N3TXy2T6oq
fCjrNJnpZtQ4x5cu/hjoRh14A/4kJeyi/lyqCbAYhifcGA/VhHINpSCnSx1HDfkQ/H7u6B2isVyU
wLvxN5xzAu/Zp0cSSDV4G+Z4xnjs4mQVoHoejlHpcCNria65lQNqUKw771HoaJYoUnaDjkqCneIa
GOslMVAHNz1ObmKfo6YDdHi1/oxQJ8UIa65m3mzfC4EdwxhnqmwEs+A9HK1Ncqco5mQyiu3TYS4l
yQwNv5XO5e+GWAvML1IllAEaB6lUdwTgsB8b2REv23rK574pydWxciNBPNKAfwAwhOE3M5hskvxL
ABNhekVR0vsA3UDhRR243jqq9BBs3/oOcIZeqMPvluJGCXHWLFfcIAACJb/7f8VygvWzYjunmtaI
HjgIXSDJU+YxOD/R78QEv9Z9pft6kg7Dcems+hn+DCUs/B/mLNuXU/PYzWbpFjM7RBfDp1tiCJCG
Epp8aAXVUImYL9MVbd5SjQtUmavx9yhZKzSPE94yTXKdxPO1Ika+o3ITDr59HqaTaqiSEtPbjgSJ
3WL3/SbVopbndwDB9j5KJdZ36rWlKtnA6E91/LGGeb2EQKUmHsuWC3ipy/qD/gIkP9V3rs9DN0lz
voemb6u9mvqe0VielTi+dF8mqm2ihNzvaSLt93HzOb63j4S44+vobdHLeusFWbX6g/6t8+TDhOyo
/nkwdIuYu0gTL7djlPW3UwAU3y302M86wLdZdD9GELOafW4zsQ3rmr2eyQm2e6Buk4QeNGgW7dNj
0butlXpTBtU2Ju/vcN9ztmBMv8L93GzsZwDKyxPhK9ZcawsoKbx+7liiT9P0x5N2uqyRlfVcxEVM
WwEBHdAwsoFOFsQB7XquU7OC15F13Bybw61NrIWXwSQWnqwDfZiLDphVhGWCGE5jg1/MdqrUUxEl
qe16Bw5o6bJkgHSiCEg9cl/Q2a0e/PO7ex8hfTPJ5a8kOEkQshYVwaNjjZoQF58gVle/ZSekxwu3
5ZPACCCCci6A4g3HV2KAS0qL2x8BTU4lyVBVh5oMRZDGDWvVupPY9H9q8KlQkX6EHu0cFlV8Xp34
uBmIYvEQLddnBFX7qwOQqkQcIDrZrlg/FVGphkInZv80wbeQKaUmFa6O1RfV6qZ4DNV1TsdrGNbl
+7/TodI41BkiiIpg0tYYp65abl2U08Kd6ssnfpuAurVYzlBfdiaEMwaQIlMM1N4GDz8oQZdv/XFf
lZWLREVMIAurL7iF50ZPEgxqsidftoZ1atttQ/JYgv3AIiNXSbIz/tDedE6HoI2KVv0KjDgZN5Rc
sTpP9Aalk/clF+EhkaZFde+8JzIGRYveVzkIRblGJMXzxObUvtH+kCh5Q5J4RyZ4gKrenxdDK51V
ZT/tTkQ4qUl3E7mCeA45nf4Ywt7adoUDTNWhaIcYxabd0eeqdtLdDtbM+lbhKH4t1WOkAnTQncJh
/lWf0DIStlD/oYY4Koh3b+UHbRCWUN36kVZPDIPUb8T95nyiH4gAhdzAURbHI5Xe4NBTR08u5mrH
fMqCucMDyJpwtoAFakkPLvtzwhSoF2A+QJhsWuPk70SSI3HAb0gKR2QnMsnSGHybrHCxAt3Bx1i1
ES5ZBKpI8/nFQ9w0OqfXE+LS6f8xBu29TQfSaT+xNh8jj2hRvSikgBWhYVKDrwfUNQiwt0fcNin+
d2NLDowWk/9UJjS3mEeHbq/wVrLS79YYurhec9uqXX9fOo79xfvPDID2g+gkpKBtMZ6T6KaMEMg4
bD6sxljk9NDUDLVn69wYO7e8ceuIT367Mu9f+7PxwbxwM3VUAJK/69IlNNREHCOICdxWPIs1PJFU
rBjQN8pQqlZFSwCiiXM9fjWaABlK24BJUuqCogIwefG7rDCPQRmdEBl2r2CP6OoQCXBgwBwgHEbY
7Z0w4bzy+14i/46X8FngxRYACaqM2tMKZAAL3E1RGQrUbNhr8wH1O9awJ5P+Gurgiuf2/kLqzUPN
Qv+ND0qnAR+yOQ7dJjNACzQby4+j7y8tph6TxeFMvK/PEKYnVHYdHVKo/X+F8sruMu00LwGa0e0j
8Byy7SS+LU6BwzTeWDBDdsuepw3RvU/IrBpRPf41rrV9OoCz4NaDyZqa3btGq1zLqYhuZhweiOSt
5XUBTXkW0/kveWC5qbgfAIXmGRCtLbF/+IURCgE5ED94JCaL6dAczoovj5BFmf6It28qTCeAaPe/
Z/WbZtr+6aMp/QSvuIlMIRfuZyJ09FB6j9EfZTR/mclKlpzP3+o3sdQ+hO2fU/l3wbYC/P5/2ZvP
WV1yRD3gkFysaQMHGTqZGAm8WFIztByfYx65Loct0O1lAJS8Mb5sHgaoWq4/Z+7wwWcPkSvWC/ur
iHng0295/RT8hzjDrCwMugpWpOckZsQv+SMu+DRXqAL2uzUo6h2NAu2ivCd8/JeqJZGuKO9+0S7Y
+3j/Rck+A9zbsdjfok57Jl8XIRpn9kYooLoraaNHQ5Zu1fuPCAKdGanglpATgTEQcPz7GXGj8p3h
Ap1RnsDp3i4+7lgHbN2ZRcOv9MZg0oTtGuvtAtpLtAp3E8HqefQEataHpF1rr0xlv5br/YcfYgdc
1WAs28uQspTZje4p9je83iVPe8XebH4Eg1nHngOLGFu84RkJzLW3Jtc8g3XbI2aaEgl9sHjl7dIW
CY5e/y33OO0VMgjnrihgk3TkyCDpQu/YLXejFV96SU6H/yls+lvz0mx2jYKaR0lX6oVPHQKIMZvU
tgBSYHijd8yhyju+ivSe2SuFgaE7t+qwkGW9QKVGAer9OzO70+fo08CveZV6cfbiI8Q8FQhmnJJB
bEjfT2/t+WH/iIQNeSvT6hvrBNDVGjWh73AQdRHNPFtXi0YI/AQXUqdSdIwB6TJI57oTzhIIwYP0
dMBTMrGsBpBkdtqarqAKTp1Myo7fZlEcTbPYvqPLl3dLnNJck8leekR70oo+pdjwBqaNMvkcg5aw
4TggBAv1DE6uEPZMsqeJmejEPxzfKDUfyTC2xSMpwz0sfdWdPD5AJShQDpSfejrcCM6UduloOH+R
Zb7BxnjVWqn1fK1E6ZISuWEj1BV9Yxnkiov7wC9oVzCvx6QQDwzCpWgaptBmcgv21oKfWjUbzDMc
2xSra4QP69ad3fHABnZbljh6Nbd0W3pXTCkg8eRcj5Py3+1XmqpsPZ40Owq2aS47o1wC6tHXfjER
vNlHxBztsDahJVNCU2QeJ7/w1hv7KFA3XqO5xrtBhV2vhucNfhwVvHZ+v/b8M5GYSNpcQu1EbRYA
BM8e5pL8Hp8ZMgfT4RMNiAvfW1dZtA4+1YCdx6dgC4Usqe4JCerkbb0u0CH1L0Tu/XqTIZFKG53q
ECdtk798zk4665imC4WdjPlscxZ6kFlOnPWn5ruBryZMSQlWCEO8KSY0ySTW/0K/6Di0PaTsMEJ9
xJfSSQ1Z7YF6RxbZWg/WPhZLqelOVWxfpaahGjWpO/IPJcD5bkSXcmkjNkrs4s+6HsMze/a+6Vks
4QAAmCjdmVUXoGXM26EHXbNGDQJOYP5rhMIlbNq8Amjq3y/cyMgsN4OLXDr/f2sSRHXXgwsAFPTF
RkG0KmXGBAIi/wkzQU/j47M0Zohp4mSSiVnRL8FuQnTQIalmvoqjQ7TIoyTTYG/8rcm5H0HKi1bQ
7BgRpRmOPk6aCH+11phAgsnZOKEz/SmbTpffTj7c5JY4BBVFN7Nc7Qda9SoevxZKvYqPBNmh3MhL
VW7OjRfLKNFD//ncivDl8bNA8osvPa5I1H1hTj1u4WwiNLmPEosAT9siq6c74L6eumu/zce1bvMP
c3trhYnBfKrNFXGEmKwM3442jU6PexcmVyA//aZ0rzJaBJgqwQ+RRjb5MUlkIBIdjVFI0zhtJVTP
HYDF7+g7PZPd+v1EuirJndkOMdlVcI7a9fx7iPsv0tPc6rpaNL9yyWDMskFDciYxCTkf7cs5R5iU
lLQfl9dD4WbFDmWQdiNZqFhPw3Gw/zh3ImlEKjCfjkEkoaXed8WNT+DJ6MkTlIFJGsFNGG8w6ITV
M3ViCkvw8YJz6aWoRmBGR01XYPH/rFRDqRBWCnCld0y3EBONUt9xm556+Z3EeZGS5C1QKiY6HSjI
e3escSSKj3xbUOSlgzvyFP2hLulSjHu+tkKNDVLfZ4D18i+ATRtnpMznkKBU7QJFQTwB8Wk2pPMP
80jGqIYgXoEoHjAYxOn3MvlNV7Q+0p57G8lyvA/4KxTUprV5z/cXxvI4oEtC2LpHmqVY5oLD4C5n
+nn22/RONYFmmT3u1jVcvHzpSsBn1dqr4kKwg41+HaukBVaVGeJZzl65JiwB8S/ar6Wy1zJxEIan
bjzJVH/LspTXuNi61BDQpy07J3PKP86SbZBlRzVJP7BvV+dKccQM7JGwLgnhdM3HB/5mtIvY1Q4K
hCcSIul7PuewWEiqzEkQioXBLqZ1B7eK6mAYxoZxCqzcRH2fx/hXApyY96zcaqNXFLzvW4bp8l6/
qNYjelQCkeJxCcnyl5LIpvzsohYC+hLWOzTpEKuSE5E3eFToEB5s4dWyJe/qG105BWFE+EAteN8Y
l3mqmgTMFEPVE5OIQzlhTtZTvly0nCgHxwn/+OxBGNbjVtoOgxySQ95ojmhSSKSqH+Ue5cnnXBOd
CjX/wSIAxFi5a4b3XzNJ63uLdllc/KlJ+KIWvlShqfrDMMBaPZ7Usmpw5tdasPblA939pACtXtQ+
p3Qzk/OZwc7Kx51CwhlwG1qmIXywrvifK7PlhTfDgfpLS7niSPed8ruuzSDpTMseBUyJUXAafCvN
BrnACxFJp/MNZP6aXMv8sX4J41Q0+/d5GgEBY/lIu0NMF9w2CsAYjOwe9jbH6jIqNOhJ1ui80BlN
IUdDqyvYOPY/qZg+UxcjqtXhTDXp7QjYkYbC9ZbalCaYMycnvr8NF5TEEVtxwWiHbjoKtPwdY/Qs
jwBlOrtwcVVIitl/tZmsABA0Uz88wiB5UNjT+t02fsx82ua1nFXmA2yQXCJGR8fGaxBwbWAbx/FC
T+AlDNtHjivJOnB/or6Bsln04MUUs08JDvFZ3MA+wBf6jxoiUdyj3wKfisoi8HGu1Q5qKT8b7alu
lGkFfh5ycI6vmCthZkQLOd+ED0867a0JQ4GLxuWH2VG5d/tqfM3maIjQsafj4rqZlId3T9mC1AoW
un7HrfbHKWpTu23G7veJ1MDeVK2fom8Nw4nd+AYztySQ/JpaXHe1JvgupHxcdo3Ni7Zlsjqjm099
Xw4EqdpTFf+JatL30pKfO2K9q2DPyhCaFOZfqLTOKRUHah9z8M9gvt5x5IifyxJmVRnbVFmgkhAs
JYl3NMXVzRa9ofcPVQqTxO2/SEUtLFq6hP1PekY5Qu7+mkLHkaGbz/JZSsNI8qQSt9gMFwnhi5sN
MiwveX1Ab0bQOkdZ+MbLR/e+YxKRo3cvyXbD/9fYsz0CV+lAfEhn6u0xdBieF9PM0zpZnJd2o6Lg
1VowuuZKijQwjieUc0gCkf7gTCbipnekAYjhIwLCCimzBcp8g/FDEE2nLAUoo3V/muBf/VO0CSmL
wBkHrCxtkQcvLFMI664HtZU0Mp6lfWEh+7Z3ymTNTfQjOeYF6srXxFGA3AUDg0Dev44Am1xEEBpF
uP+qECF4YS9josNoTatuwnboppo/JyZbEtoFcDXNSCfLcgeFz8Fkotlvj7DDkSzbBu2BBfqmb1mD
rWE9U8f6Mp7EV6bQxcC3Y7EliwJdAqXyCqSIBuNeSEFTPdtMlWPaRspAPJAbgmv4k3tDAlkTSaYV
KmZKaCmVHyOhBCYxMpKZThY2pdW5nOairOC/94MZAUvPHKDrXN8d75ZLeTpeofFt/yNbaKAkfoIi
2RBTRWmRJv/yieZaxK62IxMg/fS8tqQrw5NTBj3UlEPRZ0761qhXG75tDsCBQana7CkMMchzg1Jb
O1642q9A6EisnXHO37O0/hFokNOJoFP9zFOF4ZyjhkFDx7uSA0oo8CbLOFNvXu/ahZRIx6TBVjxN
l6PpGXxUEkhU+7++1m53/jcF9MSKnVJ2BzhaMxIu8lTi77zcyMXPAHQjwGDTSWf42LzAL8MJ+vCQ
SMK3xEPiXgPB6rPnhDqx9f+iQYym1+0KycXYA3R3sx4qEJ8b85qJ8sS73p/OGCo2v8FcALnV+gAy
Ylz61lxPCuHBa8+Iq48sWaLixBwX4nyBZXGQ7TaJxeSP7oO4wqhW4QzZnSENez7x2z/+HwZDe9ti
oS2YmL/zRwT2RzNkAzzCsivswjcVaGQx/1x8GtHqVrXXpP4xRX00XhVXRHbCsWRseRzZLdCNQKf0
3RqQvwLrFxsjkoRVoo17W8H4NngxOSNYr9xUVFWSbMFbetcwGlrZOInbz9SBFg2zs42bGmNvblzE
QKiozCY+oy+TrRxXt2cEK0xrPNXA9OXw3oDNRkUQ7Jrea7+vOoa+P+8JNdjMbD73zKncy1IkljYF
1hN9ydagMrauOB4mFWWeT5Ml+YMsNeUbP4tsVOb1Eqqt74gabY4+ukQSqjltvT+sJ3oqLZK3BSSK
6nhZXw+JIkZZZfXC25+qpxUQ+9nkrCGUOCVbqkdf5n91ZAdXPQgKVYR3ZNnQiS4k9W1UYYFq89+k
D+1mzw4+xFLyjxX7ROwouAaTwurG2yHVei/SHiYeEN55ZTexRbWAhjeqnjOWC6no9MGu5vsIvgHT
8h6FeFd1DxnjabQuVdQr1+Em9aAiTGEnZSd5ZcRNslhDidd/ZNhlKuGL1L7Hz9N32Y1WDeylkqRh
sjfns8Zt2xytUyxfLiqLe7J17H9lqa5n3zkKWHnfKu7dLZMpRYENrPesu9483uOvVcgmoNcdpICy
l21QckbUpoKOBjnT7CxFgf87xsLrK4Op1AY77IyGBSQfA3JxzWz4oExnkvwtsqaKPXC9u4c1TOPH
0KtH8sAH+TgTo9/DIAe7R1oz5JPEw5bnz1HDCIm+mlw+XnGEcfucef+pU+H3CE/cTpufcXD55RCh
XnB4cmZrRzjRX/OjK4m6iYA3p5Q6zZ7uUx2X9gjrh75g4FnCmyTvTRRw7K5kgJmV5M3BMDqAqUx4
tqz8F7gJFk8uT5uI4mgjl00WPi9/lyxn3KkSx7M0sL4T8lgafmEe4V45lYpok7qpukm4MUwOElHh
XDK9or0/ofDVtCU4lQ369WNMCXAttOYwVIz5dW/+gYbXHBrt1lGAAMI1Yr0FFIm79id6c8eQ6xAI
ahmgfCTUYDCWGLoHBQwhxSk2icMpHUbejU0lTX9TaYQd9gOFHcioOrXBnQtgUoOt4NeXEiPc467O
l8UHHoCH6zF11gA6Jru7+EY6+qG+5gLOM7khfXFFuIwcw3Cby+DjYJKUvAc0Cn3yFa50+rtYc/ce
+VlZTqF0dkI4EXEvBmvWQpX4equab92dF1N6Tkj1pmE6eFTV1ezLHJM8+pJGnTE2dLE0HOxEYyci
0ZljC4E0Ja8x+5to485WMz87M/MJRsx5bvdTHhmNXItMfEOrrQUJox0+AlrkVLHdG4wEGVMtV8aP
AE74fOOM0GMeKAc1odFHj26Vs5NeHVcVrVPzEGubok8ykmO/lCebVxpyxeNkAUboUdogVNyU6wMV
vZE+hmNod49piPxI1rLBfpzBmlEsGX5UDDiOlM0u7bqZfaVctVQ81gN245+ga7a34Ws3TnYeaRhM
onLw9ii/08Gdbeh/f++42xNY1EgDlzikvDmuU5iEgGreZcmMzh+rK5j6WNfBBuH/NnV977YRDWrP
oQ6ELm65lHnzlVHT1NJ57u4qLulW0ZhHOtbTKGQw+MdbgnFdZxXGeS+g4djwj0u8WsniJtaJdpoL
IkUowL8Y1zc84mWMCWVLH4iozPrqDkrJuRzk1v4lix9zDwqr0Oruo20K82uwl3ykVpKcr4aoZtF2
0merXPn43ROHdvzD6j60qjnfWf/YLnKLi4olY/JFV9raJfgi1zKe4acMqVNoJ3hd/xZagwcdUBGv
YtPk9PU1YDMMlFmM9Sm+uPPlzo1HVsJgUdp+erTuVg7tlMFMFOzFpzrIevfHTYyatn9v1cg15dPw
/OPFKLis4Lg4oXvRfx7LZRg6f1GK7m2ISfUtWi55fCYYhwkJE96nSsUbPYBuKdVWRbCS0qi6cGFO
Cu1wdLqmmJr8xXRNOvU3iUTYgcwd7cDHwQdmHirsUyAR3i1TPcfCSSjvm6ia+Md/c70sMxgCVMli
RnyyHvs4V8VIsD66iPmd6A4A8CyP72fmv77eiwJEtO3agNi8mUOD+Ed6DGqGV+ClF/bvrKdd0ybS
DxjNA1sbzeAsNygLTAp4nHTc43Zc090Tbp/ZdMoPTMKybeo3Ic3czuWgngv7iraTGyqeQ4ZhoKRF
bqR01j/7Y3pZFSH9a74nTi14SsNKGxovr0FukX0hID2PH8BKOqVW845LVzxtJqT7uZPYm0E0TtUl
e6hSxMsUwnILdp9oQNpJNGR/6o5DFkOs1FyOEW1Mp9a7DbdOIs6NhN0/FBUlsjm9dO0xMoVxhajG
nqLf3oINXZSPcQMZHtthT1ZUFMxWDSYTwuZsLCWzKM7nkObudKQc/o3K028wI75VSIrqkpqP21lk
hf2/9kwLVtV7vSME8xGncWqVLgvIbO2ajC8SgaQhi6l9/FNW7U/nr5IMylfl8ywsA1wJoY7XHV/A
Z3FrO/WNfEPZiqP7LFilIzkQI/OoOgJwtZiS8OEQdquu/o4xn7WReLnKz237W28b1qXi8OOXXQ3M
NsEd1OmfQxq9Gw/y7mRlpK2Yu4ERDqCcABGKiegBGUbZyzsnwsJ/3qEspTU3wY1Nm31I2+z+jOMu
+/VoEPKnbcZ3cIR+S25AIF9MlgEnzemEySxP7DR1CiZhrH0hXB08wJ+pOS2SQHKRsfrXFNOwdj0X
5L+uicGobRZ2l5ElS8s92CBM2js7gpEZfdAKdTqtXmX1LYhR5piq8a1msKl1myIc2Wx1AoXWGO4g
4nH06tlPmkB52UBIFbX5zKUq/80nZch3e0FA5tCn7chDxMB+bqjlgX68eSY1Kk/GOXGRzvNRNR0p
QLEE+d4cHOfB7KdIUm0jKVHqFUx++zEbB/x1h7tC+BWk1mU9H5vii/y1QRKdkJ3sv9F5JV20UF3v
5wzI776udXZ9fXoaQSoBb9eqOA/evDWLNNY7+dZjCLnfvFusX9jilnnx38dtzeCu7bYRRxialYbr
vwp2iQT9WIi3KvCbnYz/gWZXWOjbGh3JhwNns0IDOk1vKvqDKYv5m/isuTTGZxPtoK/ydUUacCIU
UahmO0uaDKT8i6x/5yR1U35pfJ/IShF7lQxs2EJjVreUknuydkXtTzO178PPHMxTBILCEOEEQS3Y
izU7/Sv87VcKq1ITALNZguzHX89lwX1uX1xrXtrYEoLqNnSZT0tr83k8mD1T+lPDDBoudBl9ABSY
I9f6q0p5/S1YOBi9wjNmwAitRGDkiQl9GM0mq3MBTG5F6gOCYZNeXebJSkET+Xdh467xr6dxt77J
OXV0Aog0PenzYZyCN38zELZYK8k+VxGIyHdwJyAvM8y+/nakuxj8S3F/Wjy91i1XljiBtPRzxBOe
qqN9TWho4YhCjqgUgtc95kjO5i4adYOJfnll81wtOgp1FN967r3k6MTcopRt984h/OZwbUp+a9mm
Tm19fvZAVgE5pxcRjgb6AkolpEss7CQGY0a+eb4OMnCeL/wo8EWMlvnlCSScPoPJ25b/KAAPOQbV
OKbmHfdx3B6+OILOuoyP5nBWr+COK2FG+Cg3SPkReWDDyvyvqDa1eNYq+7Qb5EwEFq2KmW0PjYpq
v0Vbdg5XjSlCdzSpfkxT4ydVO7gsPY/0irW01mMOm38Ieftj0y6BG0hn3GajdB8c3pgoXxSsykTv
KBWOOX1hUYYWV7D06b6t7/AfnjYrokX19KU/oBHM9DhRFJCDRGTA3ABdQpT8FBrbggN5GU7/nosx
qK5qitXZYlccJzJP7nvP/cDObJDu47ha4GLbmgdkLsX9cd1uSIQTpIgNmJ21gfKnpMHVW+3ILSr/
OfTEs2EqVfq7eVzF7ZjxZok1ygBngOsAlDuMSVWXpfW+HCuQ5376pc5ms3s5pnajEeZV5qLuHXiB
Ftkqmxng4DvfN/SY3PSbhMk1qCnuAzW46Lxfz9ecNbQHaRLGIhzrpqe9/6EyqMEryxan+Rilq35I
mnS9WBJaE1eMRQepoS9U7snNdnLhWY4r1f8HPu3772f0b1ybyigBjkCw1BI/+ptav3NYxzWvXOfx
9S2vQxifSwvQpuuFI9Oqr8/3VcmpZp8uV80I8YqfHVYKxw6vYiPNFivPhyzaSQNuH6+TPdZYyNK9
VWnU3CqXsvzMS0G3JJFPYZaAxH4QHrBYV+xboacg1+R+3VcvfAjad+CVyFO4KnLgll36hOKYKx53
6APs4XedE/sCMLnwX7347Yny93AfQicVS3bCezX4Ovhgc/wMMkh64kIa5kz+FcvuMaoe3B6ancnm
sc816PRY0UfZW7oacxB1nfGHqfKZu0dnSPRjYnI2gf5Abwx3Igkuf6yQmy6ABTCucQKRkhD6DY1+
8LxQ2YBT/z35O8O9hLfYA76bFRh8yF8YVN7yfSn0VbJ/1ROxaqDfIVrn/uc8cIOjIeh2ve6e587k
Em+pgcALUgmrJT4SG9s+qKg4qpQGJz0mXzOo7zGl529stqFvSfXh2j61jRQgt5HZ3sNyrzcxChzl
DvDi+lsImncLnYd2nf30gIzVqctWuWi/658zx5JI9TmUIg9M6hFCn0sFRB3ceNh3wHhrdd+brNV0
AAhKlqOQQigo9jFucfDyh6+a4hYkMS1/tCQ/ZDHcJQhRfLrw1Sp9VUsQDPh7jwKhOJeqYQ7Gz3/u
xalWcdoEEkPcIrzyirdBQm+mgfAYzkLVwEx5s6DiUYlDtlFXRJ6N55DcHZ5PW5EPb+7vg/DsjBB7
g8E8jGgGrnXR2AhuFPUsiUF8l1eki8HlXCxzSvuv23dcfmLhHG/EAmN1gU0h7Y3plJerAmXZzsLA
XkPkWECgPykuoImVOrK5eToThj+R/DR7BR7kKzpp0q44Zk130j+0pJo6Ix8NSDNLwXibC8MxSyLo
nYXnOXyxUkkQcZtcLYO3XisIQvnOHcl71/Dxb5oYKU5lQPnKSi2OkG7CO44/XBb9vxny6sv9iCnJ
A9X7smrvtnO/tifrO7HMqxMo8IR//9zGYrkVmHfTXv4zzk7tP9NSU6LpRL94bTSW8iwWyGt3K/oh
fpuKyicA2qTxDWlICt9VRz6CPc1uM4o/7n9WdTTMyB8nsy9sEXS01jf8MtqiJyQK03EajAPfEkac
RSA5qoZWMIZUqn0VnYvhqyE/FpJZs0VRv1oev3HdHTAdPa3ypZelbOlw2D8ZDj0pcgpEZBN9B4nc
fO1u2dOusWdAmshcTH8YDjZDryzD/46LZpXmmpLLeda6Pr7aZUq41LhoVAntA6EUXEDV2rWdEmx/
S/Gnjr4Icra+gyBPSPFzbH50drpNnTRzth/DzT3xgQsAdrOOB8EW9pZMkJYRv2mZWHsfzO9ODfyL
jEhDxZbSx0CFzC1CJq82lPdDaqs7TjJBAHeUWiys3Dt4+lqB7Cf2yLTZQrbv3YubA0I2SF5SM48X
3ZGV4ww+qIl/NsKYSSdS3huCCxtI7z3KU6ZpBy1gG7wMwwYjv8XF5a7E8hC+lxxEi/n94v2sxyGo
Loqwtgv8vadB49u8JJJrtvIkd1TrPkICZ+7ldxTvFGmxekfXIDia0WZwaap8sA8xy/nkqVv5gRvE
HRFDcObiSOIUcikZaeLXDN4OHYKVpOZR91ip7x0S6lDO3AYM8nG4Ni10o0z9AWbl+qctvHOy7DoA
0AH5GlFwEktLeXTo396mctS4DayyPvFAIU6kDK3urS2WMmGOHwvDqJ6d2WwrLpPnonklwmJ7bSHg
el30iOwykqY3DkY1kLwrRQ0hpioaewDesJzNW8PRyn4ivFR5vPIWWOXgfUO8DO6Rb1FZ9oVoc0se
ws6OcqwMg6NTsHZuQwi5qb5QmGBbb4mzKltWXvsyA7YH1wqqnkjZ9rXaZYUcB+7Enrin1MLjdtva
7+A2J1DseniJdDG2CyKvjs7ZM5Ptcxc/turCgfdmLXwqTKMVhSxcxg+5RZ59Vwun4XLbyzD1HRma
dZ1mL/xw+kZlvHiMMHww3C3IFzsKt7Fp8vDHhgmTgIiNGLjdVS0SAlr31a6BfdBlQMnS8Q01FZMF
/EPAa9qvfSSpJxUan6vj4PvPxM1WCrhPexJaXZRtXtwm5SUc3c9vJ5J0BdG78D0nucQRqABgdcrI
v6PUQTCiloZO4pGzgQ9jJK71NXZ57Tu5QRY7VSjJLi50+bm7NaHivmkw6Obuq6h4iNt9YW9jJ0DJ
dlioC72RwpN6CZLwBKoUw4S9O2XJiM5rh4W/1a+PnJ5RctxthrgDuxVnwCwqIhgxX2p84Rqc93R1
U4aNlSdjPlX4WsXu3i8g5CGP0cNFaYn752jAhHCnNsquSUE1gmRMxEVny6CP9jFItKF8LerxTlBw
8rSxoLrZomzzrUG+v7RuDl77LOCVzSB9S8f1JgIAAE1+TUfY5vL+W1A8f7kkl+5ezM3N/+njtVqU
5brHt0eJQBIumteE6e/xcBTDsqOd9NfwDNCnK6XFphSj8x5UghahFOjZWY4WOsHq6759bBTHJYTD
lhPbuyzRtgK2zIwuEgaQH69DG0Nhuup6HKYS3V9Kf++O5mQbeO5MskxXL0moHxYKZCwXwm6ppKPl
JU7X2WykA24MbcaAMEPM69Abh7aR5MjG5V6LQftQV31JZVXo+rbiqli8RL9q8HfH/l0RN/7FY/mC
VlmAoJFBwp8ZrDeChdsHMHeXAFRTPbMOETr9j7DaPwn9OiDCenHHcU1rzUrddAmsWszqNIi8dFm5
iwqKCbLMYFCQv6sMKaZsREIV6zGl+e2LEc3j9aBEFDBmihvswiXQPM+LNAsVUjhvANKE1tm2pB7n
r6nzL861bstIeSy1rSNnuXDMZN6jUGAFWd2PAAmapnAHBMDtQB0c3KAkcQt5FkYXsIZ/kLw5CjWV
/6BdvMkDkmY4DL/MZfGF03EZ1Q8HqLIblnxylFuGYozjBBKcYhGeiEMRrerAdomRBNCS6wdCMkZU
zIeXXs4zMbQiGL8EXtxWlt62eoVnMfGJvCoj0dD4ey0rY5IjTSSffSaDPtYHT6NyfZqaZOE+z4Wm
xu2laKBkZiT+S5/Krbd+ilZJtembFe/gFQbLjov0JesgY/jaU58YyuMtuhrdTO4EVXsUmqp8EKT3
jHXR1wPYZx0LxqVFomhSuRA6E6W7hSj0dZ4iOEYt+hz8cX0KiNnJfZHM6ptiqCVgs0iroyZacQS4
UufRrBaoc9MQ+SNlW0BQAfq1FginS9IOFROBf9NHJF2ZiuBh0Idh7hChwGVmHjVRPVw1BsxlKYoa
01eFBwhizhkq5kFdFUTR0bzvijePAE1hxCLRlbsrYsfWEm5kJSTBIFXRxYEYbJ1r7X9QQQhPAPqt
fW0BYLzMUyKWqM2Zam1PWiVOGe5DFX2GJ61VSvST5sLLUO08E/1cT1FAk4ljzQBstNkSRr7PZRVA
t757hqbubn6kcoHMyCGjk7tnmCAwemsv9mLALuYSxy8pfM2MAIleOBzoY6PVLqemtnlbcaW/s2pF
QSC25sufhUgrr/i/3vj9X0zYAENgRER/kg6wl9AUVnfoRe2QM4CiUX5RqwOoPiivOERGGVbE+07j
J/5wqLPPuDC1QhvjtKA0FVnDjdFFjuf3ACK/nhZYItykKliff3A3OnF3LyjSF8KD0aIoCYrQG6qd
3Bgp92WN5lZkP1qSkF+IXe0l6eW3PoqhP1mmBBVfi2TOPnHDcFwGp9uMquSQSps7Gf4WhZK40PiG
MkfCip/zEJYUdsx6qH7ohvJI0wCYdf9XKStfinQYT940F3vav4TJG0mUzyvzyEsHrVhYPMWd03qB
+1HMv8DOx55nOcLcoHj3loVFMyUUhP4muaVepvyzvdHlJJjWVRDvgBk13oqss2hic+/Oba9LdXFe
7tzRdqhTB3t/tNdz1QjAhzbb5oPTVCiiZL5F1BhEw8CHyzlDlQRqUQ3io1f/VfGv86xBlszUj0ub
Ih1fYUEbke209R2bcpj7SQfsF7XWfli2Oe0UVpMpSrHXdwQLkW4nCFzixLetmd5jRosqCgiqjKO1
v/wW4HZROPLFkClTWcYdkKtrqaw5wS6lhDPgH0Ldh9jEg2OLuMF+jVdfdmtYKm1TschXHl6Vs+oX
Y4RIxCliQDzWKbN9Xxfyw1oSzy0mhOFNxaOdSaq9Nuy+VGA6RM8+sEN29VZApVskvjFxOFjrV3fO
vPjLVunB6KdmNocX5bNsDU7N/FkO1zU4JcNyQWTWtASfowBBRVUkwFLNv/ohPFg86zqckU0IBht9
uF6IPEqlmXi/a0o5NJ+HseUZF7FGBMJZrsI8+2DX5ebR8hRLB2tZj2PguQxcFfGxEwt0hzkqpwrp
ab0R4X5fz4VmYWdXe50MzyAJt6/usEMqb2YFaF9FufcndkgtKOPPtHsdGLAQ4H8WMuVTgUmZCgl4
GR9hG9fdVRlHPKRcDh3tHfQtanmJAvXosFDTe/UipNePijo/0uHatCX/nzSgBORbvKrh8Syo547U
puVitP7NNsjTOYbbEsxuaueqZqbfRiOIoLu0xUvHEzlH1J56Cq+t0900NHOhaYlE5KuHQi72naI/
92y6ZK3J8ugIYruPISFQUc6MZ8LfTZBgMfqrS5/M4/7jHqLYENHPuS8m0kg5A08AZC/DzFS3LZC0
Xl+Q5oP6Ky6kywEopx/CHzRhLZqLVRAMuqc/PaJZv3hPOMOpH30PKMB9Q5/1/jDfg8iisGvcgKze
Xlox0H6gKb/e74Dzzf/lxDSTqGHyu1j9+6z/9D4fVgJ5g4KGY+mEslnKDeOJn209Rh65flN1eVPl
cyTUwlKU05l00kZhFYiEPL6KhJEAxdsQ4QCoz8IUMqUdK/7wyXvvlWNcZ+mTZ/zOsvhuouFpgFBJ
yywX4sSFuXE47nH6e0g7Pm7y7Y5r91V+SpGP88gKtIMRvEwRIW9+m6j2jDjr70kaf9RWYexdb9sz
OHE+k3PTGep/LogB8W/R1VP5c3tyoXsMgDaQ8rEVAg4sBfhTq5I1fl0l9NEp9JCwJUHI4FkMUX/v
hUbwFXypzBBMqUmEsK5IWYIHsh7x8jHRSWvQf0XXgwE6Ut58Dc0mMCq6AFALN3NtavqcGCi7Ajpz
azToVnjk2uPiEGuJK4lmMWfIEEGH+ikmPHFCo9PvRtqav2ESV3AINt2rsqUY9reUzUxVjVgR+oub
X4co5H89vquYzN+rClUlP3CfnYCwVF7Se3Ic8MurWmixUSSHh6xAXBxK59dEzZYKhDTTx7PfxgCM
aMmiwzxTNUtc4DcJg2EIv1MOy4eO+8btXJlQYnhFWeUFL+YMODu8V6yeHWOqsEBmKLpWS4db4DN4
JPPww5Ic6DFkbYJ4rNEJAYoMatIk90Qzcp0guYKqAQAUIoGXEGv5VveaLt9+RCKZJylly1wdTOyL
1IZWqmNdg6RDD9fjfBZBxXDm8oOgyTzBdo19yfrYETcaZaQHhq0Agph+ZmIxR+ubFBVKHLF9j+76
ce8gc0Pm9MvyiVpo+S5BSSKhA2uAsGqJiUjY0F8JQn9MwahHk/YQe/q2dH3CWfyHVoDmgfKIACOM
9BGjNlmsd9sr9BPp+AMx3H6JRMV8TZ20n7tUD2tjurGuyasAMCABteYxZK0CnGCPMk7JBX5uc9tV
n4Ad8XY+xiNWYZv8aZHzEDQQ+vt9Ua/2hPEYIlh/8r0VG2sVFN2XQh1oUdATTd7Gwyl7GpT8HY2B
KDbE7Z1+x9xc9x7TkjgcpT772h12hhCT1vGNhQqNUmFNT1dfSxFpiHBlejSgxzxOYmVODHLR1NbA
yVcJxpeoVvtgfIotCnH4rz9r3v8uLaR+EBGLoenaj8uX0cjF3dyMid7XjgAJacCWxbK6FPmY9HIJ
NEKRYasAtGygmBLo1qc+xIQkziKZjApz8c0G4ErtKu8/Ay+P/zY+OiF1R82FgtDlXE2t3ySG2Zlx
HEP/4Lh21Sfd0icQVx4jouTriIYFSE9N3BqbgKQ/59bH1h4D+O517BtUGv6EKmClaFZERYouNySo
aMbQrwxLNFN3RB7uEi7W/oM0y1n5fmPy5TrM/U/7ayJivtBwz3diMiiHIfU7d7T+7Pk2Wd2EfxGp
owc2dEA8is8iGiXMvsDwyT/gSHgQuwM4FZtx3TucS0GybTRbf2CRCxhcMycvt5s3lamiN9CrwrLR
hVb2Ukcv6dIkJR1DtnhKbs+qmtqY2pdP11ZANEYP9pFOmWHIosiOXPgg2qaWbbJ1oIQzHcQIg++X
KapC0a2TnfqXfHNPqyuKOWTmSP58m9XyndwaeBnjUOw3pSCaN67x2SZ1jPtejecpoglsjMnPuNUE
oAhhnuvEVrIjNgBW5EMb6+fGlA95fzRUsIo3MXmKz5HbEDd4/zm9A5djJk8DPArTNMZsyyj7WyxG
1HvZTN7w2TITEEztszSkVAJPbNXrSl8Lm8OgsvmC1NShncQpha9K4CVqi5XwHaYJJGPPppUd21jr
A1zbfyxP8hCygOXw+syqHCT93mYOq8+Y1DH0PWVTJ5LjZWLd5P4RJqxCdVEHEDKQOjgtcECLlBX5
gzXPnW8qLvXKRSy5HmUmXvqxba+wiFmRzj8PIRAAx9IG3Ij0BMoUEQCv/lcN7F/ce0yDyls/uNx+
xc7hBdaQpq+PSI39HfjN2aFvYCcejzjlQ0gb9HZDSBj1W/Tg2PJIUAsZFB6VKUYGfzGlsGTaVvXw
s+C6sAC1Pp0pyYgxnECN3lG8lYeb1aM9/HqOflAAqPknGfyn5bn31mpBEU/J4yx2OBlJFNdM36eM
CLw7eQ5F5tPeIfTHsr+VixVtg3jzJwjmJfkv9D0AOFRntrAHEmxlZk9SoZIok8TCzswWZEWEhYu5
IXqAjjLl5EARb1zH/IXOzO4XQI8MWRTIleX1+nZz+ERJObD0zqI71OZRT39V1mfgB8iYUifk+Fwv
JEAeVgLAF3t6cNJCSsePCIHRIBmXxM9C3WtGrZteq78nkMXnh57kPf49y10H4J/b9+0rmF8yTN2U
90MLBTW9KMvSf6QwaGjvBh3XpkKL8C7AkQMSFbPVIPv4ixJCpEdex6nl8zVCzNqGm8fHBcRCWyy7
j7Jopb33G5rGyt4IYFPDaGniNQQAJEKmlzpj3usVfbuPn5Cmqy+rYID6q9tM2gjWW/6kv3T9wYrD
Xa5LF83JSils6TcvaeIvwt1+zH0K9QjpWrES9RoDdIHrWfWdZhOFa0oYsPR4duLJBZXsoj9EG9kY
6OYSkmV4SAYj4XP9VbF2LPV2VplGQjENHYjeDfyTxK55IZMVjpOcI4bllKTSJaiYFdkfanwb5ve3
C+Lt41exWZBRXVtXYJBZ3Gv5xl8EUQ7Qudj3mVmZm3o3iYxf0ZFynwspQNG54lo1hs+Rgn6hqWby
i9uPMIoxSRfJ9gjXXYmTBrP+pY1CW+1CuqPV17mU98kqZoo3E/uTXRaKBNp2YO36EBuRYHX5+Zp+
Ze6+lf14rbdTta230zux0u4hONvIRjYT+S9DnOz/hL9ynhHWN2gpJW01AyXbHlH7Ae+wTShcTBDz
KhJ6PPLavWZvq0rZSxOLYtL1mpeIODtajdnWH1y5LhPPtMtNaH9ygxvSBnUpYX1+oWJSGkMbc//0
+O21dVOqPldY1cMnZrHlQwbMMSThry6d16sIDaAk/jf/eFeVFFM02gr1q8V5htNBfZXeoKZPROBX
QValb9KlpSuQivg8ZvVNQ5REaeMTl/ITrgQzJTndptpFnmGCllqXw8Pq1VrPzsVp0lVQCnAyMOE4
vLxXAYfwLFYMs7FYzzZ/FgNMCSXS2V3ya5QmLqZn0Wa660qEFPOO9XSEp4PA1ojdA0ylPGjWDBZh
GD+LcBbbxpLzlldNgwIJguVVxQ1eabZTlhOshVZpiFZasRQUlbCvd9ecbHEKjr4IsxmtmWvll0Md
wwlRc8Fzy/u/zU3ob2j0BHBjPw7MqtSdwJqXeLrjCG+SgjiVWvt+Z9435Eps+p9FuQD8V1PtzSlT
oS7I7zYsjPf8LfxG/+/9aizRttSL1EtlDPZlN0aDrs4+5ztCjKobe8onUElMbFBHgVDDidCmNNB9
H1tgmqFFjrHJtOPugexKQ3anZy+a4kbRw7Oardp6jWntDe4p2QgK1ykPx+EO16qesWUsI473bBfS
vRRfe/Ak9q+wnRY4zSw2vkuSnilg7MPBtuUHr8SMW/zSufgiPouvMakaamBTStEQtI8QyTJhBIdk
Uo95eMv8C0d0G3eRDDCXIhNsftQiPUUvZKF6AqciXWR77mdDCI31HMqzyb9ipzXrRbI5GlPqB/z2
WvE4q5GMok4KR/QxJILks1WymCDvcp4K8pLq752dBE4b7zdsynTuBAOJ+mGoDIq/+xnaswMSXRiV
OA65am3Loq5ujvE/7xANyY3fu3PXg1qYY0VwLxy3TWE7GOoBND7vBFP327S6b4g0ntMxjwMSAExk
VQcohO7HzqaNjtu299ogofJRRH8WHymzmGJmxzMaTeW6E80jrw7WXYkNECYv9O8J8k+G9M7yUnYH
97xN6vchmi2bLFCMXJ97tGwAAkDM0Tgknfe+/GYAvD6/mVx2kjzHuHPUmI99kwUSzEkOF5W1+vUw
YLP60s2pQqq+goNTH2edTWJqMHBmAK6vY03qE44ldkgKto0GtTEYkbKOZexJkHg0x69MuMsjDUlw
dpzWiBe1IjYAyEMuOU/HQXGg59OHQDYtdwp90dCG8lmDv8y3vlvL6KpiyMA3ibd+D9r/fuVPKIM0
0jy8Yib0bk0/Mjx335+Ye5PgqT9aG1wPufajX79v93AR/nntWA8EHgJa2vprFKGeJhuFAnL01INA
v81gWXn02whcxePAwnOVbbI8oR5V+0cnWfRDFKRJqnt0lugQj04st8Pr/Wx2n2s7Yb8YlFAwBAd/
Qk6Vh7nemko10XPlIt4kcQumCeNUmIa957fd3EE4+B6yajh3gixhlgwbmW98HI1ey4Ih5MKJunlw
EmUbyXJ5xvZsT3CKNmPx0u8Lia5lY6kpeigyyvxKuKtzMvVOh2MWqPIee51AQhmNwWOZoi8+Qll7
Pq5pTLoiP8v+l5NaGe0NIHDuLwsC7dEJgnS61y9N/I7Yuf/VJQtcOncPQFvTwxTh5SrYjdk1UtOZ
REOoDjLI2LhaVtA8PBD22zaCBYoMYu/CBN0q43AJH1djz4oDMgwDAVBOP8tseG20SpZ/yF3AQTvz
Hxe5ohh/rz+lZbry9v1kPe0ZhqFFTQ7YMjh74mguZZGUej/Ja3hw4vjcK0f74GWqhqCCqLe4qJqn
Q3TpQxfyvjHczPKKPLv2zpoGpETMMQrANWBO1lM2yL1vZ4GkMyQzE1v6IarVRT4/CxVWe1931Tjm
MiKQKzkmF93vUAZGgGtklFvvw2e06pwQ4oLjSvN90qbne3D+bN1/b3rYPxOXc+9wy1aXEAVTUqOV
q17sbmKp3zgehiA2ycgKHIkDzhgyP2eM1nGmTYFIetdpeg92d6R8uHqTG1Ds6RVpghETMuS3mFvn
JOVPuqy1UgBB2PvivDVrzZ/FcM/d8mYICc+dTVxHm2s8YPfY6X+Khc8zm7S3pgN83R10BIfNBdjs
U3wjn9+mVvzYJAIroQOgoPWS+Ow2888X+EoOiLwV4897HfqitgXsv2l1KBDOkIKBZGuW0AeIXOGR
n3h3K1TUSuUQKEG8W/odtL2+Xi7s26N1ZaNRVcNtXERbBe5FtKqnVRiUGC23tgTAOXxOCyKSpMQA
UCfm8cHoxVV9S00CvLVSPOi3rbrnseNY4mrAxHhsXts++B+L0RyGeKDB8c6i3eSAnzMqdU6IOzsp
YcXDxGS80WCYUDOtaJTocJ95WKXSarCuIClH2FSSwyV0RbMDacGmuZdqb4dpoP8H/D+zRVErndjC
IUS6K6xzMYyI3BWSlOYUkCviBCQFsEsvexBLdVpLmQZ1egcq8yncTfQnTqkqyQSbEE0+TD9oG42c
5Y+6iRKjuqHb/olBrtdWP88syyGUU5szcw+gy7KVJUZ9dnsRV3ztXuliUBdLQmMa3RbNHKRgq5qT
BfjWrvV0AvudUBR8Hew7jFesNCbw95FyuikcmfMqfqKrBILMcWGdmhUUndRlXQhU99IQxHjYxcx6
qINmPnKAvNYNJdiVG5oNfAQD1XAt7c2c3FPrCPn84Ja3PHNlYN1ZPwILNM8iL7L7OUmspqebrXc8
61krz5kKc3bF6K7YZoZJBRF8a6FGBM50EMOsSTUt8sHSl4gAPr+ETWMp6z2uyqIehVmxZBLY3fIO
iG3KV37TXStPioqT9ivvSvKKTxnFUDBIAH1ijqLxtP0DE4U51hsv6wlj0Yj1BDODlYxNBIYq1HgU
z9BTQQ/xKjRG+aUgjIdrRAFXBSxb0icj3nYZ7+i752TJn5wtju+uH7Xr1B6VIXQNwuPckhjV5hTl
KwRXT3VxwHO6GjCIewdOW3OgPUJrqVD7dP2wJi+bF+1py4LCVvO0MHJhsuj/dG9uePL4RtlDph7O
sWYBQ13W53MYIXBEwnog8abYJbqiO6ZoC9YwhKjHwAeKzG/l85l5hISPS6y9EaaAFbXdYXUR31tJ
sSgmTBse4jBWFiw7YSlSK/pFXmSiCDbd97EQPyyslfSewRtkq46fOT3MB84TcVf+b4/5PAhbDdax
gfZcnuBXqQ1upfgmbTAvGf5EAwCdI33bloKB4eU4UQLUp9x7gYe/+NalOlpBLLbxA3+Iig4IesK8
l4XpZZgINQBgC6gqlEv1wyMiDcPak1pxGHLQzUNzmhaGKqJw6xFpSqSlHAFHQlg8Z6bOpwfgzvNp
BbLleGyQR/AYG2WHxFhY3gT1TPZIM7+skV5DDfV7niDk1dw57JY0O0SEcKbt6QSSwNKQ2ypRW72R
fl8+IDcpTD1Btp4g+nnZSWXTJk4c1oPncuoRi5GRjY8fgPa3jN5T6fp9Uhsltq4vI6+LquZ72nIi
nwU88CM4NalgXde8W6xL/ciWj5aNzDFOMmLuC3Nu6hD30P9IVK0u0K5S77kiCbCSLZaleso14QbY
YYUN1ik4vcFqyAGuI539HVJXatrMQJDKSiy3+AoPIJh7bhnzskurG6kBcZNCfEMQEwx4GG7mo/Bt
aiY/x7+hooZIqK84VfxRG+gMI0bFqgGQQLFwu6nZLxmxDgoyjaYeHfUHWyRWUcsiIlKB5uBgDQ8f
/c5laFFWnLT80BKLHNhQ0uLYjJwViSaVg5WdY1DkNL5u7461bNnuqyfHfC6rKpeQy72xysQ1GEyu
Dc0HAEPrn0hM8NOgG1dFu1fJwP/ijl1PEFp7ka4QkhBo9U8grbQr4fuXYFWgshw1y3eAHc9NC2Es
2UHLPYc8S4wdVwZikEbiOSlij471zGs0uO0LL7XCDAUm+hVfCoMqYgHEnUhBkaSHcHlM8LD4Cu3Z
vIVSXVk1HYf+OZSbBCHwLOR1iqWxbVPx2WzXqzlDFI+Ef/EulJxduPCRD4FUfNz04+Z+cBS1/YyF
/1me5SgX+lXwirYV/6BYLHZvTL+EU4W2AX5wG9/jf6AopTJbcVdyMs0Q/wcLMf0b76LId0c+2eQK
azJGfJt2eCcusNwY0Rv0pKXuYa2vSvdOEiEnQ8UHgWS3gq/OeCUHwQgQM5exb0MvcbXCokwlIY6N
ouJxRu8J3HmYw1UMKBRzQAHsNAl8xHq2I8TRzU6VUAOaQLdxy8WFibhSKQRGZ7yv3Fht6qfg1eYW
nwOebKzzfZDc61aVcQaYlsUGbvpPJUyKhtDiZ0a+CegU0E5cZezeouhrRkMa/UslY4i4b6Wqb7EX
ldZHmKHsx+xMCWMVBOAoPEYkawSW8TtS3pcrwEbt2kDoWnRH2NGbYaEfWjwoBK+rLrlfF0WypIe/
ipmcu8Zeu/xPM6VmtfOYd5ZqSZ4jY+6BHDY4dmemEtaCrNRFxx/7/hzVEQY8A90upu5MeR23HHWo
UsygMf1a1rBEFCPMjjZqiLpqqCd2waECZ+nFEd4mpgzeaQ+aA3c+5zUnTgaeI8lwy2Rsut6St4gO
K+u7gd9xjZQlIvpvlmtH6RlwMwd4tsJrfuwxilvEWWfX+8hOslanRb2clwnB8qF3FIi2wcch0vkc
2TEFe57/9NrckzLmEhYPIz1YgsCmYwsiE7XSeQoYMPVryetQ0nhnxivBS261XuFIjJ8gg/Xmpw65
kNEY3El4aMV7QhvY7gx28VOxje1f9+7IoZYVfoLof1CwBtJnTn68yO7hFs7RMoc/MRw9trKE5fBC
fq5vM/YCDAEjVTIJjgSBnHyw6tNY5QiVo1PK9VCdspHSnrQpHHBWLoJmO5ppjVthfaZI4j0mQ5vt
QSYTAMZeVm35TYLMPh7zAWrqoaepGJwKWxuThoqtdwkdLtJvUMXYt+/3OpRYCDiH6BlCp8jmEYTw
4vCjw8idXUhNprII901NcinHrIgZM989b6MbGY7T5MESl0qZtJdiXDN7GXcjq5yUCQA2r2sQQdrn
5MHjwbyop++QhIwyXzEkzA4P73kzZcE3T0oJjLNaePTshNOILE1xi+yYYJX/j0twBi5B/uMxiCZs
4dqLNOnCPqcGW8N6/umHUwcxVQoigoeMsgx5BqW1kxTOtU8yW+s9VkX3NxLsFrHYv61Ha/N4rm/o
iiU3/uTp8Lw7zINLo1ue/1HTlyG61/75+zci6XeFT5jyU/6nCcQ2uO//BvbItrXqsOAR578B+CIP
1HW4WOZuUg/GcCf9FGobRP2nEGilTHQnBomGTN7PLKa0/vf1GQQVtb2QtIIQhT1vkEeWunwo58MD
x6hLCvPrfoU0ZZa1OGBbtm1FNQw3A3u2/OXRdASpjNepOAG4lwNHFeNYYpSTYRiILUn8yng+uYrf
RSxafDOEOVYSKhDG/ilm2SqEbWZeRH3BsjkcmTROtRnC7q3p7VN5vGFv7JLc1axH6UOxFepwlIG6
QyqtQpwmZp/h0jZVcvt1uw0pFtuw8aS8VwlaVpTXU4O1C+l/i75pFn3dzy0ljlP2vWzghRaS2Gwq
MXzk2StxjIaRoQ7gG1VCcVqIObJtMY7KK41UAFQyA6tfYre4YmyWCYb65T3OnIGIb9hhEmXDWCnb
mZBepPP6oU0G72uapzQv+a0VvKa9HZz1KF8kTSOtsOyXaAPdoQy5cSTs9hVA45xAir5Y0bmoWEL7
JdWQ/EQ/GC5E9IofyVp9Ik3j2/eENXbZzXikcej2s7aSjZOg9iVpmMOcq45tKLT1uMLvY3X5+tok
8ZN9GQfB/5BUs0+qSrJf4eYMkn/kLdNvXusuTjOpPx9/fzQAh96oY9ttkxnVQFOB/nnRTNzRTXK5
SufE6ye+1q7y+ROshz9APth+5aPbyBC21ZZEbgnEqd+fXLKJN3nlev0ZwjeHnOG2vImRZNhHkO5k
+gyydlkBgI5nLnUW20vVHJCrCLbLIhdfWFXhs4CbCylsVIqdvHNs/I63YvLRdGGOZpGBUBUYYyek
HopqPdKtafb04nMZYb0q/CGh/L1w0HMcD7UDX+GR8gckO199uia8GQcl0sQnoyz5m59P+CWEQGhq
axd7IBIBW0Hjg70L0LLLjlfvls5e5HprKbj8MyFGpWSQ+3WqwKMgup1SRTADHGM0EN0qHEPqb9dQ
hEGcbMq7mMHKKPVlKrusMMLGA2efX1HkKsWSp9zhONe7HUBaJICQOQUu4MbuFMevjT1tEAojBpyM
xUGVaz93Ki7LFmNJVuklL4YUF1nR3KVnQfwD3ICiKejGmCJ47iokiSR9Th9B422MCDf+3iUlJSvS
ScAQ15k0JRMAMMZRY8VVe/jwOpT/Ej4dyprQWQVr8BbATIH6vTkJaIMW6kiUIJkSMzle64YEIZMw
stPruY92D+dzamF/oQsDyJqip/SvZ63LeUU6c6g2g19jbPvo9MOJMaiZyzwWChx9G8g5UzJtUK3g
mGJ1N2msSRi5SrxfWQqYBanLvRlh2yHOOXXa5fPmnB1qq8aHetUarGIdm/1sA694QM/yjQShnaGR
q/nXlsNXeljcPQLYCirbeOoNUuYJdrN4XTt5rJzgzKVz0SFK2+u2nJ5pjzmXI7X6FM5FEtLnZEqJ
xqAyKg807XneNnjkWdqT/za+u3n4H+xzKmDCXwxLs84EVjlozMkWUeEa1DmG5nLM/O8eniPXyrTA
E5g0pjqCFH7Dbrje/6eDOUbuI0EIXkEzvWePHeHvSe5UK48Ftund5bpymSDFyILbVZZODi0f9IdT
OolWo8bn3LyLJXi7KaLzPUVtRWg3+NsStDnBikc5HinQeo3LiTnVIEen1KLaeR2uJGO/yonjo9vF
jL1P+CG//2pQpnla8sOZ5RlN+p7FZBL+0leTmntR4QK5szvNYN91isjmASDNsGfGevLqEXh5+cy0
c86Yhm0kMj8krxlraEOfDggDn5Em7VeYX21JPD0SwnbM7RUUXlmcucXlsKFDBFy5ynzurBJMJaQc
j2cU0n6QNtQGhCBhDHeWKKJgocHoSTpFtIaeKrvl7VSm0McTVnCvYhOqFTIzs70g9WCAOWsnPife
QO8KZ0xYV+YsSJ/TkKpKQEy8hF8KLTPynug4LzmECsmVH+k7B0LJPNzv5DxKGuuUvf5pzeLxfiVg
KK6H0WpzwFYQePY4EdsWZ8u2EM6Ojb2QiECnJBKEJtKEY4q+HXokx3Y3oVIWq1MwGZGg0p8KRJep
QOOVvbR6uYLSIvD2uutl4pKs2NDv5Wtc5yhBOTLy8//feBs56sm0zwkOzxCH82FMcmAHd9tcKdUk
BITE2MfwcDUU7a23wCcdM5CJFAiXJk/wzh13zvy95Pv0Qq6+6KH9y9btAr5f2z7VJIaXgxG4nbiO
XQwOr8tFYlWFOM65/ZgFxwyH1j3zfUfKcrIz84q8jYC9ifydNF/+Z7m2srI3OBB2++R73gFobe29
Q8LdTFgBThLqRD43YNYRQ4AVrTg/PZv0WZ7e8yWRRkNez+OPit0sMf334eFt+Ane+fx7YTkzklEW
637WeiUh46E671R9T3eyPHv9njORO/Lxhgd+iJMUCIW29i8a0ll6i8T69B95g8ecvxtdZs48Bf/6
OChBDHknnVisWyzCdjr6cgOIwEUMSFfW8FJtAyeguVmxnUVfRIbEkhsxsb42ZcytLbbdwTWFt8RQ
KNRXwKHEKdE/eWMD9oWKAaECWUMNXQ2v0wAd2ICIHh5ntbvohkFyNYVDNlq4OQ34cWqbDyZreOFO
u+WaX9XQwU2/mbgD5k9UKvHORPnjuFovRajiI9nDCa+Q0qvwyCdBWVyQHnZxmV2jAaPtQ8NLBeh1
OnbDTBxHoxTfdMC/LpRUmZyqyGzSmGrEIPpZbtLGCMoE7rmdZfeNdt9Zzy1HBm1qjRLasV8s2vTH
VlJHceIkPqTOpCzIJLv25UEF1cAdBEpCJn8H29SR/QiHACxOcNLnGO79Jl2kpd3C5CBEpPwHtEvA
pOAfQjGsRk4O/hztgPEbDrpNa0OPMXWmgqe+a50B89c1Zlmg7uMVInwegFfnN6ypucilZBk9DwEn
iAr1TLHUooKbOfhC1cnA25I7KceJ/xx8Dd3SmFEFKK4RF9ux5HurqaaVk/1FUS97wNqKDmkn4t2N
hzEpbRb9pyISy6v6xiFf9IUAAg4vo0NfkaZkmPMtg41+48lqMeOzSXCOaCkhoqjibFTlG1NTYxi+
yJCLvDPxAvjvASO+mVMJsP/CAQ1y7DNV6Bbfu8DjoIWncEUFrIdJyeweHGME+hDirEbbp/LegBZj
/3sRJms7nn3yJ7DCbAWarLSDPX7PKj6N5sXTjau32Thf79XbFPlf+iWsUT4GdtjkQzXqleeVrEPk
l/3oydLfPjA5lbpO5bCOjuT8ZqlqHRPyiZhyut/qUQ2XdOrjTxYgAo2L8iBFcqS/W6i++Hp/qWKW
ISNW9mBQ/WAUOxyQXtRVroM6tj7kR3OHd838scygTfNmQoRHw+fae1Bzx9YnPZuGzUfPTDAvur03
xvtNWBsRKhbpJlMc+1gaXNyeL/ZZW8l3g2i4GbV79NDHqEh7v/Fv4e6tnRKfw7ay62F++IR4k2e6
jUNqVzlUf/cP5J6b50/98Pk5UK2+8pBxXG/p+EY6Yls/ll2++/Z6/iyc7JsgLNqkObLNEAQXq1hn
LTCvreQBeilp/fw/SfNjnYrhwhyYR3SaIPkfytBApEVGQJ38z8r1b1abJ18ETiw1NnaADvuk91L0
e99FC1oqL+/9tBdvEfU3GkfhtxhC+rqBKWIYyAzRWla8FD2cpQA/h35v7OqbhAlFvoVL/x6ajz+O
bU1tfjLlkwcnL7TIr/8wfM1DvhXfl1XSHsVx71Zq6XP5or5Cuc+kiPby93jLhnIXwj4R9sJsa7vJ
e3uMYhtCIs9V5g9RQ3ALqTZsm7Y4PiTKMTi7yAksZJfcxiZAROoZ6fgr/w/resNFyhUPLGlk7WUg
4ZOvsoXRUQAhsizzqFaYcWiJ2CWhopG9AV/97jXGY4XEn2NHebI2HELtS4UAIOitje/f33O3cDHj
tPRwpLa0nmFi2yUV9gKWoj97neMpx8q4QhpR0YTOLWQr1gotvJHmDpxmQxdkSOjvs3pNqLN4ygcQ
aU6TO+6v/IFaIRWviirWRBVZLYZmDGGj2SZSHB5ECwBxvlNP4DZVso04yAufo/NCzRjWu0x91Hwy
ybL30m2vcyjRBC2hwTvWgkCigWotXfKAOjha54PPKRllSVvgI9kM02x9ubqN0H4j9mdwK7wNKpWf
wpB2bQmVunMwWkSNqB2gh6DEgmgjzFzmOc5mtj98v701xhXgarxtUbdxExznBZBern8tQfdpuUWI
P3Sjm9RXe3RB/vaQd4CS8wqseh7t7QNP6pkmuWCLiZSAOwMAM5oQNdqzCu9JvOmlqLNohzZJzdqU
1OqANQTGDJlwxaqHJuioAuwfeD0iOOcIehR9A1FFT+z11zW9gehNzYLpItZBKcZTKX1eU/NY8CtY
iiDF4iYkXs8w6rz4nSp3ZXcTN1YRBPKV004DuZrU61iraUPMmSn1yYhNi+ZnyuaH2EhCrMMsyIMc
rogfNBkMGlKE8uPTyDgVcjQ+hCAKti4A6RqjxFfRC1p4dFFbUHVzyrjLuyU65uOg+ClZ1uyVdMEf
YOws+dKPwWbQ2Cc2FtQgHhp1FVQ0BteZKSvYuiORQ2ZqWzQuaQrpDHbpHWprmHxXekpHLwBsYS/D
efnniKh0dJR3vX85Hu4GUrgNRzDaeeGNP7iuR8giNCl7e+7Y48IePoYQv4ptDv38xQLkffMtDH7Z
cLT/Ib6cWxm7up/j+SwT6la6WFZAm44TDajuPNqJLzJpOxvs8LahSj5W/msoX1NAX2maYiLBvQIQ
JKPD3euHGZ7kRBuHsvYGGXU9PuLhFg4Gn7+VyrxuaJ3a4BD92RKP87HnKtYJL7RPgdsbpxHEaNKi
Xlhnku49JKf9xzpGa6R+F7s68/ef8HiktehdkEmk4tHBjmLTvawen5DXv/IcDfN2RNNqgKNwptp1
URiQtN4dXUND8Jju4UZCYCOsYqDbFzlO10e3M4Ou2aTNtyJacpL64GVp8OMgfqZrLt2yZ90ACDyy
s1etoZdsNOVLn7RgYFvCw7O6iRRzoRhhfQx5fZukQn9CFL3JLtBqfvT30QAwz2S9rDpeYs5q9ARp
75E9BWE0kR8baQigJsJTWKOkI0JPwwiUrsNfRCzbfuAlRcydFbV2lTAdUGg7jdxvV/L8NafD9cBw
Z1gaw9XEv4ageVdVdGLxXnbuFPyWQewbw9JZsKJTPPcAmKpIjkMkOa+J4HRk9Nk4udgtsaCNlLS0
oO/0wunRnUU3RMUPd7dICSQLN0lDGNZuKB7UpKXQBzG1wzJvh4x6kSUac+Ztt8Uhh03xTS2Nbu39
B9yG7Sj1nOyz7YGgYczo/0bv28l3r62eUUcy/0eDeicUyifn6nq3cd9u/H4WlQlzrNNzbVzAtCca
6wnrLylEAarCPKL5Yd1HoH+v/fFCHXoF4DG+Pd4tEultPxLkjfYudUuCB/oxeMWB+ehvQxQIG+dM
DHIMMFuXGKi+jgB8nzIkT28HQOzLPhYPSAiKUX6aPjtd7s0/pdvpIaDcDHch5QbhpDRvidhXY3IQ
2Aq2b8kUs8n/T50eYG53ab9w17F/FHG/mzqAXrPED4x87PyCZ7NT30fMLZY/ASceXY0OsKFQjTn/
Km0rmCk0/z50LAirZSqbIWSOMzn7LcrNH5PjP3wtcxa5O0TN/OHflh0BhWPFFHk+LrIgn+zYiYuw
gVHyGc84act2SJVFb0B7p4k+T6Xr3jtnaEVI/raaKB96tOafmW5fNh1kxdgLrhhavrtMEbUY2wHZ
9QKFYO9SN6yqM6itwHSJGpy1hNm08B+FXE03h3G2RXxnQT9cyIz5sUjTm3iJHoSxwWLAWqrp6ZrW
k8K/lAdMCfCoYCutc+z1fadBfvGlzOimDPDR6qReOWpChRG3D8Sr5Kgfa6qkKK8WgeXpGpdB2IV5
kns7HW+aHa/88ekIf2Uxv60iXQ8HR876Soh/d/bO2AHAMii0L9xhsWaAW5Hc7MbY4J0cbWMnLr6Y
+0iDHmNajknr/Hq/LLlkevuUIkvCX8nsFktQqxne1xIPnMLxaPyykv6nb+sBXyaEkXjPWzi+40m5
o4Msg24ff1C12PPWHocLQ9jqA6Q6uaccMSY/NvqfWylWSkJcvU7F04OociT4mYSGW1VIeqipSz5E
7TaiDgQ1fiaTZ8eCip5H0T+fip7F6cuILZuZ3u3JBGCHJcwWjmGjjbg5Eoczn2eLO8+b2wClMS9I
UP4CbwobTH5LBSwGbsVp8MvZcujgz8AAb2Rhr0VY8Th444SQC5cvVprrEp3XWBBGZzxkbDaRGjE0
9JM/nihmspbW/B+P82QcLBHAIAA3KYIWXka8TJUUExfzdA/QaaMrnIx5l4jEPaVaYk5ubj121Ujx
9X1BUV/dYcyJU9Y9dLsvVcE3oXYNdYil+1Hf3UmyLu+JHiq73fETPQZZMITZJOpjMFPVUZ7ehU6t
hLeahpyZpk3U6mxRP9jPgbkZ3B8OCg92T1m47T8kZ3CIxlAgI5ZvXQhOgZmMy5NHMcOnbCph/WMt
DAp+8bCkaCV/DZl9VSQ9PpNaXw0EgJv9lchiF4d1psZ4O2uWCvxYz/xYA/UMLOx9a3p/fedcs6JO
5yJMg2SnVdvn83IPDlNz7Cu0iLHCm/tyY48q1D0L3JdkKFhbZMqo2yasteWYVc8DxWJqNUEsMCVw
qgIj2UIm2eURfllHhio7s5ltu40tu4po5qAOEoZ5CyzfjUG3LHQgyYsPcWc7ZhegnWCLgQTmo/3R
HJ8pkW8jfRYJB4kadbzEo9g3vqHljNDPZbvgLmLTtRwZJKai9aVyfGiCuIevalG8vOulV4mQJhv5
HhYuasaL4JmqZCeoPWGp9ak27rPsEzNbgemxuASROiz6FsOU2pxKknxWvuVOGPb+hYV3/CC8peHQ
iU2Y6C5hwA2CYyylKDCwcSWixKrSu6EDmWtwIsBzzZ143LTj2XvbOA4ZfhEr4EFcW2/vKF462X78
hzbp+RCCHDncYuvF5vRQnslBYDn4W3Zgk1ImirP/CGg7truJBzKYMAy0i13Wn7N0cBFjfNJXGbvg
CrupgsRnKiucya8ApNQii0XLrOlv0nThhA8zBk0e0zTu0epzbESAy0DTp6QAW6SGqRwwl5qhFN/S
GvI+aVSDvJ47P//conIkrF5Yk62nE1KeJkexUIgQmr+ZwTkryU+GHL6xo+eR2rEbBhY0QVpDCJKX
pM5R1ZEUBFatQKU6zEoBPnzn+CbeyEVmwEa76xgt1iryulWdXf+/BSCSLpGARKWtXjaSf3PPbPyi
mWRhwOH+wrDJeA62cb1MlJPwx9xnYbBGa6EOZBVxvbpLnjpF6Ps93RyMlqt81bnKUw87RPijOKZd
5gH1O5wJFFjRsA/HQ/nUN7Ix0oWIz43szq0ohl12BX2HHsKu6TkhAYdLWfP7krfqsa3JduNi+90Y
JmdBpTnc0zrKrNOQD8q3SDtpr0z8icD4XF2Qn8katC5rYY/YUPhe6f/MXDZLQQsjMuXNRZ96f717
sSorpqbVedihoGW6F8ikLc8ns4uCBy2elLhy9gTXZ3xpLpuONhvUo+9P/kkcZUYF1EWSKC/WAl6N
gYOCnGL44DBCNvEYOerULviqKcec0a05yePAnQ45iucSP5RA8e31G9FYFnINlv0QfdB36aHoRSXs
fbr4CU8MR13N+ixx3bf2afmcgrecYJ/kuE1tbK69l3A3CyOkYAGKlux9HFU3q0PihZdohm+4dpu8
Y9hDRfGIdz7nnEAeAwYDp/IAwdOizFApn3F8NIO9N+3XhGhmHsusi1+OJNqcihA+U1/5E+dPwA3N
S/HLgzaYD4SXQ+H+azm3QTIzJZP5Twe9pMM5kDNcmkN4hx3FPQmg2SREmSpkzSjAyraI10T9f4qr
XmHVxxlIJOH51gYc0cG4NJTWzz6B/qIF38Xtc7ovuMiHHfIc2deoZzrQJjkvrkBI3/0yhGrZuFDJ
tUMejfmVZxq/qrpMpc25vM6ROYccTKCDC+NNsamIARnWWuQCp8nxvpCZdKzbA1g1geKSG7NL7fdC
hqoAICJLNSitEQR3RHsCmtEJ3gS8b04tugb9Eyiin4O5JaVxOvgbnXLPJV/MtciI2VhlcBboi+uX
OEi0xMjw6Ib0oYnmKSdUtzsukw3NrNKy2L32GLkD5Smj5RzAj6EjbdR9A6MBpQlAZzuaGdIvMgKH
1jo4lLzOUVEkxTtBTajyTw3cYx5Q7JOvzV9gJUsz9oy4+8/cn+aEtdjbBuaqwyfGIfzF2wGp4RsN
1Rpi0oLqAE98Pb9QUwlStIo4j9gNrClVLi51MryF4f+4dDHD1fBr8R8jwQxse2syH9YyPrtExsvN
49t+1yL5hNZOKY962DVV/QuxM/KrZEx0wddts8TylswImw0joSD8Uthn7Qq8EL8sN9yiJFWUXDWA
a6WLnNJVqqNi4nYR9Sy0dV351IHxzq8Gmp2w06jSga50gaF+f6HOlFKHmDwwFjaMt9nBXeEn/bvl
fOOHzrT1xx7oWvTOitOlCLXYHyRqxcOQxmxopML+RCVecOraee2vo9RJ9Vrz3U4JWTYVvCrX/PQi
juHwV3bmaCbYwy7lsOzw1qK5EB9iII8W3DjNTGh64r10cTkiKyqIp6aWQtg592U8G9hHEWRhTFR0
By6rIto4QBQoh0Y6TGro3avFebw3i3hoSMwqkh/jfrlNPrI8duFx50ajpYbYN/uv8+oEBWQxDrCw
AAxjv8LZYn0jpunLEiZ7C8o/Lkf8yyX4Ei236kqnYH7+Sr44hgc+GVGPW+KGQpemQ6GYDhQCHUu9
xYI3JaZyodMIPdXboMAReOorDI8ASFtzoE+P+kRlBbkMwkxCyq8h0z0qFq67Kk045Xlw0WXFdPJt
r6dVMsihjhLsx5IssWb/dDYSKBG/wXFXFfhmHniGWC2J5tmjhou5YNB35ODgsOln3mMiiRk3w3zY
DI9eGvvjf6zge58mvodHGZZQwbTFdr/54tYL4Tre8XH7JdzQaXownhbLZDIcPXu0kDJnfux19q48
waeoX3mAhjepAbYiXS5dp1HiuoWyyy8SXaMFMI0HK3rJ8Uhl/OsbTSp/Z10OF+e0vTF0Z9AmA8v/
8WguDpHiqU2HanhyfJyrxkusIIhi8P5X3fahz/4j4+OAb/+3Bzu/FoTyeZ3pA3UPIFiOAK0JkCJI
scB0jHYAKZbYe9Bq2iQtC5qk064sU+qn6QfCim1tF6THySghhckFQ04bVIUYTyscS5Z38SW590wH
NDtdLd4rINLn40l+FkzvRJ05UjpEukj81MwlKJq6OWS9gWXLFzrzPd9DdzOzbK+VeQYjBYzCYtMw
pExw+CES4yGHJh/HqmEwVMty6JLEiB4OLG6Vkay+YyNbdKOV2Y+63++/7v/owBSHBi99ah4aJDMa
Kg2K6YUvg/Dr3zVv/rB1q8hqVpQufhdLvMvRkS/adi7uzAa+lr/gH9OGng3xGn8VH9N7bFoP3B82
GiT4tlQfNiiv/44vo/9jSAh/a53JkOCaJ8TU3gMxde/mZANeGz8p6J3zy49KE/iOMgj5UR2L9Shq
lwgO9oZSY3jlcyFx2RB6EdJJDBV6HDVHckZ4ejzYLemjOHGzTgm5raJvaNCrpKk79DFevid27x/N
EJYCulp5e4MgfoZ1MMjYalAcYuXkq+tXzqlGqdI7XqnprevMc21yCl9SOjcYhWLipO9b9NXoelNQ
m8PNwiL4nZsFFv0uRSjhUS6eq394I893JW9HEr2gRzFJynbnkNgM5VIsdq1hSU0va+4WINvasZMS
N0s+RYttv5LArvAdUCVgBCSPo971UksIXwBZWihxJLZ8TrC+hk9ZK+Hr7fw+QlnZ146GG9vI/4Or
OrhIr1a3SZKjYjWIdxTtbMuErpnM5ulKx+D+sloGK7d5D2GUHp7lVjnzerREKtK4nmCLFr9zJEV2
nFEXao3mQAteaO1u9LWcaHKQbm5fDZZYv/xJJNjLzm4DuC11M5Veb3NGqkH2IiQ9TQ2jOHEjN+FB
OULfmv5ub4VRJi6TjIu6EFt5Fa39BkMZ+gwsnZIzts7w8PRhsjsa3psAyi6pllWwAb7I0ZAEbCSh
bNli1LaHnz8Mhp9YKhGhCLCIkBn7fI/ZPlNSTXQWUd5W4OnJLHAsIAMP2PVFbXVKUlAdHlctALdc
bIlz4KXNHxfu6cRnXHLYINzBsiMtLeHyMgB2cRnAq5UKqVYHth8R3aMb673g/eRPAFzoNo9/rEUx
1zFHamxKGvd3hPo2og4rmwfWl5hs42q74gXc9d6BWhR3+iFbe3/c4iEuqk5rXaOd5FWqtpKCkDfB
AuVWGt9gvb86GmZ8OiPhIG4uVdNQEV3c7AMjJ5Df1zNzE5IqxqNiIHgxJLlddFN90WK/h31YuDjj
4g9FhAZver4Ngz+e0ghNR8C2MmfEHuxTGizzE5kSEYNi5hhmNWDJPmAaJg3U61nRHgIvyit1B0oq
8IF1HxV2agrisRzVIYqtli8MDdfvMooJP8noUFwNrAM9XbaV38dSVWgnfuRSSeW723+3Vu0XlnlI
JFA37HiJP4sI97qhzoHAWyeu30oPlfveGQMfkZ6i4a+ieh7dAgoH2QTY+HPQgtfsV245SgraLbPT
1PWkVDK9f8YgnsNsWakP0i+GBu0A2eofPA12dS521I9BZs/uhIe7EjDlHK4OudqlwdRPpnoFcQUl
+De/Cgkgono79JdnSnH1PmND3l4cQ0Qd2EogskYWOhMcGOcyDuZ6/ncdR0f3+vo148mGtStn2W2Y
vxq+I1/VIdKRbv8lsDnBdYBoQt0+8uMkaFERzeWGQuLILJUviBVHUpN7zZRxpxSBbpaGM9+n8qqU
0sANsdYFznfjGp5vy0otdtqPropQlKcZSaynyNQ4BJCZczLyJYz9vOlRn4KS6pkdZP7ObLh7aB8e
aFtRXXI+qRQOm0Cnu6DxdjyX73jTYkz1MDgKmxx9J2U9geeMOfPLUJdQyKzspa4CwBuAJZlpNE3W
RFq1VcXXDNastIQrR6lsPaL74MQfveMwZUZKTU0YCtZ/IMlyOgrR65MJ/YMJZLo1sO3yOFPGSvNI
gdEDgY8PB2oojBk1CKQiEcjG7e7flsSehFYJub+qtqCogRHyDBJiarhd8lcUxdNLfIQ+XOfTpQp/
rrPngzpChOgVJwYVEU0QbuPYMoX0Cf6ikwVyIM9v+kuhTFwpiNLxht61gi9U/rSumJ15zdSSAXZV
Y0c6r4KWCjQZt7qd1Ce6y2zHdECEpARW9qH3LA4cVhdMoaPTPlOL7laNirqxXcBCklxjnOsBIWSY
hUULaXISG/YcjRPKM1NEtElgblIVv6pfQQJkQjL5Xlsew1+i5WZi+cVKgQEBJiN35dChX0SSHnUg
wBVpeSjJv3ptwi0qCwpZuVdhjNIWiiDkogbzU+IhgXN92MzpqgAWaJw3Ec2q4PED/dfjr+k1V79N
CFaSJ8rXusJPWe8SiJMy4sy9xHuFuZ1L/wEyxPuORNHAzbLo5UqDxK63oFITToa6AXDctvZAO7Ma
LSyzDAFy7wgerDl+DfGDJEmrAQBaBqkT/hIEktcIjLt9BZqmjH64F+nugfeXm630rbVS0hyO1+NM
ZzcfsKRDlIreU6/EdAl4xer3H13jnldlc4kH81Yf1iKPkOson1QptMcWVw3o6PAoWOIETEbRqq0+
d5pYwNP5yHitp3Y2j5/N344pxmV0pajsg4xCvzjoIKpvNjdQuDxOHggHL/P6adLHyWDmR42MgT90
jCdlk0yMnyrD51qaPpydH3Jo5oYPJbQ0eDM7LmNkvYKApARt010L2An/xdW+CQrNOAdKZ9TlfiHd
3xeaNvo79wYqKrr/eY8eBpDuDXM3JVCOHQMqiIxgRfuIWa+du/Df22YZCRNwaX0TaE8WkpPJXTq5
pEAN9Sj4kvh+Hf+kabCmoBJyCL8FTgWwN8cRBp0+tjZlL7FADZiaPBbW758VuXa0sh12oqbDepW0
9flcXG5YFoXZR+nsNpRaDmj1z95yVWW/kUqu/PdkV8OFTcXFLTQ4B5IBSYkfB/B90+298uvRJHb/
Kn0Pwe9IkA7rKZSVh6BpfAZM5eC+D/wGI3xuATXfpQbc7teIbZ/ezDZ7mB2oR/dWilOOSt3GSSq4
6WMqfFbV/IYSp2W8snjIZGjA4JCze4BK6wHO8O50hl6TKntxn587BemYcFS17u/rrgggpSu8BpLL
EVrA4uPWlM2NAy9oS/lE2iBeSL9/8O/fhbRWUlbA0uqpmpBd5JBRAZ8BqpfXi9S4e74PmwlKhi61
hEgTgiQzywUAd1LyG53awBTrzWzS0PljUCUavWBqFC3GBtzpAt/6rEtOG5PPp1GBEyobU7Wf+6rr
U/HQ9QEb7lnrnsJKvAj8H4JZ5JwCjIEKVkPHmMC9TFGEd0Gat60zu1z+euJfyr2Kc8QkSP4EaCPH
SMRR5oWpWBHsrpVP4Mzt3Duc6Wk58jgi6KRpakuicIxhTRUa73+/j+mSFxS9fxM99oyqseQSnh+f
HP2PA7qyoxZE/VXzVaK4MGtNTlohDQg77bgUiAL44SxMi2LGQSWC4ldmje5qMavjpLueF8TyT5YO
pVTowowFgO8kqbj6qlzGcXCbCb1CHGMnKhavgazPAXOS/TrWodOQyAACpRYiQZaT2wgt+LIRirn/
KdDkty3iy0HG8/Fcpu1/jv5OYhr5GOcG/SZI3Z+LI5+S6U9qvJmwjfcEK0FUAE42RORt7Q0q7G2b
zuOWB4Ix8H+mRPfmpejSuB83pq9UcwSHqbn7DlzUFGk0JrApWTY5E2/nQmJvtZE41SrJB/Di79t4
k4ZIfmyhm2ZzxoqY3jLPt0RR8EQA1cIWTBsN2ohEuWaA4lNs2TJkhsgXdKj36XyMIJCxNWxMKDeC
KlvBlpFMYQjraFAPeTm1X/G7bZfhlmg6gdbWqZ4EQ6x/6LsRuuYLx888VFHwAZ0nO5KqLcWT7/JD
xxI7+I7hWkhH3pt/TrlN9s6Op9N49ozXEk5YjCekBKOR83WlGJb48g1FkKgXiIJoTlIf41WiFcza
+asX9oOiucp5vfTTJB/ApO/pHa6AIjkAN+V3epVD29ae3up4I90T213cGmT1Isapq7vH3r8DAfXN
fknO77yXvPfCv29Z/YbUOlDwTSX4m3/bI42Au7ocn9/zcq+sstM3+uE69n/XqAOlRkS/zXV8Fikn
92rM4k7Uy0fdwDybqGhugyyL2N1w9ywo8EtyYQuyHiCoMedUm+uSJn20BODFHBD3T72zP1EOxD7l
DtcxDmF/WeoU22m2pri2VB54V+ExCxK5q9Yd6uzbQAeJsH7OyKFJUYJDkkh9rDNx+daIxa4VXAWv
ceMQMtCb1lL4yNAAN2ArPgTDWhB0iNTGbk8i8bH1aLDLyucx4O6oT7fVlpGB1SKFQSt0yN90uAMZ
n9IvbHg7Tpr8HKvCHZgizHD97KsUH1HEMvRPV6DBYW69BBMR1YqKF6Arf7aUtymdQT2UwCQ9perd
08Xyz4OY7ifYEEUoU12PPABjxPPnZ6xHxTzuSdLQtVTXDLA/edtu7o0BhL+U97f5LYuGYBzdVwi/
ZgsOJc7rFPtroLnKRDqNCHdbxBjIdix+pm3phHtBtkgYTXbJ7Px3qID+coy0GbneD7Tq6b+BTOqM
Ms0KUVfgJ3q+dRsrHjyM6OOxgVibhqD2VNIxgzK/Xl3vk+S24uHzR3Df+VgD+tCDALBLMn6yhdkD
iCmoIa07nWHeFjyWiDD3lxiVd4v9z9BxLBaTtrpnvijopfmCFBSny4jCkUNmHvkDa7c1jfub2JTZ
BWad4Jte6cnbDvhs1zjmqU+Ck3TILSuBLiC928FPr2OlF0zqNdoLIDoV4Y6FgpF91HvKMTWE6Kyc
HQC7unWdHVGJz/p2DabxRgW9IrFqB6IjiEBtrd5wHHO0Sms3o1aEKCg23Y188al27k320/2vt34+
K2ZNt3MO5AIuw/UDIvskQXC/jcuDpgm28lvm6XniSrq25QlUQeFqhQA7JrI5/hzQ5u7XEQeAxO4A
Hi6yau0Mqx99sRFMThun+1jJSCqtOVSsBmRqSsGuRjhic/yZ1wjyX4yZYqnHbkooudxsEF+11ls/
hRsvMgNExEVp8GSq2WVjgv0Jmx9PlT2s3IIF1HzHNt092HtYSnx53FGt1KB5ls8L80XKJxkxcCg+
Aqf1xOZe3P5cn5xRB+oI7b0mrUOYoNYY4fwdY0Xm1Vvvul6E7Z0S/Sr7oLyXoSR1Z42KlEZpmc5N
mPb+CSm9KneMK8nuuWw1HUTT6Zvq3VYbRaMfT8skzuqMGWoBlL3Z8ZxdWMhaHVi25maeZ1C3+ont
EBCpTn8wl3Z0SXNBmW/SmUI2SkAhbheOkKNXuIwE+A2LNc2kLvH91VSOhx7DC11MkoDd+c9ImuNW
IytvAPFbKXr72nceAM91TJbsBSOVLkpYHdHW6TWsZTQwW43pDkvqMd6MDV1f8NuzEDrmmPB5LKJ1
AcCH/b6n5REfHQHIDy0UKpfWb1SarYaxgXI2tjAOSvII4Ou03NuGLgomWRyk2KdMwmj2MiHnt9Af
Zwj854OmyNOj4050ck6zfqjDTgwPerGdqWyKkuOVh9FSIydYUmXtcDNqwJ7qwjLNQN4MVgFdgjwH
lNYmtzAm9wyoAoDm5+vJd3aX54lYH81E439Q5xVwZJf0Jwtz94JHHhWFnptmwFAHA2/2yy2fHrmF
x4SFSFVKqG4ZERz7FwPGsXGoaqmcWtGjZaldRn4z0V639K5N/NgrSdH3icver0dU1XebH8nRTKAt
4MKT6YKg5pkr+3Geu90asoW+bjWDjUGjbL++8pqOutX8Xrwhn+1qettrzXMEdV9NhYQfBQKKIH89
gmJiVy+laOjraxJeVwWUSzs7har9PbLPAxI+YMv64f1kcFri1+TZwGyPbwKhy8vGbAhpN3v2Fdgh
vXYBOVh+eVWg8ay/Wm5kZ9F4BUShxnZxypAh7McjZz3TjoN3GI9XbX7vWs0ReTObF+S54Hkww28n
0kRMA+5wfoTbBrx89a617teILU4XMFMRTAUkHDyG6EP9Y+kmL98i+33jcPZNjYGo4JAitlEwZy+R
qcZ+/DXowj54YRh3jgSEUXrL5LZx1R6xzQihFMYcgM2nvXYavBUlb/18c0PFMOJzlve0JmwQ4RCL
QJhvFkUruzOMm7VaiqAoUQGw+tNpqyy4gz5xOD/uZYla47/EnXj+cadwYglpcWobmRY1LI+nO5FH
R0D7S4sZ7wdGsXzCBdgCK8Q8UOwunu3skRnAmC+SqDD9+xbPsK4OVz+AYnu4E3kb16bk57upyPYx
jUj1X4xpjhmIfVOXSgeie6T6aHNYdeJqUFe3iozIz7mjNcZEUw96s+G28jGWE9rOL5GW4XpdiGc2
Z7oVpMX2hBN7oC3uLTDNkfE7f++lqqH5lI9NQfrg37OOvyIRQ5ynzesmh4FAlBflf2EtMOkeEHlu
LoL0EFJ6HgkNfcFjiajvb2yM6V09HvQiXTwtSgv6qYvR2Yy23pD3BmubM4BJPUu8dTYjkQqJzKeA
RFQkrJDYGaf6p9xcGJ/FjbVykjTHsKBZVK7wr56F/M7UmD+x5AuwZ0r2QMlwEeaSxWbfQLgzzlOe
3PY8uvrcPH1+MYl2m/3oAQ6IgNgnLmi/TYW2cKGNBFbnnmyvf+N6KbwSxLCe7QGMvMqvFijwn4dh
PxndzI0Mhhq2/Py+rbfWjt+IcLEehIAGg1ml1wkcNB8M/irn3ufUeiZ6sBGy6dh6theJW5ax5wOF
o0EJBgj0rt/XbKXlNSXWYXTScZiPZZh7ue5q3CQg7lGCXl6Wa8eyRK9nXw2HWzh2svLExoNjGlZr
IohwXM8KyVBVkfgebg4FhDir3EN0xzkeVZwq8H5LSUvFIYgXONHMyccS/92Kex8sQeW7EOe26R+u
5VWBL88RB14iJ6XuALanbV2w44Q3zojCVTlOkARMfUce7M0BDGBWm8NXGJ16C3UleCGB/0EdRLuE
XlM46o8zckuBNAHrk0XvcrcTiBeOcK2/0ymEoFFtH42OFC0Xq7XTr3FtwOEyzaE+goHkrlzSJcWY
t8GnrX9T5u5lPSMXxZGnlmRFMZHuYE/Egbx3xNC14NgCwV46FeZdvrgMUXJ6WR4PDiu50uw0qX3U
RIBiGY4V9Xm0agQPJLiAKYsxuctM/+viX2+AfvZCcP5ZI4qUsH8c1XZHlS0NzHKg9nADxD5ymTh4
q3e3k4DqZJYGwm3m/8zzUnfLQw65Bh9JCtN48QnXJY7iy8LGy4R+LcmnG44Lo7xbi+sUHU+j5Zhc
2gTuzypdyrBuhrWQC+vKvxo5l3Z+toO9QshRB2z0eZw6lZf84TS0WGajbUQfRnXIUzXRffArfFTQ
PVT2tvWDU6CWC3bFYSOZ5AZ+mjnNf4TVwiaOFAvpQJjq4gEnaedc5ATyyPjFfV+W7dEAeft4G0hZ
Lf2uGGyWmb88R2xFUZ2TJYX9upankdE21Dq+aDnjOcxMiQ7RSSKPB1sgRkP48kMfYsxrj35Rt3Jr
VaF4v03P2Cvbx/FYJt4jld7I5zrCEH5Ky1d81P9e77EpT0bo9hVtsuPS/Bg/htvyosytYwGYzhzk
GK9CfvXfVylA9Z6Z6YmUxSDEi2YN2FWAKOht33Letf6oSOJlKKIaS2kOxC/1ohmsYIuzxU+Lw83h
FCY1pIvJ7tNccD5LZ5xbPah+nAaDsUx+PS/MCSZXHOC3q85q/YV79g6OE3WadGeUYEIPrKXXf1J4
tMEoDS7Hb40dsyYJ7XGkA4J2hzhsJllbU2ITv8/8mM9JyCw3TrXNt/5CMnRRpxmvzaEOkAQI19yl
o/MXzcs9n7GipaWks5nSHF8QPTOdlnZS1LShLYVkgxzF6sSc36HMurBrZXc7VWtBAiDbxI2Z1z1+
/aiX0WglP7Bz6s1kjfGv/i7Eid7keeDaGqXokN5EAEBb6EWmq9e7rQG8uGmRJqrOA/AJkPptyYAH
bv7UL0gdfc5MLY6ttlOVvtfW0nQ4zr4SAnrJ8G2kJvog9jDzq9UjHtrXv6qvhA31kdeaD1ujfNZA
mJ2R+IHneTlTcO0kEYpt3oM6nnC9cLs7dzb+guBANAMffKfGwwvuEVgDsXTwlLRKHeyM2ITKtFzp
w4J9AEQczDsDM8Tw+maAr12AaWrOCLtc1lFh+8HlL2kDEJHvGhgyV9Jk0VrzbPcY17SNzu6KkarL
3Cty2COr5gUBJ8xtKypxaI0TnH2GU+aTjqO71b47L/SkHu419m2yEfDIRpXISbo2AFEKvgU0WPwa
iQyLSvm4EpIBAmHPeahjzH1EvF/wFw02Oc/hqOfeWaXGfeNO6+Yobv9AuNq7aXAhyAtw6bE+OIry
pbzi0ntuf/KXUedLpxOvREnW4Hjqw6srTtJoOT/PvZvdDjQJIXzlbtgekIr1Z9IqLeUhMwcXdy2a
JswgAo3vul7mDNoJQe5yg47UojaOOVBcj8TaetWj7fLlptqz7e6ZGfYlhci6n2I1LxWxSj81xUq4
L7k9WX+0qvK6mfNfhEFYrHsGKiovqS2mFAxky13v270eHlqnrrHvBccOPHPwHiFbSvHoaf8we8Qg
Cpak8Q6wKysqcQjV+ptFtUSZhYOpN/J2DU+Wp8yli+43lTryuMBl1HLTEgV7v0Uco2Kd8Ma754p7
ezMOOd32oSpJ3QJdHZMCRLRrzFLjOOIlZ+uRDjX4ZWWqIfG7ubjtjT2wpsAAKj9Hft9guF88QLRS
Z1SGAK1iPBHIPAiidV9QV1/Pww7IDl57eh8f7f5Kb0Foa/30nkKUtrDEXBZ4VudDbTmXC2w0lqi2
QAGSWd7i8FN9dr23WcPeVfahWMPmaa0e6fLrrAH/CTtCvoOoP1HwqPVBqhirGACFF8ZyduGNJaw1
XLkRo6VEFELsoueJxLa2sftyvtDYdgHauZMIQcYMMqL1aYgWoDtzUPuRf59YoptMdx2pbIeepNOp
Zx1iAuqlMqvZsl2sBcIVQza9GLhevcuroodHWK9ZJk7W0vzNf056lYbZSUFeM618nTQNPkbuZz/s
0NqUTCMvnUfu/OEubagbDrfbII8rDXcLPx/V9lt8XyC3lEoqrB5bMjG8RThzXISHQqOS0ZTseiIj
33WTP14BFRpvqe2owIpjEkviBmrw+KzMFIVfP8YWTK/Jw/mimeKSG7AcTMnnb9ZEjRLsS94yGD15
C1ROWeU3SYHyTGR52ooTQMIQamGrVUXBFkVCIHITed2PzfohkM13QCQfW6IUmqRhhf2bzsCAqRZE
tbX0cuBQpjs3SPMxr5OopJQ4O7u83t4WB/g/5tmpJgXdwcrx4M1/vMxw3w1QdT0aK7JC2FHPXvq/
XKOmNC0xb4Z1Dwln7Bou+BzoIETGwv6Q9vwvEn0Mti1Oxarkui8OotxuS2/G3Vhkb7pFxgPK05DR
3MZT8KnB4HAb0m3Ut8N14lUR8aW6f3+2G1v6IqB4GW0WtYYPqMDWRsz1ufkr5UFxbPR9tUWBq9cv
eEYPJM4EqzEFfPnYFH0IToTcU9KE4Yrv1h64SF7XCJ8tdGEcvRcdrH6zOudYpCerOI8rw7sPC1mf
pAggXLsDOiOwPAdh6UG26uradW3v+S0kAaSB5WpMVqC69kdXCBcTwtsrwzAJWvA3V6Ra+6rodRV0
pz9uPjAolkNOFTLMVleBlbei+q+MMCphNmwavDXH3y+gAqcK7ka4OsppbHCKzZAAiFU9rkLfVbyl
yMtcqhP46ruev0HI1F9AKykWA85hQ+RvfhjjUBXrdc0TLqMWtjaY/FOJhM3ujx4vI8EDh/+NWE5B
bMADDWIEam2Zy+yRPl9VGYWfnKVHOYRl44SFhvqiVYGXSQTd2Xrxu7QKVvkm8gItfXSIPusse3EK
G/4pnUgflow4LjzuNsjEQG6rS9c5kSRw+HoFynpM5MbbfEDIWwuLMmtkWgd1lrp017boKwxjeVa8
eWfmpu9cMS2OznlSMse/J3D8bc1WXTV71FNgVkWqy6QXknbKHvZ6CW/3qpT4vZxdqgPZZJvBpPeC
kLPhKqasEPhzr7yM4l7cS3CPI1IXwJkCBYXwT0dgB9VtLChEX9dSD078h5oZb+uaJKH3kb8dripL
YEoMPVO9i3tGZPtqEIVof4RGoKYTioN7U7k01XBuozobqIgb9+qMHNSMwbQHzxZuBjgu7TnRIs5M
KaSaaJyQIMSH5N5I3ytxG/bxfNVfalZSNv+HtnR72VsYBDjMMkQJ5hzqA/6PS/JULCupsxs9L6dR
tjRjfUwB13ESFRrcteBPKWMmGLl+7yAFt0pWnGwQfZjscPFmQ7yg0475lmqJApx8qa9l0/y9QUPW
yOjicdIRYKfT0d+LqXxQebuODQll6IdxEalqiOnRyUazM+3gDT6/nFEsVepwioh6oK+QJ9NdqqUw
crqeyDEpdXMy3NWLOD+vEoh9L7Q8/2DLzFjnRmp45K7kF6Xxgut4+FfbLIpDpV0McXXADOQkOHkg
vSb8Mzt3Y2J1dZGZ76Cg9tf5oBlak49ede80IzJZk7sJY5j//qkWoFeVfLLeIwW/UdcO/oY7oj8X
IMIOT6wUxzpo9s8AcLJ4WDYsWAEObAxL85+gzTC7vddEdkF/8R7geOoxo+zNlvPnv5K1GOYVXLnJ
MS3zRSiUgQyVVYXpu2A+EBEU8EpmjYJ5mO5/zpr7bSksICkCVQ8vSmxgu0m0ZxvitLBjTA308kIi
FfsSKh/lJOu5yHZm2lVre1tQbzAzMJmee8UCxc8hJJ+L6IpNlT62xaRj3vBxb9btYIvygSko2NPG
u89DqY52knkLC724zOBUPYwQXa8AAC7q72J/SJz6hTm5vxZAxu1/d7vFo7/aCdoUNR37th+Az167
MNDDZkyef+okXQf3B3YclEihyF+WwmMmoDX+JcH+EtNAsz0A/xsQ6fQnBgPE6seoPzRN6YBlk98T
1Ka/BHDLSO1vQLL6udVE+x1CMmPDvi0LxreXGM2RkO5hGE2/iCRTyVq1O0rzCFSRAuJOs1czFKda
13NrdBM4dAcgBRwzj0GYkgFAXICCfriBUldCNGlKI2Gih/u5DLdUZpoJKYYn2sP4TS+/+1zFTdjV
Z99ga8JiNZTdfsMq/wnwyeM3krvqrfOeAtNNve53zyLxHDSoZHvgY10+nCDrWL69tgYtvEJEL4dY
3aHuUKc/maKLHSUfmFp40O9lx1zYBTSK4rhX68BYApo7HF9LecE3YZemXcUsrvKexw7FlwbpVPSq
76M/kSmYfCW9Q+JWrIo8OFSD4V/qfZS9Ejdj+EvYTnNdBuo/5wbvxhMp0AMFvF9RYYcbLLpQi78/
jjJEAO/mHqvNA9iT9LTjYe77gNPL/SmKYcyYa4OYg1xJQ+UuYRjXju0LHQBWC0TToft3DJUCo/s0
Ifg4bUASSVTnzBYj7iHFsRCEGKxujgvxiSG1qRAtGIxJaQq79DvI+59o3I7sf1+6jg1AxEv0Rigv
4xFhZdr8L+Z+Q07dyZmp0erJzKmyv+wupVAaCCDVfc5npbwwe3xS9o51kywC2mnuB1cEm7R/Z0rM
Nrt1tVJvOfTCc17R0TbveQfIFJ37MyWnIrMzm93eVtW9qWfHPWaTy5JDS8FGej2ZntSGH7iTKMb3
zu86/Mq9uv7iCnTLwLEoyuQd1es4ibE/6uFN0GtdIjtPmme938oIxhRXfWFyCizfzwY7KDdpPM6i
J5ZqBbxcK08wpT44kIeZ6v1p54qRjTzMF+MxRbvLLynZZ10NwBk9q8bQ9+Z/icTKcCn4vKKMyYoe
af2h9zCa19iSN1zHQcStG4Up1VJjdDbtkxyHM5tUwdTs/p7Xx019daRWYSWWATq8m82WD9YCGoDD
FDJRk6XeRh3nIvzEk/1vyBfrvNPeax/tflv3rOJM+f5472SiBqMdupL850agt+Siaz31GSnaqTzp
iSbBMvRTqG6cAIde5CVbJGW0Zjq6KAoN0BNZfEmabZfGjNV3bDQtAGdv0T5RSqhZEhpO+RmjAsut
yi/A7UGVZL116tmockI6gcxZRr+eN4mdzp2MIBT/hFl21ovGRU3+uzLjJ4Dg4/i9GhNZnKsxtqF1
OwnV2iAho3U1yU2rN44bgDKEtcBuzrH3AiGTKbi4RiyoKdK2jHWV9QRY4sa5NbsRzxyPYnToGIPr
CnVtU6ErpKCL1hEYc037jNzMbL/zkPsjLFrBTLYJvPSRJXqsQTzQCiy9EmgygiEsUP1oQnzxUUH9
blGYFpxrY+KWuhM5xTRpl9n9CTUdmTfFlKxXuYtKQkv3Xj72qDxGUJYb/RPalGjVbKA1a+Ze+ONO
CEVEO5UkAwbAQrUdnCXJ2Z0+ZIGKBGH9xdzdEGn+W9V/mp3BDLIoj+fAlt239t+DvNQqrhDsrkV7
tSjQRyBCHXGXTIsFshrnRUtavKrp7DPp17w4kadjm/gZP+J4I8s3V4ZrYNiJLNw+SjQ6cshKvA1p
ACTJ+aQ01t7WBKKJv+uSCX0qHFtGbijVAzILNKp/QatjMgERCAYjcI1+xe16C0lqHQS3z1vF75w7
/amHls2FGUIizcv+cxgfc1ZHoo7/KAbSPWkiy7jT2JtiLowzCvpzcytc3RL8isb9jwF0LVh1Mmrq
dtu++p5nn/ePkDQcDrZADSd34XovCYOxGSoZSRZNHErMVPasneevu8ytcgxu0ZcKwM5bGdo1/W1g
b0myVRCA6fSE/e0GIUfLG46kKf7v+OToHHkw/MCkXMyzaQji0czeQzNtmgz++8C9EP5wFKMGcY9C
VogI25IoxQhT/L3CHnQjRUp64nyYz94LAx1r3KeE3peEEkcBDKp1CrgxmNoQHObkm0QHcpnhBDu9
dUSUlCPobF+X8uY68fZLYGLAxiYclXngEhSyIn+oAttcy1ekn+3tWBw8Nkc257CZSMaM0LxBA197
y7gLD/rNkbkmGpohm3zxh4us1/eWc9uowvueQh+jcQBOaXVUcHSQA4yjV2tXsLVqK3yQIl4YWRXm
9wEly3K6p6l9XKNJCNkR/N6/EUms8rUBE0Lj0IyElHeZj/NgC68SoH2UKP8IH3YIql+KYEGUF5Cr
jLTpY2bzIb+ydJZ1iCuQUcaVbgior21YCkFGp8D8qK7lXxmKyR+MICmmCod+63PLmdw9DUC1JePc
78ivY2NtChCLraB4HfNui1xyen0RtVx32CY+tlVVbx/xojRyBjZsjb+O2q6J5n5FixjJ12EeFkC5
7CJwUbyKm0RVuha6T+CbBiD+miGKo9mxJDnuly8HzQyOBlNM3JgeOxTP/OySCFlqdmGgMT87nHf8
tIhirFgQXvoYYU5M/hQVjtWe3HYRDyJ1FYw7mg1tO/PNpYBRn/1ppBqCLPsFhPXav5EAOoyBdsL3
nVrXCqnmhwqZJZTnvTLibLNtH1Pm6f6UTYy1HV/rESVahOTh8ZKUYbMEcNwXyO1m0JM+sNjlWdgm
rl/1nJGq+UYwdCg5uoBqBOb38705UfX8cIoi2bJ3x/3RpQBkZdjgbIbTTwUIXJPXj3CmGkGRe0My
xjFYt0BmxI9+ytLDff6t1yEm383BukjbiQNT65EE1fMxZch97Roh76YZ+mkLXYgKJ1BWfGln6z5Q
oLaAL0pDaDAQ1GrKm8yxZvGsyosDperZDEKKjkggVK8sH9oKbPJoh870Fqoof6P/60F99mhQFeKo
42oMrScJuPDM0n1yNjDVL7tyHWGVFEmD85w7QaXNDSer6wSbV+gIrh4jbxAPG4ShyssicbVPg2P2
JepZx7NWeFsBaQLp+AQ7uggnURflvpRaHf3KGkg1ffXK9xve6uuimo2yyAbD9hNTh82a+wY2eCEz
X6ObcL0QzZp4mZFoHaRewLZepiprlPbYjvCtgT5q3y4wcsCHgDV8DHYnOv23JEm1iyhrjuKuLVha
AVyWFnlExmYr8rXo3q8WDYDn4LV5DStGcMTquketNIXegXuadSIx8ZdTSREMYAnkOwU601CXNkLz
t6uxsZkmungBJj81NGCTpjOt2j5Ss8Q4FoJ2PH7UFDairzPp4QLfjGf5m4wpm9laHeKa9Wj6xV/B
313eIlq9w2PCpCdP6Dkzt/gDOZHeaPToBmq1ncpUPvvx2MFl/mvAWiPdBwYzpYU8Jj0kPJSNKXPO
FPumwqAtig3JD/Su8TWZZ7kyAH9+2EuVZcowQpkpLR8APmhf5YqTKExrE8XaRxxuwzHTZtKM9A0m
ZVKcYXDOKSYpR39mA6RHDvIslHMImDh/iDr5HwWXxbYeA/eYLG5lTqm4bXzeiShqCfs2KFtjid2T
BMz1EUvLYhNFMcMZiQ8whdrJ0p5d5gatcIQhhNcNepcIGDK72Yay3qMwRw0D2Jcjood8hBEZ+q9W
ajh4pBXUbhcn8T6dIYsid/AN4Ik/z6ev2ClrGtlp9+LPayCSNa/h+apPZtR2X655oRy0b4fpWB8Q
SVXNcN4VLG3S31xd0nP2rlL5SqrKtJZBREpWqGKnH55s3zOIxpYyHkE+8cXgmgeo7AUFKhTfIvnw
HA5mcRNdwBNa1BbN5uDxaQjYfLDdSpc9VpO9YDvRhmbApoobwjc4cxkPvPYvelwNZY3CNgSsn3OB
FGxC/8YHTcPtlDHNE81F1eVKD+RsSOrLHRokBvnkAKmOHmLOkcpNuWPv2LgVO/hp5dFeviQyHoNt
H0smpivzxTyzndki1SsJEF0s9fyDedGJoUhADHBPXZW2TG0haFIhBg+ZsTWm+jOi0NQJgHw+tlq0
uw0bE5WATCpdBrGKrf0kUnY/XnEZ5OcvFTUE4LoA9uakr2MZ/1Mi+HZugNl+31RQFR1gtGvCuGj0
Shas8Bsqa6cNjePrO7C2OKfLjZU0SouWrPAkXaQteWoys2A/Vks8QC0NTCAILXQDsAi8kApRFJeS
42/lmGn3A7lI0FLyP12Kt9XD1JWxJesVSUyAGX2r4kTIBgW1gL5a///L5KeE9zb0zg+UwV77Vt5H
dOlT7yyvFaN7Y1FXewSZ+rm+zwR0pnqm7NxxTbWv2LoYxnT1izdtr8elzND5a/n/QvdN0NPkuuG6
wREs5S8zzzYZu5LehtIzOFChlNAi84JOJhnlqN2AKL+lxytpadKy0BOXGnh/LPvHB0dXLYdJX6tV
e82n8UBdsQwY2PjLIusmt4Ls2vUlhr2DWDR3+NUp4MOPJUATaxRjVUt5HiBAvDXYCtv/f5acvaoD
jYvBm8TT4rf3TwEAyaY00eUlrjFofQZD0ZRK8/BTxUcuT3xd35+71X4gSyL5eWHRgQdp66jHo59C
xBUpsxbuw+i80z1N18cfk90Rtw+2M+NWSvqxmytPtIcFf9wWYSrnDOK1TnOVjcx8PEZWXRxWtqCZ
FX4jmZN31+9tMxcGG+kAo3ZIYCcX6ih+l5/hGsXcKLOVQkFA1VRz4JscQkujBeKqoUqFIVHFwul2
hWC0kRAMmIUxZDewd/O3rm6XB3++bwdAC6qNgYDSsZ7hnU74idnJSHPRewnZv5kf/0RWN7Jh9HlW
X5Swa2ofDxlH503zKFazOREguIofUqlq+I1ENHDqt9YfYmewAYQcbrTXSCQ6D9phzr6WH7hyJ1oM
EHANhvJKI51pwfGSfijyUIyFaiZXUlYFfsepqK61XFVPIRLCnAGeeW2/EyhMxbMiun4/HSMO3cFG
z4dmclupTwXIZW7mSwUgaa81mrnJMDVi2XErh3sSvcqwN9VgumUAfbFoRjzyaDbp8uDi84mJzl9L
B3bWvUpBGm/S1WfgdURDr4VbdTN46GRUQ2iHVOR6gYbAv6bKALYa87irqXsh6UEQrq5wWa8MTPHy
D9YzLy79/L/oQA4LAbRqABt3R6zqk8hjBAIZGKMMYKbdNgNkps7YgdvXcqXSZkeOynFbmtGF6tkU
txARAaN2mw8oEOZzCFXgviIP6hbldnw5IWpgyZjRRkPQdQbLzra7ZZPl7U39tEwmzd5NvltMJyd6
8/pFX2jK/22Qa4R1bHMLoaUGDkn7tkcSd0qpF8Hq3oX2OwBJL5c82PT5agE3LDEqY6jRVKDtVMCK
XGqmykoDOFJyIQRwz1SzJZ758zdHP5LxSy5ZQI42dTD/Kq90Q+YpF0r3/LiODC2bkk+TB8BxHFdC
ZPZ8wndhJEaNSoy0mRjQEo5gROR3ASiLMXsdiZDrxin0mpAARZqhbR7MRkb3t8z98+JziDpIVrrY
QPeH5DEZq1tMSv7XZybXw4TdRFo+nELaGS03bYX6q7hdgCzjN+NlaKSQEO42VBkxpFiajf8OdChK
PTiZsD46WIUkCRGSZzBeI6dBkYx53Knl8vUZg4CRxmRbVJ0Y/ncGfwD2HVci8Ncy0xM86FAjewV3
enIkddtzpVX1aKkVl1N95yCNYPmHN4evDboRIbp+d+HZEG9nlnewzhhIABIQTpGmlZ9vIkF2SfyI
4gYV4Ok/l+CwaUL4wpIgJaIp8k1n9wsVR5C0aada4TmoJrzLTnw2y8up9VkCfK0QgbDF55SffDeR
yvZTMDGYIlWeQnJf7w1JIuBQ8H4Q9XHBtLi0ztT1RxYUeW+t+xJQKUyptLBzt0EnqDAbU96AFoeC
dhGsMTrE2Ku9+9QPj6D2VQ1FKkwsenwCHYwzjgt1sLV7mpA7r9rTeWJ++WP8I/FsnAY2/GR3BDvd
4VKzB0ASpO59cCBAhnHFsjX3zcEfAjXkewOujzB+r+QCKcJfHPaFxONdCUs6MdRMa/eivKraELZT
asqX/9Gp60k2Y8feyy9TcqtL9nGPTm8m4aZn6fm/Mw5n/AQw/5/Ye1+6ko6MofPcQrX0l1+509ht
C8zct7t7gKS/OKNnSVUrbV75uitdj9n84KvYAZJdP8GOjdrHOvS4QHSKkOmlLASN5Xrt+sNv7nhh
naRXydR5ooWfVh7+Ox3V6hfoOEsgcYSQNw/qvsXarfGpQyU5cUFun0yobhrd8ZVR3M+PKBcHPVGq
gZhnRlB3sQiAQgHY/kMgo31xbcUV0xEGIYy/Qh4nhcheB97exeMHX0QrJtOrzH0+Z3dUMQKF88JZ
nbgRgCUUr4Sg7DW7se7rOdow0plzh930qrZF4N3jzQ8I9h3UnWPXTYlEoSucTijWWA4rnKxvvYgs
+jaUb99RttUgMMkOs8pYRPgm0QbKKy1rdO19Js71Eafe+86nGjnfx81Ka3tHGskwHgnrcPO8zJ3T
4uN9+RX436TAXX/DCO14HCsWO/l4wakqfAZba4lWzfS0sVYMSnc3SKccVdD1+apISpZP8dh96EXr
D7brMTdyIG/rhmKAxnwAkLo0xdUgcUlblQsuxPtNkccCl2qIiOaql+iGXh7c+hXQJkp4122f7Zha
Te5j407GKst2BmIEJKKQQZrFecid6IVtVWJw66cf5TsFrSVGMXhz6A3zbU4OgxIchNIP+8ZEXiB7
uDdDNTg6eUl20VLZVf3qhxAzPTQxjaOR6tdsylMPaZd6BIWBTWWhoB12ly4DrGGLzNXK0tF1/zFv
qCOuns503K1qFzeSSS5E1/wkisdegrIhXecIbAvlFx04/oDWlAgt3iieqJvoGwph/fq725MJMKu9
s9jyfvBxB38ifZnPGyCUWy2wdJnzEsHx5+zlvBxn+8VY5LGLlssMyiAkCvgfVqvW2mMqK6R/+RQP
2uDD8KB4u9k76acGw/DOynLAjPAjeNiQOydeOG+R0PPVwFhOCTru+otzvBrsHsMg+9lzaaNHuKQb
dnkP7yRdWMppTiT86i5a+ZdOfck00qhYdcyIt26ZowHM5FZvVilHepexp9Lf4AKAy1Z9HQDp1r3p
HLWcH9Cj10PwtKd5BI7SSd2j9t7wCB7fZuz4i7nu7VfAPeyytJp2jW/ElTAKNRzyHb/P38dQtaJZ
INKdevKoRDLVNS+RVxMGwSAHQMMdfH7JceE5ENFaxQZ75BS9tE0O4SrirqRDo03tY4f7DHwOLuiU
5VElFKg65KEWxURxMb4SpnUfvWk0Gk2VXreFtuF4rFyW5jLFrNpG2RvHqGgQPyaJy4mkX5vnOTfA
9VA4RPRm2swQlR17RH5XvpHSnJwBeR7BoFIi1HE/jSpADz3Q9LXovnubBF9qW//5e1QW8gbzU/NB
ZjxWa4KgN9HmakKrlsfKN10mLo8CJ2V6hipdkcxrNN0+gC291BvxNlMee8ggOrzhTnm/rrIHuJZ7
+ryEhP7Rw6iY5gzRFGyRPrsLQxZLBNXCIEsDipxPuAaH1fgVQ2sr9sf4Syiy8BYnlUd+WRCUbDrm
V2lO337J1uPmH5RgL1Yc6C6T1jugLF1868nEgSNbZxvMoQ0OsvFEOEbZzrv+9XAbF2blaytsvK7G
wbYW5BIfw/iRjE2bTm9aj1BuPSRp1ZUIhoeXCJz7tDwnyXmYYqusvRZe3Yyz48u1+F97KxaeaCsv
+SK7/Dm0mlN9sxhs5WMLAz8pFjkYr3ICpBSrY+0h9P0FvMG9Q3tp4jgAG7ohMtXkYyc/MYjasz1S
+yhc7Lq4CCEx99y8uQRceagc+GBJXE6w/hSmODrIcHtUyLfV0WDi4LXQ6RersEX13iPg0AltMr6L
i8Yatrd7ktPZW8KouizkQZIe80i493owW2Vafma7GaaE++tCY7DN6halYYJP2QadHtFfbw+Pw+Dg
kw58aEVLEO9hACkTyUsuY3jMfhzKR6S00ghExH1SuYoXDSD4EIHJa2w/B7D01x24GaiL6QnqoyHP
NC0yaiW+56i6wxkQ94ZPFxDo09EvvaKhBGlZK6vYNl8mY5zpbYj/WkavTDm/p4xZ5CugFm0+ytdY
Ba0YYqG/78Mk72iaJ5BCABsoamusemw5eQU76OIgdrSo8UEWKgoj2ssnyWjQtU9Qk5l5cjWpjSxG
O04Y4u6qMEjsXX4FFbj9/OAdlzXMEEO/ItRhCUr/oXxFOCJXDG+PUus6M1P8EBOvMjMM0lH+eFZ3
W4YTdHZuCILuUe2E8tw1VF21gd3DN6PqRFFNIrpGUxsEDQJmcS5CgsOaoh/NTU639N0weubbDLxO
Mve58h8PHsasfc94MAvtlMk5dUSBsNsyvodB37x5iC8S+8dSKTNdmyvqpa4b0qGl2kP2/ec4p/+Z
Ehhu1TCqqH31Wr44HsVnU0IEDEpTkdZbj6keZbuqoSA2OXyuNtV1n0LKChe6EOvK+d8hRn46dVba
f/teTRJZf50cbAtnHcYuz9H1YngMSg9M0+Y0YBd1UL37bHA0+elnVjiqfFLBPc5LwDHtJ092uWGx
qTkbMud/FNqQvLNjL2k9rte28JXh66kXKhbeEgc7PEzYSyBIParZyT+WB+7wM/ONbS2ok3TTuOu8
dA1CBNAlTjGS9Pz6p2ZECMAIL+npQexBjWnyO33MblluP9gPccTYzYD4doQv0+TdnDwcY2Xh9WWA
T3AT5cnYP/QOo1Sy8yUQ88KbgioNszlxa3Ew/2EY0SxbIxTR9fZRv4qyDrLqOKXCeEsybjYNFc/9
wBvCMsNpzAVOTQFJIeR0QN3sneemZ0SQqK2T1NK4ddgref64LN6lDhA53cxgiyFaHQr5oR2/ABZ9
Wl0xcVjXSkhC4746/OePZSO22RdzlbdXSxHmFUXYj4QehiudOzhBW2QsunbHoLFR9jlo7BNdqW25
WAhomYBT/iAPa+Hi76DVfVMMQWZDBgArMy7S4FXkNEM6brB19hBXqFySDIZS3brS8jDCsa7o8sCO
GOORaMjD9xRO2oqvPq+f9LnqyDAGo/MtU03YLVa+krXwp+FCYmfs/gjz8IcQlaR1tk5faX604kh7
iZKZsiO+Ey9DIc3GOAq117SzDYQcS4liqVutPjJQhgwiIh8fYuNN7SSThKtvG/hJNNpdHfbaj4/L
hSF0dcbDHjlwAPr9sUQGxVngrGvI1iAAxIPA/3XKRlNB9ujtuAU5pn7rY/5eotKacptVmIjTlQQZ
bDxGWwHlO93GQ7frA6TZhpsHkpegWTBlwrnVnamVDVbIgXpvVD82gkEFRylY8Ej85BoFFQFLTMr9
5sb7f+bJy9VllYzMJLSk+qz+HdSqxSblTSAvKWaGeom9OrFWcsYQfX5xMO26ArH1LBFjai0iu8jG
VmT0+m21lv3FJVg6M75eUIV1YQvD3kj4DGaROzY/vHljTQnT1ioLTE0R4sGb7DT9kSDd9wioyFUD
u2xZYoRZDw4n0YqGvTo9CM4RC40q1//t4kll+yJcj7xuLsj+9vW0FpvMUpDGC8YpTm9VScxMeb0R
9ccrrZ+j2sVoA8IpFp23NgGUr4Iy8Y7UiQJDjAWlFpaTPq+DZCkEUNstLiHUXB2YVJcBqVgmP5ml
7pSB55hSNzq7UhBoUInryOGz+eJLK+HNKC8G+uo0w3RFME61KH1t1ONJe4K3DUFbrnnRIrzUweHQ
WZ4HAPQUiQuhAZJ2pQzv3jSjxIjfpIY7nbS9T8R7+yl0bLYNhKMa1MmS6CW66MH/QQqx5V0EVETj
ZuCNsWFc35TYC3cvhbStWxPKSGqaoX494k6DdsIStb2BVpeUE7WjMxQFP7JF0sTJpU6TNzZ/FtBG
hzL0OC+pSX5nX/9GZdS4YuW/GG8LP4XpwtRmsRahnmHK6Vh+g6mvcwX9eYAjUgPB2ot0YEOTMTXp
R19X7cSTRAT1Q0Aglz/BteIPjNRaBJ2tnqyq2s5zvubCP7P+ILm8qTvpoyYBwdldXLK79srPXWY0
bAxA/SSwz8WhbDtpz9T+xxPdhop++4PNoSVIs0K8KxFDrqmTaE2nNJvGDYdcVTK/Dieva2udO72U
tP5XU447GboregIleKRA5GYvvb5p4+ZH6XeHQ5xk39YOrBRt4j2l+gwDe6ueB9Rjs8B3Ai4nWAVy
Nvh38g1apz3D2w6rT9N8lA8ctRy3ihpLqW8OUCAYEvGagVEiqJ4+MY5hqGDTyD8A405s3FdXunuk
lkhH0hKGu160UdV/Zt+/TnHHfcXTqKvxcyl+LYM5vVjLtBIKgjzKRy9iEFQxvhScJcpzpJ/mb17H
SntRMo9NmjG9RUGdOrSAkJvoxo9SEvtuTLLSARM6/+Sz1QtMp3nzzhdHeqwDQSriqGHtnGQWJsW7
t/aKd7W9ogHK7MW7k/2zg9PId7y7oekFWYOwKFJ4oibgwLLy4s460kS+j4V2HG1RuMO0LpdNpNYx
oVdEPj5lawyX0qhdZfxZSLGMHwLkN/EKl8vgBnkw9XQHhbKKyNbBgCYBoaxDmqWuJq0KT0g6sPrK
cezEhu3j7crIxJHdxqlTLLJaLVVyz3TcvJ+pTfvd3eA/wjP9ru+UckE//ZTxs6IC9tYyvBqgXXtg
0nZhG4orXtF68GJi215nJEDFtpDUcwqp+o0v+l2yC8LHKCZo6Wadmc4a5QZ09UunV5dNtLbcqowr
nr5m+w6pTU1299MAM+cfHck2Hh85Pq2ufpbf1ld1xjuFtj88pKKrQpVIk/JI6GjmxCJWSBfLswuw
uh6OTLNWDt3aJJAlTzvDJtYGGAHp9T04DOIEkRIuUBg10fyOf0PTcJEEgzB+Shzx2lVjaDfWyjii
PEGqbja0dG8d8J7B5F2t6GuOUZHjbjBU8JqbAmpYxmivkMPR3ixgAhmQkeOZHWnRAwRZZjVz1SYu
mHhwiJ98rrL+NdBh0l6ssalJ+2u5hwsyuoj2J/XE7vsHPLQEEsUvC5+Tu/oG+FHMpOrqSKKP8Oke
p/YmO43ikR6lAddiotpZMyHd+7dum9KNoH1fg/B3FvaUePH290XxrYnz6TZm2SE/YVn1MsXMHgyK
6Tz5IV4yV/+5IBan+VdrDxk38TMUXNn104D8mE4WAVitgp3xvrWZIug6ti16WBdGBqUOW+71dQfn
ijzXXzNAmbYoqU9TXIgd3+VvVQm0WfY2781DCdZG6SX0brn65duwhbz50ITrrVpgzrR4QuQfe/rS
fngn+uXdUDuMfaaSdV1FWYyEwNK6RVs4kqCMTCVPM+N+5WOljWJ8Fq9Nv6yU6WD6u1Jd8hv+av4T
9VrrDvevI9ZJjNmYVO4bixhE4+A3J6CnTHYcOsMSzB5SzmwMQFG7ZB1oZeakUY0KNQX9gmA1Vdzf
gF9JQINWCIKbIDo1nd5UDYnkDxdK4l5KgG6xk2MJImuaaMQlS2C8w7rFwUEULXB84FP8ADUbIVrR
TQ2KSjjhG3R2WbyZ9A4IcxhgxbVFIL3fAqCDhZl/twO7gR4OYx6/zAU2BxQGoHpKfZDCTA9MJa5j
TVfrzBf7UpvYVibIj1Tav6ccJ9/Wf+4taRH1B9UdJ7dZcUdaQ4O/9Hl0N01teJog01w5EXFej674
Ma/UZcDCbUbQ7f6FecUkCuEebg0fIVL47TjtSvxZk2RTz5ALewTcpv/E/98lCXwOO0VaL1A8CHpR
FTsEw3P4KkKo67eFp+vs0QzbYEf76Y/00bZsc4k93/qyuWWYoPqMXNRB/Rk21mrvTWWB4SpB10Wq
TSAknO4JNnNWMuVFWLgz9bIsTl+iVXfH3yEn1Uzv3syLTYZZdQjAir47Irx2+fAruPBu1FC8tjHh
+lKMoWhVG1UDOuqGBHnc6110cDof1YJEa2Uc7frqGwaxCj9JCU3oLCFRsk0tSrZf8nG50XRXZpa4
F9gpQIky2G4EDFHzSV+QbptAFapsDT6a9vpd+00bec4lWb7cpwmEMIbdncXSMpbqBcCxMugU1je7
l/hMEcwICq3Of1AXQoXpn9itAFxDA8GoKhbbvEDMPHkg9vnECUKzdjptNI524mDx4jNI5mSn0svW
q2DGoFtdbpyDHWH2Ncce2rKJbVy8W16OacOv3lZ2nl7NfN301wll57UT2d+oUNEKwLo6iNQFzaQ+
jkolBbr0SKxwZkLAvzyd/e44KoSIIDv7N837KPGiB8zwGkPjZqHC0T7MqKiiUuwk65UoK9J7czYj
dHPQZwsbocjJgFhHU4PLjjYYWK8sftxXmGkqkaOQ+sBvIklICt4aDwd4MicXOE0EeNaECOQKQNT9
ngeOyEbQ6KEJ+xv4f6ywgB2q0MGKLNaA5FWhevd7r4o+g1Hf5tcDq72eE+HeGgIntV+tCphjqac/
00OTX8ou328qNHHNIZVJjjy4YTtjKVi3CWxooy5uAF0muDPbPVKPNyciX+r4/Bn0GcibPoEvOmAM
nyw6iVXB/8etVqRSajUr5yOCf1CT3IDKi0gol6Hmg+rciOeGKRKByHZSjNVcBrKUwF2upUTIoEiL
W1iJTey0miurXUZbDmh3C7+YHYRwwwzJRu7K5/GNZL+s6LF//8/OWyxfgk+jtJ1H0gugEmsTJain
pWKA5jSWNUtDWwXLQbES6nhe4a379xY3f6Yhr5cKOigZeiNdqMdUUnzQEyaVN/B4VdZ4TZXQjFk4
qXLWVV1qKiNMPlNwtzWelV61+Z+5smpT3tinFb//gUgo+7wZph4whsBDl3sN0zaOjeJOmIIjWrYt
H993L5xoBsd29JTVfNI3CLdTblef26SD5XBs+RY2rHW6aau882clzWHPE8233gZcgbueUylL/b6e
KdgEJj2uxdV/88I4C7LWAVwuDaLpIjHoy3cUCX958cnqmCff5ICTqcLPDzzFEFAK3Lg2mhlZnjpM
fa10D4i11pV4UcxP0GBL+hky/dGS9dUHbITzEuExaTBPszbRtBWQ3W3olxWWgDBugId3sK+Sd7g4
gruxjTD1U7pDwubrQBDR3suHsr3z37B2FxDqg/Ds6hRgOXZHaxJWAek3meFDhrGW41tKWUwhQXcD
MBlm7Lj7jsmeQR1q6qOFEvGxckrG5EjLdoZKykU855Cbgwvyl7pF5Cj5lc3zd72/5SbQY9JMWl1+
bNZ6wWq3e/gJC1QZbM0Qr1x2aw2yFf5GLd7RamoS5xHS86f9068WUAyhBAd/hLaK/nlKUvWNrNlh
X4hGOIokjCpEqe2+vVahPw6fCjy5TgXYgiXf6TcgRHUh01mkfIQYAU0Sprt94G9V4277+xka+osV
m4stNKLExirXxVAy8imOMNmkBUwo1ZBWFjzlP/qEC9wV4KWOPd8Q2lGlKqG+YCsA8eCRp/fZzSyQ
KsCJ1uRJXIoZoYgyr/cM37R727uIVarD8YqnCsyFKtFThguxCqlob/lIXD5uQrYG+GLdQMXWT10Q
aS5u5h4trjz4EWQQWRwb+gl608m9gMGUK1PVFhBV230ySlLh352vxSln7WlF7ESbhF7w2ynNnIEy
2nOKj8CYqLUqNJQ3wD8pK1tc4YpmZHskT5WH4V12D99AIEnJ6atvliHIw0M6ZRFVFVBcg87qOzwZ
n/cGE0OnOtajDrXI2qnsecu0UUIF3zbRoiSAqvkAxssyTZdo1CNgODZfdbSqCAB4qeNwYPTSUXNd
dM3mMtjh4YVPO3lIv79dKcd3f2idoogPB7ZoAnKGYvjg/plCUsnrDo+2m1T/UsMo6qBZgXJ+6ZsR
RQeIQ8rJ9p8FWrVcy7Ckbrly4Vi7xfPiHenYp2MIq9kTYAiema9joHdmhHaRYk0uN2igFILH3pa9
xJlHvZvQd5zFybZPd9CnhDp0Yedd6rAqfOpN4fw4oJ+cikfKPPkDeXL6++IgTaF+kIYQg0mCeJ9n
1clTFIi2s51zsIWGqvbDPYKVsJp/kPi38CZNbByeqTbZPTJHTu611U0jqDVezbcWhYrt142BBIY6
Ao4SqcPV3BZkB07gKeaI4ZYvVC5WMuhY7kVCC2CydcR07UanDiIZzNhrTA0+Y/RfDsOrQJLvI0dq
LuNCohCIYpa3ecGZTQE1chafv75KrEugYvLnx1rgjWeaBDNNKYcUTNd1mR9BtGvDWOdz9Hx5x+wk
HghRjU88yVyoH9htPAqrLNTpWv5teoxYZv/Ypos/cOWwMfGtl07PYqPu8O81XhRhFidF3iUCM7nD
C7apkjNErHN3HneffCdUmFnflMM1NlmmHn9AWkrxeuZaU1FXS94MhtBZxs0k9Jdq0E8DwRgaMmwl
b91qpzyEhuoDWb6SpGfDDDA/DSKS95xhYXaQ29eNYo/5fOPZ7cyKF73knEcdVRU8+VncyBd31qZ3
muYB8aOMeKML4DmjajMZUY4oiDMSEVx5OBxG1uTIKcVlRW0/aeaxaaRT5mz0gtCvUgGBSuCPfa6A
QE34dGOR4bgIm6eEvsoCUl3n/PADsSniyjLf1fDDQHAfy8byWKY7bF3bU9C621R6OMvcxuRpjeLx
7kon2YV/QhjlIXiGGqNaDfxJSpCUiBu3pm067oqXGLhwUfNHaSuW0IzExxqh4q3gbt98CzDuHaBd
vc97zs6Gat0XLnY8eJGWDdhdmDcvbNzxy0XjyrvbfIpG9aIrgOea0+2hk2Uiz0Yo9c6+K6zxJKdq
1wFRWOST4goSOeXwpNJKs/2w55sd2VfIPhEuo97tW4CuKtpB7xLlM5yCyHF8RvhrpcMMUOuLwhvA
OwQOGu5QFmTgdLA3rOrr6f2NWYbSd/0qnAVkdi9B2Hxk2nGHsWEbXwA0KuQu1JtISy3a9LlTi+kz
8gW80FrlAnOrMhsb6u6HzOP+x81yCCed0gdB4S7TPDlAUa7Zq3Qk5uqb7ITO13TIWFs/L5fujW+x
kF9iLtVPoEA2l2l7p1ln7K5/ebT0bx80u8nlOXECYM7svbVWFcazcpTBq+RI2ZvW68OvwjIu4yZi
XibBhJ6C99eB8Wef/nSmuG6DxSDQDEfzPW4MnIrx2usUP1Sdg+oyzoV1szIuZyaKUFHqBqQV/l2A
rglQ6q5yiefTKnQ9kHfl9gXv7fryRLRHQWjPnE/OQwQa8hsWLQXimCF79rzdjNVuj29pHQGpnhRb
suyGAl3u2CTDQDoPLP0/wyakx7cfOHBY2BwoZUMm4EMlL8UiCn9Fjzt7o8ErFPgK3p1VhAW0LRit
QxtPu/Ysl+D3eq84QeWthuM87/kzQo+LwxGbVUGasP/7cPnNoBvgCLevUNRVgjK2Jrxs1fCscvte
1Qqwzq410UBkhjVJiZSU/SA2+8XEWk5yvfkCVBKSEAWK31qY7JGSgFwxfEqWtHRtWornTtzqtpk6
Hj7/8G+ioX4T1pH7LDzUq78jEcU7DiSWXxIwo8AhqJuy1g9Kb3nyvtPyFnYRra898iiemeb0Il4O
hZ3cHW1UnElitcLaQpywAC67Das9j7sADiqlw9Q8JaN/LdYVq7+MMo6VUIdwB/4Tw2oOlO+/pfeq
o12uJqfOGj6/mR1zlqlwJTVLZjzBA8+Q+F31Pcqf14K4TLO+prEZjbgHZ0n8dxDsVLY324gRPkFJ
sGPL4P8g+NBuAYlcxXsbBZoxysfgc23R/J7Njvme5MPIzz0k42hY7nPpm42eGBf5K2mOPMv610cc
QWljVY/7VTmcCR2vubXwJoCf6fw5dasUrMvT3QkOZ8cm5wl49CiCtkcgds/dvup79h3QTpJFtx+d
HTXQnsXJ2Aczss+HaLBDSNxk04Q2lMA+ZVULasUZX05os0o/FU5X71bhnBhz7CEk4x/E6XNE4pqe
TJF8xma7oiC4wCaDKJsST4ITW61/w92oD3xMmqQPpxZQrNKx/K5GI8rXA/OVr+tzlZ1TkhFwb0WY
xVSzTG/5b9jznH+OcN887ioeDbixjGYNyneCt4q5qSq+1M2OqvahfRQTUAp+szN9YJ1RBPWtF3cs
90jgC/8t1ypsoUd8rWqSIBSYLtpleeLFwc8KgVftX9rEUqlBH0k5RXn2CB42Ng9ep6fwpo9e0x5B
uauDw3DUID5402nM1VC1+QWMNmHbvEftEqIMQm8tIIeGCUIgutkbM7Nm94KFoa1TWVzkY+9+pc4j
xergylFfAJJViGTjf7I/iJ10QVTCynfMPpUVvKLZmkNsOGEdRrh9Ikn8NurPfmncTcT5LpARyqUt
9WsF0NRGI29hCQS6z0NDDmYMYhm4j7ehnOYj7xcy9sFqa+2B8bQeErylaL6pWHbPDU3aBf4V4MEl
OUROZJy+nZgKUU61AB/a7anwQdaYjfnY0bvG1p0D3Ah0CrIA20ggf/m2NYj2T/mSaTEA12c8r0M8
xhGUpm8PcIcNx40Lh3qngRwH3U6i+40gUcPiizLF64XDIMZoKsAz+oThRkbrT1IIsEeDhw26Ftcy
PhVbF/8V7yCJ3ciqylCZciS6Cwy8e3TezgORERGEb0Zt+cES0ps6+aXE8IHjJK/cOaWipl7AuZfN
V8pbmER914/JZRo9pK5b7QCvfSK8GpB8DJ8qnOWNy2tyg8HTj0mIFgTdJlPoMKMmzkvb781eEl5B
WQI1KuNB+LyfOFgcoikvSipssJiEM0uw7yYfFGUHDOMJ5STVHKdnB2F9OkoBioSzfJp57ybh9YZf
KaegmePUYRs45gm2lKjuV/teHvXNzYduCVTP2g41UOBG+AIk0ZMC24CNyEndDj6IsVR5aZ3VfP1N
0/302oJnrc1+KdNbCVqTyvZ4IKQ2cCJ4Ow7tQxT0OM3EG7mC+pjXVrgl9VJuivfK/q3mXRdKjfAx
0R/i45rpgBOn7LIbWg29xacGLBIkxMcFsU6Et5pXxAXFE3yXVe/ZAwvANX0B9+6m4sVemixMhnxV
0c8UMn7/TWQ+upMqyzmtI+JslyOIMnmPNs/dSe8jGnGRUVAC10dfnb5vJ7IlfSxf4eO0fO5IysIS
Xnn9RNjpOWxfEZAndLkGJjMG19jM4X/1i9vxgQmMvA7ZtwetMKTVqxEB/SwRNsPxnnac77QBb/xe
lAdORgEqkQqww3I23ATN6e7KttwFqfZtnh+GyvIr6+8KKk1kiCT9O70YHCfg+erXmE+tBil1CE7N
3tkjoIxuUqtOAcSlZlopYyl7v1er6Y4do7eZZrDrYGo+TdwqTdNodM7iuzsRVwWjJCWMQsa6NYQ5
P9TR/ZqA4sfcPaWEeNsJfDtwJPuPcfgfnTtn5q2Rvir/8cLFU6znLS+yElWQfJYEA5MdZ6lZ4SiU
Eq3U13xj3HNRYklgPPea+xBSDaxC7atFQOMc6Z7K7pN46FpQnzmozscalG0Sm1lahn3loMNJwaUX
8bNzb5VetEHLE9ZfI742trHjiS+ZX08CCVrmiJVb6MOvpkJfH+Yw0lHwLOGcGUwBR/kIElt4D0EN
49LZjDwLMLVTUsoE5ZTp7F4sYLDvQ88GTMpId5OnPZXi3WN0QdmRiUFoiVesiQkk/JPXFO0JLqTW
O/r9S7+/LNci3rXYZ2MT8ik9ehJwCrbYOUXPyRF0wJmFg/x6FyM48lDb3eKYB40A9H9W8kYxcCRR
SwAmVP++giL1aV7+ulAGxGT43/x3bATm0ZsR40AQaS1hez9alvc8ojKTRk6pj8SrmUAcVrnje8Lh
+FEjEmJhMfmicq+aUiZcmc8LQ0jzjTk3wwxr4epqyLXCZ5MRmi+WaQ1nv2s80cSqOvA0LYCf1Q16
DuUwuXnf9fGOU/bmWtiR42N6vxRf4kvMnM/nu+1SeS+HpsLgivF4+w3+iL2M575UJ0ctafZ6PPG1
VshHyfi51I3DudibAroY9mK93szjcEvemS8mXF1WUrDk/s6a4bNL4ZWNf9eCqxKYZnJt0WAxEY6S
SXLo6hIj0vZ/iGtyzoazFIyqWrswTl/CQIq1v09n8ic7kBPJ1b1hemk4PGpZsD2EsqHaNtqjXxqD
giBUjDR/C9nuFd3laDQCJ2dTUYZ3FYh0oMPY/T9ru8tpm+wpARn30REd1liqIgU303LA3dG5WW26
O6jdjtkwyUJ6RUyJgp1ml9RdxyulQEUiU+NN3zuxhQF+GjvlqFOB3ITgXEyQCdU18qBc/0nfnnhe
PNFMhO32MJEtMe7fZzg5tgX+HBfKVkQXotbQ/RldL8mZNC8jcuSiFC0CeAsKSdXBMR+A/2b/ydKn
VnMdRMdCOeRzoDGr95xiF0Fd1nGxpqWdOqQ/I20aqcvyCok2RDBxzzaOzhcHDeKp9wPhTNnunOPk
ZyB2wRaMODJ3quQem/xoOUy8bBpcL72cjLlcZAWSy2ol/SYmsn1abMv8i2M3nz2yBYrqTN8cwZho
foVcKnXxcvkzZPXLI7upgbVdjtLJCtDaZYfUXXx0+cv+uDAzg/DK33nGNXbuD+9w4w5qIfOhGxw5
ElkAkoThDsP+JVyQWJt00Xr9Y2Zc0WQO87hl1VkL9IHluFtC8zBa4KfGYGFmIHTQYDA5nzKvolyE
VbSdWzxOzaZ3Fx+dZW0LOjywsguKFDqqy4d2cP2aAVotVpA182JQDBQRraJrf1wd2OQdOBWAqigF
eLPHqVMb8ZTe8iG2U2qb2qyak5J5AgNftMyvpgigpwlzAIVyy6VyoWllTaw6Yxcc9YQ6Ti2jnwnp
6Sd2DNbvXppKa83LW5XX3WdRKJBGHmQTFgDNVNTyVLS6CZ7EqoTIAypvq5g4VfuO0yv6Y+5RhE+s
UFe6PVyt9inGnI10elXMe6xiRoAZvD7FfyygB0xbQlW/Q9fYtQVxjxg8I9JHUTyXnw5ZpF1uLRdk
HNWRJzWjOp501/b57lvqHceflsq4VKHhGpdpI3qMvdF2bjXA1+WTzTG1+1EqEepArrNBkiw0yXaY
0/hRNX6+CF3EtXm8KYSyEVHrAvN//fd/KDWRUqzugw0TAwiE1LzfxeD4BfEPRs08YBnplq6J+G6x
8E+AEE8iB1F+acSRwKRmCH2F0a3tQ0ZoZ7tvxSWDVKE3+CGan1NdxBRkgaB8G/6BW6C0SD218nb2
01ZWm8PkXTHX9gCypyceXW5+UMKpa6T873hx85wHeDVh/zSwV6Y6HJvpm00D1eo+7tfN0qh8++gM
sL2+U7GYQuf2XxWAKreyg308szxPA8i6+QrIO/dsgEsKADQHTT8D78VqI4WoKpE9NG7q38anPrn+
OlyU8fvvLoiep5iBTNUSbwmj7++JGwnfJx0TlA5bG3yYLWl1fRbS7A2+ZEGt+Fo7OEXqpvWnK7s1
8kmU0X9TaHcwh7zA8ACCGt5XMIAZsqQu3kYl++Som+ATB8d7zYUkXXiBNiDBXdMIrs8ztPagGX69
QPmZ32LOHLWQEBAYdtzCkdZpAYxmhwoNFoxHwA3jKuo593K84fZzs+uVNsNmpejZkjN0IbQrjXax
059LvafNLNH8nYRM0MROFB8XvBMmJnVYUfYe93B3oyUDyZnwp+a1ovoRfsjZ4ftW4XFIsfAO54CZ
mqjDZLd5hOCA2tQF1UnW+buVJDTcj3m6HEIGjaivp6LieP+MnfXmTQ5qVefCJX2CDgCydTKt4vxL
SZYgXPm6m1QGtpE1BZdCZ1HSTASDXt0yK4RJNmQNqlqCzdHr66NwWJZKXtwP7y551KlXVz9OzWeO
zH29csJDf2ji9W1mn5ph39RUKXRZAj13whxjSuugp90tI1WX0vt4E7k4WwYsB0EKap/Wo3XMGOTG
y4OLORNISJwS7+0Y6tQrR7pYQgJzFcFUUZkvpGap790Cp9RTNYzudHDigzEuUjBwV1W02nCUJIFM
erYcpRCYSjsnML+2asAIvRfdQcJzbOA+82eeoo+fRMUzte92phYv7C64iVFt/jp/Itjqg1Ho8tT8
auhCD1E7vKkLndPFG9WrDRxNavCMQ1O0opyPC82llMCWupLkSVVtksx4PdHJJTkDSc7T3vNL9KXK
GBIGOwtP7GWtDzay0/SQyq31z3SNG21hvjFc9slWlHU8yJXULKPnb68ybDcjCQsfG40nPAOlaY8i
mARRHfQZ9AkC+W8g88SZBZbq4gxJ4R21ZotSB1z4B84MaNt/TrSusy871ENFAy+/kFWdhYsGHmrk
1W6Tp2Idu9ihlEjrmk06jRkcnrxai3FlEvidJUmFeLB3710ps8uJ+o/7DinaGp4WETBp9AC2HOdX
9b68pbtN1mHFpn9akJzA3U+ySaAOFyMUc0qKJofWwl5Kxuk96O0h1hbkjDSB7OyZBNBa+6jIYh/t
wmgEoHloJ01cPWxj7yw7JjHsX9iZbFgFBPAoucD5eUSLEpRIDLA4vM8zBPlya5/g8l0STm2rs9ql
aWfZ1lnGaTvElU0uww8oUoGbeHm16zbmotQ8kPzelaO5sWyDgSb73pXg6fTeGPIc8PNmJ1EnRkwR
7LeOVDmNgoF+tMFiemZyNwfigb6ep27Fke7jM7y7bdbV/9Mo2KyIxi/d1FbSV3AZw1SU8MERFlvp
tg2/hlHZCAXLTgDqor/MBDPc4JCj+IaZwV7a/+oKI5yJoRO/zIQgXMb+aitcL70k+AdP18Gpjfed
MNO93Z9O0H0LCDyOP1iTFR2ovAdq5htIc+rgaFKl6AFeYp7QE0yWkTtW8uG4y6xci2YS9fvgTGkU
3RN0mgNedR/YIPQjVQhm4BThAEajpIvE2j85wjhNjzKnGl7JFlOfhtarGKnnQ2hN9vr63A8e6Xli
cN1Fs+vgyJk0h5jeH2yMVzZArLz1DWcuiLiRiSrWQ24vmjMQiZ03MxqG/YKwlNsAcC00pSFEBoLD
LRYGmDHNFgS/Ox59el8T8DtZh0hi30kkCH+xH1Vv6XMCtvyncN8IeYfZLmR9DmqAjB+omZlchzeD
JBW5/CHMQ5U1llOB7+IVHl3oUxyjsAzWLwK/W5/XIbXLYbGyObNv4PFF9JtOdGQMb/5ed59V2MMd
nTJkva7SaQlO2j/AhoT5mCCJsn1A9KWaO17t0CXCmEDmSC8pX6MgvLHP4sUFbeRks2zItTSYaqyF
F/5dTk+loIv2G//7WdEp8e/XB6743Tqr22mQWN8UiPun78GMX2gh7I5Mr/C9XdbnAIkcbNAk/o1i
DVFxmNVLj1AnoOHSwwhGAtgRjg3ZhQsywqXKHX+zO+WtcXEH6pfRFSBB1+kNAsM14FzZ/GOj9I6A
NB8DRbTtXWgSRn4519wq3/z+0RQJcwyVtaRiMUgc9vjIsPI2Yf5msbPLoC+rljdXsjvf+cmlMQ8t
Z6ucuxxZT1ky3wimnPoWMwqY1T3eXtO1F2imufqtHGP09ND8mh2gI7NS4luW0lFCycoYlyjOZaak
02N6a1BlV8gJB20UZyUWX377eo82VDnXKFDgsZFvPsuOWcFVPqqfEg6Pbbd/s53I4XBLl8VWhsXv
tPLFl/jDLzuhIIQZrrgU33g5HZW2F+Xbut0dOoON15Du9FaJIHOjT4448SkmVi0Ft4Jh/qSlBjOy
5mEuhwSzBPVqhi4P1h62WBmSjky+W7HPrXQE8DtyaXhidL4aII8EPs8zyAFIpl3Aizu5DQ6YTBVs
AxQd0msG4EMXl+gqsUvzTOzGJwtF+dGfmHYW9JUhpC1TnIO09cO5ZnAIDT3Cx54zIpnLzb4D0j06
QwAiFBsbKHRUp1ulTPzAzJRR8NO2iEGdkYlzlk93yws1aLkUOomCA2HOLfN2CrMC3S0qgV8nI6/8
GHOcT3+sLAkem59QEhpX58KNm2ZR5KhVZqVNgj85g1ZcqdqlUmlP1R9PudR3fkqi8RhUx7/+B9Hz
EXbt7fPLam2KaXVEH675mSvvluNOmGSJ+MBErZZAGsaTZYFLdSU7QCW3WuMmdnXdZJA4hRfi59BF
f20mCJPe8fcgJzg8wfVsX89sZQ08lAjfranTu7YIKwCnRcuLrDP9S2xc6gLlfUswuwc1LLt37NlA
zse9fME3of0YKUEAaaJaWCmJRJsTbKdTGbOdVxPiS0/8+k5LY1X3Z9F7P8MHdw5+1c+0pbUU9wnN
HbDwHGQy5ehy+exfCvzh6XxBBDWnGQdKESHVztyRA3uDH2WquDGhL4SHZqET+HH1BJVdH0GvcHg5
OQDBxp+NYWzvlrfPoEUI29orQQIyM0t3LR4qZYekztZJT0inIIt2EmKoUsE29EuqfKppZclaHNhq
l8gShUrUadM4TiPVSmIp842QQxW6BtxYstHP1pu29U+NqRuc2BeXilYYB/vf7SKg411cJtPN4iJM
OsZF/gBBUbPtRrYQt3dbk5nWhQU+GP0w8q1AkVsTs0P4CEyZyCFnI4WTuaUAZpQFUF6sg7T98KlQ
kybJlJjwD0ZVx8wLLRt/XrhfWSzLs4t1E7UF1AGRLl0VuwE8rrcc19ov+4cq32OLxVGQgmZTwvOG
OIyxrwRk/GlXozFToieyK2YPf0evIkF8MlOcg6Dd8qelibwytd6XewhYjE3LPbTvntc9IKvXxtna
Zy5BVkvnPxO6x1j94wnzjJfEgWNpRqA5HP+MC07ps6aOF3b7c2LScb0pjHKD+ZNH0PfyBhnX0cxR
q1JxJmVk5NAi6cExzFsi419sCFV0QyDxWk19jtF9PjfpZ69fTc3d7X3CUYeo5HT/Fg+sMKNgpMCv
MeokeC7FdTpKjuOYzunUvt7kFq1ebgCRuw7BtUSfFGHO3C9ySTIprOExiTPg4QgJgNcGC0jN9/Rs
QlvBNZcdIAc97tGAGlZa7vF6VZUo/vS8/S4/FxKvurH8uO+qY9KfqXyTrtDqNhAYY3wcpyMpSMo6
TgBl7WO4d0K9Sg+BjFT5K8EwBWku+dtNwFtxs9dOD+ptuOl0ByMxsJ+Hro5nSQObS1j5li9Rg1EB
Qek3EvDvrMNl7dbdSxOmDAIKAkjhuWbsZWCvVJTmVnTTL25NS8M2DXWHBXH9Vi8PCqY1TbUWquBB
Nl0VAcXm26Tomxtu6ZXRqL6v/WuylTozNjDfzLNDTyFNlYFlFfV/FuraxRUJiyU3fyQd2mBRvfh3
+uNzdMgX53+SYX/UK8TYJ2XZpRTi/ZSRZBjAd4OboeErBIzeTWrN1l62c+8MGIL0nfEf5/xMh7Xb
fLv8CqhYzXrDm+RNaODAsvKRLOFtQPH9mbBqJ++aQCFK4gAqI5gZBwYXMl2IHhLMoErYWCrCIAKo
Wx9MXGONBk1YLuxn/wsl64FWxq1vAWX8KA9hf28BlDv+HqdWDgn3m83U3Us7pg5mhcByc47gsZ0n
zyBUaFGySze1spgYvx8N81Mp85dicCO+go3bad5dun7RU264ya8+qNnMSUV9csQ2yLsjxKn2KWZe
iDhP0P9r2UVr83W+HQvUpruUc5F/2A7lHKXhLAjfdeexPu5rZZc0hpSZPiuFgmfKFaGgwsLgC3AE
7GGD7XGntv5eLA2LwlHwJZ2oMUr1mu2b6CmsAfwis2/mcsZxw43FjyQ8yiEkHYoLKrVPNFYVVuQZ
iI1oFOV7rAHocy4umbbvI0UGQ3btzniu28AKcTbByZdGL/b7Lv+gjSDJpvpVlV3ghhawMqnLYKY5
EhX10EheFY4qwN0OIibxiEiJgV407P3BpCAl9uP11MRsbqlXJuRJwN1X4tO+VImyidEXzKJYq0Hy
C2vWk9jjqLpkuCmEaT7Uj9quUhYeI0nLTx/cAXT5UtkDtk3/LH7+z9Ig4gI2g450I51H3wCOrotn
30WbicKYOq3FRD3fLb3jpNcesvJan4FXa9+KVcVVRgBhjYbDwYk6YPmSUxZL4jY9P/GP8biaBEZV
fWgdLPa8ntw6ntVq6lnrtcEKLQwRxMDWpcXIbS8EShIZp8J0q+zc3FcAhPOkYbcVrFVZMQienEHG
XqKoeVo8fL5oYKWVcN7gNO9ogqs6Z8Y7V9sj1BrjRSXeGsGT/IG0WYRTmGIldH3J7mzBCa5wC1Yk
0sc0LFFY3F8+62b2wZiLwmWjEOzKN21QPJMVfzS23CQowLcnpkolxcIDOocsRfy/8cSyvO2Lt3sM
z/1NfJaBQ95GzGC+HxqP5RY9muRvGigg4YYqYED8J3s5dcKvL3u5L5RzdfskcgauvnnnjOUSCeE7
qrM4TsBqAKsiUbHnEgYaKvRbsx8WEe8tHVYfcSfqXRF37q/AcX2hBN7Q0wDhl5qyqN54F6DZ6ukz
bYuerWnrDSE/utaBAI0L42jbDkFy1TzNBftd8MYCbgMc8mrBioYLpi/y93Csg3vT5+HBr4n05Vz3
3sUsFUD9r5s/mGUda1hvG5lXjmf38aEvy16nPkj5YQEVvBtYRO7sPBsiVNDnLjIVdUOVOWph/233
ODC1u9cSvSwCXDhOVKnv/IQlkQv2R3VUFZ0mAY71pEcx3epvKmO3GNUoDQ3nr/AQhaNNu8/pt+CE
gZDiJDcTo9k1fuLeE03sIOOLQrUpaLGA0V/OppHzZESP5dUxSh5RdHFCIDya8N58VZAI2j1rk4Aw
Qln9uAjTYnua7nFK8SXkZhspATP5RqQxYbYuLH8AIyONNhRNE1xWRuMNuKVtKVZUNg6OqK+cbYYY
94X/c0pwi3iFCodeKFnPcwDdmLubKf1rmELZIk5s42foBGw7hWvpf9jbe7hGNsWjukFOCN0DlhQU
Riv2a3VicLb7fPHLjA2mioTIcZOWQ6ToPwJUqjx8RATNv7CIr71JQcPR/j4f4hXFEaA2AJcIl2gl
RjwhLrKO8qZg8fQ3RDH4RSi5BVTZchK+tBa6eUXO6CRfbpUgnfb6jzHlg1se4gCPTdBsE4d0WzWE
iSrmvlZZSodN9rBMftSDghdmMqB+E29a2RLMw4Y+2wS4oVsV/W38Q7s7+yGUDaeye+ssZveFyl68
/gqO7265svQ5fikJshPpHhx9OsXQnf+nSG4Os0n0gEDOrB9hM26KzOtjFHGlATNeaEXuxsAG9MwD
b59zkJH4OS9yF8i6jxDN/98cPN4ZgKUtbvXLGXJC25dfmgWowZNk98SOzRn5zdC+sVbdMlSygJPu
UmUhqbLT4vBjSHYjrgZLJ7PbRTwHWrrQPmlxu/WNpKvp573U+TQ2D0yXSg3ZSzM6x/BY6JEhswUB
oKuHnCBfDFYG9XxEqCksr5xYVOT+0kdN8jmkp66il6EtBDqj/UYGMh/qHluZNf5rRcTBIDKqpkzD
kKNUoWiP1oaOezbUGYTjLam+vNIKIi87dgpyHSSqwKTGuTbNmxdt1ZuTAsJgKGoodxUdDB0gCdME
23uiAk0ODIXhAyHB/rEU1JtdcrRYG8I3FvYr8sq79v751ZvKGLXRYV2g2oCaaoTzzmERjaZ5mRYb
wHdIrELRMGooMpgPGfWQKliPDore3haHBeHyzcM+YTV+wlC/BxPtr4f6UddVmWqM2X5rMcziQ7ey
YNgyNEUwWEVTRoepxEXHj894vaOqRFH2kmhCj8hwjGO461MXDCM+1TjNvK8dLsZ3/xkRBLwSULcs
phvj4/ATRA294jo70lDogMv5jsKoyPBi8EwwoQqfrgIAbfFN4pH314HgjrllOh5tlF2YJW6yPEt2
0g5yCBVJh7QvK36+lIrJp25iB780Hqroc+Kps6PD2fpEYxHLx0Ls46Z3e8R56d22IdAS3MnsnyMB
EfbHAazWiCIP+uf3VOomG/vP5++cu3FKxN7eu4y168T/RxN0/6dyy7cOQEkyzZECO+d64J1PAkwP
43hrsBfe3nNSZBsKpbjH0rXy3+ZYzYVDF3WnAIgG/CeMzEV8as6ET+um9rbahHNXlkE1gBxjXO0f
utMuKG5BJ21uAWMESAQQICzBRYmRHA/3EXoBesKb/tQ7b4dnGKkU6Gi17vR0jtnUCQTethZqgkND
lv2xEeK3R4nnWEXWOUuyvt2FJ/vJmN3r1CMgE8nxOhOulxFM/WkDrpojZrw0+TXwqyupL9ig8rUR
hs1+tj4ZCmBcTmRneM3BOV/AJeaUUZXe5QedPcNXM6mlmjr8qmWkUhz0RErbe7NmVkFp5ATMVOjP
spl1iiskQqSTbcI1pmbnAAYQiV0MpZFZarASHoCCRgDxTdsqc5LxQsw47Ct2QLLzsb9gIe/eKdzz
d+E2OAKk9UmOBMjarCcPMD0d5+U0njEWUmjpcni1VbpDaO9W1q/ByR0hrDfhlITNeG0hxh3PWqHa
Q5fuTi1uEm5tcTgkdHLpThQvnF4x87ZWwVlrh/4sjZQFM90iKq36Cc3fHYGRtU25mB9pGbJu40oq
XTtM6eEX4RWH9eLIGzQgaHxRsMR48sxa2Ltin0+h/xrkTPfPcs8PYvAdxGQchv0vC/xKkzCGaGF9
EZedWOQOOpd3SH8G+PuKY8dg3GnDqBqp70bkRr2lxXkUIhC3EZxoUR6rzvQPc6zz8OnXIRDHMjxL
fsaqUu+3kJvdb0ZWCn8D9LkwNzaXXGslhsPOQiZfrSr/nIKBbASep8u3FGeyV9kBj1Pdiqv00CkH
V2ZGNPyu9Fzjr+YOOIyGch7bZV2w4g1OqNhZhAOTrb1CaRp8f4vwToZuvFQZmdk2vaSahuaAmIgc
ltlp7hv83t3/TE8aloQb8nDhcK3CZTwIqYx5oL5yAxa6WZ2Qni9wZCrcdse9/a1g+52bcYdwtp5F
9cmmv4iEmMboLBhGeOr5rgn248Df0Zk1gr0NAQOm9QBG7/nWUWcXkt9SjpWos6/W5HroAdbWznhy
lOvSEA6BLPWe8JmZ5SCHvwVDVWluCoCPzLEOtsRjnhLJjg0dQEsupAMTG2WYUKNb1NSuaddhRUOR
DCSqPkOBQL+UxhHL3saWIm+FJ2QntS12FLf/TSMVKDPjFzdSxG4BPaCJq1ayQdaUbC+y0310JRvl
taMb65nM7PrRqA9b2OIQjMOkfG7TC4PGd+pAmPdfWxbQxhtg3pPwkymUATioQdC06VCf+373tFZL
T3wpEz49p0edTAV8rpLTHGyFWaSGS0CEgCoqMMzX1FEhZVgjHKcsddQ2SQMq3I1szjuGNXjQmbgw
VkIHmO7orIQ2FR+aWxYkZ4/fsZlpUuAXgr33Lx4KZ9d7gZeGcibbm4ss3qW1OZQRpPT34ypbZvHZ
QeBRw2gtkz6BOMxHRCwI3AUyVwdhyJRkvJ5M/Zdt15hztKurSC70vgarydBK8VfVlkqV8aU6FBaf
l1e+020urYXv+LSWDSjPYbhSW21LXN0MJTWu1Iu48jzN3nk1gOiiu3qKBXM1P8ndeMJgngxY3DWN
U0tEEzIQz7pncrJ9sXh5eI/akk7AGdy9+J7pnO1dMIQcs/oWD8FblbLire8qUKFSYxmFXwlhryk4
jF2K4iTmbVyTieAmFAjzchr6DEMRzpnoVM44IoNnxSOcpWmbF7K1qcbo15qN9BJneikaGRqjMQeh
xCitip1QtazrcegI5MxOVnqQD76EucsYO1w1gGnUNpHhv99JB/WL2W560mB4aifBuXG4ayO7nyjc
/ZEbug2hl2/0i3V3DlMhrV0B1TWyCwQrMJblLUH1+u0+w3uaBkr2oGl37CoDSywL/85nwtOXT+su
RiZkDzV2E/FRkrXqG21aDr48rr9Ywr8YzGujzzQSoN1jf/B373J7ZSk62YGnURGLwo+TtrRRVVC8
jjOaOTriSzbfYZ2+HGJ+bCaTLwEg7ls0UcAkgQC3VjsrolqA0O5dyX5pt19BpeG4lUmnuxxnhfJf
oj3kNK/BuOx43BZj3J0sx7bKrSISz0ULAbcNyeZ7qzliAcQALwChFkXhC5+S4ipmE6YBy5JOFnNO
Bqo7fokEiQjdCUWojV8ivj4D7UbsKOake7W+W995w2HHyafyemhJbO4FfgpepfkJ4Nlw6CAsB2Mv
NJzfqsiOwarYp+b9On++e5ZYSDgFel7Gsv1IOn+eD3YEIgq5+90TpHEd9bIsGXyzavD3uQFovoHJ
CuoOj4+B1Zi3jsppnzWifZNV56boOLFuHaIcr+ygnWdQU30ElhfpNkDYsW4IpVDX1bbaxUxEEy48
MCnkmW3y5YzH3kKBGxXgqmJULm5RhTDtqyxuL1v4UxcSbnmpug9BfHsIHdZs4CHiX5zcjAp6hP6M
F2HSbFdGvgXtGvFjLCWREE26hdPQEWA5UY5a23Vjx1oP72TOKJjer55jgULAbROTQjlHFLytP+BO
MGip6U4hmCAqtSRCjNDcXIoBNElDSAKqUaghhzfGPf7mKhNZDCWfare69ln7UZ/ZD9crZzBbypWo
cQmJdDR9EpHNhGP6ob3DMIFCyh+aT+oTMvM3sFeI0yd6XyCxVlwgKQ8a0wluB3EI5ZknbrqrllJn
7LgYKgcDNwTsvFmiEk4nPLXxOXPk4jXaWM1DgE3dnqs1nnnS3ef+Cgv1WEOkGzpYusoIdBSS7Vzl
gZ2tC6RbqM/5QdM4XOBUFwwRdXYL4sZBNf67FyHYFz0vaZIfWbWy0a8SrtiQkCUGanrDPNTLhwMN
gdw+agphW4hDWb1joTbKsMVGbLJOWo/Kc8JlWYegAFPIdpg17CjUBvWvy/x8oC6O+bvyQVET8d/z
r9mXbMXc856CDl1PB9p5nVR6523OFq6IABuESU15SDm0H3qGq4qePp3Ia28VzIyuJbEtL/3pLjhz
ecEVKgkqOIevE5mciVYA6Da7v7aEBozwjuSelQqmNm5G2TmfVAxagqlyBhK0WSx/nhE1aVPTHbul
zwL+3ZVby83v1dinTxMBF4WjCkvGMj8fyWMW501r0Vxugkkyog4fq+KrsiS7QGfkQhWGcSEFoPAK
SgZ50gakzn9gBoR01iSfWbtfjmKyzxtMwYKtgrsMsD6R4KOOxDw0PDPMBw9vrqHOgULG9o8MzmTA
Xn28rn22k/RQ3nuGJwrh65zXnXGqGi58MrFN8uqlYYmYXqRlYLQvpz6R+6s15M6Sx7Ls8Yv4J9C+
2DvkMb5/ytyQroP+tno6TfNMCOANKLStR7pwsmIItS8zXeQPy1oOzzd3pUeLxvN5SYaLXfObuUYS
VLpb9jjAF8EbqF+vyPS/P3bFXrOXWG2otfwewnxH2cX2PfAaB93XaACm3CONTlcrrZiILEyUh+fD
iVPeDhSd4JzuBod6otVItpC45m1EFW4GTcetKufavA7B5Gx3JkFsf7GHV2/eBPhAKgT1mASoTKXN
YKmQ8xtWgK1ps/kCzEN1g+eJAfJJtMg7S3RFO1V32qIOPK1YZXMi+I0JiC4XmlXcfF7n81JpC7+B
h4MTC/SSp5Y0EyZ7bN4qt/HIjDHmrd82plTuW7yyj3Iff/RMQExfv0AGg6NKJzyEBLoH5np8ILHO
HaM/KJBc+EfFITAo3Q8Mo0UR1TDWHK9YAUNExkw7cSwZw5AwY8qXqsO5PSydFL+jw8Iih6Z9ZxhF
Tc8cJTGv7f38UpApaW0u/VnH6e4NH8RVpcpz8HNmb0ivJBcIgR20ezkTIwdTz6cd86H5EV8cR0rm
SiUGx6I6zjXRJDlIj1WLVdadmZeXminYYW8cwECK9pnyGbuEj5v4u5wGs7T4AkZCW4AhvBJ7hF4P
uu/pfC0vIDahZFVh9RJNUSTnD8YYNiPTPjVM0St3pDPkGtNhwggaUFNm3R38gf6MiXgGYRAF7XuO
daC4msfxcAWWEhl6XXB5Zq84SOhNAJia0WDLpvvXLSoJMm/1osCW+Q9HG6PmF2dS/Sqj40LN3leb
6OCoiKVKwdvL98NvG8t8q1LnmZekdihzvjz+8TosZV7WIOUQKeHLB+xu2LW/AIihd/cnxzNORKJ5
x1RlLLjmMqxI7dUYtjlwPlu5eH2+HjDnVVZz1l6dPspMDfmOLYQ7p0v8nhC/dkkxs7oK57jKum+e
hQaYHHelz6m767hj0oheImOoLxxtXVTUCvrha2TCOVO+TrGnFOsl6HhhYiO4FTemdBJb8DIqSZ9z
yB4mB877gPIKJrna1CTnkGw3bhWm8DFmbbzLhBX07duX0mzMfCo9kEJ+BU2bCGfOAwMc20MpDUhy
3F/7fBhiwbuye9DSWkhxu9evI/devUytDv2SgbJrfPClbXe2qNJurGM0KBdyWIFuh6vi9OZY2ZWE
Rs5tMmeM2u3rU8qeAP4N+3UsG+47OoaoOXsQPGvUT5+RbsGCxcRRScfbAH4hvc4knujPQXd29Qm/
kNT4zmXAOyPrMaIK9Pb/Qjthnq3EiBm2zjsOped8IbMq8VzvtyAf+ZYhwvPKTWfcKSBbc0cN//Lv
fcRaF5gSdlMyy5h49fiGV5n8GdzMgfc/1511pzQ5TzTvtIxuW+L8Heji0aDo/yrHYQ/+jWJNq+Uo
e+gqT3nRaX686uwMc9mLlvOdmD6NmAhs6SKEakpejzyW2JE2CyWh/ax8O2McLGMxvguJ+4Vf5Js7
4Kv7C0YNsShgWVLD9bfMqOFMXIFby6q9qVX9+HomREjPiaQYjmhDqRMK7MgaTW6ytBlsSTcVJWO4
oicT7M1kQXDuSQZHEx0SJ6sFr8a15qkrIjJNgbzABV1XxTCmQ6T2M0gpEohQgjrZTLXGa0b++XQc
6NEt7q0n7SfhChkB/nPZsKMxk0vyftCnXgPYToVsI8VUIvWtBOKCmIvsbZ9jtQx9dYOLlxBh72IS
ldAEFmQh8FHj5wTcwsdDl0cRg6YhSn6erZwB3kw4Nkg2UbdCUhv6mbg2nu24jGDS+CJme0zV9kue
QAp0hxSQGkYunwNcs6VOramxRETtwqBRVpUOP91xco4/YNySTeZ048uY651/NidDCtT5L0GWiCta
mJlTW1Z5AaCLfifJnSAE5aiw1YblYVpwPQqa+dMy09qwkxTDTiyNGLEXUqm+suU43jkQhYDd/ZFr
MaXqjtTE1frlzZNp4qOXexe59EedhTEa9QdclZ5URkhgVNWYX4sDghfQVgZKLqb08IZY5olh1IKt
ZMXu59PwUa/UmZlegrT9u0j9ZzMlWZin9c+3lbgf0YxVTNH8NXnDZO9JWEW+yp+FVPPzFZXeZrsd
k2Zbx9OqDc/1IjPJ/24erq+O6t3AFzzfwguy0JY7FtcSCNi3+hcwvo8lJZOAIFlUnHssfyE3CstR
XBVcZoLG/b/W355bqGaRtvHSZKAk+MK2TxFNgsLqRv53Fv9R49J4exOeQVtQwgQdoaLS1amijNUn
+oFGcgYW60FrSG5+CKxhIXUottWdxClniKXioy/42Qfpu0wXsJMKk1IUbB2mrgrblOy1PIOkhpWL
LXKVc/fbkXIuDq+0oQb8TCAXL8tbTHRmO02ARcOUgax1Vr+bfq5miMWHk/bXzg8a2QsShGSY8U9F
koQDCI6RjcAh8dz4wjRianIwAakbhLUfyKtQLCYCY1X47Rk19Pgy26yKidU+AL08X5Dpum/SknAs
wISTC+zStmpTsS/fakNs8Zlu823k6LtN+XxpKhzT8T04tcCrJYKGmlkHQn0xFHPPPmSvT3w6hVm1
ZnrQ4qzHjcoRgvXSwQi7vc7f70Xp72XFjJJwtqVJl8laiZR8VHcc/6NOGK2HiVRgOyErVPpeXnk6
ELD2WZlLec68VHatX+h5GFQMNSoZkAH8oCsBGMX3KFXwNW2aGO/MldhzPAu2at9fYRjdHNyy3+Ke
pngyBr2jby0YbnxgdW1udhqepk6YzMcb/mTuUNylcElp2sWkkg4QXym9asUnr9Aauqz20DBFuHpu
BchsRdJo6LM4n1BVVMKvyLTLd3hsHzir7TpTJGh/gbQErf0L6mTL34qhjc3xzxmr+E2mPEBpiMgb
v0JTFMBjnE++6jhTw7lh5kvJ/gjlyjCw8rIEUTKiEHFBXsuyZBPUXPVKnk0cqdaFsQeC/Tm3WHEN
TriH0qtz7SBuXELiUN4PKpQPS82+oCtYImGH80mRT7y5vHObVMsb1gRAy87NstJ/30BPJMApcd6N
/F7WXTurLu8ZrZLZ/raV8juQFJ4zXwxCVrCGkCw4MhiWcpu7OF9cbYTRv9ZdavjvxC0rwtA8HzoU
Efv1QogWKFBtHAYHoQSvMqylodO0foOUBmQg+nmcKOWvkqQ/Kn0NyfDiSi0oug5m9VbQslMlbT+C
hBwgsJ7BhI2mj5PaxKIZ3FqvED19GvyWyeppDJ0fX6Xb6WlCkEAEbYANXkr0AV313ZXipSGAoKjF
S7okkHpJOzg/twbHZ6PKdWIdEFqv7X9R6baFrQyh61J+JDaY8ft9wetONBEEOypqtlp3N29KjrVo
VZBXXOoYbbqPZmCCr+3Y0CLkXw5LAzSScWNyFpckTBQOcO1PWVXdboD0r27FdvTmT0m7Hp/ByMXw
998TeZPdnruRQ75jqs4xdaHOzOdSwCZd9j6kIyI8s/4UC/3zFsuvnSz4obOkzLHfYMGMgYNJl08M
Snwe9e2l31ORV1ZhzA0PI9AtHQturr/SF/O2adK5u+aVxpsaj5euT6rKRAfZGMukDOOE+cd1IkfT
iFNVyM7JSqJukJp3fRL3yfsTqXMqOwmYc+s9sz9GcAe/OtJBMaaNx+N4cb+YBzVXVA5n7PQy6G1D
dVc2+PfWEhRSg5Gn4edJYsnYq7zOzGR/UHsHiZhiMohwIcCJgz7MDVg+sGr/+RaWd36aThfwB1GK
tAKjLEJvAkqH6jgbG+6+FPM+5HmzFW5wg7tejId3gnoY8bJSh1P0gej0X7FaGdqguHTNzxVI5jib
VuLOzTOGCEhvY+F7t4pFVV0kuO/+P8fH3/C1rO6/JEluhcIxrtRYM247/qWgnXeK+mYX1/+I6L3n
LP9S8WSkmRLpJlqclnpQS5X6bZNGiDJitgSdHYo7sDd3yTEMCMIcb6aDTCR10Q80a5EnsZxNlYdC
d8zzM1gd/gBOuwt8rbVgvB2OsMpRhwSfzB4LT8bjch4DvzW8qbnbe1aIynwTURX+sx/bhy/kcre7
Ghp6u1T9jfc4OhQYMwRovJB4Tgfbbpj1CJG9cyXywRgNjae636U0lV91NN7rxCwi2rj4QIJeoLKK
lQXs13KTIQitoG9KiFbHBy+6XtJYJF8cqzBHsNjWwpSC/6v9tB9N01pe6pW47udU6edT2oaieGpv
a3pxGdaKpfZaXoyYlMa8NiOeVhxveQJSZcecV2Voo6uT81qBWRgad7YbY9bzayDKJuqKl9JG92HS
M7VBMWXqYI2pRkyjtm79qkLKZAiRpK96ik+TR9ocuB2W1W8fZRXu28cSo8s6+yVTQhsAN55MQ6y9
+edkOeGxJIMyPHCSY8WfEfsY8sp/AZVicxeo5P50QPIifkhnymGNzW3yPXHGtxfK9DPfqPp0FmpK
GdTHQ5v86m8PK6knaZzd9ipMERf8A8rXBMCBmpmZV3uYLPIl8XbYv3C8KfL7cO7Zto7GM8Nsyuui
g1EypInnXrHWXwQf5K1tr74416M6JGimbaJfUmwZSsdoFltZaquzDyHZn6fe/Avh1sAv9MBXZuYj
P8oU+OsGVkrjjf0//wZOHencJiQnafrZf4I4GSLLOvCtS9eHL2dELvyaNZw/bI7QLCBcMfI0wduO
Tjdo0IDT3PXRiK+71hrQjufFVoylLyYGshIunt7ScmjkR+xg8e6KUUagQNj9P2yOqw6CjUCWUjVX
5lGsuv/RKH1Fse+cUO51I8CWyBI08o+n2ZP8QmXLxaSLISz407T1cvbxpnSbpXUMWzNzjsANQ43Y
yHrT3vXKHzvf+3JmZ6tTmEMg9TfelPgNO8KsALUmrpsIEeln+NYHzoB+2P4nP6UtItbyonbpVYk2
mRk5hD9hE4RUlPBOF9ThY+5y8bQriT3kRVtMJiwMjYcrQNUUfJZhaN41lLln7RYJIRv6xrqwM2JC
ilSro62noW8SBsI3sH6R06UTnJx8/vBtBn1Tk1RL8HDwYuyog3664MSZxsIrEdqsBa6s18DETIYB
KfwhW/dExfylNEGiewJpI11Axmi4CWvvN7pnihwYoF59GLso9Hy5tL3nfeciDa7jbBAxFHFWWgM7
IfRjV9QtjabaA+Vrg2fzba4pU+HDE6S5e4f8MEGZ1o8ryA93Sa3QA53LGwKB5pdlSmG6Ez8tlfQ9
WKE+0ZJ9pAzaeMwknMss49NdB24uEsEEc6dFZMZGk2IqzP0ds3wzkxDgK4oHgxtyRadX2FfnVt+l
h6+zW2j5Rze4VKUtGH2X7aRKCGzFZnOtjjJPE4b3uFqWwzRuEfein6pBKGGy7L3JAEg0nGWV0+I6
1pRaBhrG23rxAp4ZLci8WPfYwda866RhhWzsIfyuf9UYXTVa47l2/WGH44+etgOiOFNstTYlNT3N
OPY2r62zLYZZs8pHhnw4WTRkNImrNsRohERPDJzr4H4ys23oflEeE+QLp0bzRZi0If87FlGt4h0Z
d03uvhRiUpQV5BcQkFBLvbofcAWhQzXU+gXQwPljQ7MWLCtbHEfbsUEV8KaEajly6Is2gjRgL0ZG
dW9dwTyFvRA7iyWoOpr85YboslAlmi6dWZQDO1/fTVNq8BtKdRKb2eAwsEzDd++KxkoLfi30nghM
1tgyuSt1jQhpXBwevx9zcsO1jyyQITbU6Z/o6AZ1th/O7D3MRmu9oub/67DiTJJtPceINKEwURWj
n2XjKCLUsFCJXethNCw/QYTVZXwC0emGrp68dXj94q6xNdlJQYFslUjuOAgc+hHbGaov0ZoiEIBy
JuGBLwXFxMPE6cyTRldkDX8kHaeMiIc7zwE1pNbQjmucAhge/ZLXIVhdMR0qQR+n8zj/VW3FN/1+
Q8Uml5ltm76A0DxPcCpQWmTwu+w1WAH5TC9r7sZ70Yu3uilqyBJlfMfse0c0dkMTx9oHcV/LDKKN
HnWwAe1XN7t0ybiO45+S0SP5T51+AHDainJ8XrYohwAHl9S8DXU1IfMG1LZX+2xMI9VOgkRNyDTF
5J0u6+2UHAJe+BHXTYnMNbZe4dwleGg37Oz9zJzjtUFEMMaFD08pUx+kIDpqcwoi+12H0rTUy+b+
TJbfZc8Ex0fCz4/Ml2EhFh1ghdVodP1cPs8fuei/Eb/03zKJ85h/U/0HNbafjcQJP10lW/Otpify
E1CTdiaQNHIJryDbZuLZmUXu6UoWCs/2lXhlhtfOqpecbXktDmPIQ9Tw0WWT7xIP10Rt6Cb+5ym/
uyECnNAuMts2qDFX/bRtD22RevSYlV3craCHB/xUH68ElYo+f2jx3Kn/Bfm5d5d/M5xZOFIYFfCV
Vp9hBuTmXGS4khVAL0bWsJSqYtU8J7quR0jldThzZSw+PoIUVZ8fUsOHB+nYyjKPGP/9FUdBXgJM
LNvLabb8TYABvavzmMzyKHvAZTQWunAacLuT2YTIUO5LdbeQ+zhe5alGRsmo8kqNPAzE/XMpI7bE
/ZumwTXAhPwrXRYHhi600GTwd9mb/SWKr/rrEMWtbW363WFTPPYuMTaYP+Jkp3FkR7/Ao7A1Pnbg
PXQdvs5uHOdeTh3jiK00CMrIJFNDN9uSOA9dBal4z0eKBLfLq2HDRnGIc9EZUjr4xZemmyDy7mc+
effNiAgqqVENtgq6L9RMYXxtbG/som2ADt5WnRqT5X7C0TCn3foMxvNwq7E8eb2GAzJYpvkDgCFb
OJXvX80gPhedICy4iUVTZ06l0hru3PHYf/qkAWlPXoG9k0yxVn1KfptTNPuW3iHcE4mc/6deLf2e
YUS1/m+3+ZbCQa5wrgL2/L7miwc/DgEM4eXTXCPLGiWEpGMnZKRlKYwlT0cg4dZ3jacZYHV7IDnR
jxIrQ8tHTvcdwTrJFT/Uucqz+ar6QggYgCbEJGJE0klXElKO+NYoPdpxDsegcZ4MTZtu4EUAhWNM
6mrFra/4cF+YsMAWZIuAAQADu4dlmnzXDVg4JMgZdRLfkiUYZFcdjOeNFL6ggsdMnWouwzZoT19q
7JhTqRUccpPVp0PbTApoNBo+kQDt1HciLboSjrGbiUhnsB4tf4TPs6pNR0lScBvmMBhMZaTaFhtX
x4DEndv5wO9e0XVIVJR/K+QYWk/z84fdIcWniB96lrfOJqoWnELbkmjPdWNMVg/RSg89EBZ5GFDI
GiHAD4TlWnIlW9ReoqsS7MXG3KmKVyCeHK2HPNuMUWEQncIT6ZbIz2W2CkmBaJVjhxaDau9ADZZt
wXqhyrD+x6gbPjE6GD57Mx5fW4+t6csRTpPCOR2Olp5utZX1dVd5I2A0f8Fs3LNRfaoDona4rHBd
wxzlMRVOMf/MDipHC9xRYh2O/qRjbL9p8S7yhIMeLEpaoCgz+tqMap2srSQqa9uIHlYlqk614Y5J
ysN/siuPF4NyPQznNyWKBgG5fEcQf/ni0dijtl7xSS7seWh9Vmjr7gQISoIDbU5tKEO+8I7/OdSS
aaOQMTyuslo7aPX513Z+dxrf8NVQnZYT3GQFMlHKn1RuIIFtZJc9t8oP6Iyga7S8d0JLG15z3CZv
hI18maYH4VJVCsh34dzsoBmM32HMAlu9UkTWoPhjQomqjlp+MHO0qhAZczSX8E/U7igH9aS95zAK
jJCVteeSzyp79cqYTd3wzCHaD7UO30FJpDUB2VcvssUgrkuBM6o6QOj/kZjzVyLEqhskuerq59yX
TToPlc2zstO9g+RTh35Wkv01WaxrSdIgBrfjbLmixicYIxnnc2LNgz2Gm2o+8OJlubHHwJjfSFOi
jWaPS1RGFyEl8l3rL+UaLOE4cCA/sVsXor6TMlbKAqreWSkk6EWOuRgbpbSRg4JzBkyXWP/N8FjH
c2OPUDYbvcg/QDRjk2NpCPPEpyEfGHVoD+kOhuY1RdR0zvV1vOnNkulC/bjM2bW2IIRYyU3gqDX3
ycRxvx5oFCv0fPPEWo0B5IOGHDeOfTpXFwE46F7EMbmsfG90J7Bybe5lQz+oCypECEVXek/Ipg8N
CNHK+yIMExZ2HRiV6/2rIu07Gl1aZ1KDs6qP1+JI3EwbLUEE4ozIvfX40p3n6Qi5qPcR1w/EIB7u
67o7Waw/JNzSkPuMI//GG+LcAcq/X0XQvuvJt/u+exbMTSnvXMhGiHwUCS48/xMSjqiOcY6Um4dS
hWWdKUbp6fT8xMfa8AnzDedX5BYIfkxoG0FxN9HnYzPIff/pveA9OFsd6GIm8WIamlyDcZ30MLUy
XH3yHAay+zDj0i7AioAamz5E/gWeGpn1S3wKWKmXtyk/Kp5j3exnIPJx7KHhybXK2B9gMI3ujtRp
vXCDyExGDXu9Aqos2060eKSNE/7fNsssLsFVAtnprYlvGTEJ8+dH1U/7JweF9okZK0HZRqYpa2Jq
fnyQsIKASxk9swPx/3H14OjEyn/Yz9RXmz/eiaM/WdD2nGMc5exsGtYXd5KxQlZE7a6x5cvJaisl
WDv+r0T0v4dF+hDi8K6s+QLWqNxUe5uBh9miFP7KlThaXmexWiAPge0QOz5CHT6/hvxypGWyL5mO
qKgQZlSxurT8mQLQxZZLWmFrwa7QQHfMNorBt/aM8idHxlxU9wPx/6VyrVvGM0ew1GtU0zHQHz5E
965LQ13QYaRvRkSnIso/jkphZRJlJCxIS1rjtNUTgn3kJMyNqiJOjDmGQtE6UFEQVJ2IisQL7UtS
Yxa12cO0s8z4Tr9UlsP3a9dTEg3tNsid40rH2vvB7WTcb4R8k9z1vITXcGLgqNm0Vo1akcXNEXoU
lv0sm8QUkZzjbC1s/5lhmFZnx+7+BKt2U/2QRN4ha8Vi0HGiy0/4/E4/ibBHor/kEE0BO+ZLchsh
KQMk+FsSXanReNFXnzQmjj+p7mLYivy8GkXdJ2LQe+1fV8Tzc+hng9qbPIjoIv+t9RpPm77sJgFA
J381O3mPLNPzMwa1FIGKMvV9UhATWMk30HYqkGcHR1DZ2UZMEXclt6/YwW4Uu7OOmMy3F99MwQOw
x03acr2wBHzou79It+jpU8Bd9DR4t3Hx84ZMbXuX3FA5AKGOny2QTmRe0dlvN42oLPm8Pj1Y/oEB
bxZPo/CNjLNTy0nVKhEpVbtq/k19Pbj3UblnDbYT/jCjK0cx268JOV1cCwq7GCg5QIECqaEWFrmG
LEDyYTWWs875X72XxDN1ffA8xtN3D5iICmjGO5ya/trwXzUlegvYdGQIYrVlH0sPlHXsdVzkhMQJ
QDwtWAAh2d1NOQcYxf3J6E/UzUZ6N+h9vRRnxF/HGQq0RDbJFTRssoUMMJOesZGXOHNXpKmTtGWr
H90gG/h/Cm8nQyUajd6pKgKxtGzBGwO2VG4o5onjY2KowiHyXNQcmTJwjS08FMqXjrKTAmzHUMEV
BjDJPYD42x/p4y2GgUdqluXnLG5v+HJTXlDDwG0ydRwR4ptmvYnIHW6kL5/1QBhbtU/NkxAXuwh3
BXxPm4KDZByZMF/v8cLOmgRdGb03POpADEMPTspHmBNpwtt04wyK2/oMRDEfUL0I7SbtQ0HK60je
grGd0ovBIJvVhAR0Q7LqJ/uV1TTuj0RjaJKrIRNGBLkPyotshkF44k7w56ohqK2DHV/f2ZR+BOYX
+2dlDoA6eIO/O3F2/XF89KbJNxI9A8ZmFRvKnJZYhz6VpLMlXwH7hzcUU56dqn8gn1E3YD5pcXhv
wjb9ex9AwMLqtSviPpniqzXHbJo+EAYf/yPkQAP3v6nQhbMJU1DtfknoUcERQOAi7d+1EkDosbXU
3DkIpkAGE8mwbmEFDgJ6T+mxuOXXpVLpgcBtAmGEkKLYYTsQyVpkTaxGxLJuWA/nZvIT8KIVxeaZ
2QZWxeGAgDY5ean5V8qgSiyHd1S/60DjRO0pszqZg5LfKfgbjIRQmGQLEG8j9PwppqmD8aISeQTT
yQQPAJ9sijBRDXI0zMZog6GMpGIl1ku6B3WY0rNF/tRfHW2y1QSRDQnTu+05PvOMTrrzd67iGn7U
a6bSUpMWrDRbbF6s0CuHTKK9KfJj0WUwMZzysC5soeFLF1jKkDskW1rTfKKQhHSRkob0rnG+tdnC
c2HQakRU+ikCttLiX+CnKmQOy3PotV50Uy0yahTBblo6XiCTRtDlD0/PzXV11ogDTLHX6DYK4Ppi
2Vp+l3JgX6IoDtKE/Nj2vea5xKI9aTOO8xMRTRNGbG4Fjc0hosasTX3GGLgZLPfxBGQve7pqxwuE
ZPLXiQoTcDlOZBqXda4qb2ZLAJiDiyuUek8wg5mDUDoz4MGX3vVmEogeBUKoX9POF1OO3G2HKq/X
OkUT7w1+0Zd2tTC3A/b8rulzC9ujkzJXO2epljHSXLkUyYYo3VRgeZarqyuwCISa+inWZ6yj26T5
KLvsI/l8yfxyYQvpI15Y/V4H8J0dzTW7Ttl2SdCxGlbztBllLq71SHm5S+T0uYLxc5gYe8q9/mLP
M9u8f8lABGRhuVWwqxnZfaisTc0631trJvIYws2E7h9+5jPmIn9PY0yMdoazhDlfBbk9oXupVNhF
v253+SQefm9/0WTbVkHRMuvRGeOQfljlQYusnf/5gwQsDgOTjH8LoNcBpGmob7tHDrpSZvIKKCqn
uZmxrd28EsqL/m0U5jJr4DfddqHkHfZDV81/Od/pdRLzNnAPVsteEfonqY6xA+nij6ZF+bKbZFC2
V33w98Mml2x5eUy9LObd/AtUc+4JYlvsbZ8jFEhYrVIckoJYzaF/tzezNU5Oq/vtxZX3epjPkVnW
PXfghtZB9ijRQrSIHyLfQNiHYoz4UkRvmz1HBMiFqmM08+9XDzJh6MIc2vwf/wf1pp4opZiBdLGx
NTPwyXBlxspLlfRE1t5hd4j1G5NrE+2eKDxzfl5bdeTXizGuOx1YUpjFb7HMW32mjY5IwUz+KHj7
QcfbROAgfEwnQe36DMOd2WnrzstxWhop+BiRaP8yp16ScJr5V2+Vww7k3nN1dOMStevolnkqw0wA
Q8Sgrk3Xn8acIsALZ/s1XfBeeY8gRKBilqBCI/k8IGZFshHXiNfLH1BBCCzdArmjuDgSeaDsLgz4
ZAdI7axtBOWO2z9ltLRGrpwvZxyJG3cokldCyGzRK5ISApTnAgaeS1Cb7uKmfSnDzZ+ih/jfT4qR
F/28ymJaU59MeG2P+r4xtzsiv94MHAvtsaZEWqPDzJ53ZC6SY/IVnfJQjxb2C6epsgE6WZs0cikD
Hqn7xrdFFKmxt/0PV8k3u/XHQtxGtRxB7jE/pWiHjIzPdd8X7piImkqNanoe9kcRNauW4bg+jlKU
oxBh6NIqJ023capHu/ce76kmK8TcxTO67aF+POY49wiElaa/cCwRixiA9JWTMYIXrwxf4KEpav59
7mhuk1E8+Dsf0WAjqOcj4suiDeQdrhLGwE0Eb/W4iujiIGMlxE7ZuWk5kDjORMoasB6iWVbmedWW
8ycDVomuLtPwdtIJzSpQ0TI1qbNoM1uTdas6QIjyR1I+DIxMhbZRxnSN2GKWL4zb93pW3kBPO0H+
hfhlKVPOt2wARmGm+cO7wOxkIlD161LexuY7v2lGOiGPCzyP5URcTLSF/QF19Rdg/RZ5AdcFSpcr
LsRQtjZ+VmYkS85cHzu1gXpcRqG9xcM379rV8yQpXDb9vbr3b/CBQaRinx5BEuCMPIuFGgv65+kC
6Jf9nhAOYcK7M/gD9lbfODhmSvgQd3aglIz7pt7ivnbU+t27+pLWWNLEphlTfklm7qMj4s+n2gIO
tS4ZOgMKr7fsrxfvMooUAOy7+RUBNGB9/PmASXSZZjr3Dxq4/ai3eeWCdeUP2ydrrcfZFic9PEpA
FkuxPpuu3PVIcb0s0ep4vmBDutsneOsrBxsisD4x63WLyZ4efhZjyEExn+mIk+z/DHy0m0mqXnpI
j54DMuL7v7221REntCDw23oSg1EH3ujft4Rk00kJUwUIjavAmhtlwGLB4Mx6wCEnIXGKN089ptWS
JoQqIlOWoZXpyOJTy6P6yQf9M2AIxBTer5W5bS1ATaM3sfijansFcq1M80EXFl00xeo5YUyYSthA
Qp+RnQxD85MJ78wUTVQ7tbMIOgB46yXvqAA6amY+DbZNA8VSPAoRdJN9AlS530RmB1lA//ZT9JTn
obr6EGSE4o72XiFTvVHqFM1jYZSPG45p5CnHT+/gUKyTaYe8g0vRPn60MSqSkOBePtqXjhk5FDnv
0JHabzOP0h5ueOD7IFo1tjeeSelTGLOD5St0GftpyGbz208fh1MgSKHX++RnCUooz54+HbpwfsH+
UGcBoYkKmgBEmg3TSftJX8Hr339cJtD/op56pLIyWV4NeACJxo0EkdymQ3dwDGPfYn5rjKkqJ1by
p2W1/hsacTKTgAp6P3XQYV/DACLfmOB+BzvzMXiCoXJYUMxVw5PmBDVFXKhuw5UpXTl3NtJk9kmJ
TXHdGrQob2oZ89VPIL7INA3PLLVd7dvhj0Y329KnzBnr+aBGEYsibfGiInSjQIVEYfp+pbDvSyrD
nVQ5aZlpg3dfQNPlENXXoMIc3FqYoa+MfTsB/3Le8sBKi4O0Op2IdDkHVohPMTdEgBQnYRvLx1Lk
CCq3wC4oQAHJL71UTHNZiJjNYU9RzyfHONAD5k/G28kDVncIFVq3jGHAvA5OOSJJuhT4gsi3i+U/
oXsD3seHg47y7/Rl5eSIsmIXPKHcS+8BxWNVqihObpPw9AhzH8qxxs4zkD8jpzPtP9QWwDXfDcZq
V48Ztyy+x7rIU1SLa/Eb2s1OVJzhQ/7eoEUpxsjb9LZclZ/WmHrE6ckARqvULgz4bPm7/TNL3CAz
7bzJAhp4U4T4U13q8lzTQDC6xxqhBUnJvs5Gg4fDNFxIyQaIJKuPZyZxAa11BjzyOet1CqYsJxNw
G6BOQE1NSVd8GJCHLHhICwYZdqss50xVvsAtImIVbmp966CdjIKu63papzfiOldh8AN6Hf9Khi/I
AzvIMKnfCFyD5sYC1/FrENF2M+3E9BlF7UMEdhoDqv6riNSl8u3tYrOxFX9mUUYIoYLS7j4Mjqjr
kmdRdTKLcrQy9i7gWZCdW18SgwjiQvl1JASQu6okOhlciq1k8Qt2OguSuiFqLsV/XyZ6cUaWvcpV
OOg5YYRsLcD4lhlp7wYMWBXhulyfzHMisJDB5Rre7r7aQhgA86y7F6+EXPyOc4zTdowt/jLv+D5d
f2YZKZXP3v54CBaXV6nBltuyHW48Nu7eTmlG/wm5jwObTfTLEWFqlRFQvyTSXFFb/iQKVvbsdQ1K
k7caIot3bmOPNweE1BkMgWTBJ5P/WNv46rdJ9Wy7QOUBFqbFBUSPjHcwXbyK1V1sKXekXXE+UkXm
GC7PEQdyIrey84dH04r8mZMv+6YKF4Iy1RvIliRNsnrd+qiXYl06R+yJ9bzaCFgOm6IfaqR3ingL
EKyhVTQ1VRLpLnR8szqlC43T73eS2wpXM+2n24efhNai8ImScwjUxtEu7ykUzw3/vxzMTNgDhGSr
HIc8yV0Ajs2eN1H841GQVeieOrAp7dTWHOdVufeifTQrvBu9/YCKLgudmtbg/hTGbnLvYn0WTTDc
tu1Q01PzKBa0nSc1uwCcM+soRH5UwQje4b89kkBKAW3ZS9YQXxXgF0hsVZh4WpzSQw/Fk0q0Wukx
xjYp1+0j3kTZ293yXGaj8tAWhDU922dDzvV8h4X+4eWh8qF0C9Wu2lIJgtgrnOGH7E5MaFtthUmM
erfRf1+AJFWdNG36KZWt+WRxh9yTQbxkPrPpufjA8MwKmwuYzjWiYlK/HNb9siKJVuHwpocqinIN
bO/wOoy65++McNkAfnGv/dRfBteuua0RwBOgaxBDLg3obQ6wt8rrt3zNapHotkDqe7Ks4Wb7yb/H
GgD8y4tzDWq2NOXdjQZNJcczfR30F38GSz41vUKxX72GqdL9axQLpFVQIG/ESTtJnJsVVoYqtZQ6
Y9oSrpwbgQwbCK8mKsKu8el+5l15/RkuBpKRh6Xp0n1gvkf9AJIbw5NIMTtAp5HPjgVctGHR/y+o
LuvbVW/fSj86BEsJWp8oz33JTgjlf4MbxcykJcR4+erxZalM+RAhg0yuLGD9hgmMSvnJ2XPn6LQK
g5pLxJlvNLCniGWccSH3y4/PeUAo7p6yuz2d8O+fSVx1CqUgXzlQKsRpevfA8R/tbLTthdbEoGQ2
9sSLv/Vm8HyijwJh5iidW6unPVqQYVby1IVN38ncbCVQ1znSmMVxXJdiu5zNp7RdvCUanI0/AMhi
FCPrWBrdMhn03hTaB6gYXOag4AKX62TiB8RqfklRJjYk4EV9CJm4tppm8l2EV4vwZjS1j7hF/raH
AToZoWClxMGFEGUxT6xLRfIJscdURoPfRqNeJuWGvP3sWF4LQE2znnhSNHU0f+El5UPIUWx4rcnk
0uE0kDxMy5LZCU3b5KbtCC5OTqZw94RkV+gYekX3xRhzevfCnOjmeSSM9xEvOqLznj2xCKtAJ0R6
foXimJ5gg5W2DnjDWtWHY5zWpUlULD8NUB9DIgJNugzMsejwrAIjG1ZShx54ZLWByfAEMCP46Xxh
Ujc4SnKG9pcQrPFrFGgK1Qub3nrfdNbmrLP5sBBpd/2lhViF7MQV5R1hqmUjtH082Wn243ISXO73
xzhOH0bDP+2xtA9nVBMsEI9liVuPEAYnegvyeB01DpmN9fY+huOACzXrDcKSwcXrbAMVNh917Bwc
4hA7Gzy+oZsGCdlxgm9XwymQ9NhPyEbe4tTlsDyk5qyT2mjUtXkgxbf1z5Qz++j3BbmhEGVf3ToV
TqOU0W0tAeFkj+ax0vib/JEmI0WXZf2/XtJDSc9DGvII1HwnZfFKpS+kwNIKX8oTv9KlmebIUiha
+TP+L6rVCyVo9b8XDypMAxi9vZ2+tNNcd4I+1TBLun0GLjmjXzuw+2HMuXmsSHR/O3IWHkSJ3PFF
qi8360LK/ADxsJd68+dOOsNyGSkU2WazWMDMzeMi3YOW8wJfB//CUa+sUYz5XLeNgNSR6y4pLjmu
sopB4XGZDxx+CBv1H77AopH89ZiNF+odI9gBCP8Bj/leSkqT49vbyCf6FaQj/K9A1fof1dm/otOU
pdMK+HKQwM53N+yP1IFSyfgPP6d+k/PV+nxFCWThHykJfexpsf+/2t9n1QD9ENepzsKQ5OCqlvBk
OCUTjb49u/dIO9KvSH7jkGVLHB9YIXErPoAlAQ5QMDKvIS0jg0d86MfTq2Yub+Yi4oJ/Dj9rQi87
Tuu4cO04djYeqCtrp4iYFanUtzDihT05FsQN6LdT2dyxfHmaKYgiOaKrr5Aj8EIX1O9Tr7wcAgIF
ssdLZLB3NH4i450XwP5uY4vFcEe9bYWdjS8Ess/tJjS73VuYs6hg9j2yLhj8LnfkbQLt0neSuMjj
jqBqiqEgVgzd8BjFTRNDVPCbg3Z3cSvaNoHL6K+8vsqOavC986iSxzJwb+Gx36XI+9gKE+R/+KHt
0Yn76fnVvPK2jAZR+xSm5IH2ULjPdI/Rxo0d9XP1TnD0VyL4PoEyv+G4IyyBI4pnRcp1OfvPZeeS
6WLNbOxJSwhyfsHcdcwgy/wXWMwRN9970VOBzc35weSOeBOWK1NsJVh1eRXVslTMws6n6UY2GcX0
LiX61WUTG7LI+YaPgz3dmKGb4d1MfesBhqQwf/NM1If/BvNAVyrMoRyDifY0WYnPvyWYgzT89L8b
VN031LuhJz8i+f7fpgNLKRn9TGgcjOSu+gYi7Rtn7+TaYisijL4hJ9lEXV2VaE/VU8r4/TUTXxCF
8eGCGuybaPGwlPS9Djv/bSGHWU0q9KxREIaxpiqa0D5AY1i3RNbqWU9oA2VSNHBQ4wnF841MDX0m
ybPlLUaIIO6pbvIieQ7Jk1OUjvqxZD+NAvaftAaRPlyMMldhTUfSI7Jknb7Pg7VygC4VUUVXu2us
sk9gbeE9aMlrrJAv+omjIS65eOMTGeDxOUnFvta+jm/im8C8R2zv7BEGs/lMLIooA6M5m+x9uBJM
H8BmSCHTEYvCyk3UZ1L8fb5+7PYiYF5n/zMF/Lm4IXcxVv/f8OWEFrfbwkmH993XJWfwVBLT5Xzk
aiBqEWD9NOg0Jke2j3BWpzA8Gt5pOBxenGhDIRLOBoGsGgvLQss4ilrO7IvOCPFQNDkgY88CTsLH
RL1hzZR8CvweORiW/dA17rIpmswFyoXZ731FLlSxPdXuM3u6FiI336dH7JMZncwRpbcACYdmNhKF
HlMNvoZgLq0FKlADFiejt+t0DwMrgg5EOEKowpBt/T5753VODtBmDZBwfGw4xK+8wfSp5ZG0y5kN
ku+jhvTN0c/q/yD/N3Tn5jxeavc4KkXwUXWkFKGEuBuBjJdrr+7S9ml9PK0+Tt+px6+ljVmDb+on
nhwCATHL9hjAyuGLVcHfeCXiagTglWb/pLoVNC8zkXPeTOSvA0rDgMeTyGYBjNd2CFKrgxWDtZ4q
oDryIaelu1S1yIr2zGR1iDkLdVaTAMcuSzB/FsfnEwjXagThE4kqjUtyne1kr0rNWtsIWpwNM6Eg
jIXs5BGAD240mg9m1QheTvQvPTDGpgNXXZgGZ1tHqCkBprHBl1AdwELix/A0IJ5ZM4WnzUoHDabC
IRLTvwY1LxZBeWn0wqqzYsPyoiBt7Jf7Vpmd8R5Bx8yP7yn3CcSPXfcPwyX4XnVO+aCCwPfRTbSZ
5kgUuKIhVA0NnfT9bu3EkpgGv/Haw0Aa5dNCDPPOsCEyg0Gc3iIIoAL7hRYCYBrW64kT7JeGBhOV
mpWyyNA0b/Ep2Cd0Jv8TLRns1piRLtitoSEeuKMkR/EwCaBm5Pwbsp1TSJ5F/DjY4HFYjTVvfrck
PxZp3NTmZX5UYVU43XfeAn6+PMIZHBcXeIDWMqUFY9sKFGD7NUGpkor4ETuCadKw5Gi3UTpH9V3R
AevuAhYTIjKM+vTnLRjVDQRgxnqpXJo+au1kNWczgkUVfvkoTilQTKkn865AJlf1QbdxBcaLW0N0
Rbgi92Kk7Vf0hWpLepyNRjJ/346Ebn8xQIHJn4kwN8TjQI29h9VdbqhiOJ/FjkVp8KJ89mxjZ9cN
iZ+vt8X4n1+/e9u07E4xX6eYA+wisTCpALCYl9LTjVq7ydOJ7T91sBrNIPn46u6QJsHN7IfJcN6t
jfSUJpiSWU/wceUEtWQ26YcIC0xI2OHccNRgI3TMg4UUeChvX6CVap8ifA3IfteVTUQ0dceHmvcS
XgW19dLB/lQA1SHWE150Zfk12yyhvXaiEXfRe4TQFlVkfNrXjIAq1cLqivVpoHZA7TxRhR/4O8t5
5OCWgdRH6rJ1kDNcTJdH9Bl69NOqc8bGiTKHqucm8mLID9eQPWEg+Zh4cEblMNHoXEzJZcB+5NwP
F44rpn+Eg+DbggozzpAgf/pfT2ckz1d5jRDeW57/MT+ql+CyWF2i1zVMJHJPm4cKUyocUXGX89mU
N/KVSJc3Sm6Lw78lL4eX0HJLxU0XJlPOyThZOBmh0fhYU5FRE6kx966ni/xJG4pvbYpFgf4VYMJw
oFtOECzdRnj3T2f0hjgGsiBeoZR6YRdQbiHNY+nceEAjwVCY00AuNCBbRsvkcY7g/8GoIM9J/n9q
4/54mcJZ/hkw+2wwtKR/J+fdQqNEL5m7PoVNuwLH+M1BE0rsh+09EP/h9/p2y/h74d0bsXtFPKrM
JKnsdKpm5jV8c4KKH6xJl/waqUVkzGSjyLYQpzCuAGFFbxoalOO/0W91IQBdbhj43jLJRaPQ4nbj
2hE0en4hXaH2FyQMlPP8LcTf6no4dpdgPUOlmqzIYq8EnCycdamew6uWD2xUJZxeWCqQ7V7WnmYG
FahRHtpcyzgK0t/l9tH3zPMjCOW3xmgGxfm+XAM/l259pz3ciOLkCgBnCCT97sZukgxa6bn6LJo8
VyUkfUQp3ZqZcfYsX+wSAVMBbxJOS3ZJnJ0eNgVMXyDK+FegmuvBzccaObMaoKHx+D3GdvOoCeWn
6+F5kAommr8AzbqVLJopgY+KcvcTEpB2yklwzeiCCoXtMqRnSEheGJPHZzRb72ZjnXSIfGaa4AaF
qg1GSiTIT/u3Doqd4f12n3jzCDg0QZHJWGqpG9agt0lLvpbn4pbeg5QO1D0OQaOGxgfNq4/Pe3oy
ngG7SgGfEzH6/9UebtwaqasbNxMxobHHzTm7lW5NggmUpEA3QBmre4BqKmuLW5xhzTBozFPjaM77
xCzeURttznU20vR+8bHf5m/1CiRk9ebl+J1qPqXmbPpQnKEklD5iQ2uZzpmGsPgi3bCzv8PCuqp/
WpA2cnStoKtLaDnYxlKIE1qsN51dXqiFRE1OL1X6X8Gbp0zdGjUBF9D9p6dTCXMpR3tsWYDsYn+p
MpEsRAcxEa2UKsp7ll6Hw+ekAQkRNKeKPN51pQD4CTYL8Xguc6AOt2CUoVeYi1kD+E5QyLH5I+kG
bg5tIIfKdFW9SdbvjwELai033zkODrMQkN25h8j+WYba1C0uxa3FQDfX5GWBFBy+SovgPXaiVr2p
jelEQMjCdWk20nSEBtG8HzWKIZ7vvjlARRdn0TSMv44KZZ/SaPerzDF6ftiVAz+dF3Zsf7PPSCdF
WQntdEKX3aqivUCUUdcjcNtt8s3h7p96N0Cul5E+cwkTCXo9ewWBJYB47fLHcH4G0awA7hY5BjSM
z4tte37XFe+5SEbuIdqE2WeGiYBHZPG1Q9QDpEzL203VzCJCc98frjxEkavetlNTr7u201ev8zHD
lq4SwTast79BCS69z2JWb+u1rjTskmjOhSu3nXdiXbVSE8jkf9ebEkOzdUnlUp5JLKHC2qkQA9sw
TlPn1l9nu0Yw0kdwabQDHNRPPSXQtv0ZZqmp3c6u5xuJwKJSaKp2sTRZOGbYawV50z/rH7EPioAV
z2Re8J7MIV0t7WRATAxcDuItvKVrrSxY67ddMZIwuZ0kETD1aABScuia16gWzdCznfOa7sIGPsX+
jg1w9I+avM4CYL8jJB+gY5sTrcnB5vHY9EccHZnmIv5lnhNdgbrPK8duqi6QexlWYCYgbfyIpISh
xwuEvClRyov1iYGjPdf7V0Amqe4REKXZPWVLG+0xfwVDc1gbqApEKVCj02KqebAlrhhYS2E54K6x
lAw0c6bA/mFWZDXWhNJfZaBmapzg224b1RVXVID1OA2UelFZlMarNDaWB4i2jyhzYI48ilonKiDz
4ousoBdr99hL+vtXrDTgGahulgfPFhzogJw4cNuJv7LW8WPeWAMeKNcf79emQQ00K8lnNA9Y8D15
wyM8oM6kBlqCu7/yPIh1u/Qk771Tie9R8DKTEh/Ce1W1SlZtBdLY/JEZerva/I0H5ne/01d7yxzS
UpacaKwyuQ+bENHIgLdqph2bcxTA+NpgFgf47dJBBYvFxsy/58Y5azTvQht6PwyEfqyGCvZHlGB7
CDu4fAeidEM9JzDku6V6Rp83qpAUDrfnHpv6PmoMPCK3k1AIAL6ihU+1muVLOulRjg0LQXhxRlh9
/pChmq0cZbO0ZdWjk5EYlL0roMSMCWx3L2Pd4Ulq9Kr3UwrqUgKOuA7emSDmu5J4pnAjDkU/UvKQ
mdTsTRqj62KY1UEXO1CNIyq65NoiunUi6K2I9i7l3hsUXoGUTDfqd3L9u8z910T89g7039SR+rie
99ueV27FrxqdFQbDcSjkBdbn75/ZZSAdqCo3zT3iT9Gfjrps2OQjxEFodYnvDoGNAnHieU0MbHjf
uOvVAC7GtnuD6292svRUCJgKBBKNiJCBI2nFS3eP772/z1ddWoGYZpEE8SG84N3RaGv3tSmgcoRC
Ddj1NqBQXrwQuhQGH0fp9BAuUMCX4PLM9eDktTIn+Htk6PJo2iuvuTNmqNCIbhYGuMcen9I5ravM
CB6OwYkWA0C5Ryc3oCYSdXpD7u1RX2hA4332TeDIwI67/we/nx7QhKTfWcY36Pl5E6nrjclKx7KC
ThGWFB/dZZCWfOtfPvG5emFBXEbfw0tzx1G1Qcr2U9IxKxol/uPw1ObvdlQrZP9eY9uAgKL37U5z
qCihfbZlk9rgSz6P/dZ+DO28fOJwFMAzZ5WqZl935oKkXQ4ND7ltEYTpxLtL82f/kYEFe+ktGzC6
F9XBxaXE4K0VizA8LEJL4kHCGKJAE7CY9HZ99tk3evbFS7wnqvTeK1hsZz46rDBdzY2bhPU6ApR3
21EXzrcknkvoAyJsaYayr+vI3xMmHkcwxZJUsqHaTiAqrx5XAQqEPRcqgmCVUsUqPAO+20tcAIr7
8eekW10Vf/UO2SqeJsXKtZDGWjwLxJ7rB8DE/8ZAieegWj84BbmH43O99yU6oEa7r3v5yvaT9rHX
zOC7AV3mELjPj83cTVJ8sGLPtfNtj2TkRaDC9iXSapzPaYGl4QSWmWiz8V7vjbRup8l6tLc2seIz
3yUmksCGge1Zp6jwjML9ZENSLto4h7DpFb41gC9yBw/ZOmimLnx/k21dwDck5gAX+1d9fKtsl8/f
50PTSCAmx8/0LjzxBW4yrNDkWI7qU1EivrTwu5u+HyanCpWt26xzIiTQ2RVC1Qcy487Y54Effs0Z
3F2hLgBY4BXWe2gjusjLQXicgCQOWwsTZQibXzq2WJ4D4phR5XiDGK5vITmXw2k00Epee/RbW1Uw
1mEC9x0h5cE1sVqxj08ay4oIPD2iWz/XbTxDxmq3Ik4aUo9qODtElPXP80vpMHK+t7stjQnBNlJ2
HsQ7zKZTKBVHPv4+Sjb3ucBSNjH4WNEb4PK+dtMgkI+MzYy58YKGu1Da/sBAVvDL3znFsbqHsdsm
MzQPwoAfgt7UMQlvObEidarMU2huEFo71gQumm/SJSVcDJ0R6QN1Xy+pd5TUZxhN4sHQAivFxuxP
ggVHFm4SJBSQgfsfy582wCjdsiMTUrhdWdUXrP5CNDF3ZD7CmHNC7+OC8HJIWvmnIziLeV4+Yv4y
kbdTfunI5vZNMQe1MK9XIYWPRUbmUWoHUb+3ENPwrS5KmMjeqn1ZcG/3SrTYvvj3860yNblprAb3
odvJX31Blng0Dag+MBG2yze5UifBiM34yvBuSBEdRmA90woOunbkW4yhia47yT+qIQetxB2utbTj
/HWbayZhHvBBJxj/hfiJPoXNUZseK66nXg/3QsfgkSnP3Y6yTgxXEpU4NahTX5HdshtR/powwvRe
hpNI2oWSSGFgs4OnMBGc0orbSGRvY9cV3+Zg0RNjxytE5StH+thKE1qnqXMCcUOKTJkqeSzGaHAU
ubKI1nafziXQH+5tD48h4/b/NwwtBD4/k/VsAP1aQO3wKyaw9AqeJgBopwcxtGZ74w99mtg7FdUt
w2zr+X8pMNqZMWPOGRfRPMd9gLFWPQ82KXMSsHGg6gd0/6rgB3KGLXk8dKdW+qctsDKPAlVnYhDa
K+x7PAtuMP2gxZItFQKhb5Ai1s5tX0UgNv95pc8dArXn0EccuJr4/iL9bFduJaZM7Ea2YksRcS5E
kQ5+pHOk7iNnGymeKnv3bxtSd2BEs2izz7CvCdRGifap+m9xVRT/8nnnsnoo17y4vIgRojbFXkBq
KDH3km52EkDgBtKnrvQB4AugzseRJL7QB5IqMHcO9JtBCcDuhOE01e/Xm9w/dBEmrmSxnFK6z3pz
oFjhSui4Whwh7PXU39K78KcRlSJziOoDZjUt8Df7/1V8E8m7Ieodj5oGFRZ062nkwRtQsfWWrcSk
BaYQY0pnx86tSRX2kQUOk91OegvR9jlKq8gdo1lZOs8rnHPwa+XGDoV9WnQUMn0ahpuTVItVbIYX
26/Tw6FeX35dqeF7V39NghjJ3T+DEhS6zpiFd4fOJzX/P1ByQvgLM0WNCru8v2F8NjEvFUdCBBHd
qIc0T+2dqgKQ1VI89ArPCvGEP/hcClcM+HzVvLsgLrUJgOHELAbf2b1CcqV2g/sHYKgvrsLcUA2J
gvQS5k7ip0eVvPVutdLgVWkG25Bw5edRyjBI3n8bs65H0Hfhw2GlgAemQdwnLRj47yFGxrzOuWPh
jwE5fvKNbwFO5M6bMSe4VuZnV3EzMjIw9VNnUsKi80sZ3y6BCMxX6txmV4gVXVUmWTut8Yql2MqT
PANHXcb1YKDcvT0OEYqZKCN1E9hF3r94Atb2tWJiNBD4eeQl7l/dUB7J1J5ObX2XS5FU0gSgPgDo
3z7Pjc9VGiOcaLfRAn1UrD1riPcviIbg4lfXsPgP0sp0dSUKPrRS66cTY9kMAG0qAuxPu2x8QK37
1GcygEGqVm3PpKjmybOkei3oMYgEY1pAbM4j6JG99HI+2jWoHD0QL9uBP6hvNyI2f3w5/0WMVVco
UB/fp9hT7IArb8xvSiMZth/e33duADwlnunrUo7OXSoDQWMCtuIE+MV2fQU2q70bMQ+TCBVZGGh4
nNfczwzfgLkL6Bfy2XLL/9ru/2dJRomgJR+9GQayQHKAEHTR78gnq9+BiPtQiQojKOGoemb95Zwu
LGOPcemKMshReSAytdccLlOkk7yg5EAQC7vDzDKK96yYj5OQRgVjs6/WKOb0S9/JTYk49qSCfhsM
Oe5p0JaecXql/vjIoVMja6y1/RCWuIrT7tidibBwWhLktcSuXMWftpZiLJW0ob+28a/EFzKS6GTa
FXo0b098bige8L4zAHR8XR2cQvBJZjZ0jK+Ywzss6lG9UWn4HCBcPgl3jPJh8hxSDAjooEIJWJYm
zZDEGbO5p0ruuplhC54Q/RiyCjLlmoXaV5Ienw6XfwjqC9fZ1PDN+JThlRTxiPTLVwwoa7knMcvE
zm+PhGqldJGgt7nYfYaZ8vJ93W6ZQTKVKN1M04DJ27yUuYCNw179wDG3cp/juozBqrkDgsgq3WFe
hCUFopJMWBbD493wSsky1q2Eoh4eHScG9aK4/6sdLTjgN+8F7d4+tbzdsd4HePO5gj81WC9AH/U4
QZGSNKBA0PlitJuFyf6mx+9J+4jGSa/XnbnsdlEFjVhM0L1u5LAX42wHQdrE4J+G5WanpAGFpI2Z
GHX2Gh3r7nxhDa+sZYAMvEhxWm+ssW7k0JPVpNE2VQ6ZsI92BI0p97irQTWWC3kdkUdG/PRMZ+XQ
VcP3IrHdgrCAUL3EP2j6ihNjhoydaaXV3ynbns8s1Vfy/zKA1+gWlnbBI3Zbu50R8LOP2Weppaqg
6SWsAdoqtFOLEmD5gZAS/6v34bTlN9wuN8JP+wrMwGcbAhfth88RNwKSRNd1EAK6eF7PjiyFD4L7
OuCkdUuOHFFxyV6s/CPngUInf20H5IwInf7hbphNtfBk/DbD4kDvkXV5zZ2cAg/07M3h1dRxDgdU
XAcPLSVzmlBFkGQgS2by9U/w+m0jt8ixw+XAHFQHVKvxeZKBoyJ0kt1CtdYWicTBpTXKiuYaq8mj
tRZV45A8x/I+dXUONaOQr+EWBxWYTOmNSYyIjPS3QRkQRHHhJ6BcvA/PEx6rZQ4XDQwFJFlu96QH
tOyxBJ/k7qFqvNh3u018OEJOYy/+1N3TcbXJCtQsBI+2QVPbVwDR1mOdUpw7XEtPHr+hdn0eQ6wR
4BVh5BrMaqx8ogUaHsTky5Ohwuk59h60la35JpZbtZAqg3ngmqNp7W6W848eSPFm8S2Vuw1NK854
EPlXStLz89lmAZHfoxJtRs9EX4zq550op3+ms1J//WcaeL8j8kknRmELjO3s9b9SX02i/kH9K+Qv
6xl3b7M8Zh+bR0S8gfAvOJefDh7UllXhyPx/rehJYmuypD36KCMN35azWChv0lfLdVO8S+rkyXAb
X1gY2AlONLMcQAHFmjLajXJPbMrdMoJ/A9DKpFJVlOi3x9b6Tmr0opDo+uKQc4p7xhbP9i71anWF
K8GDrAfCgzLw19CVqoe2Et+OKc4dgIIa2Ws9jFUYfVIIa7lYo8wO9cjzqMsD5UBXgpWEUVy7S3l1
FD+Vdnhicp4+cTd4VASm5VQOiSgxTwhVota+EqI82p1Gzo+0JxiJVS7oh5E9hgzhUs6wPhnE1fPi
XThrCIA+DexKsTjzVk+tScPMMLUV/RLc9+Svb0zmtZ8xamP3Bdz+4q9WbQ/pM3zcnPEXoL27ifg5
y4NS03U7vhY9VG20e9lxQIX5z/QRKJjhTXR+D/5ISgxg+2vNdj1XvCB39t0F/O5OZ1KOwY46FNwq
6u0vaNnYUCmsCzKZDHLqvUp1PKhbat9+FT7aYb0XXfeyJ5I3eY3dHXHqjRkByPjIK+XgZbFo2G2K
kn+o1BuOVHCOFMANdeOLjFJHQwNIBZkPE86++bWY/X4E8s0CTKMWEFELi3yRgRTaEa1QRwHtJXrD
ej1yR42DkJu+42j34p//zD5rLnVdN3itfE/eHn8VDQFA/9c/cP13Y7XWVr9KV8ujKm1+1qhlXLKe
We7iAK3LxBZVQ696cCvrWfXfGXdNndfKBciB6LfadfgWbmbO/p0g6dTZyjNnKPSM5bIfecWKyHfj
nmKiXHXWSau7RFGWsGYUzbVF6mMx1GX6vmi+jYX8IK9zwk0ijU/bvFNf6CECuj/LGnIrzEf8K0ix
nDUZT0ZixSBXL3+9o0qqVbQ/HRaT1JMHqff61gaqpaa01yq9x6NJYwoj83/OS6kQ7e04n9XgUQee
QGcWy4oF4jQZ8aia+XzLVBlYKSKDGjsk5TsKJslHtZ6u3hRGC8V7Gt5bdFtOxxTh2i2UmnmrQa//
zukuzINptjRrliSJEdTJfTFOTy7YOrcEjEZMPMN42P/1mQmJuTl0ATst3Ur0tiI+NCJupZyoti/b
NsTua7ak53eWKJyVyLncBIfeY8tiVAnulTtKYRcn/j2nrvJfR3GLjzXzGvly5DERyF22F3FGcRC6
3FuyNqshJ9YT5qWPTaObPtoz/Htdh3TpP2avXx1xsTkruOBrxlSri2eAaImLDZOQgbdDk2O9k7gE
Br27uV8qagIAJcvof3LpixEuiAm8HVgFjSQ41g66fhjUaG+ojDpUL4RzexXAtOuCSVVUYvqxpeg3
QDKAo6dxV3gYgF7Mrj6InXKgMOlLF4Zo6QRnSh0ggihmGWO9PdiwR//ecFf2EPGJ/46Ry6P109hN
48jaoiZhJdZ7mmRLq1s2h3o/xqH65Cs5dP9xIBfFNtRhk+AWupsEEjcDT9190pcSWBZkoeg7Iq04
yFrDYdkYpp6/l/A2x+tFOh25UrxZwJ3m+p6yBj2xvmnPBQuzRR/ux58b9rsJV7Bw+sx4C/AOGwpZ
MJ7gXazsZSAJi81rWjpdeUbFV2EWz+tX4AfU2AaFY/Ub6tJXNi6dfp+MqZeLVZwYa0y5Nk5/00IO
LDOz0y7LDMPj6a4j/oa7TuRkh2WBdyTnR45q/WglzQzyVC+Ydd0B3uKNmrWLkmXdNA1WoMSiLO3/
CAPyo8P6Hc5xx96tCc6qdEeI64dalRK6f+k47Wfc/fxvYQf0m1nk6xW73IzIMzu31rnjKRamYgAd
4FNExybB4xRRMeiIaNTUZ6XU9Q3Je26kjdUHzRvwvdUP6E028XiAJM2ZteGsahkaXMzz1QJOFVQV
/Lm7BekqFOfpYvfhIgftPbAa8f4zInFm7uRTC9oiMtt8bY67o49xil2DZBA6gjHqHaKl4hWrQKQH
zCKSYTdJ2pBhsW+qzJFMbQcecWdKuFcpR4xcDDU9HT7eL9dGYMAdAl/Jp5ktTIN/cvyfVZmg4iIP
UcMMKitDpunRB0aSei2IFxa0Iw+NIGuhh8Hf09oiK45Y/EJqRebLLq3hPcwFj+ydcL0ivWr7MXMl
U825XLAMXytbgpdkG9gNTX/s23I9cuBDqmJ4nrjNW9Uz+D4+xZHU+OyjkLrWN9IgEcjjpsx7uYhR
ffmQXsv/Doxh4SBz/x5G/f3Uj4uHONe+uw3vhpEnLX/HXfMdM/jTA/oK71EfFM1N+Yk6HfR6jxJP
eeRxbCra9j5UCPViTRwV4D+NmmHTGFSYjuWUPYuEy2HZ2rjj5Tvs8DZkmeIyRojUZ4gmtDiG8EFv
XcPjTpBAWU05RJP53K0V+/HC2YM2RvFPZNJNE/6gPRuV1LtC4Od+Q/cEOZWgXAGLtfPKSUnxk7ow
zMcoQPNnm3NnQKQ4a50ixR2bDFMSeIskCUNWauhFaOF4nwV5yvJOIe1/YI11BX611OfK/6t6/cqq
bXtQjUoagPDbgWWLU2k5S3QDLh0MC4L16nWPVmKeqAKZZ7ibiQged8WGWZGeTmbk8dANuqe0KxEY
e/lubP9M6/TZpSvBV8jwBip0vjAsGs8v/yLI8AU+XqMggfXCEmWjNGFGGXs2brzDyEzfYc3QvkTu
OlrPmV9c2C3e4v8IYLam/CGHB5waLHKFreD66q/zEmiGwPzS0uwRQ1kfzzb8fGpMBsAuFmCSpeN/
UwM0fp5ImlR4jXBi2SuydviQYNYAJV5SUSMLVDXXgZe9rIp5A6+eLeGgwS9MRa7GHPk7tlZ63I5I
QLlZXoIg5yz+pK6JGcxh86zulxT4VPIneGuB5YTFoYYZCd8TEKyuVZc5eCQO0Z7Lw4XIlM4/loix
KTXXBi1EjDKMis2yzfiIK8XJ/AAnIW7ICkWOrFxpzcNIinNrWXfPzVi+vpcam3QEBNJI/QaKEw9v
n3vPfL2u1rcgOEFILNFucPt/OoPdDQnYma5hHEFAr4q2+5m0syNIuCFkRUwiAnjqWhCQhAk1hAFb
O5wb2GXIRAUvvpvCf+dZzW0OPtYWNDHD+TNfuLF2VtN0MuhPK4rkL83fLobwciJfyoIzJLImvV+O
ersp1MS8v2V8UkVsofXVQQKgCEGx3t4hleqMjuJ5suDWVSU6Sc/v2l4/tCObcwCoAVGmNS5DayGV
ZnqZY5mtoj/4BUETIRqTsIuzfXLZO81Ic3+Nv7pb+H8zd4EwpAPN1nWBrjBim/FrHR1DOMGLcoGj
0iB/SWCw/1TRbWIcEG6ldk92haThjxb0F3duO274vXYP5VaiWF5fGIIGdtcd+dhAM9v0WsV4JZmC
lMSuBuC+uam6WJICzxioQkA8uZEx+QZLjjsDziez8qHiMMWQ0B966m8wttT7kCMnM1e+J5O1enSi
xKILL3cYwMHWU1FWjBcZqPM0Qsxd5S7lFlT4MjsW0lri14SP8S6mZjpC7su65SHJztiO9DgEw77l
xi2nJ2ueXPMeWivHjINzKvda1Z7HSPtPs/EdmS3eceQMMDGOO9AoNd1QKe+gu3zm7A3vaeXSsrto
/LDd+VGg4k3zNtsEedniPXiacVW3V84AmzsG0tIvjtOE9qC8vO/rmCUtxnJwogDMVM0+Lu1qUtzD
ZrZGct/ahcEx1nv3E8Z7VUcgON+k1MtLzhyc/gbXuBPLLwGpmG/i8awHfeBKaXhY5X6AMoF+WkRd
4xkKjkftzHtrg+LotLe93eRM818Ql6OF605E6SoeNO/PEsReO33ox7QSBOR9UA5xkiAQCtTZEtXv
Y4gBaLnWlbOAOIUBTQC86Et37AwVQAll5JSMaOLHXFGnDbJL6/W3aWX2YAeJuxjRwo/cj/JTZ7wR
wpq0ch5OebUWBj4RMYzuvnKEhcj0sbNh5GS8CedRCLseTS34P6NNEcwNRu3K9fSdFXYbwBsz7l6V
V24607uukzEWCLyQOoIoazNr/VFVlx3VDATjNKSGSGYt349kd1YPuVATShtb1S2y8NTmgLPA/uj/
1t+SCBfXCBnqZGztbXLCiRdWOHcvW20+Pm38PW0/6/riCMGt1t7huQBpbFnXrd3DesavVm0+l32M
bQSjCkat0J5+vdAf6vrWFQDuI3w8Xps/tq9M4ZQWSVGBFpw3Q0DiiMxA+y7Zd1QhAbTwB3X/XkfD
zwvte2pMgEYXFAx+Nt0wueoVj7VPuEut31bsju4pcuAsXUXjeNCHXyI5sj7EGR1T6+QkBL5s8YA7
DBB3SrU5xGnNOEexQcxnapZkhaZAAkb4777SSxBh05rYMb+o3MzXk/UGYWffpFVnqiQOnMrBGSsw
KjzV4b1BwdXD2uTnhgHhPWmkbB8R/BuLuHBkxy+yuFg7E3th/ZYvLD4oQxIdBWkspKzNNIoqgqLo
TkTvcI/GD1/WLDGZxo4DstnxXYMVhwt09amgwK7grjtJw8zpguvdC8jDCu11ErxP61MDJiJXdVP1
3ytlrgAxP7NtGyN1flHlSxG0SviC8rkRTqKMUo8FsZWZ0zNTFV+/Mryn88f2y7HHku+H3zm5LQ3Z
Oooz1x9HFD0Z/PqSTt/+5IwrLos71b6vL3E9O9AQJ64YqBt62hlgfvAVlJL006Dm3etwHkTwA6K6
omfRF9RM/nCczjT/M61ClAYZrc18pBDb6jYIsG+TgSv+2KYkGEvMt5s9TbFo8zg3QpahVB8LSzk7
K9GRfBl/HG4mZcXa5NerpW9OKwxD/Y2KXmT4DPpM87IU413fmI+MjnpT0sc8VBwM0yZNLFLjxIij
MttDM0DriyvB+cf/HfyU05MGv2iowmMqLMX4FItia1JkcfboQCPONl9a67q+8lLWw7m71QfI6+bG
LRCoVEOmEeyRO0C1sJHR2nmT1OeGZacgVmkPZXT5CHSJGr76Q/WuHSm75qFlkC9kz61jy/2wvONS
3LX0ou8l2Xj4WyrYEbHQ9We3i4JHOaLqGO58X+FGsn8mVUzkITGirYiytTPnaixlffja98wp+cdx
z/eyZ5ANipj/NNqyx7wYH4JeIpGEe1+1dDVQ7RbC8fPaQxGEtCVUoxsHcj3oL++2zyGVyNOyUTWL
eZdpXIJEtafnY6Opas92gY35AkwGlnNYrwhDg/ZmqiVbixcVu3lXmrge9SXtpbh2WoqhqAwxC0wQ
MhCDEJMGvQ8hZB2kmQbRZl6nHYrIvsD2hmkwOAcLE7+JBx7P8cucCI52AjRFCq0ZZntSDLBYjxQQ
66ZTLuYDdKGiSrEstsOCsUZyIUecyUDzuaTZthS2mX0dDt5X70QlYVXDWZBDWzRwS8ZdAYLhUeEm
9GsAUfCoLF4K0k5JdwmY6WJwJhT6epPhpv3FGtFehsn02SHi/lBwZaCVA7I5D4FifeLFp1bxiiqm
FJe3CDZpHZh7fhGaN6PKbvQCwSM7+upzvwjfggQDtVyYaHXDuQXxUd2E8c+z7FKvZW6/yaV6DKeI
J+tnQ/jg3Yx1aBk5GnuufCN0yEfeBqaBEkm75yamjILuVaJ7FTgAfuVigi+WhIqIuyK/KvMRvxZf
bePoqbtEUE0HKzLePvEIVwJzC+XOls+TuliZgDJMMdqpECMU79Of0Q2iz+ZNaCXiG9mXvme928Z3
sSTNP9eSDthsEG82L1SugNsJIKpR+Bg9/fIrl7ye4fICA2aPeQ/XHhPhZI0kVxjQBahPm5uWe2Jf
oYdpuxO/GfEHciKKnlcy9npt1E4H37Od5j28Cov6zoGzFpgKKEdQ8t4Sjh8FxedHgIdah/62Xyvg
wXjCNjrRLVvI+mpuORXr0fi02igl5hoOOsFeBvpTD23awuPn2CHvlBfvIXwtJgowQVgjsW/y2tY0
Nud5wn5Y1aV1bG9cpeZa0+hVzO/TExVe47Vclxx0DkBGzC+FyB/cmyJ9lTERr5kDRjnZExl0s9lG
BJAIUu5KETEs3ezsNgyLK3/3uY8jjfhbhBHTHfLB7MYkeI7E6h+Jz9emUI+lKA3gWk4fce0XwhH2
PVhx0i20ILYX3NCWOdTsXb69pct7apeM98CkJmbfdW2HWdPuPDiXii3VIsH4vHAQ9k7H3bWGlmbR
vWqWSYXqkZ+mXe5PGKIVE4m/R+4hSWQnZ2aekVUMrT6IGAPERC1JtzyCFFw5nO4yCtssml0Y4f1x
QMqLe6vFjkkELESZcSY8NMLyomhA1Or9UdS6ZuIMjf7uivtp2IMWkJFsa+GBVxPjPXY71/VAvssP
RBvu9vVog2hnpQrotAig6AgJuQijQfiVkaW3hyRNbHOLDhuzTm+f6ZN2EsaiVmeLDCGRse+J9LLx
X+GD+ZaD01TPdMM3L3WAAvTvKGrFI9zktIzHCU4TmdqXul7NFrLgAx9zxZZxGjIC9u7LohzmyFuW
m/2LV7I6fIEcGwFAvAXf2GCEhzEixlDXIFadTT845oKmLUCUPrGeWh1G1z4uqkNB3m3ZXVDzM9y1
wwX5JP59hm0zUs2YfZf4ZnRCqyokPAkSh4SbJJdBD4Uh+djOcGk/hmHbr8LTbM2l35bv48URFHGI
Uzt+u7a76E9jo2TaGDP8JGi3A4LCmU4V57ghK0t00IdKfA67i3JQr9KEY+39d7M/xHR1JGrbY2Yr
EPD3k+PT6HZF8dMy3WC8OHyPNQIz1IvwPBpKtLnfp90eL44wc6yo1p1cBxhxcH5D1ZedHKISLdxG
UTheWjVMz/PvsWSx5PZq016NilbTMgFsfsRoGk06kaYZt72opgaAjrUXm02Zy9pli+4D/kc/V2J9
fOoQOwQJVweTvOhSpSaIQzcQ5BFK48qqODCf/XBsF1+Krqp00sw6ZDY2CNIAmJ6UdRPsRGOLfNaZ
07f0jpkDKp1E93iQFNvx5Q+PtCBddkwCdo+8k45nFQwgwg8KJuzvljzAChvaiU3KkfesogdAIZ57
DuuyqVoqaRXl9aQUEXeiQi6MvmCjl2hRbBVXTje3jctGA3ds/X+VQ3UX3f5nlsiwFdd65KVK0Dxz
dh3sCXpyRCO4dMJLfG7FRO9K2BrLofRnIu6YhBaFw3D6JpB4NpeDuXlcza4UFmiFpKVFvwjx4XPK
7Y/OhE0v83Rmi4uAh4p/e965gEF4QIr5G94gxeLCPXYTGgkMSqMYjqIWwvfVnjDjBc5S0pQkEWMz
uznAbdEkfxKeNgw5tYBRFY3qbvVYOYAgnMkVgmKNH/baAe5i4MCvFOaYKHGh1KXdfKMhH+pmCGkE
cX0xk1DSlfrkgavXdkkZT5oqJQg+7YXvQqXyISDA+HusZRAGKSrDYbXtlBqmX1AJ3IZ3zigC/qeW
+ey3B+/FQn5mNKgxdH25lMyzERRTROy7fYLskHd3kHtD5fjvez39stcSIfnysVc5PGdDlpFWtsG5
UiXwo36lJ6GPTnhvYcj9GJaO/F7O7xCrm522OT5Df2JGnuhb1CEULb7eY3QL7UjB4hdBt28t6MwU
ALX4c0DMeedvRIEISZXHMVhPbbJrm5nOOawm3lDuJDAN3j3s82yvwUaigqx0CNfY4oLpSJVVsUwl
Zi5RpqTCM+SOCo6UMNZGyvMK7a4MAVZnhXzjYV9IV4MLxeu/aJB8DGk8Ca1kiSuAGXnWXt+7I7Jy
SGCrvIHA0UZJ+v8tC+YD3Q5hEe0DX39Cph93Qf9jYyXqhknl5kybBM2V2fz1JbQ2dz4gKz8DQ9WM
Ow2Ao7zBO4x21XMm/7oIgOAa4B8BIgez19tRILfkbT4RbLnHPjk8ljFvLBjFFrmeRRU8iwKV3UXj
4N8n32lv6EtjiMEiJG8CAUmHbHDEAfvGwXPau0OrVHZasTjlepL8X46lB0Lb2vAiREtBOcbRL3gH
3cOweoHPAdUnd2PmsAut4M6bX9sNFhCDKlyf4xUdjZkMY/0nPOGqED+t2CShNcvi7dY/gY042Rzy
lbK8J37cSeXpxVqeoVWJO2xGsUkpDdwptB6Ut1WNZ/VkhML0tFJvKqRx6v9Soe13UFToHC7or4oh
Krl1tfnqlPSfUHNg/CmnEefWgopMDtThssy289p7iJr901YX3mxMOM+mK1cUUMuW6WRLg1E13ls8
sCzmhOk6CLpKoYCyJrjCNDFrUtuxN6SZ3TPqQNtn+2XSKsebOys5SEilIwIqI8JVWgXyAl3kaEMd
Lkoa6XEXmqM0jm74ZM55rMH3FIU1gx8FOXbAa0y3U1OgWS6BxOkiVXsOGgSB1RFEaG3MCpw9Ww6U
xF99yJ1b5flh+MTv9ETO6TUbLshecW/FH+OLocqW2ifJO921vKhB+AogV/EXHEGcg258QjRek12u
zcViXI+KEfhw0jxXTbhRAJd+5LJ0QQtYGUNiwunqUT3tAYIx5mTc6maacIeOYnziXEewwcT/+LDm
4WLfFgQZ7Y7qfFvR7SRJrIQS23ZO0UhGDhLEjiknTEPebZBGd27Vhu1p3pJIEHDbtb9+SvveZaec
VHkZfTOZYFq0Y8COznA3wISdY/myZs3Nr8NJXhLfgY36AwogrCYb9tMtlBqbsOlt2jdezy3Uu9MC
xdniq8o6MXlb8wPvMAOfRS8k6J6b/4vBPYZnqYU8CalsAAGOx1r3eUUVnC90fYa4toXnz53iqvYy
QUt9Ci7LpLOITntonFGE89F9518286APrF5FSQ7+xJcn7ql6yGuWOmcVNZQrok744YQtb+ziiCjt
Yb3JHIcrnDfOGEIl1QhSsOrf42lbifx/CkiQKqWfnLgUTuAsAqtnBZXKL4XMiGhLSGru78N2MEf4
C8tDFHlFmGGO+SxM3R6vTufWkmvHuNtKspPHCuSMi7bxVXEYhGKJifibdIpjmoYQm5d05HDLqlWu
y7cB5/JEMacFV5rT/7gkK+2uMTCQc/a4gNzRv02vf3ZJVpC3iZktL1L/XwadH62Nu6gZp3Xes+16
f+QeiBkWb4YLCWb/M5yvZLxGM8oPPtz4oSS9GGP8rz/21azqklwq8fv+8xbGKf+krlyJY/lJSbkr
ZdSJf8KClguzIA0uw7+htvuml+N15w6UpWxD+yGJLJv8kBrl38zT2Lty7ceIA1bApZPuRAQs7h/2
acWkD0l2AAbY29Pla04+XBBzasVclrgsG0LjzsDIhGaeK88CGX9ep58rhnJO6Kiz1A2saClVqd79
D6NwyPyXY7m0SZdLm0hrnZoBkYYICovlCTbO3QcSKARmLq/kdtbebu0YPIJKHwC9gNGX80C4+phi
eK64+cYUpGGiHMk4tx67Umq1MFawchf0aC2yLQ5Ayaj4Vb9rhW9dmhSPDXoKQ44cwzIhnINKwt6+
YCE3EpBIoWX6j/eU2/c2LgdzYtZO6UEalQY3Ah8wDnra4k5XB8E1RtTMQtLqfEbE38251oVsG1/U
ZB24o3/rySUaj6UYplts28dHGJwqbTOajoZoVlxdsrUFlJUv5xr9gQ7Q9URKQ9OXcwMK9RgsmCmQ
QYHlDzauzoXhMma/aUZnqFW4C6mhlSepSeyXI1sA4nLtuSY2rmoM4D7GFyOPx//4asQFp+EOVAUD
8eBL4T25v8xoGBIp0O9I/WHJVuJXIeiDr5zrKoVzHBnHyhJDRquZ/qXLOgUF8GiJS/p4MqVapc37
ED2zVkHVRIxQIBTtS0ccFkE9exs2mp1HAXTYXrXKKEOGkYhqBCXmsTg+0USimwzlHggNcyyoeJVz
eIh1KwzBIJuqjVgGbJ1MSJYZf2S+dlvUA/rd4/NR+6wsdbzCM1R1qff59xxyKgIzNNLPWvrlh+Bg
8qOCJmHesqRvJUoOa6rPh2l1jtqPqlfaPrJ6F1OvHOndYtAIPg8hxXt9JMLrVRNonOyCALYIlgTf
uIbUT2kt0z5A1nyJg3ESCa1GlNEjGk7ptbeRA0sIWPr4WqOgV5gmHEF9hSyO7cIrNQP2bPeK2mvO
S9Px0MD1roozoQh2yO7pF51usXOzaJ/shshLc2QFtx2TGDR8vuEdPJVU9pjLcy36Y1LnfptzsgRW
UmwVspWSCXUeIuXJ7LVGygzqhW+Z8T4GAN7F+a6SlHXT2kBpqiYfL36CXfN06qbw9OXnOKFOml1a
psrzVMqW4fSWo6Wp1VshjeJxI/2XsBBpn75ItSI8Yqt3nsLHLdMfbvN5/Z6CWJIxUlp3Hrmxp7yO
At2XbQYBxBNXrJggTSoBkObvLRyxU+V8DWyJmHpxjUYHOFKoxzeAEKJivsQzZeE0GmZ39mzg5LOJ
QAkLa2tk+Tq/xDzHGFH+6BpcFeQ95U4rzW8ySYvlsL+vc38ERXrDZhi61ER1L0tPmTXCPOetCF+3
lO/wl5zMm4x+diNLs7q9036S47x5lItDPrxrJOtWcBcfKn/mT6nGhQXlTOuRv7DHT/GyQliF/QAb
XaF6GCJOBD6WpeuPQTXELq3yfq0s6BhJVNnw/ATD062BbfH0Ca8IUYq8rS3kAG9vyTDvZGb6Wg7s
ZE8r0TRfbANbwjWhIVicgYHplQW+76fnKD5TbuQdUbTTtGQgAIxAwJUdLsNBdG5I2eCSAdGmW2GI
SccR+4yv45KPE1tqVfX/DmNlGHX8WK6ERptIMnYfwASfhcOuy1PD7ikdh+LgY/tObFpEl/eyyg4H
z9+/Qog4U7cfMAV+xTL4d26KRB3ldHOPR6SrmMBtY60Q7m/Zae9y/D7/LUDv/ZZhuRaexGIqM936
KBm4oS/tgCeE4DDRK7Nwh12HE7GrS6P4DrB4cDNyGN2vrJDxs1Ljyy5NpCRC4FWQY76dZ0yHp2tJ
lOPdlsVspAC/IDh/qmbP9ezfB+5DYraSWXXw0Of/xoxYScBLAUBVzxJJ/GXojUl0EVVUelBTh/cs
5S72I2Nl9Ihh6nyauXMuP8pxdpOFetbJfjeiKHj+M+tyEhraIGQdPdrGhFG4YblI6yZN/APUR6+Y
ecTd9HT7nhufOX35NGQKUt5owsfPFrzKuRzdhjeF3E2qTCqEboFFUNF4b4I2X4+W+GDiGmMAFisa
3bpsQhGnkAwLYrQW92undPBqxk/PeXsovr60MNWagGbOE9/L9vyNgawbdfrfWoynUeBDxftDzq60
xUtI/VlKdrNKwPecMYQ+DdBP1N73TGOqjDy5GfdbeQ/DubQN4b1UF4fK+KHyYFDFoWmSBjeFFJik
frWdc0GK7PXeuzmsO3UT4y01j2EZu0GYSVvk58HDeCi2Xy4n3SWrfsLYqk4/gLU5jCzi8OagxTCY
E4dNhNIIwRmgT/YUY5Bjo7nG5phWXeRMfZekuUlpW4X+2ho8joJvTiudMeH3nMcBuYQUpH9dYkrZ
G5QWfRaspS5+EMMokZ1UgrLxci6MB7ht9ydNsG8b/xIQCkUNacs9oJ4Vq9+SnQeJXQkKmeasxcOG
uqdTZ2SwltFHNAgmPK2BuaQZ/kn9YUPUFagneRXBAPCi9swUXh6R5YcCpToTAN22D4oQKi9hh9YW
XLy+mANmJThwPrnbJp/KvH/9vJs3517AejF3ufGOaPI1ztNGEaNovZTdGGue6JEdiWSOxgy8iJny
O489yFyuA71iUxsgHnjzkGgNyX4ns5lwaR7m4mbmGWaDNlf48vKP3WeiYuQhg6frdfMDxE8hoVez
pg9PsvzhJD5kfV7GVGorkrYLI3LCm5cJYeUl2cbZhamDvI4SOI3eQasZTvGFPICOvK3MjKfkSkR2
HHpKxn26JYMlXKwfa+xaIIoUp6XIK1A8X8B03PX0KCqLD7lEERxe+0whdnblh617y7VWGfipqDs4
s9GykNt2xbb98A7aCAtjJHwDbgpZAqRIIPpgurDuNJYFw+MJrIpsr2QTM7k3r/XccDIUYe/lFAVZ
Pn2zXIihUwYXw3/qPvQClWT+qcnBUP4VW7n0NrHImvG5oBh/b8c0S+2lNX3YIoJrBNzjqebReMUa
lctInMWmpUCwxkX1zSPqRgUCNMqejbM05nTe2nXGKhgqO4qVnk2D9qTwfr62PCBAmC9IGJcmFpFE
nAsFR7kCtWf4FNFLV/6+v2yFJZnMJQl33PTV0iF8EkHaZlQoS/DRDxPEdVA/mprgl3pJOQsxDZpL
iUnbjeJbvukha+1mwrqlODm0bXxCA603Ghb4dh6f3jNMwTX9Z1acjh0MUEL4CkIzpa18FNVEmmlR
PYVaqcCZps+2OhsFFVcJw/Iv7RBhyYoHU7kP22VgxqtgwkdQEDtKz3dDZucsP2bLq7fX4et53dqC
nuGVyceZsrM/wf09051pPtzZCfWBQWWmEs/PuqgWpURHJqqlbUY2p+rSaJ0ECebO6Qqc06/6665Q
WOaWiu71fu0ghEXEYlrE20aAL+0lsWUMYoARQfxKZtZJj8B0S9YHbF7ym+2Kzcsyo5rov5OccMXT
fgA10bD2pjYkCQLuQJYQC29V1x8muoqXxdtNNbH2+lHAR82i29mF7uPN6iYLyEuA+k64qIWHsBd/
yR8FRCoECKGn8x+XKp3T77cCyLAuy8xKu6LOXYPJOp4PYgSYCMDsMzwAeAX/nDzH0/g8LOGDM/uu
5FOapvXd4hRXeti43i3j9ypXcxTMWPcgrgt4Umqe7j0ZxyQgw1V4GsKuBjpyYF4Go7WEV/tecg5w
JDFwoh/TR/cPI6hPDfclkhbu+kVCvMtDiqsGJMPn1e81dAZnAU9/NFRNTDYKtQLlO72b/32l7ZM9
AGJCAfs/92N/KshqdmaGFTy+T/EYZnrUyj/kieAaTeqapiCWOIwsmrWN00t7WHFGyMxiu3zJyToS
XVuUlMH+6384CcW5xndEKmBL8etQTvv36u2vwhpzdzy0Ot+i117Ht4vA5Y6suADfPT/0oWq40MZW
0cN6gkMb1CRZfRz7P6mTbrQb80ZSZICt6TKmehCFJqJFI3FGduoNkRtkDRmuAsOg8NaDl9G+BuWb
zV0sZUYfqZFTi0Xyot4rAbW+nQTQwlHgM+I8ke9gm90ZDNPmYDaxhWZySbLJKztkEn0NaY/99Au6
p9AmimX8RHFcNaASQlWv+dLD2fhtgaSVNhsMqZAiCaGi0SYwx+vHX1580dKAYjEIVbv5BH93tt8g
+OIwyO0mppboN/AcSO76wfWOb2gyutUKiffGYCM6D3lbHZ5EABxldqzbSTAz+b+BYNqTPEDOdMxY
OKaASOYMQvOrVmw2kqg0q5Wau4R7h8j1N2poL4lMRqkdQ6DahPg5SA8gArSURYRIs6YjM6KbCrGQ
HNBFaUIfv01lRH6J/O4jEjkgTYCT7mNpiuvV4s68jZcnEJ3gbbJ3KBSYGSl3f0v8dImOpHj2/hpT
hSHa+CHPWKY55hRxm7pef93P0f/kFhuDHnXuYNwdi5yKMLXTy5G3x+z9Y1R58wQ4Qqlus1Otaol6
ArxdQ+GXjMxgLSDwbCXhIBuhl3o5oGXHJBkeCsg4U4iado46nyA1syEPGT88JdK1EPkvLPPy5UuL
gNe1dlOle1GFYSq1ZgfPaiSZVQBhNd5hv3AlfOESNrjsNXIO8utm/zXqgr+kHtjQNQfKNGiJcXS2
9YhqmW1PA7GCG7IOgl1A6dBVja/7X2CNd5h01wjNSwcSROa4RspJtstRDJXYc9CU/0x8YxyjjKWq
vCVoY5hb5YgHDq+zHE8R8cfECcpgDXDqjwcg4oc1XK88VZbMTk4CvB2ck73CUn1XVh/ApleAalxW
LpR1uDAYDiNg5BtlpE0YH8q7u9AQj2RGO4j+P8ETj850zYEF5CqW08hFinCjuIVYPziUG1uukHYj
DtUWG5K81phRiS/xDO6QovGNDxnNk2GJzlgD6Ojk8covya6LyexlyTMGRHX+Rs4Q5cfw6c43hKby
tL+ypIR0V2g24sAqmwTAhA4ZKSJWyU/VPW6s/pGVHiNmPlX5fbd+vXmAeC4DDJ3guqHnHia2hakt
kwNQQXyGLYliSru71X6OreexzMr3LEkYm5i76gcNQGiQGWlsAdauOpFzTKmCZmyrJRigN49Jgh4/
PC3rh5AVPR92H60mX8PcHyWfV8xkdlY4quPcMqTj1cELaW56QXzD/7sUE/g2RL12ISjuN3vVlgYY
JXsBYd+0JyfBJVUfUZ0DtpoJ0TJkJ0f1hkKdLLmWUUANxeyBWIbl43TU+A+eWp1cPkw8f2hk9O21
XIiVWt/4pH25LpyRVtSJmtDj+w60W8jQdnKBEZlK6SQE6Mxs8orsQtYU7hNVMT+J/BqecMZsYh+c
i7oUmYk8aC37uhrqpd1hbANGGY9tlQykl1CQDfR3ULP436JIhGzSGpcx7P9QmEXryGDlthsiNvUW
lIzzgmMnh8oSoQvHTC7uq6R1mldllJA1adnRqqewR1KTq6rGqSY0skKyQHkQR6pyVvM1uW8Dnee5
TiMPr2T7v119yPkHvvecg8wwuIQORaXs2ssT7zumwpq/CaXdEuCWeETlnzdBxtU5W/cO6s62/NzZ
D4rd+wP0lgVZrdBCvYSZyCwa7acjzHMyD11zLeqTXLtLPws5fHcSIjZsQs9qjE30uQj+uz+OgYYs
w4gQIOcTS2X8VDentx5v7y8B174J+l6xu0N8FXPmLmKiF2XLXaiYZnBzrtoltpGuj+6+2Mvu1VoD
bP+MsKRF9CuryrIv6/OpRoWjOY+4mEcjiFFL+Ky3K7OaNJ6U+grnsOKU0TTXe7ez3s+htMElOucS
vPhHNdswN2jp9qcU8wQ9zmLvlHz0liyJ6igpaGiKQrekSrZ0SRmwlTZoQ7dVpjGbm/P2Mmq3iQVC
GBNOMM+dWhDjKou28Pm3HfJcHPdwtP/egwCUWj2Mp3cZJli40MxSTMPgJgUxhxE0livJC9A7vAKb
07XJJM/wgAPggp1VkXhyuHaSwZ0wBf9Tlcu7g+Plpsx7P52l2i2KJsdScNbkAJ4Vj0rfpOooEq8W
BsaUa7wQITfhvqQS7oL6zJd37LbQjxBX2QaeCKMeB2WAMD7UWoZ093BJalevvkDIz1a7fnFEGsL5
Ml5hriXToBDKOLfcq6YQ+7lbqPdrDciLuI8Lg/hQ0ApRIKd6xxjSM0E844n72LlywMfD9cDsOHIA
aB1nR5e0PJuSSwkARJdbHn5TneIohf2S7C80YCISQU8+tBT90Jbvuv8pleTMb7oZ2CLXxQDOjlaV
i65P7eTrjhkrOkAkxyll2SUUl+/J6wkrGp8WJcSl6VfJcSNP4VHK5bBhQ8GL66C2dMmgAQiYyOay
xvRH52O4qmuSDuLfPBxwLep+7YnMqVW4lY/WZEjNyTIEn5KZO8/xMCE5WOY+ieJ6QoKG53My+eBw
L2BeOxEEYuPREm7mmZwnsoCWzns4RFtvGdi1XdSzL2mz/MrekIIRoHi1ixF3M8w89YJw+2WetTFv
oYVHS9jPa9MZUr6BtepGSYs1DrTzrQHC/U/lCytDFk6t4rMeKLWOU7QA0RzPoLeTxK/svguSzF79
N95kDmmyY647RWzpqIZYUqavW0pIfAFtYmgBTc8NRj8pZP2iMHrePI5cM5az6rkvzyVe+40HNVwT
nEOgrqOCW8qfnHpnomwGoiZXJxqfQjaRgfgTpgQSwk3AbnTqf2FXQi4lzMboD/xmp/FLcWK3xFc8
D0FhFK2nsnILlJyrbnROHTRldlu/DBzzYtNNI6PFIUcB3rcFjFjwfwU3P7kYkgT6WbjIfvNY4fE1
lhS/yYAl0UAZ5dlgdpxE8My9LLeJCVWmcCvqS7UNX637t1zcoZlnp/W4CYP+EZRCer6gkaHqdDt0
uReCb7hyHAe+i54GoFgHf2OrN3wzvJeVB2CJeHFqojwB5uLBZnOEw1tsCX/WmbGpU+YOWhO64W+a
N8sY5K47awMAMg13jK68elQH/Dtqw6mZ5ixnznCs5Em+dlFHt3yWtl2fX5syZ6TCebyUAndRhjL7
3Z9S+tnZZFsPNMXaUR8E4c1je5pjINQTyXueG3BvTMCHcKRxu1iCAl4IC8bhMp4yrVhjx/huKAV+
TAiBX1l6VO6wIn6j8BtyhZxAUKLaZ2M0/S6Iie1CA7garPFJbWKKMftYsb9gfuHB0SSs9ZFSOgJX
BXOai5Ki0nS1cYV2ysqylIPYLACEdB4Ua0kzqpljQy9SmVvajDymj4vMm479RGv3YPFadlVWguen
wLb22uOoJOqWnKLqLv/9VxRwjCcy56Qz8Qmfy3h/Z3tEAMutFJfJJbw5ZJ2Ywpdub9bAnHyiUlNX
zW7XFOUvZThv7rzecyvFwsehLRVSqE6YO+IQ4B0jcEEuP0d2Go+vWqpaQuSGu2lih8BSjmFJTZMc
vJumM+ztjVXWY4yfqFDVqQiaHyESBwNzuvQiSch1jbHGeSrlXnhvhuaAuCLOtxnSNVh+vWUmr53a
1dROfyS+4eVbIl6qsBfJOXXMfbCbxv7fFTMqv0f9Br+S/a0G+z6rf1egb6j5et4f0qUV5ARenfPJ
+weycTTw2dAFor7jmsPUf1BhhIDrK6u/5BpjQ3sjQb13ga9ahkgIYEqJhgzVc77JntT3MKyJnlhH
P3ZWo7KLApRjHh4l3Cpt04xiZrydJqqZWI3UAZbND+vRVBO7Pk/RZxhnVFlEuKxpM/DWfhtfKuGp
Mg1u3+B8aRt1oJf0mLpnsOo28Bw7PNpg16kDgX4lf0s6qPtjiJ34UTcEyeUDvZyl0mnIpA1hN05c
Egd7X2kQdSIFDXR6R5469cX9gL839r2oBjGMQ9gWYrGOMPcD5SUJ3AV5z/FTuTUgaQYwkFYBoMpv
HBhPDkjfAqDYyvQo+FjmccjxVywduCGSx/AD3h1KWdgYIUyhHVUiEls4lfFO6Ed7xiQVLCFUiPAW
0sBhtxFlreRs7zNOr16L4Mn8hvc7e6QiofXtyviKJxVZypLySW5f2HzieXvv6Hx8uGkvi4zPY6ld
ROXEAvwtlgRJiNGPB9z44RuFKVXuX+vmBp0IFWaVMVSPkqZ1r4FRnTGTUYekVBCNxO91VRyIjgI7
YLChtJ4WCeSfuURIjRcyDM1y0kM19eStwnfmMqoCdi9P6e2NYoYvKXHqoIdmtUVm5S5PZmZxbmg7
wHSvS4BNHSfbeVPXKdh5nlqLLr9DEGiylan7zsHrtbgg+/rXQi1xJUlP0zjt374MvuTXGRxn5Pxb
4QGCjvm427/gEEU9sDRIyFPD9km5DZO+DlB4ltjH1isyTylqSwNOqWd2J25FxxXNPtSH81aFZIE5
kTZF1gkvw7Wz/mv7PlCkfc55d6w2up6XCqAJs41jq81cBbs8YkhcfDZ2isZsO4opZowCrJkCl9sv
REMV4Okh0pdQPWPDGpaXXEUR0O1nez7BCLRMsM7qw6n0POEaIqqQLd/6YycQEGZE+GiYrxUpe0Sv
oIUvSUCvJh2oNROxCnyez/2TUV7QArq+SyFR8FF7G1KpjSmzYe6VwITE0QOyVxSG/orGZkGTu+9i
ui95dTxcQy/EHQQrU0C2IHY0zRXpN6oDiD/1KCds884qPL5BVirkvbY7+yCloOn/nN+ib3c6ncCW
T2484HVJYjP5SCvrjM4jXMzRxwQDVWnByT68w1yh5iLD76ZURWalp61tRUwuTUM0hkbX0b1ovWw5
bHSHBCPpGHVCDd8UkyHzEFAHaFX0GePpcMy1UJXP/03+Vz7IwCqI3d4ZMUNPP8IeNsHTDIJuF37i
Af7D7lL0/zkczTrnsudyulA3GcX4o8SazxR4agEuCsw1TDuU6dgZXorUN2W5TraWe07iWCxRGHY+
tlW70usLb2bA8jQs+atiU8PIyRc9LrkXaTKvbgurglejB06SsFVbyGZGY1eicW+cHEl6dTjJITPs
LXzV0AHhGGlQfPAVSajL1MKz9zaLiP0QuPF/83sLASIHCc4xSsR+aLcry3aCGRb+BQPOUTyXQ0BY
E/UWwzhAadtHHL2MWbaVCJ5OYd3Qu6KeAsKyDJjP+YgbAMBQMYzVFHzTJxphdwrVYYLnAWxiCjRH
h0Yeoj8Z5n/krUjjCOU9cUodxQ+9kJQGTHFeRKle51v0VGg22czCqRiW6u8B2byW279DxF+4McX2
CVwrX7JUoA8bzhxDTzdqnkSH2PaGpKghj6ATcX0fNNs0jZd2lKJx5+T5dwYmQf8u5c3uHNkYDdEa
yGO1hLzuHIy1cGCwV8xPiR+mvW7xuG0wYhffj8incGhlncX/IJWLZi1L/cZZRx6oRlQhx1lvFrEl
x3xVSEp1rgIwkSurAsdhDfRxAnwGBOdJ4NsXK2LWu2q/zhODRuSMfdIw+Ot8cYNVr22utZ6G09G9
oNUAxQlaLiYkwPiQB6mNhKZoDrdbFxDie1VJ7gxy2xjj3o2jUkBKqDxUgjuinrJF+vatMvhzhXGB
51PggmXdID3hOg5HQSSOW83o9nG1gSMvjiUkNbgHNw/Qs/97CvtaPkU4FaWcJIrIpt5/PjvW+xRM
Ttv4XedLZXyltJD/+8jwjVgLGoC+i+hDhbt4uvTwySRQK6eX/h7eoYyBRRNjGnS5iX554Gd6xgMK
e13zS8/MYgGYXxcxB6BTlex3yu0jr1FCprcaJY4You+ezYrhIPjz2c7zgl0DYA+DpZny/p4185hj
JNXBNiCuzkO41JPClr6JJYVOjj4fto0X5mJ+nZVPRaSpqEpNFz8lxYqZl50/GnqktvZnj1mPJXHs
w5ZCAIrXCvbfleo0dn7FOTQSHU8hhTr6ydQTFBUuBDDJLNpq1aE/bar5bkepNIS7RagHhTS1eS71
l0XA4GOtpoYo+DULb0PYhUjv0BZ7QAX8YgNyTzQW+/9tZlu5YGAg/NxhIU9EloVb/+E6rsKsQeDN
Fil9YP65J7TaWjaFpv8B8MNFjeoT6TDPzUzl3EZ5WWOHVx1Luzx5lux0hHGE1Rcudfhc2iTjwDuS
Q8MA/ZA7hETqhMiKxoDDP9Qr+VHH5MwcUvM6EOPVS56A9e0mdZNRZeThg6AISh/4VTxeur3F0V/h
bVxcQ1nNxIEXUBapA7JCV+4hc3XwYQIrIABsjh1QbYwPSb3e3jr1X6p66klAyWG9eu8uQsugBKqU
YxCWl/DP4hUTuFsFBn8/n+1+xw43PNU0HCWYXwOLEb0mbC2SOfdzVXtJ5+IEXFOg6m4XDfoJWF03
wxmloNhDrak9ucO/T2QYFkWw85xIFSqAQ8zCJs7LGDCoAKo4dAc93LwXVizmZNRHNJ8TWiQi1xUT
GrPgvhTSiAq3xJaNjAGX9gasKxWytWl5TifaDuz7n5sdcLza5mZZ4JhOV2j/pwaUU/FuMSFL8FeJ
gKdC+BOV3YHBLjlxCks5IwRFQsKfMuvxJ4hewGt2Kl/bgiDbv2RjhtsP7efP9+IckqMgOxqZc7xx
uZBgv4XedMT2cimLpZktRdT4Q8xtFahEeAqqhckGY6xSxhOOztG4zmT2vdKStJ7K5RmOcUJKrmvr
6lx7Kk/lT8Vrr50XEJ2eUontPzE6ZrKDbbpAaw+p1oJGY5pHJ6MFJaqdtSZisJc7fW0z+nG4rrVR
aCyzj4Bo7y+7BD+9pZCxYknlz4YPEoZ1VD/2SUZnqKg7WFrHi6cKv89Ucf/WXccyQTBBKrjMZ3KC
heCaOr7blbknwO1yzi/6WG5t+jR9+CibihscFRar4z79lpy53avT8RuvdYiWymnLALL/RmQ7YCxa
IC62oUu9msRZZeCh14YE/ouxjMq2Q+ZxA/uvFNHC316waVViNs3Oe0DCSy/scw7BBZEZjKX6s52y
wBT8TIvrLRvl2qSXa1prcUstDwEZDiwpCPLoHWE7D88gl/ryU+7jGes8FZCOE/OKBW1u60wMsfQx
tDIO/lU4ZlViG39XU1GKTETJVjlHItJsp6BWBuGp8KY2BbfSX/5L/tqSvRJ8UMEpES+5z7Ovjcwf
UCookakwmHxbUHZg2Twe0rBag0plELz8SI65u5I1JWKNq4tnLEtz1hXaiLosgureLFxuEhsZf9pg
xBNO4iGbUIj/O9f/5YnLKhiUktaX/iCrXuqfIKthAazwf25Tto3r8Dggotik31Y6glH1CCXIYxAI
YT3RYPuutA7DIDIyqOGz7aO+eUqkzTOFPZVvc3XJ9jqQQx+QujL/R7CrmpDJyrHjntw+Byc7Lziq
lm9OGOhtAazAwu0dn8tkp+Bx1fncgQRVJsro60mVM1YKWZVl4pTJgw9rl3RbwuZzLm+btBLIjCAU
y91NAr+L7byuJOZ3NPwQLg8OB3grI3h/D51+oDO8xLiqPzieOmnTbktaqj6/0dVVishbZS+clVmv
BLYpxpW+t3OyEsfIiI5Tg3tLiKGUfHecmlYw5JDkKrzJQA+PqH0VUcDkgyEFZeHLLaGqit+KOsfN
ggI0OCOx7qP5whP+GYan9asD5hScVophCjoRnlFegbGT63QXLCC22kcbIh718Z7EZHHGXw42LJ+g
tUPzfjPkRuIMzZn1zykbNpTujkcleYESjI002qHjNUz8zY3XzV0TB2PrfNbzl211ZxOA7k+9+xPq
ylXf5nB1Ucfg0E062VgKG458kx1ALDTIblES+/QshEzVpGsyvko3YsakD6OML1fZ6LXzcjKTQbS4
e3LSs8geLquJXkpVnQE/i0fEsZeViMYYk4BO2ye12a8Za9Q54EafBSYUfrT4GfGgpdvbSa0eRqm0
SvxA7JEW/3vkji3HMfB1bbottgtg1nvgCPA2SuL2wu9xBov/kAVQCKD5lnTSqwdhb1TonzGiXm5i
3mm2kJjh8UNeTX6yQTY+HLXJFEoylNCQcF8uLjrtzseBxbLc0tYbVEU4UzJB7jjE071p72HQ/zdM
HcZsh8tp79CHJ5kUIkpj5rL1tB7kEVyP+GW1/tXq49lR+5jXr3vcAGQ8Hq5dRv4qi3G5zXBqbV3v
aj84PnfL16S3UdIMNXhqV4BvqlGJFZHR5BsSHrCQa0k1Oc2cc7gajA36KvFnxRGLgN5R4GktFUAz
xqMUZW8Qig6CHHOnjFOTXDrDQrXfl6Ye0KgvCnSubaFxu7EQAcHmZuhtfD25KRqj2/CpqiRMa7Lf
cmxeZ4hT6T7BcyHy6hZot1roFEi/STgUhkjyd2U7VrTPfUkxQZHjM3dvy7+PvHxZKiSlLN25Ca19
f/9jTTsHVetA81KvZlVk5bBFNyNzH0Efdh4mTyditctao+ooM2y9Dy88jnXBji5Mu5mFxvZClwuL
trwC4XIUOjQB3pjKivGGL41xIryaWakmIFZzKjLVewVergAm3RMdrX/1y+MCMxPnYyDBQAy/ZX4W
Yl9bo1C3Cg06LbaIKB4b0QmS0ZGBAQc5QBbSaZpImYRR69T+IZ6+7D0PZTM62Oj8BghVdIX2Spev
cn2Xekh6Z4nJ23zvE6O9kSe+96/9y4kVOqtS61uMdF+l/xzYV8HWeP7c07aEQ9vJVPIE29LM90VL
ew6jgR2baYorn7XKqguzfXUMFgLhNWV4WaX4hvHSHtcZrxsrhY3s7PGXqbYEZzTxTmegTVTsSvLl
ujPBKcX6QUPL9A6Z/kB/lBGiG9Ifj5t0q+oeV1MLpg3Db4RDgteAdhmh6TaY1mw7C8awka/CoTA7
YDKYf3/3VYv7Qb686mvXgTi+0fNkaY6X0PDYHVSHWleiPvYa2fvo3cpMZrmPptQ3df2Zf8m198du
u/+fifUvLRB6Y3yiUOkK5f/l28koRV/aAy4KvxaT9i3jQeS5qGhHVsCn9bU2beghMwE0D6vks8wc
6fEzbgUiaLozSrVMNJ+X7uzrCTXTHtXGfyPFwHygFM96EnqCzyJ33hvvJxWRwhaR+LujLOvSesUN
t4NiC6kRKcpJt/lGynMpKTZKYz8SCKCLM8t8TwQdGvis8oqwFYI+AAi8FB2xKsnn5Ow86CSk9OcH
1IEPo7L5sfqJ8DerVAqcHcGGgefzuVJRoWZYu5L7EGrZ8u9Edn8gSvOmw1HWEsTRgWX/KjtMljJ9
sB43rCQrVuJ93EeNwCr/KxD1dxR23hQ/4hHGLVpZmvOTllMD27c8qAhTIjsE4KpC7QdalgjtZVXy
zcOLkXpvaZA83oQEDGolhzlGnI6WLMz23AjQfvx3TOkM6D4VLWgEA9xLz/1IQktitQgE9i3rH8MN
+CamjG64VUHEzZqnCau7AYv7po48h4wJpEPVFLMKp/jZUFuWQMkkzVO3xGs3ZPAk6xRikXKyS51T
Cs8wkKDhijgUcmakv8VnVi30lcmvGxmGcTj5+7umqQ66nU2opjHA9+ulLW4TbgKkN5Zs5zSXKKFo
yk7Gxp3dCi9SHQ9oiLWRM7mvHszq4bCQVAAFurl4m//C4eRaXppLY81vAAogcsrEU6VQl+fxejjh
riwZCgnC6/kvvCZurZjJbekwjOk33Kpn7ctfZO57v9gkcFOPxDDsyw5//kYMS7u+pOhLsmNRp+BH
+1TBSys2f092ISwc3UkYjzcLm/4sJ0Vzvb/cRtq7gcEEpg1v28setH4pu16Q+xbvHE7dPhTH5G8f
aXF/xR82ONgZbXsb618s3ksT1CGY2L6vng07HyPr6cqKq3di/NP/1/y2AKbRnTHuStwnhDPY4sh5
Z63s8WVjozuFl7L8zW/R5CB8rFKEDRn0I3L0yYpv8tzbzdq3d7rgEE+e7CH7yxgRJC8glge6rMNd
Ji3Kr5H7xwmvuvDWJhbMpvIA6GBsmibSzVSvFKESqQivaQvn8H3KZNdwjTwJ15P4RrPnYknSqkXc
vq9DsKQHIdgV2XYFyiHRoidfwuTyUHIAngGUkD2qM65SmFDfSAKm1xGG+go3wZW/36TyAfLMCl5o
yk1C+vVmMHT8wKe8RpPjxOeyRQQbNQjXkriJQFm1y8XlK+RYbkztI0LAL+Yjp3X+8KDr3dO+lx6k
a2A4WpmLX4DqZoXWvkxeAlx+YMNQl9pL0P+vn1aHNG8Elsmw9dwUzS312kzk1eHNANO6NMQD9LcZ
MG+LR0KKvTX4CZxhadlOIXYoBHfFKrd2Z7ElmXES2FOYgOgq2Ozmkp3WOvqFuBoR4R3RUrLYjc8d
3cvv61bUZ8DXsnnN+B6s9bUhjDE61GVOEpHIPM+PiI8ItQPhFnf9QwH/Y3/hnxqqzytuSo0paFZ1
ku4Y1l50vV5lopxAA3qrKMNNCKz5RDmff6V1i1UWNhvWmKiZdRTIpe3gsV7Vqsj7NAHKAgeJVHCc
9SQX8t5yfck+9bvl4lJuBljtKifCKqMwF+ZST19jnUvxhcDTQoVTCA6m5nbVH/8qHgSlGdxLX51d
vXWMuGxDORCt/RtVyCMRpDYKCXX6GyMsPjy2mRbXksLjiwN38HXAMep2M8WocjIHYkl5l3bm4wl/
A0ymD82QspW1iKjGZyno0usN9IlwkuRjo/YgYkg/KnVcBxMW23zckgI+1kWUkZTUIj6+PgsBgk6c
vMXM5RJ7vhHrfrYzMubC5kYcOHk6ma5NPhbGv08fBhgs0q2rEhfx008IaojSMVOhYykjE35eXcIt
yWSDv4BLYfYtzI99ZLPYLBFjrGEZqBxCIeFbZcJJQV75k3GoC7EfdKm7d2NKU9iGPBDZvCZgvJw1
555LmGU3j7gIbU6pA+uG6TmKNdHN2HMdPQVZrlpEOZBgSudsBdZyQlRoeoYOocD8iq3ORwT3xY3y
tqNUGazJDgHhzgFZxMJGy3JKVL3AKvScXKxwKYJ5iUM7KPJvqlURhpBJZlEq5qYljloq25h98/o1
i/PqaTGStRDyh+svA9fwip2wyLVIm50LZ5lKcNcYvMMdzicqlZUbhEpJ2ywebMiw5WGkcXb2UdoG
bz/Bs6r3u1t3eMgzw8McWdgcm8L5O0ICmnvNhF8SZVB4RxqXT7kRGFY8Ue9dMvXHZudR5hEhO4eJ
HSZL+5abGIHcLU4/xtAyO4MCIhpnwE8QRGS7h39r9gDsHUB29Ttw5CvYxltp0RF6mvcUbINjAPA6
gAcveETH7e1AHMikiXB0rBdRUeOP6RPBAVKCytaJ3Kljjw8p7mWeu6mKkqpH8bu93MEDvvS0rmw3
KUvdK21kNRXL5odo0ZHZxBmoYYPwVEaT4aUDjhxuSBlUfZNCbDEvjzSdHHMWundBGCzAmfiABjDM
3Kwca8T4sbT6bNkmiFUEDj4yBJbndZuzO4BsJcAUSCfwXh9npWzy+/vl6sr3pMcu89pYcllipM05
KDfeldSvKxSwv8ZaaKFjXH0tUn2BXUp/x4t37ecHLRLJ5F7/0f1/bfnbe40qtTOQXaIdypLcFtl9
HW9Ip5uy9a2swkAKN0n9iR+99+L+xtB0AqtWazUbnBteuv/+HpGQXg8TLLJZi1F3d2XXOxFRiCie
ii0keJUayEd0yJQ9MVBcY6qTMrLjzYTSqKO8gwXWP0hHSAhLGW/moEa+ySTvJdhkvW6qKf074aCC
hvpMMyeOQp8xapCYW1B3LkjY+O7PRNOapQrwpSeIplUzkjfSLrTGe5po/pzO9RAK5mzTsAvbx0+D
45MeAsPXgnAK67KNLm6x1YCWF3yUnSNa4GQvqn7rAbIg0AZZi9Y5QGzd1NnUhrok7jUuze6g23BQ
PUxYAJBc7TcON+6JPscRbaZtjBhrMryYRPIqvkB5mH6lRGMbxfKCQ7wRh6vKtYRL3dbviyrfXJ1O
W9HHaPHx4rO0C4coQo8M70u1onlpQBiRC7nKDpod9VxG7bMeFul2nRty1VdJnCuhaf829b03WZUp
JuP1QkP8cPIrabqceUn17ACDZ9xrkv66sfV7k52uy5ibv6uWximN+vYMbdC00BM1Iy2slKLa1hCL
8+axZGiUH8FlQXH4t/4eANYI+FZS6p2o87BFI85mD1KMiN6UbEqQsbddesJ5FG8io5aFQ5hZJCnz
jNzKZvL8s8XCowdjaxBuQ7+bZIFjnRNYjrkcLq7MXltgvnrIAtQYFKw4GGe/vor/SSt9+rdlymzU
1m49ny/bipDzagghyp0Rv5h+12B04+N2DoH6yFqcmJafl+OO4kCCAWKD7XJsiTsTK7Ii1MG7+Gkg
WWmwooAL6bFrr+EEOOaippkBH5gaOOxtBwEXqAlOtItsOeR9wVIBo/5D5tckUEtY3NGSqo9VStwB
mPajCw9RcpMwDMR93Xdsuh8SRkHLd7wxErQz/1dycVsG6hO8q/u8ZNERu6XNFWknQTOwbp49BiLq
l2oeifMv8bzViua/7YoClEY0ec+O2PRLiBfYN9p3Jac3Kj6Ex50DUsPpABz9cQRSXsNrytQkHig2
/H9/3cbCbv8ubERva/Q90Z2W/rrO0fwyAztW9TFkdl7jZleCRH0QVNHhJi9Vw1nktLPjTuIClKeK
Q32IQ6mIKd0Ry2UXZ5LE4AMooiWpKW6PvBVGoQi6w7UCLtf09tGkoKML40OxYa4t3eUHKeg0pfho
uW6VvzgZP0figBnkF7Gmmgty5SjoGCK4616UETSuvF9y9Q9PMoY61yEzn/mAwmMD7QkknzFHHz2l
zh2/Ds3Xb+xqjlvD51gnHDUWZTQYdcxhv9+kjzGB73mtMK9ewOcbFTNtRzOHDJb2drlNJWLu0KqE
KD3q6nEgw2os4A/YNB37Zp3lkjfFFAVDVQGHGA5n2DUXSq8vFIGjRXnGxdB2v6JtILQA5SbdNOsE
jJO53a1/BBgt70E6f7s05sV/nQ6r0GuInppjAM8zUGeFBOlHJLayPk5zohVoeqByLX3OvUVlC7q/
JKSfNEvmeudKI3wSQyJdjR3y20u9Ajbm1JR44cLSrjq4Ygq4eIp7MrFjlqea5WtoOgE7dkh0VjQl
LoBQ09/HjHcSlSMgA3inX7/jeHeFxZvkjHnxdT0z28c+b+Pe3cWERwSTuOWtUe43KWKs7rJ3HA6w
LNDXxrH8aqk6dX5lh3lIaDL7XFDB11gFrdP9NRMBpFzgRBGSelOZ640cpoBBAnoq3ozCjJWhRGXc
ZJLyYhOuz1iC76yR2rzwIwCVIdt5nUmYE/Lbo1EryWrBIO9rwAWdIFcmg1+I+o2vAwkA/2ZZGOSt
xoeUPolOgcwYbN0kuMYvqoNf+1hOFMamXlUcSbAfcsvx51c3696caGoj67Ck8lMX39x7Yh2jc/Ib
ja6sRlUlHfrAw4RI7Dv+B9tlS7tKiRdriad3d3fBJYne7ZlLw8Rm4MNnFXvvr1g9dC90VW2LOygs
rjX9QJzaC7hUBhVKYA/INjLEbEOmVClhPSlC17wDj2KvjNGJJA6EEZx0lETeLdCAwIFKOhK9EOVn
J29h0T24mZjP9cMz7bs4w45Qh9LqYPRkBzYMz0FBUA/iiOfhTouDpdhOAqiEqBO1s+ma872mid0t
99GSCcJ2NtdLFiF1MRwdbAItsNIrvVR8U9RzHcGjuwmAyEPdhEamuQkW2pvRddReiZCZ6Rlinu5P
XrIkMfy6mIrV50IYdvSzg7870N/5nPbZLS/V8A1BzGJH5uuU9VOBrtu471K4IHHYx8HIonekwAhH
cWnBGC5maSZN+dITjS8kc37kUCAYJb9HFJOIRkLnxXf5mq94Yyp+oWJq9mAVMNIwwKPu6gRtKrAq
HGJV/YY2ioDuDpnrKIcm54TmRrA/21wb2RNIWRf8qO4hUS2we/l0v661wx+ke7VnoeCWoRP6MWQX
PXAe05JrlOZNc43jlAYJj+WhNYM4WVrOVd2y51RyfMc9uPQtXR0j+gDaeuAPrH2hzpGsHuX5phF9
HeI+WLAm66PvQQkxKzzfWPZJlWz1ujxGtxnu6pfjkHUKFTzwLENlTsnq2CqsCk2LoizWEDUmrXJY
lOlmxuf1ZWATGbFMIzTGYkC6OZUoohMeMny1fdz8dupV7hpM+WEdy4/6OvWkP4DrbQoETmwObZu6
08x2Ij/2TNmYk44dr04FGeRU73WjGICz2k9YVLxmJRMin6uRXWW7bEyLE8F3MU4xsuoIxfw68+pN
/VUfNp8IdXAk+v9IRLWw+F0SacVWUBpLUPIcj9QsXMZ2IxoMs2lFxyLaYPn7EfLa0wnClqmMV6I/
83kzG2eXlCCfLNj4CvE+Yv71llMvkChOXRJbBqcjxEcRMoWScaHxlvNIXhyyQE4yCIaF4QZTJIj+
2NYcK2q74TssDie4Ddg5Dkt5nCEQAWNMV9kZqRI7oiOKohkLnfqNXHJyK/MZXna/QQNEnGPVI4Nm
ToU38TW1HcB58MjgmF5fcg2KF4sNeF593EHzCPIjf0erx+7uuAI0p11nGODGhgMHAnm8mxb+OZJq
fZKYyD4OZX8oNnmmLMlvgWmrY6goAGSdbg+k0Z84h0xYYJOpmWEyY+sqlG6KL/69jLBziTxKxgZf
5n6yBQu2agV+4aKEVMWk26W++Tk+MirhCD9sdeGk/h1tz+3WEbbTGX37qhLvMbShz1x1kw7O+U8r
mn//Sx+/XRhWEDEc7sHuMmwaVOrk65SaEhU2ckc6Az+zWDPawJ9uRi6zJHC3aCvwk3HhJcDYqd58
s6F1Ll/ROpid9smIoVCwcqEGKniaJUd0AKknv/Rj2aKO4eaMX+YHOdqGShtiaZJiwFyoWyaooMF3
c4w4ki3wL7wPYljM5+ewNuLDE6xBDAPfGS1NBv69m/ZvFKAzIhD2NRORDGontK8t/hnyvMFEhG2V
DvuicqwPlDkn5yyy6eqlEiN9wNwo5h/pJJ5+Viant96AEfFlo7Xw0x+qbaqqI/O/mrWKYnBJgekm
7GOCuJipGQF8q/0dEFyPLFCm8ZN0LsQ0WPAIx7W86oeLuf6OKToWr1TBvlgpnqd8ZAvvfAcwVisO
lvyApMsWIE75xDJTrtwYwkYlaVj0ryMGiWpWlXV5pUCj4J/6Po/ys9zJgKvxIIUuR3sW/PQfCHba
JB8kak3uGNk+52+eedbytEaLt5jC1GePkwcagqfXzBNNOgXbyI3cNNrDiNLI7aXh5ZRkuiI9bdXf
T5bOZfvIa5UvJJPhxFN/mMvvCMpxCl5/CRLl/qOVMEgAvbJoAx5w24gz1q6xdqoSrl2KV/keCabO
gCt0U/DORyFE15qLVuWUGedVNjq4zmPiqrR3r3DiV2soNhIMG+l1LyeD5XsnodQflmrfbDnZPsZe
MRZyYoGIcNT0givl6yAhgmelbOMi8ospRz8A+ytkF3g4V9WfS5MG45w8j57+J01XSZEdzh9myrIm
VDRvzvDxhfwF6HyxwJRlqNK31ogi1wu2LV7vDUbedTLVBcbjcSeuSxXIYCtUk+xdcseuBtFw7InX
rB9+U8Bzv/NTJDKEK+fNRaUgAisyRksHC+iV51pMq1q1ogHc5KDElnijtj09erq0tqbsBmiIAxOt
A9HCzcZ5Fc5qsMgB3SKrepuiIlQ+7ET9mkctNqD7I0pZoCnQ0S+Hl5C7wVCp/S0ktI57KlIYwunG
YV8snV05TRoUeFdvvFh/X/kqXV9wMs1imIGDTMxNnRoE62KD1K2LfyjwRT11VpDTNQw/nu2EEtKW
s7JfotqItfrNaNalmiJG6ok7GAWBqZA/+KC5FwZZiPhami4Cx10nir0lX9NFmx+R47J+9c3uVPXI
FxMd4Y9aQDWzv7zYpGNCz/6ro81F/7y/fQ5IyU2G8d12R8u4y1GcK+DrhD7eI/iZvKjlRDrfwQ6z
KlSNX+57Haq/+qz06QTFv1obm+HtfIjbJ7e/LjEYFPJW0hYRsepsMbP63FObu3KvWQb9A8UFHgju
IqQdlqAt8ZoscMEFs7KmzwFN55aIKyW3p4Jh/Hep0++XLR5GDZndLQONk0ZeD1pN8TaFnkB5qpcI
W80zgTUeL8SNFwHh9Sue7Vkbj6UL0NYK69/nyFO+4DyNysIxXIpxjneqUsGWuw9nEtkVGmboZqSr
SuI/jPMvkIAadEmTYlfogleDETIxDbRw/RpHRihgFdUwj1EATPuFpUFrLstobF5QkWn09NMy5203
djdknnCfuikeCNoI0KW7hDI570pRe8nmGmRhOO5CZMrp/vR9WbrKRcxjVGNkfw2F7I7slp5Tvt+g
DM4YEYha4SMcnu12lCH58FHTFkI1rLdQSC8eyV3xe4qNu/S8ZQxoL6qLXI4QoJ0M53G8eICj4/No
M81WDSdCTA/cYyJhlwnwDbvyCf+nfplIAGphMeKrBRg7jtseh4dmqmfpn9ny2H5ciZ7zVaK8S8bA
fGQWBYSCbObeonxz++LR3XlQVskrRXpbseo34HX/CaybmqEr/d2D1ltzXRvDuLljGOfLXHFlFvMA
28qnOtz2CLNgvbuk+Z9eyMkx/afW2fNAQ0UcOcqh4HuIQ5q6d4zUBdsiRDq82SU1fYMyuiRa5Uz5
+xmDhzFSwB9P0uBYN6L9d56gi3rp+SHfzy7/jw5PsudRuSlzxWHt4mzeqD5CZDfZMFF+86oMyRgr
GFc+gxCgXKTLC0naBS1LVi6KmtMJZZK/CpDmCySeW9S5bPiRwhqHmdVh+moUQJWC7aCOIo87VhaM
eF5dBSZy3QVtlM2nQtBdapz0Pp6eFjOV2YGEz+CUwbzFHZF+QItfmTTQTs1fCC3Iure5t/y731f9
5Hl1mCxQ3qGX7eso+dzN8HH2rcy9OzQ4NmfQWhjCNPj6YBq2fdvdFFlq7WdcZ25L1b1ZZWtgZHDs
PGvPh5ifvy2ew3BijNVgpfbQEiqg6v4lk536tkZzQnK0iYaX0/uKO3J5sUKvBaeYTNoGdPuEhsSD
t2+5qm2NmmzwCa62dEtQlNlq+X0wViewq6x38WJ4sPtFytmCPfUb8r/Qj55kyFSIeqe7wHlEkpQc
E+de0+CKA7vURmp4m9ln8ZA+GjWz+hElO9lKX1N12NPCBpUfZdNTz/7TV4Qj+waA0MvM53P8mjoD
P8AVpofM5IcnNDmYe3vYSu8q4YI1cCMf1ZDMiOhyWTchNnu/qC+NJE4BvVExU9d3FGqom9f6u9E/
HwO+LPGKvAes7hWHxytLDQiyQemVg3+tng87hJTwWrTSBneo2Smb6NTe55pSovAY78M4wLZMZcnx
10wMDMIgLt9aaKjiy6j+PyLuqvU9j0UzANlCijqpqliQ0RB7Rj2+w62spBSID+dabFFVcfIAfHQu
QX10ahTyFHKPWxcK3AcW/AWTpehfiCwX5jZrVuK2H0F+adYpS8OI1OEtDvJQ6JOJsN4ta+WEoxv7
uPdYniOi45mEdGeE6hngWJB3h/crgr7GU02qzNigRb02shbv8GQ5UkGKQvQiPezI6/1KGYp+MImj
mhRZynunNMxBkZWLHa+9pTx6vuAZ9wO7EcyBzyLNwoegOkq1olTy9xW1RoTQo5q5f6NFEqqoFdxi
pZ+bFl8DeJp3+gGfVt/7QtBsmaOHGIWHqIRUmmwrFXvVvsr0090jpCEOKrgx6nmdCnsEkbkGhxLf
3AP5Y2NNF1P+nG/p9LttMqPyp7vfDfUlHEsYBKdDnpRRZqwdzh9ZVR/IzO7DZ0TK61X5FkN7Z7zd
bXMC38k7GTqgCwLJSHWD79+6Zkf0lmdi2J+dJXZ3KMJS47usRvcft4MVqfyc81Fm901khppCeQgg
6FjwI455nz7zLIAyMbusox2R3fLx+L/6VtoAqRSe+b5fPyzRFXKHgzsB+wEfs7QfWGLiznf4VzLV
OkaQyZ46BQlJqNLJI5ZOUQPSBDXajhkbzO18Ofh01viScEFAqfPLguj57Ra+/dJyxcu45SMdtRpI
kexunuaDiuDQTxTlrkvVbYnF8Wqto5Edu7m+1h5BgDmFkcX9zcO5RoMOWIg8CWLs0D8FLu6Zod5y
WQ4oEdEy3zy8EQmSnlXf6o8a3balO/uYplRTdqUv9eY5Q2/IKG8vdLFBcpbbbOwXFvTa9fHejr2G
LsNhGM4T/YOFkD8aYfSO1ClXdH6ucPbXyuA+qUfrVuS2SnJdYLrUM48n6cIra1SVqG2d9Fo2oOll
YJdKdt2xhXsh4c1lNF/HxjT9UhqZWNo7HNW8A7Nfw8UBAAZiBS1VSXUZZ5yTeezp103a+UxWlKk6
UXcCRcv55ToeR66UT2O6W43OQ6yKq7WTDP92Dzra/gXPJj9JezhRT5tWtyEIuVT2nQC5EiCn6992
cXfoHwm4E4AW9hhNCE7Dc0AH76iHtLjPwczFxObmrMfJlmeeDNPFkOnVYGIy73l/Ic4FWyddeMao
xFlHzyyCDmYum+5DBJ8dbp2D8AsYbW5B8K43anAHVX9OSJgvZivKIswrP65PIxuxHFimaFFR+l00
lW7Z0gO+8ATWevY85P1Ptf5nmBXwAMU/O40C5Y69UViHnFdcluM+7aeSZVL7Ll6Gzear6EOVsDkv
nOF+UqgW7Qk0kovbnj3R1GQEBxq17/aab76w+RodjfWoMzjD6Y9w+Q8cBRKeaakd7LSWccsNcV4v
ZFbo4yuFbEmvFTOJ3wWvHkWLrxKX4P7zks2MMMYx9rQFzcL/F7+Z/2kjaA5Vlvq2aeYK/XXhWufp
muia5HizZYoybA64hazfC6SXxpDU0h9vg1PfwowulxAeC+gbZdrafhqMOURV5k31a5qtpK6DSBD3
vAHaKgqs40r82onEWiOri1Msy4p7Y9mP/URe0qRjR+5yBrH83YasNujw3azlMDGLnUhHQMeegfTi
tzw7bz6rryuewS/5AQrxbf7vECdZS1NjZiKa3p9rcXKrCR3P9DT020M22fno+vJGlJDhhRPFiF4i
jc3Cuda8ifUp+F1oSDDhjbXjfif9xL25wmubA179lyL5U7iWMbjtyk4mZyZ+fvguzvIUX+FLrqB8
sEbonzZHxNq5w7DJ/75oqVMuRFbR1XJCIQZJKyI8I/Eah5YS2lXqDfCrtgSCtwAtNK5FEWpJ2WvT
Fvo8KV+ogfaF+iaSIg+WoYgIB/wrI2UqiwEZ8lL+6U+7Ay765vHaWswdqR/UUHhViPosVFm4f/Oh
br8gDCBxqkGG10NFjMlEQUGAENZe7rCry94vxPqnrJE7EfBDEQitFtZFaf57+0kBPUg1mXMRFFbw
ImL9h9Uo7AWCi0isAMD55o8J3s4Zrc7gzJh/QjWu0CHAZGaPFyrQGbxHGAKRr/PS9bz/HHvlb/5U
lGS/6NCn65DxG75c9Jq2aGBeJ/lYoOmtVtRv57tg4PIzcfJJ+0Cu9rzd2PLwi5fR58viRn+1lWEO
FeJE8129MRiyajaZKlWTik+qTji5guhKurNG7UD2KAzLtoh4eb/j0Mch6hKtunHAR9l9arTLT0GK
Yny/e2sJYwiGPM7XCrdz24QURs7J5nu0AEiCL2E8DaCor5OtB0/LPrLvAR9KBZYIlOB4DxMljN56
p5UY9BGekguqVPtV0iPclRRcSQV29lNXDQblCcx1Zslk/FIyeij4GfRvg2S/CA+jpDWWm3p/7BV/
5IXars//1aZKF9MtjS5r3y68xyJ4PNGh3Hijf/Q9R6E8YkgccGRliDZ/dy62HdbMY0xdG5i/s3Zm
+Eh9g63kP0dvKpZZOpB8vETjQmww2YuYeIwPlvrY9uhBOGxciaowuwro1l4amxeGlKB1Ds9D2v1Y
SCmlxgq/fKTSNPCeDi1jB2ri8WUqWrwrt4GjoTBMaYr0D6HlphociYoFXPPm/QX1YFMNDQj+Rdb1
CRjNBWf394JrBMRaSWB+dT0ovOUZJ2GzfCsgzK+2z4Ipxhe0I8NHC8PLh+aSmPurUDEMCg6ILMeE
ftwp3AFrZ+RiCKgcuTSNAmIuBV3KZxnM2+cmmRxdMscPRhbCCUdWWsvtVwtOhVOEj9AVMMcZWjrV
5ao3tSynN2nfc/CGxR0uOB/zFm5Eo6rHGB8PZX/emEaaHOVSzddqxe7iUgzvo681U3zIMnRyZV1I
S+0HpBobvB6NzE2kCuOXQexol0i46kCuqz9N2ZYQFi2g7DQKB1/mvWBJEaZr5EPdmvtJs0JGoCxx
hmAPynFmFDBx683LmX+oC5N5ShzyhAQVh+QqHiNhRpTduD8HrFXJpjQfzN4QxjFzLHTxMXYipBQd
cOtDq8NMLzTnrESgW1Wj4/nWgqjj5i/LOsF3+x/TSpsoH0piyS7q10YWoheTRvr/VCbN+tvSAqQp
+1G/EI3ZT6eZfYtsIkdNOMGblkxvQGMKNorejt2dscBHFfx5gSP2w8PHLrirk3AAbbJlyHKvJ/i5
Cw3eQFvlv7BFDOl1ZTnMp9hUXH25noViSN0XZH+Ytl6J0ayovcC7AV4SpALewPcGqlpWiP4/Beu4
PQl17iGPidTDeU/hN1d+4AWukuOdc3mTsy0R2zaL2wFJsk7fQsM/a9zwheRAvTvlJblNZtRIzeqh
quxXUEqo7DYyvaJ/FHkm3VZYTgJG31WOR13N0+zf+cntWDdQofHBCNcuTt8ZsKwbw+c95UcbFNls
EL6QaB30vIfpqlpgDrusGeIg8DTtROOmu6q4m85gDtICaCtvrgUe2trBWPDPtTNrqoqPVhuD2tWr
hOmJ1SI8u+TaV7enjJYea509DpDIfP14N2gHoDVwi/FjYtNoCNbGP0Q05DuOdi0LfAyoK/0JR2If
at2peQeMH+7Pt6iu0MIHJljrjhWGXRhocXGC2xfNF/Cg5BPxM1qS3MqeiR79trUXOrpCZ5mNKFE6
IKOQmKkSd598pwAcfiECFrDylMGpzGprWUv1B0SBt7mTPBeyx9L3PM49dMhZ8WKS0b9RnvR0k6AQ
8uRKjoj4TfhSl1G9QxSWkh1nxZ4qZ6AAg3gJqmxG03p32sw6p7m4O6p/rHKugQlwpgqYpWOoJP57
JDCR6XagtC/q9WI2OSNAhyDCzL0lvCIkG2bbQ1RY1x1nHgcyhZrgbrneUXdfAhJhiXcu+o73aB/v
eeFMOS+o9/1xLtdD3DaMywgnqwmOjaMc6i68XXtYvToupr/P1VGM8niBV07CFyJ3w8ZnbEgm+mBb
NIyZQ+lx09EiMgeJPBMT4msVVi684Pc/JobZpstbJMcTsdRvoPSsgRQ95g8zf8UjPHj91VHwplAy
4rFdCdRvJ7TOV3XEK0D3aKtq3HOgWYwiVa1axnMKeMPwz9Zp0MIhtjaYM/xP0rhbF3r044bjJmzK
YaUzwelQckjXRhoPIWct2ySUPQBYiXrf4M58q4bvFVQm1TFZCyt3Tnli5SxlrU3kCiC9R4YHqxyL
aIlf0IcvIgkfcY4CCKOmHdmccku1mz1W89ewjBH7x9iQl83ABpmvZqswV425jMTP1uVtlM6FnwGD
jpYmXkWMfPWb5LDAkisTb/27a2gA7kPuvHpraq0zSPzrids1+m5rN2t/TVtxo7Hw1ES/mGYbrPAZ
o73O3dseazRAMoW9dBZC5aw+WvKjCQD/tNoklgOyelC96VG0pcfUtBaJXBBlsq/K7DY8WBzesE9I
3+4hQUEfyyyoe7HRlPhe+80gb1YBDn++VEFpn2z9fG7jKh8jxyXKfT6v0HJ39Ar97VN7LKVxoqHX
U9QNoEDtia5QYaZWiJe0E9KRVBBBou9RhoFtQEWVM+tS+t2G0acbE9UwbzmS0RayxcOroUrU8l8b
Q2o17bcdyrnOiJIOPtsZBns6c+npfYPdpDqzoO23ULGG0VGIfk1rJIVlct2SdbZJ5dBjxAmM/guj
e1r8BfV9xajKIL34ez/SYPETchRvVtgPcOLoeucGr9uiRBoFIqt+MJBuIE2lCmqWfq9Hw8et5H8b
CpJTaCypqfAmVgH6e0EhuMlIfpQ0F2jeQCnPoA+fvVR4Pjm1ybptH0bpWjwYSxKS7CkYVc8UqcXg
nfMQMLRqmzwsbbLdMqBo+fCpoo1HsmRmzHL6JT7ZS07NyvcuRM9fPwWKwYbiyfek9lh4HMSFwr63
tCKK47wTOVjLGsWGnQfChV0b8taxpqg8fbYdGQ0kBfoulhZLRxRIiVFxXyk5gC7JSU/9kVOD0B+o
znn8KMgFRCAtbl5o+2tXIDQ93jUGrJKSCspEDHkX5ShBR2hPJUNUdc4nWWeLq8DUtf6Uppan5ZVP
YPkpitTnSMQUYx0pc1FsllF1jy1S/Rff9PAarCMQVX4diRiFzudSQOf385rHCXstXILQCSFshYzZ
6DAQcHzcs8DKkTLjqgJCgTouGUZzyZWknqLffZNTX2NGyjK0f04scGyUM9xH1reusm5q0bl/GwgM
Nqxe5DTbO1K3qil8JqgZqXJAGBk764tM+iB0eJ3Pi6yrsvJMAtBxFhVzgpU6SOMYPH9DPFxVblo/
eVdWcSQtct6TgsZgmR1WSzQ2zjNjlLrWbsfdBtZlCsx5pXN1XoEMvuo/F6QJrEl4mAc/rSpAUtSW
z26UOW3MUkizn3jVub8lUYxvpNOOTo7I8gLTKHzYmtbP+KUrfe4mfgpOx93i2FaoLsU6PqvCZjsE
heDQmEIyNTaF6VLcwhL+miCSd3HoJ+sRlAY9Q5TcYjx7zDbpLDKJKEJw8uN3cBnjKdMsF9AhHe0M
vb3rv7zrCfEnI8wP7uI6YYvs4TjcvOwnmvlre0bzB7f85Im2JhPk8fWJ4ZalR+bJjlt1ENssLYKs
ocIv8vP6L61+E2l6rLJx7rid/iOT/HLJ3UTh5UmZPF6fE2V3UyjsilkRWWJ1n9vPP//aG/bVBb3A
EF7cfdUYin2FGbJah+u2xCh7h46SKKtwCE4zkze7D5C942WuG3pF60bAhNUP75Qvc2UKG2fGFLA+
QY4s8z43I723196gyHFxdhwHPBhBCOlQ+2EpuosvFyurq4YvZrFtwoc1p4l4gHTCIT7EhzLQexO9
TbKl4IW+CnylWMR757RasDIlcT5+hXxxD060w7zMgtpwHd9+ymJ6D11gWs1WK+aIk76IZ8lU1byk
rDQlfxyzYxXhsy44tgLQdoEBij4dLlbsWIx4TCu6X6UrRmwCspNH8PZ6ne0ACsWm4t6ZFr1wo/Cn
v0llFifs9bO0IU9EhfgtFiRuxz3OvBLLQg+d3nlad9FPhr69SmFlLNZBtrzeApYySM7QLRClnjv8
s7inorQ7+ztd95iWOWmbHbndWD/uSD+BKjoIX8yr7Iy/x0URyYCdozVISlWut/lBWLhd9yjan7ws
6tvTU67VA3u7n4fbOX8b8GvRPT/sd4ynF+K3EHuhIFvznLeTo7Kihc78VKx7np/tnm5s1oDwv2UK
Tbcn4ujSfG0NesbrLi7zilEYwJPt5xuOyv1HTjU2GnAvZ6hp/GTJGikw56B87bMDrJLJ9ZbhZsCx
AFMs22qaJzOKkUIsTO/0p/DcVDjkWVf0L3wGgAsuqtka2Vtilvn4yxfJg03QZlPv0kVBqiKLQw5n
GpZHdbj7w/W8yZu4xJQnyzEgY1qbXEAJW4zwV6j1tqmPiJ5JrwYSdAXHbME8wase6ojnJgvR9ewx
+JbvhXfZjG0dHK0Pf3IEKo90UrjZZ/EevDfu6wKa3IQovcjB3jv9cJ16DyzhwkgJlVuJp97ykD/d
IHqjqBklX+87k2FxbWk4JO9fJvkSkmVZUrMFYc7aFBZyZqRJGn3aGipUAImV7FZFONg/BTFUArj5
5huwgL4MBxua5yrGseQGLxy4ppv3IzOtw8v/Z2Nr94MukSuG6bfDm1eh2qJp1I1RS96lAwBo6RUI
ir742LlXMH3+oXVfPY+fLb4HuNaoi7ld51e56tDlxIgZMB/RH4aqESOXlIfgI3r9mgXlvnflCUO8
rA501NiufGJMCuawfAa9JS068mkCzdHa1p2mly6mWiaDf4od6gL5FWdstVOsUp+RAuGYeIxpg7rE
1dVgTV32ncU9xiRujn5XfaZzdFJjfRJAzb5if0V/3uD3JYNsQPEx10mn1ZhgxsVQcAX0zBLXYlvC
ngfcwufvmVTx85z8gsPnYb3vU02rh0bN53scG+4GThroohWbD4eFD+VQtcmMKDN4t+BJm0ywzIC9
KqMKtYNoz1h8/kUNhdBusKwf9C+nWk6gliZ0dgAq0iUQ9JLqzf9lJ+cBUxOjL6IRtPSd2QQlT0SL
G442n2R7wFzWbO90aT4GPr2Ly4krLnXVgvff/QlUUWshWQHQbsl030dUXSb7N2d7d6baa4Rm+vXv
aIo0M+HhWmxsoJ/gFmTkAdOYCPPFkKKehaVNt9uOGiVTzCIudt7OGRgAAifm6xP+8EyF75t2asAM
uQglft9X1DQaYaO049OX89QT2k4JODEuglaHnz7pDlsZZmwcgFgQhpwYKi78UDGYfqvDwzMEcXhQ
kdA5VoXd8JVp6cLEV2JWguQGPTRF3yVbVF+T8q3/2AAf59cV818R3GCszJfNxy0jaxiol+FR60Bi
Zcao4KZymjuTfbs3sWOBPb4CGT7MbMtFz8mlDeTrXLsJ9uFFloy89huzI6fO9GyE1pdIVz/sck8e
xp2z/S5RbLLW8oYlr0uXIyjFEe+Y88nFYKCeMNjKqGU+iq+hmv/ZXjIny+WD0sdhMJvBlv76H+x5
Yid1PnB0SIJuFI0YM6jZWPy5OI5my+xSs6EZBLEyOK78FjFWcyHyZAwI8ll++QsqsHIxtGrIYRGO
ZM7XZXJUNFVtHdF/+c0T0ae73wRrM9j4AtlMzEGnpxQDfFvOnJLwAGnVN/bjETW4AS1MOUE6CQUb
T4/xh3C9UA2/FiwYT+IezO9ze98SJ5ZLMZHEI7KhSX0+o8HBAetvYDBenTfUNQ0NtNufdxr9YYXS
68CqEpkO38fSF2AeWPAs+BRSZ+gDhSUEspaFz5LD3EOOpR1jR5E6ljRrCfpbwGQ9eBVUKAOZ+yVI
b5+9dLwCDlJxtusG2f59gNI4M5EvPQtW+tH4uhCeQbMraf7Cozv+QcV0J9fakaZZNkcEm1MG1gOR
tKlLQvWIJDR9jL80OqRyjvGEVgVTlA0L+XIJtgedYA/aJtoOG9YLTKw78FQjn/08T+rRR4AQbbbU
kbG6akgKK1GrBPV9zLswaTwf/RfMVimpalywJT7Vm1JI8pQZ21gtPYuEKRt2uBS3CYop2iEFwOE8
NQKqqq5Ea2RrcOMIgUhU3HkdP+u+Es1ZelZf9gs8qYf07EzDLhsy+ber1acNekx1FGGveD+9vMMC
gLJCBCN2rmqgT91+P21Mg6oWdHR1Ei90CLdJC+cZ/jQRCa4FefdXVvtM9dZYzDMiE7kjtxNTlt2t
/ljl4qLifcbgZoAVb8c1s/Aggu1GasIO4FMqCbVpkInYsladIhxGHwRiMkHzrFHZ5fIBmzxJWsBN
GIf0E4hg0Yz8BW0FSDS8PdJPBEgs8Z2z5C0nRWq9Z3bdJuUkWA9g+5TByRh7bQdpqGXQTp/M29h0
nfgrule30r0jChOjdeXHdIU/1D75istG39tPJeaDc4qP2tV90H1iXfTkoUyvlf1d/c5nj83uabzN
13TVw+s+QGOL7+TbTqDXPlxWH+G96vUH2DHBbidBBBOv5dGmzSeXdRPd2Ev4TokPpL6Ay4dPvm5l
Yxri0Oftcu1HWnIwACe5Oattf5qFpsQPSJGNODy3ak9eFGT+qokUz74qI/viPKAZuzczhznmGHnV
XR2ncojNgzByXYVwhD7w2ScKPMhJIkVKPKbgfyY0kEB6TWnYPT6S3ZMzSe4Wfs5b/E3RFgFXSjrl
7rm+rs8glHULbR0s7IaHZrMN8bXZKpNNa3n56f58JnUDS4HZEJ62XAMGsjJvzohxX9uYGfri0y4W
fRlzfozgtVEMpv5Qoaugdu6huOTz+a+6RqVLY9ioRBMqw1UnZGGVoLjVs401uvAAxNVaqybPLG24
lXa2J7PkvzZnaZ/0sIDeRtMWe9SJl5d0oBj7ns/DbYBLhPxFSob8pC+mI2owNlHhjBfbtzBdd4N5
J95/xSAP6f//xR7/0T7Nc2sjwnuM9sOMApMahq/kHLQsNCzg9ROiGROn+I2GCP367sCaz7YNeMQf
7ZXbikBNWgAMYggi/E4JlPRRbRnvDMNdAKV6JlozJjpta4tNSHt3yWMphU0o968MIqVH9apa6yQx
8hcpDBZINfd6lV+3upx2ik8VdfAgh2fI+4QUiWJkEpr+5ALCwF2aq+PnFXGA+WWisiA4S7p24qSx
CLNgmPcc0MAuuOYsk6aJdTWLIY1pYPcjG0NrDBUzFMb0eWq3QZPhW7iSuyxXyAlDUrmk9KjBJmda
mt/wCurrkLZLUni3Dz9+xQosd4yzLJCtb8+jDDOV/X3bqCRpDTYOIiGGGqIac4M05kg3ap4H6sMK
gCaclhXKrIjOCXNjvzya4YHPZZTpMfxG8pZfOV50mg6d6QsL7AcOVFZjhc2Mz8kwQq4SxyGHcNgd
K1FRPMtSiTX2FSXdAeOhQ1s3AdV+BJNzj88iB1KORO0BlaxCoF5n/bo9XMgGY/nPQ30MvBSCn8no
zpPNSmNUKpXLlDbFRyO2BifK8U1YecPAll45Hawo5K59fR3jvC8PDcRjTjzlMrfa5sH6ctMNgpxx
51SGMV33u6siMdyw/9EWcq4HXc0rErZdMuILw2aWjfSYQzqp2Ys8JsqUfyBX+N90zAXwu+6K3n2X
i1BGg6CMyOZmzjU68y7aJghnj+6NrfxWIoQiVtNsAPOhsxk+luSPHHi5ukANy9pvDPb31RtvDweX
i9ZpUWKU3y45YsMYKmi+k/U8vsmRInMRIq7De3nAcDuWTyJ607ggyul5oBfmtchIx9s7RLOoK87+
li+YpGueQoCtAe0nhS6T8ttQhtoJ8evnZZeo8fZU05UyBi7PU/gTze/fudBCu+sr1PifZESUHjS8
wWX47h4h+Njrro4pgoRnQ7FIUFEK40REnBOIIErI5pTZ4uCdB7Phsb1i9zlyoMBeIe3ocu3VTjbB
Pg//21oQNaKJMr7sbZEEz6K/uxjLuuiIL1lzCq92AG7w1X1A0ChtuW8MZgpGbv8rwGQ5DFBPal4I
ascgEQjx4Gu28K4aLqNzlP0TseO+JKs4cvp61PxkiDaFyS+S94phN3xKTLErlNud4Oh+DASWg6Fl
CH4XxNglLs2+K02p9lQr+tpx1iCSVvkXnblooUats1iIHm/GRT2TiTSU6HMf60G41k1DHY1DrxqV
Wl0qyAHXAi38bkY9HkKr4JIfB2LnxSYJSgwPcdw/IQcVJ6eH4MgHbBsvcZ8GQOoBdYV5El32P0VF
sP0nno9kDO+usFgX76t0c2TcPIDCQk+JXCZ8auvCnbSLKLKFHdqehlblQz88nMNSt/BFyRNSiwyx
wiARGig05Vtjq6KjTmU3PU3i80kvXwOeterQxGk0NASoVsbf8265/fdOF5zxH3gGuGpdO/pDTgyj
7zRSXmmAUNuiENSiXM55HeK7ghyhQLBxVuw/YH+A61sgIeZW62tWsowub39V/vdgtppSQYzmZtpG
KxsweAb9TWGGSrmudKYU9jixfRg68NBwKkOcxecTSLEzY1ApIdczWi7m5hQ0R2n9dJKiu1aTGnUF
H3MSmTU608KBsoMj1I535gpI1jGkfHk1obu3w8GTsIpGOxBIqzSpnWmhuA+sI4b2TrTczwcu47Eu
uoi6M5kDbC1BnnWrWB0ZOMVrKlBrwVpL9vrbr0iVh9CmArXtxd8/Hv9MdWHHti3QTFQ+c9UosnCV
kASZufVZGwCNiDu133uOVECtTO0pCu95YwkCK7rfrbepe68ozg5FLIjCH0Mca2VP4EVjGK0d7MIp
s+DvHxBXb7HAzNt70zZmTmwrS0ZfnPHN3gTcLul1AkLDT5pQuYCOYtE5UolG517qZjKj086j1frT
1k5lprVLPLAibNWE0Q8blihpYckuqxQFK72x60b2Rr17nRHz1n1V7CWWsKFst+FeicNJGSavKcR1
BdVEAKTOrPZPSra08gOdyjPYUeNsGQevmV1uJoUNNawAf0ZEauN7MaktXviTwooj74IgCSy6KlIj
4jqbDt87NC+swRe4xXR+LZU5mIBisxxtMxPra1Oy7e0wFc034DUztrqPeWhBLi72vqHZQsxGfZkX
0tqZ9E7gKE0oOWkAsVAGM1oxdB/vgtGo+IX/pZJWZCVeq05Fg6GouQvrXXc71qROdI84fwkySY/O
li7cE7DWcISX3TYOwKJjQyOG9AYiE+MiivowlYmGUifoGgJwV9VhsXhs0rA1i839v0gnkZfNNqRA
sqQ6wTwomlaOh44ZNVxU3tfThnc2b/tVVM99aTEBY1CL82OXII7Hw5FYzExomLu+Bo/4cCmsd+WX
ODT8cvV7f4HqbnW4OSY6o5LHyq1nDkFnLdJHAB9c+6wgcN8qYYtkE3G20YM9vkS6drCpuS9drRZN
qR3wNokmKMjhImQwu/soAvIg9HoG59zzdJhe/WJVWwTFq4b4Jjf0mhG97wvV/SjZXgDJ8Rx5smad
YXd+42aomdEqEpKGKC/Hf8D/p6hAykcrVTp6XqGKQM/xAr4vwwztNHaxYsFV++r2EKH416dJfMXp
GpXcSl334kGGhLuxG1CmSBIxHmq8qscnd7QN6F7Nu8eKvxq1hVMElMnW714U9fSF/Lx6nwWfMOKF
oIhtOmtIO3YpHfYtbsMEzgPXtJ52YZmpkp9jf5EqLlxzT1P3fhbmamUmjuDPHP2avNZku1kHA+jX
DAnOuR/MDbpti/m50ctyGS1nqTvtFti4qIPLirL68sc7u1zg0yaGlJGsUdr+3sxJdZ6wIe9bML1w
ALULNOjSCcfj/LOpB+nbuzznLSQy+u14zAEGYww8l53OAepwJGlVBWci+r5y3Mn9Fd1puovmIzbq
GzXJ3FjZ0Bte6jK3Es5G5J8/vMpvgsTwaKpIPfRgz2ibHn6GcnLJgCExI0N9mEgxjIBnRrcT0Gvn
jzc8qMHAU7zBdzs9mQrHsPQH5GQQoes67GmavVkND8cTsjZ1cJaf0en/MkqejeDe6CFJzD4OTA7W
wdSUstwkXQpswsMK0WG2wjHr4aU7ubDCkDRxEc1+hIZzZNUuLgWtNAQlrCzqsNfumDkl9ySThtjO
jZrMAJY55+qIySMJdaIG2iNp80PvKDHsfi77eddxGNJcEPa+YeOTx+IUnwhtIipWNSUzpgLLXGRd
fh7oZJ353PAFMgap6GtAkvnJQu91hfk0RU+jfwmy2G5Q06bXUC+OVo9n6vJX/8dPCDRu6Z3QnZdv
4Na8hBipdrI4cNNbpu6YZxJp88x+xAkGuTRPKcxKFuwzLwgfzidTydjksvDgngZUWw2EKZHsydjR
X5ao6CKt46UYJisC37bJcJKJ2Aq5xe2Fbh8CwKnzCZiCZfUbESqZh6zh6l2ChuutCZ36dcBOtoJD
6YzOdBHeBd8noHgdXHWt+bN7g01F+224eUj8lBwdlq9LhjtVoVsDJ8NXZynCSZ01IULcGnP6e1v9
CiLRlKZx6tqmZOv6N0h4hNKs6ZM1JQGOuJbd/UM6uZ5vi4wlaeYTuPn6VUAx2wpjJQ0KKe2TQFXx
qZC46+PdwOCNjm7UXsX0II8DiksNyD0NJmTCvz8a/OVLDtNc5AFE7l8tVqV3M3nb0u7LMvGRS3Fm
ejh9xqc0sh6c5uY9ZPbFAn/R/q/+Ba/Mx3lKGA1FFeJkGqZ7dNvztBMcaijM4XbMdBfDleqTuk9c
XHCO82Ju7S+NwDPx46Bli/HyggYweiviMRdQnDMLb/8gyijrybJUwyuCkHcSAgYIo/8+UHYrGcXO
y1qRaQrgFYYRmqvdVt7lS+UkLZGC5K+QyI4tt31ewRj/OHgm1xwkDQTovSkOEVm43B72MRcStRsb
uoOkRNz/XaTRjculkajT4pxZnejU4/Wtoa1p+Pde0VAiAiThmo5gC2ZmzipZuzjhyMtgFGacMWaM
/G/3qUGDDXUQPnRDj9Z90x3Y6V6M8IL5AjNggNJbn/jbMqfFIsBNobZa/f/5099EMvsGx1XyqQLH
eIIZJ9nTGU5umWhA7yWjVSru5Z2TLLSnO5oXlFRgfUJfxdX9WPSfeshZKK26JyNgS30iWC6uxkzp
x1bHITjpTCmJuTI30zz9yy3Cjmy0xuZKAdyLpQduPpXQ49j6odLBrCd0CSxNchSw5boC5aRtFq7l
DtGSFzRFzg90wf//uUvKRA8aVQLThKKyqM354uA2pfef2QCkFyhyx2hBikwP7SmJiblsj2YntgwH
XsKuUsh+dIKeEPmDnhK7NetOa2NLHjKQI7KiDuS5IwHEXw/7wSoJzpZQiX4x3bnXUHdZ4fxwd4Mh
vHFUOWYHdLWkMdaqLL6r/TpFkXeFjvvAW9GiJnc7Bml37A5KR2xIoeWZtyX2EsB51GwhtccOuqEg
LbfMjA106/apRBoBgMAfyqEESdWGyTj1a1l8QCBapc4ch6xRhRSFXpSVGgTZ6FG5GnmFK8Vley8l
w/1R3LkqMM02N+gq+RR80bdixTbGvZUmOP4VhOZqRAQtytY5QaEyJf5lDYcWKqFtKx8zpuNiMpBR
R0lUF/pYZk1pnf0mVX0zL7XYbgRJkKFYFfC9yMmhPfpSEssQfmucMPN0+QyaRCNWmsBofB537CAc
nIyx4chk40j59ZMYGFXEKtTZdcxjHrWbdZFENEsFSsvX30LD+8bpCs5tjufsKix8nS+hJpYZZ6T4
r0i8qGIEhYE9coe7U3QrvhtOGmaZ02vZKXzLtoy3DP5kyAf8SVdfhMQZR8AEXBTqusCihv49YThR
CaqhRYatxXPIy8l3vnEGW7in+e7pzDTVMzIvyt5r2FAIrOiJ7uiJBfkVVD4ecDHXyFSGUJPYnUzI
IWGi8vRQqy7bItHm37FATR+noyj7UgK55jXvHKtiT7rx2FGBdlvN0HSEpFWnOCMadu0Bf9AQDttE
8VhQG9j0CGpeGIq9rPzscY9bg77CvzCdWXQMsvyqyxc2VT22ogdNEbtjTq++A8ZebUxyyQFmseuD
5eiMULMFsq0S3UjhDQ2Jl98hrgDsRAJ/8lXLXvlXlKo4glmQgsFnj+iLCa+6iYlLqf9H1svEEZVi
n4D0eLuWdJJ/88tHoxqgG99ETjDd5dhyeEF+0kCHsjLA0FZ/vwSNC0VfpGOJ/IX+EmdB2Q8kSny8
IKyA3M44yM77JiE8DfrfYOQcNPam+OG2qlnD8VNE/NXek5oWPi7vKJ7ba8VswjwzZGagIehT3XDc
P8WziONDvihmNvlxcMmrFwtbBrrEF/SWBnHLoKxu4W94p26dk6tCRkEXRm3wxR6Dz9GS7lhNgyiB
MdZxBmskd18ZhEgNRUncjQyZtoQP2veoicABBfrL24gYQnY1E8NxGBjvT50FgIqtQBESkZP5Nu3J
El6KZKr4A0X+JvGokc4ZUDK9OeEbhMdipLFQ+T9SNgVyiplhvycA5kzCXQfmX/sDHh7oHycSEJ/J
wPM392+1L2bNlPEiUeeUqs+yuOs7xkko8A8JugmKfAEptaFG/WvgiV0GQI+2kr602jHJzwii0wPj
dhkbXveYtHMwMFEtf5jC+lgvNd+nM2htoh0NlV+4nR0108e9SG6d8UWC6nj95as1vhjoH5zuwmzG
wOINBp9vqlfqi4taiRxEwYESP8Km07+mlq2h0rKTRCkFQAqEN44uUrmpohK/VKBocw6LuDHfHtlj
8oI6eBkymmxPHP1O+o9RbPsj3sz45k1VGIpzSrN9EpmWIJ+R3LpmjQmZuuzCLYGa4/z3JpWqwaQY
IeXHTR9dQ5CyczfUSTH6FjsluZLFPjL+Z4k0rbBAtZOX323oK5qdBA3pbQAmu4HUZfwk8uICENG8
v3QjBaK8ulZsueYesVXNofKRrmc7lQDQEjp8NUN8UUE/K0dbw2MrCeVECtjkLCprkhw+YkBAMCsj
H6bpDQ29rP4mDk2PlXMhgFfkdRVHLKHlAXEAT1T714lRrRpE5FzAV+ks7pGROreLMLye8W6Ki9dS
CiQShHUEZViW9jEqed2E976TV2AmVwj27X5hNcu0KvXKUM577y2MLPvET7KDIDo9LT4EWCMQ3j+Q
5yA2PH0P4R09CFe86j1GH7Bea1lB4tdEwSSC67lW0RCRDeHHzgz3vihIFLBIXGZ/h9GK9tknYcNq
2nmKUy1M8ypRwVsszJPSNlgE8S6cqWWOd+cTlzigFC3P7foZRottj8UN3cG5xini7sc1tFigus5m
6ZBCHQ1PIUYBh573BFm64cxiDobkjFSHRYSd/aVtYFq8+ift/02t5/xqmMTbeQBVQQB4zpXX1vbl
Wv1LsO7iw9pKd0P8h3eIsD95xODWumFaomWZ1HZR0F2AXYo6gcnTw1e2jArhDOLGZS5A+AwdpV24
8SaiFdoNTLoCb/rR+22oPVaCOfheF+ct1ZslJtQXDGbq/WmGnsMjwuEBU3M/cY3NbU1a2kZ1+5e7
8IqOzxIrbP7zaG6e4vATXTiNjxNBE6tb12SsZYRBMFw4wlCDapC8xyc14eBRddDU5zHizi10rDZ/
O2CErisAPrDtZls9/T4epCjgSogaH10rsYGvzPC7qj4msJTVskRH3N0hPdP53/lYNdiqRNN5pJVq
8nQXtIcwMXVIE3HtG+hcQhWD6EKX+MB7xR35nprB9ZII4keuE6EJasGpniQZrhucT0ofU8CNIVul
5Fe3pfRjV9lSEk8Q+CpP1bampTWLhs0+E2w2RCDn6zi/Ho4q5ZtTXDPbs1K2h8sCeF3XhEWhgxV0
3WMXI/puArICXNUiu67tb1mt7Jtbhl4f+d/yXfubvxKAu6he97V9WE9tMmUrFuAhonSMe60DU45o
94O0lh3LnMPQ2oRI6nTfLqkuEzNBa24swddeZOSjzfcuGK38f+9FzkxNlJeK4Cw6kSUUl3dMfPgO
Mz+IEG76qPLfT2v1YWsL276n3QgbjLjPDMJytvr3udfUotzHbxE6XtAOS584TcNA2FY4yZotAuKt
PnJceVHfX+3S0FlO7QJVkIUNs/r+dm4coKMdIvcgYE0dwpbilGODBQ4A3G8AdTL/CeLa0e6mVDWj
a/Dor5zYJJ3OSsTTR3z8xJ9Tm9xrhYYuyoMePkqTBhxR3yMyIixzHeZ9RB9TbwsRzSE1aTL+TUNn
Fg7EsGD7oyTyw1OcYm+N0Rp04qQ5OGTTrD6THkV3DWtImaqPdWyMeLKnl+esRtCh069RaFFdIciN
YruEE2Z+Jcjhiu3BJ2plJkDgRl615GuEmWcRP5rwLp3ZhPvgDHtd2USUELlUPZ+zwcJKixJ3xlMp
NoUExxux7R09fwganhzCZ6N26n3bxdHfxEyCuooTqeg+iu8sH5frUB0LUveOs24kQE/1Rbx62fjj
yeo9fSrwxL1+/xi4RCLhkvoVwhee8d5vK/VAPjfyQv9mVU+MhDeEZdHAnAz6wfaArE2XlOyetPkK
ofVavGeynpldGCdzJjNaXzMZ2rVMrkt/ICrYjpNCI/KEnFboCbOdpiOiVe6hUBd3nfkAN1iqfPcd
AJCbqCwm2r2wQ40/4FElcJx4UHGdAqn3gwsnMbdhv3XOuD7IT4Yao1BQC/H9ev8OsWdflrQODmjd
eKzs0gP9kwPvdZAIsMNNmgEkdzLUWC6LuP42st76Cy5EOtrQJJOuyNP3fbJTMuSvLHhf8RXivEtS
bXbSpBfpkZJiTSsfHQHU2yhyPEUxCg0twkU+MRQ7YEZr/I1CVFbwm3t0dwXAB7Xznt8JVh65J4Ud
2dKFF/u+jeCQ7ij38W2jezDaM32ss8plTzvafM4yZUzfF83KgCUhnl7CbuSgH4nB3Ai7p0YMTIPi
FoSdzDbjixvO7n3zwKOY7C9y+TCib3cdyLtjLqSlbTJ8bUHMXwUaW7H8vxedFJJQ6dPfkYerFuEy
N8Chw2wLO0/camY0L+fCJtfi7jUmRTFLxJ6E03AD/GV8/X8ADEurTAZtGuaGbGHLjHN3rML2qQjv
ghrFRC38JceXC9gcFKmuQZlbUhR2LLZTiYcU6yhjW5HiexEBtZZdtZV4L/4q/M9DlIv0kA3JMmaC
zaWWzMQNEkySajhDzT+a4xCdalnuU48lHlY/Td0OaSiwWgD4QEEdBgkpsQ/ouevn4FVq7xQhXkTD
gfM7lqYg3pL8CMT7HCJnVIrnueD/8fK7OF8IWiSol2h3/MFfhaJ9CclYTzbLbi7WshJMtGe494KX
0lsRJNIkOOKauzB3gMJw05adQEHUAai1gUHEixtSlFdWI61k2WRlysaDTlsQQCJobBtr9AtWXo8Q
QE2hG4bpYpA6NozrA5VVWRWbKWQZy2vpN6rPfmMG6GvcI6PW1Roda/LDBHVQJe7q7m0NGJ+xvncL
/nM7IseSNGqdWd4MYGmdRe3R+K5E/xbutscLsH3veh2IEBZUDZv8vVAAT0gP3bFO1afJs2HGB2O2
FqSV/xNf2vRhXfHIqeqqXpqHm2Oy88fudr3KY5emJhdRvJyi1BHm1MMZO6CHq++Vsplhz64feUms
jznNbeifyi9hTEaD46H43xXPcF6Kszw29ka9nAwIib2s2GVXxoO2CKlx/UuTQHbFKULEvpeVOiXq
FqePH5GKSQEOwCllq928pjogL6f+2K7Vw/Icr6hr5VA1CexTbcdDZEMo8eHVjzeHPERY8zyywbAN
zSy3ug/8nhtT3jAwa0BfiHvNMpbIE9BHsArxJsV+OGVIApVwccxW086F2l3gKkrUppxDhtm4NXOv
d7N0j1fI2vpZ9kpSBEvmraYShokkaUS8gA5Pv984wuQv9IxRhSzev7eamA4vpdII+Nu9pvQ9+jnL
dEpE/Dq65gc1PTlnmao3kth7TEAiNGNI+kTeS2jfOQQ8bOy9HOQfRPXIAexpGCWZ8nQwsXnXx0k8
um6rKUenu6sHPGX0mqjoBTAaB9yTHRju9TlRqTPrbxqQx55qbN3JIT4QXbmIXw814ykTV5jJZQnz
4uXzozFE8Ag5+DdUnKJTWH0XZa3cYCNV36Fan55wTfNDt4FS4ujc0ecEPvQhgZJOtjhzHGlAc6zD
JQkaDeYmo4GPI3Qgjr7T3wUGMdT0JCOVjUjEZQhaJkfA40XY3kti/lvfNo4tTbHyfa7jVUIveESv
1uO2C+djtOa0nw1BmA0XqGR89UqO6ThwrzmE8IMK6lCl2CPQ26vBXFDBFIdusA8jPtOQc2kqMMAr
02U0MZOW9s7SS3gz3etufMomGPgoJBThMDLr1aCR9N/zqLUHrVfO937H5RzX4RIzSEoRlCL5Uiwa
bTZ/6vQnyL2qJlwe/ZANGvaHm15ZV3+n+qpWUjc1ZfR9JylJdkc+gNuceqxeWQSwFoehgmXeHfya
s2LQHC2rPISDm+0dAfDpaL/+PafS6NIiZxWwAXNB0ve4K2qQTeUuocJ+nWj7ejPXXHNlYIcjAiCd
2GBUyyNgmmByOj9xNd+YbY6JLMpqRUgLtxOtJOYBZJouI8JtvUlrjTRQJ3VhKLbtbtuMK/BqgKKx
U8422xoiQy+ErvuyM0j+7R6p1uTiBGCLUlbWDz0+MhmZQLSbGsGaoPfJkcyjebgSmVVtPdhp1Sqr
564FqoU/zi1Vb1dMdxcwatS/Xc6ePVjadPxzS1cyrICRE+A33dElTrLMBo+P5B3lZldDHPnu93hF
bUHWXk+yWdu2S3y9hh3fbcXENq/+iqlhFzBb/Hgn+OQqry8EcFA/kRvBYEIWpFBCZn0SgsubpYht
9NQruRU5VE/is7zidmZhtHcrzPHEIocEzpZOIHDH5Oyg+YH+DoVtBggYcmsxhcLw5Ekgkz0oujls
xPogRuhg46foZzxon0mcGtUAr6JF7RAV7TCCkHsZY3R91YDp/2kYMte+J9gvb95UePgh4Y0YD/9y
FKqrzcGN05vjC8UC2N7ERsyYABvq9MdARd+V5zcv+NQSzIqJS8b9NEcllKpzMrduzV/rP1XNDSUH
gvTiNiiMex500dMMPN7hHej/5pzMbRAzKI2MbEkx9TWMvncPnkC9pn+w2Xh3EpVQhrPeI1FPa6lZ
OXofp2v9YH/v1AaoFvfSar0Ur9YmA93fD/H2speX4coXYzjfnS7cqWu8waZa98wrTRHE0P8tWgVn
XdowXVx3KunI2ezHa09SAaGYD9DpL7EovXEej/g3p+JAxDsW0F1YGSQfBHysf3T73WEosjilpK+w
4P+7+LGdAqchTqw9tsd9KHPdibliG24+WA6eDdjwB5wFfrWCrdQ/YyepGLnuAKVgtGC7BJMcyQ4k
Vut8AH47yo7xi6qwGuXrv6jppg2HxldhsHVwaJGjFbBptDUxZSXHYn5/1oEAFWqYbe9TVX2DSVsX
16SuUCTA3cmRMqD1nVpvPggNHhQeGrQwKPzyIejOe0505xutT6aIM7N/Ldso2K6p5zJJqnTwwHqq
qtzWAWO+Pl3B7dYajNDMJyEIxnrHue/+OcnaC7RYC+9NW3WuGKJM/S5qpU+62mBwuWdjqIMsk79x
PNi+JaXy4CDLk8n2Gj/mNYA+Yy14vrNgjvb3QJMe4Gco14wGFS9YjLBWf2VhvD6HAaXLeF/BX/uJ
r2NGAWX6j6iefjfkFZUErGzWyDxrKahAceeRQEndDc+MJ0uHYioj288umuO8N9XHAsg0u9acueY6
0u46ei6JvjGbRaJZihYObvHmkjfnidOb+NX5qLTjksnFbO1qBIuHHd9Xoctd0OHkj5DjGDL6VgEa
kfldO9XnxUKKfOhQNeLE86XaVrrOokA7hiLvcU/ywPqyJVKBe5i48RltUhcyUVNErXNbjJAhXhMg
UxGkWtHiO67E8YGY+M0ARbPoX+CNQlEhL9jrQOv+tKbvcZuSuYy74uEQhsbauA4oJMBGajPe/9wg
Yoq5V9Udmwo97ScS3q3EYVWTBSMJeIoT5Rx7MHvfLZMabCJU4ItpDKJZo+t1jnmwmBEC3EK2Kd0H
75Kwzvlsydw8Cv5Ed1LxW9nGNSrlG+KSkwF5sxSKGD7kCV8MX/tLJRSWmMA8/4/wuf2Ajlh6uW+T
EnppFs2kF+36MA1Zk3WVDLI++FgXvdf4w7lrGZN3rZ+2uc+ULL0jDCCjPoIYOTNcGwQ5PD3hEoqS
sG23xX1hZdsFWA1xgQrsAnHyBnCLsRonsAtfhVqAti5UcFtl8LkSLg0IOUn1dj2PjuldHkYFVyP/
RCC8Dtp2S19n+HBhTT1ZotxvtDL5QZhVeb+O1jhEPTZJdxEvuu0+gxj6nQjuwSY96FKuKGcl3r4+
pe1eSWF4+B76im3QwZqwM5ZbNbKZ63HLZFW25I3ewUcWZIIsoVpXb56dkLfSIuy1A5CuaPlO3kJ0
IMVpZRXWhf62jCbF0aumFvdj9ekgIf57Gv2DVBFzkguiYLyeiMt6tmWxOtaMAlgvxflvMvNQZSdX
r+lqWENs3PdByZjM4g7OQJzSWqGxyBuakWjACciPxSfso5HbRV4MnhIECbBIybUhU9tS5X8KkgxH
vB9Mndo1mGbTQBcosGGttcTSEmr0PYQQinLTBATTvELr6wIN5bydeJTCsbzERLFk01nJ7J+ZLHax
/xYR5fDL9jUcE6O0QHbRJqyasak8HWVH1bEJRkks++sCYlatIOUimzlDv9oR8nuQzAshHmZY/Mu5
cN19A8zl9JXqPWWStBHOBT8/V/6Mf8R+uGYycRu/BcSJ1YvlVm5jhU2QmHoeTSRzVCxXVW12okDK
L9O/ARp6eV9v3MIEujenVEMFWVbWNAzel6hLixS9wr/Hrzho1y1+XP0FO2qLa0UJXFERQLKEVKug
CVPYi+dg9PEHSLzhiIQ6aMmoEMtNlyImMtJfzFCQjpwxPSO8RPQeli1b3XtBPomvIR/yttjivKPw
WQMmmoCZbra9Nv58v1b2NvG45dxOA4sSI6mcnIkFeZ5V6nduACYTeTVk8Q8++R9YfX9iyOngIv4p
pYMLlxVevq6qkdRe2yYSo6Ch5qL8oxFn/DdAq63sYzRtINPM6pdHneFSmSl08hcmk6+cq+GiDIfE
UL3flcOELfXbkPtmGbSRm0aJUpQ/Mcg93Epy0cGC8YrzS/mZTNwAqnrWCc+yA1F1PlVLngquxvkw
TX/KoeBw/oEv+IHbI4Z6QrBLAO1EZyA/WPvPdtaHneKIhH9Wa5Ew5O60d/ZvigNQHk7oUvTooCeH
O4IovDQi11gYlDwZEBlCjqTZ7o4p3ixgCUx9yKRmz/42RP+qfbJToLxHiZMCjm/yPTlJwg2SoEvX
4IhIUEZ6Zqi/uR8xYZ3DOgsQdV0r0w6EOWmXKFqUeYTS9P2xVnmWuVrPRheKdj/ajO1hwCoun+dj
wc9XpfiO59FIeqCItWH6dSQp2U/4OI28vjtzBcTTzAsa6rtgBjGIDPBt/jHAIuLhz91KM773bwBN
H6A3NIml0Vejp2S+McwUX1AUdez6WuyfMAjqPNo3A/ZZnfS4LaOvgVPbUgTSceW7UZZWjYOImpI7
YkwzJd1fq4qFYRfIxUoqqhzjFZtUe+qAXRAKVdOtUYMpVEK1KTN8GGWzk9DUggc1BNWkLLca+EFn
AJMb4sMtOj5E9hEpYcNhyPB8JNDtYWwYwRCZDyIDN56lcZH2qS5/hiLfzOkbln9+Xjviy2MZcUEE
bxLMY4V5rEIBOTXzQuDYGpM9Cd/NM/uaiJawG4RG6XID5zZWMNfF0V6DlzVGSBEyL2XAe8V+N5Qj
CVBmEBMpa0aRFZROiDvJ9GGtsLLle0yQGHYOgAB7xTpUTol9mN5FmCuFA1xvjCxuDA8/zSQ4qpC0
8UZhrvVw+3RL6JPvAC/K91b+d/x1C3/4/W0Hpyx4gvXXwuG3dVYpvcfl4HPYgFI9VJFUyTQelZ+m
chMNPIhZP9DUjg4X4f7zicmFepGktd4v8R8kfVG4BKtYKZY8kXXZ6IHrRUpIvckiG6TZvz5ps6Cg
CbI4HJ+RytB+eurG+CMmx6ujjyxqY7UnjktbGhyIkCoBKtsdWbsxO7xcZrqSWV6P8shMUeg1o1u5
yt2OLT9ATj56XXZAuFlyBdhdEywOc7i22qeRWH0fuR7lvaCiPPtjW8B0LTWM2rhbaqWT0azVWrth
r+mlgyF4b8XRW+qRLHfD48uOIAOJ7eYzRPCigzgOGZqUIhLjIu20xGqNF0ldyBdQCBbilSu5Pv7a
+x8Dk/QeavJ4Hd+1pkMuAtTZ7Nmx+9gVqGIEqypZlF1gF8Q6ghRNTuNNG4OFeMKKx3SUjcQBlxT9
3Xz7QzrPiAJePH3ZBHhCRfa/JqKdvj4S9U+5x0CXrwZ/BKCF+SF94P9cW/804xPcJB80SoLYhLw6
MUGmpddkQeX9mHKDx1HrZeAnpd5Z+dezCU0hHw/Wc+GLekyAry76iUxj2514ewbjQkWUGDR1QWIP
yvszIxddcNTrKIWxcwO/RxaqmfrXZuhM0HGGRCLEa1aK9lA07Ys0GdSV0O/N1tkLTrMzS1+ikTv1
kqT+5wjqwFNvaG5OPwhiFVUYAXm0e7UA5Biquy/kjkgwQAtFg/wCXIEGrRGEmkRqJ5UaFLGGVXDm
2AioURdoX1lOksYG+ubg6Mh2qcazEkHD7HSvMUb3+jthAAG+g9cHcfVwS0fYZ1nvPx84N00ajAWR
h/1zuZ9OmqhGF5gMysDqGHXSdWYqiZ7GYEZ9fZc1Soq0m7S1CEc1iSuWOHjeKMZntq6KsrFxJy48
0uKEHbuCgRJHDSjWSxY68VjV1n5kMfhunOwNzTfuMAerKd2tn+c+E7+bdXQixtQoKhZnajrKYY9I
O2Gj7Bfnzab+M5UX3E8LGRSKbim9bOxO9KYirG2JnF/N9LjBcwjbDAAzb0fNgYL+QM/wruQhq7zk
oCf11riop45Mkw78OEUaSiRb6uRdp3mSDA+Z3qdTfL/v/Nf4uLx/9mLUugB+71LlsFSF1xUlA5F5
/QCSmWH64JHTf/gUDpAsL7DPBCckdamcomTIkL+iX7pACuXeyp/nm+OvJLKzs0P0JhwV6/DNLIhx
QOf9VXlipXLr8ZieqaWeTujfp6X8L1tiVYIGu7Rejdi1xeHRrGWpfTeBzMOFHeAYHXbRSjZc7+7j
90C+RvHA5Nq1v0BlOOwxfFW2TA9r0gDFS+8dp9KQKsd5hvxBbln+e9h9tUCmw3SLgrp+OnMwgmuj
qJK0iKVHUitZSOBZO44HlpQxtWZRMMqsY9wduA3M/J9ap9kOQHidBiZ5Uh97W66HOiR+BB1mJhUa
dHa8/TDCBNUuKjWhlFa2pRQ5p886CIb7WQwRGYQ7E2zwGH0Q296kKVecPBw1GF5ofapYXrVknjY4
NKTuQrGCapqEQlV16Uv/3YBNIxwzXT9E5etsYbakfZRajnaUL2u+P76UFu6A7DYkjmrOtk2Bh3av
6m5porAu16CmLd/1NxFMjRNDxiF2YedLtfd/O+C4L7foo9cn66pGEGKtTjtIgmvjlz9tA1JIah0W
5VnYMjxrTcBKYI190YLPRXS4ooqONoDdI3fvmvaezX94nIMYsQ6SfqxrJ7bghDPAk4F9alyqdro1
d7OaFU1QnbbV9gslJ9qB3rpvrTIx1V1U/xSBsZrBFvcsQ+4eDli72uAdCh8r9bjIjCCJEsJwOyYf
MQmDX5oHoSI7VElBgDPh9GxZK/p9x0s9oRXowNz9kjw+p9XDOAqnxZwkPFbBNt32GDKXLGsgOs2w
1oRvHCy1Ci+PP5n9952TIvhUoEAQcQu+yFwNJVGEibmK6N0/XqytJk2P8+fhP1SuG9Ka1+2EUAm1
cW8aqK54twdq30CSkY9PGzBAYG85OCHVcvlyHQ+4dDR4JgsGTO4FzpVXoJzlgJWYz3pyA/jNbL9z
vi+rLE2YFQMch/9mETEhkWxyXaOhlKMH9FvG86ZFr8XcVKQNcTLdihy2tnegfhLnEoF/TfyCjtxV
NATaJjJEiX1sJ7s1tXgJE2kYyLbp6Si9M7B6qqcqV7bP6XIUA4l9treEGfAmNh8cOu5ZAxuD441u
9EcsDrDtLR59KqfPPA5KwCUNSQYkbu6z/vJ021sHnBfGrQPoSaQYpwf54gIABUlPy+lq/R9/7XmT
JUreJtrk9ARcmO8MxDx5LWB9+aRDOeGpoYghpOd1Vwm3NhaP3Ke+rIvmdWXEO2btpVqIeKwZKI4S
U+c0fd5vXZiIOGtJXVtpE16OY05WVBJ0KmbEMQ+oD9B/2EvTaMjbzHkg8RtFKRguDu4GbnxF6U02
EqB4xzLoLDpSFGmHoX3WbadYmUyfWDeKTQmGuDJtBRUTcYraRUeicceGB54zulyKCudsoRzBEhBT
BYKEF2HtE1xxrLMb/x4F8if9QXkIvwGEzKiMLF5oqZZYq/ZJ0/RZs4sO3dmop8quZMchnPvDbfEL
NrSlIjtoOGeIZUEXS0EQEqcE8IfnLtWxUnX4eTyTCJ6jZ8MH93W0osEBnZG65hhUJbMtuOjVRsAx
scrpxI3BPaCmfbOTWWZMMjYgiWJRymFVv5b4c8iR25s2++0ch089pBlwfcz0bcSRLXoffxlB7IZ8
NywFjmxiis3Yea2qUATqorOSVXpL8rb3RxMWha6Zq/KqBA5B9S3frc5ymHMk+GvNXKFNgeKkHXqh
avSkkTebN3QFhz/GKJpXrMwUpiBmWg840YSN/5cTMWZ2UXfWVdQMvJcB5XbPUG8mSgbKfg/6zA7w
S4vvBW8yTuXyBfqi90vmdQIXrFbaPypnqfwX0i3cQ6JzxPEPpeppMcN4gp0EL5Gdb3MI+EMF7RVY
Mshg50Voor7680/pnbH9d3gbYPK0fQ2c9/7sm0IUnxJ86CX3if0gl9Fxrt1/trwwUL1YT5dUJ2LV
Z1bnUfbe97tiDSecCGlfnXZ535MnWxpvCZ48DzlpVvsxBa4mkFqmDCSWBBTEDIO5duVos9wlgzlf
Bh638sAZP3Pn53iQrcmGXGx0+pZtWPwSh0nQ2lKehcTjEiP565qpRqdM9FbbNF3aETGzxsAmDYj0
zNjnF+4SLRyagZuK1PAwKI62G24KInFxzeaBLIKNjENeew/3AOvX8qfEKSFtMn8g3S4DQ/vvWkzb
ijx4XZaWgR/fzOExEjSgdE3vOivTMqUFrhedLCo9WZVxNnSMX2nriossOTbHl/FfchzL/dsSdSUF
yeJB3dMMWvthrtikVXSx3wLTwvxof5K0C9fOSPei/1vonlPHhqgBXfEi7ODAz+UucWVIm5r5Cuug
UcAmwx7q+76ytzUpkrkibXpOOQZYZyYZy1XEf0hXvg1zjOq+WTRo30pTqoUyb7ue6Nq4pbZbeV1d
wRPUBxIFOD+fvjOPAQQ9AXTIKSrxMVTxYcMAWsIjQlIxcgxlVXXdFPJ+tAtV23ZuGACgExww2Ezx
EhwPZYjf1cyHblsM6UcCIoKQudxSibxUDGv3DMjn0C1R9oB6K+aZlgbfPE99nFrVonl9GJ/M+I7g
rJMB78a+OPivhcg6u4IUm5khwvnB2fXGueRWDTCISqAlox9Ncst4k+hiciiupiLo7sy1KGTrOfCi
uPI/K4O6o65eFYjmh7YWLXNn1wNSCZCVQ81RHKZZZGoV/ofaWlMAd+sJiUq+eoGNZBvY6kOHInTD
t8j/wwYPVwsgDw9+bJ8sMCsMW7BERVKSmZzEqjR9QgtHxkUPJ+9AmRMNMm6iaOrtdQ2ZHkppLqiW
GzyrZD16s4Iv3yOgGXGUquTpNJWZtDVQsC5qJOey1cFB3HOYWuRM2hNWvtGlYO1a/bkCmYJQZ1oU
21tPpftM3oa5mae/MNpTlq+79+l7d1Fz1kAXTPhYVCukJtEGqv0lT0HMVJxTBtJwOniIVrKCOBdI
c4QZ5OKCNzGgI1Lontoz1AsRaH7RCWu65/LCCOi50p81uDX9ONfveyaH2rBi44sJxGqQrIMdmbr4
Y9ZrkCAH5qK3ohiD7zlgaS/fLvcPh3bfFWnq0oaSJjc4Xqn210NYQFK2boxLyYYT8MTYWs/fMZ0S
LrzzvhzrDIn9qnWO72uxcx3o9xXvyoEhlcgR8JcsuSr81/UyMryvfd58DrGaFJ3dISQ0X6I2dlbg
7JPjkUZusKkyP/YT6oOEcLQFI70FgER17KiekCdEx3adsevgqBvUb7cBs/pmJ4piXvqZZ4le9puH
8f8PrlbODvzFhSK4i4//kFmia9PLdmzUHo5N8JEkP7Gbe9dLXgIKTv9D/iZpOnqgdNAVQ4qJaDYs
sV6Gd72jhkFAeRwvtd00vH9fj7gfSLR+kI5d7dnvsZSlMm5Vv2djQYQv2rIkT5eMPuFjrz56G6nP
biAkY937MD05deWiCedb1zgLII1FMmyytUGjd9iBpuaramC7npZGyKqOKknyLrdtaBAbArlxIUV2
Frq+6eKRixKDw1sQIDODv9tQ7IPSIFdJzDb5e3duw/ej/xJRE9FkjD1r2dmbz2M1IsTbaBL6WhcA
hmX16vxBcfRZ+KXS1VttYzdGOyIaI/jR3Xu3SVcOa4i83sSWM5uOgo48/laJ4i24l53WParSkDTo
d1GXSheepRiDxe4OpQg/YFhxAK6TxV4dyBHjyRSYF48qZuxxC6zGAftT3PFYk/XepvO0oPDdEOEQ
t4zQf/NsIIKYTDVJseyjnx3StK0e7J8Xk9nQlOChvtPr9yFXPe6e0AZJ7g+sOFOa7SithMio0u1y
/OtDsxGAj9dC6IF9vnY1fYBcaGzOYGTc70+pDFJmTlFDj6FJrKOicqBG66/2UQh3Muj6e5zboSPg
BxND49/z767QtSJlp8zHxkRC4CN+LaGAJjUJLmp0F8vAQ6jNkt5BZSrus7MrQla1qC0lwjmRu/YJ
2I+yS8NZZiUx6r8McOxcDaPBNXYMoV+eZfM/MpF26eCwVxOi7S6XLgUa2nAdSe2UtWEwLUHmzknw
u7JtBy5LX4V6bvnv9F7PJmMntJm36MaBcHwnD5yfcJdQiSvxAjECtZQPlUOTx//1CIO1cH38dFiy
c7D2d5F6dr9l9iVMFb0PtNUBGnIutZuKfYQdOUR/zK5H9omHVIu9Ue3ABsd/wO8SQj8j9FnuWWYf
DCIhVAQ2TIFzGx3+krXNsVPm1n6ck0S6svopU0pYQ3xTssUh6dftiGP1DmUgFgUIf0rL3uuOr8aW
HmfcyAWfjv3OJ9j8cL1i7ccFV3hU/GRPPe6vq2fulu0TxFh79YfzzETv3uJyn5Zap8MImdv2AYfl
SZTG+aLzMjQZKyOrkNC7Lxe1bsd0JHJa7XucpCRlW5Em6SPAMrc0mmpVoNYDkQdlOlzcF/rl6NJJ
Mt7jsTwld8wXiqc0r/7N1uYkl8JUd2GsGbMTdtaBGM88oCWyMplckxN/YZHjzHrUeFCmoF55RwW9
KX38zr6FtMxwvzCWMV1Ck4cDcbK8lp2hzY9ohOlkG0tCT3VtPE92SKvCQOQWw+MjRGDE8kHvWwd5
XMo+BHLp/2A2YNFTP0Qq3b32oQin3gDQ66Pbw7vxQgNMDDUuZ8stISjBDc0AYnOMeqC64FgSrbtW
19lDnv3ZD0fErk4sx/3FPI4hBalBiAdgVVBc3N114voxqAKy3kydla7R0unpq9uz8JBaOK9TjxqW
fcpVGE6/12apT+KysjySZCuQbJTmaWWDHAxPkS7m3PuOuC4WHUY5iDzTRqvNLkDo87uVxi5zqisg
M9JYqHNRim5jei3SVgujqMF5MM+TWqxLGiWeVOwXdBfNpvI9Tqaf+T/EalXJHi1z78gmVIRGRgVd
hLeuPcLREQZ9ijrolPZvxqcubrSJ28K8qdV6isJKGxhDdR4g7tNXoSTR2xEv32TLo1zRDEoXMvQI
ep1/SdgsvJKWI5oGBEYT8rw0nunqZFn8+SikIPOd67IhpgONenNod+IZdXBOenBXYgIRP6tTFVvA
BtcDYUHDSmguMpyVZyioELk3YV9CFYPfL8MaUCUt+4HasrmHb3p3QG+qdHrQy7tjAjyhhuOIdODq
bUg4pNpkwwdR/WWYEBAb40o4beApilPFpCHuzDk77dseoAIB9FnbsopcLac7Uarqy7XNBJR3Wix8
3W/r5acEr7cv2K6zyzfasyMbJHslEOIJuw7voXLT0nJ4UfIeKTHgu2KCaU86ie/dnZb7t2YytPOg
oM1pQKNgugu5hbdWtvNLFRqL2sFiQ/M8ltFX1H57aAOz7ognN1NNxC7uePtl9La3PtlQ9JgEQrO1
ptNu8IPYM6t9XiozzL3hftbnxkeuDhz3+D4bpPmNAGzO50YzIXekl3zHcJR8hR+NZgJK1iD1SJdA
RQdudUP7o9f2zGltQfiOFqXDON111nTgNJB9b742B/1FTiQ3IZBAXjopU2xLPBtgK6Ff/4Qbr5pE
SzIWyE64gofxXw5W1XFEHXFsPwNdnmE0Kqy6OZdBUAsIFEH7BaEr88cp6HNzSyCzXDuhQu3gmE7U
OKEH106chTOWIDUeBqa5Zq1/uL2imu0BHMb7KZX9bPnIna1CHQF8oXG8EtFKOIv3P6ZjcfPNIICq
KIBql7+mJmTZmyNnxNEALxJIlrZGSsLRZZf74dh3QvRNEjkcK7MPDfw2GMTGnmtA8kz+ao1KCcaZ
bLaRLh2nhaaqOLGVYbE4HKidmwpNZwiEo40qfiYnCaJrKav0Tvt3eNEtybjIOEe24UBxt/kSOF0Q
lIMuJA6mjHuCwychXtz1nsyC8wVY60JNSskN6S+gL68ib9gMnwcCnJJMRA/QFaWMHdGRUzB+ZL6E
jdn4bxRu5qv8oWTkMtHINGpNLbjgp4kEjU6YkQ1SQlYX2M3Tx1CXySJk7aXUqVh6pFjCdxbryper
RifGnWIeQ2H1xtifm/GrM9mhD8tmW7k6uSpEDwsdFb7EEB2eDLea2LAW8HVHjF7c1zyO9ZQQF4o5
WBR1SAYl4KbcBzizCbK9+67K35PlvQZ04RflpNX/S3lQTecwMQ1TGLh8tM3t8Z/lkXcR7F+RcRfJ
/G/ivpZw/Ak9rE3SRJeHG76GZmxnu4k8FlkwE9hL/tgxVtKbj7mUez3BdPf8YeNtc6XyaDRb3QS0
YFgX2fZQrJ6NPgD1ApwzUDutUEIliR4RULQeDjNd7vsPzLT6jXjyHNKxE+5FJ86hcgjpJ/VT5AqO
KZ6wEepPXB4h7qZZSZ1gkxndlhcA4c3UulwL9yX3giIqws8kbn9n/t7UZWxsMb4u4OY0tcCRBf36
TKTx+tYaFz2JXrquumb0r9a+GFaqAdfGDM8GKiPQOR1xegjy3WYetlokoxD6MUev4mnMek+suNgW
1S691dO2W6Z3UogwmGGPorNoz1EJB4NrkO/rPk4pwWqHzlioICq+NiKYFjU5H5P4SxY8LrNeuoVr
0MYLKH2HQppRxtADNGMNZHds1IY2nSr3Pvd8GuKyApJzV+G+DOVErgf++ZQ7q2TaKD/f0xXWiXn9
eMVuwSY4aN5DVtYFEx2m7qzV9Gz6USesSkOrZN2TPepY0HZYjFFH6X1ElPl2ZNwle7PkjX523xmt
uiaOu7q9pqed1jpt8S7Oo7Y5DqtPqHTkPpyBVhvU+8SRLcEmfNdzhiaIj8rR5fYfMEvdemUXdKDA
SA+ISSFbaiIT+urWahAK9OeWgVkVpcKGrizjqvADMhBbJ8a3mZVir+kn/a3e1REY29zcz61xjI55
31NKOQ/6L8WjIhFPQ0lZie9CBuKVwdbl/1ibJ/dAVdrfxqwQB4EwJwgfuE2Am2Y8a5BJclIRUfxF
ZcaNwqLT7yevzs59aWuTHXI41Dh9LZB7ojaTrQJOA3i0IF9bP458SMiJ6r3df2nmNBPU3CfJPHkA
43YB8WGPM+HJ86UsE5BstXLHQ1DSW5m0RvgXagMMkMIIgm4gvI6sYzHk2hBTFAvmJb6zP91T2MZ4
ZWge/dOvg0WRdOxoXXyO+L8uvG9HtfLQzKsRK6pPMfV8cZ4z53Yx/mYm8k87+GWQxkwEm1Nz0aSQ
pDP00E478Sx/WaRRdfECmgaA+qODSNA356QXVSkNJX3YN27hQArJzZkTk2R0mQKvzxri3ym8Ojc6
655xlrMuwIEntUtGl6peIvuqEY1/zK/p1S43yLnaIZAHepvGn3jbaeEi2FVKwXGNZ48BnZfveY0V
iE8LyTrcAecbnnjLLFV5CJutjW2+ByuBkZp3a/OCKthl/BgeaKkihyF4mqInj85y5EP5LZxXVyhn
wp4IxvbUWsxXyux+/2aOIorC95RuIJ4dVG3Q+7geV6Acdbe2PqC16Q0Ms5pGjc4SzcAnzrcLBZ0u
6oPr7TY57FzWUMqnavOaP0QJl1mvXovXYyuVhgapn47RDiGSQDmtowWrHn8qaRnL4K8r6sMCwE6Y
Ng0QME2yOeq/7Wf0WIVbJqyfrDNQwdsZxkrMJA75gy9R4RrEjYEI0mfcxnr2LArFnGXt6Ofck6YT
nSqzPuIiyHee9u6XmIMpupTlimep1q/XLBDfAWibQ9uJsIuE0haY4/lUkMDg7mGEKcJBXy8OXh7u
VtiytpnMgJVLFIC6F9Jv0ginhegy5Zs7+5neQF2jvs0XGm68eOQ+VWC0ctEU+IF/NWcTG6PPIa7S
2L2DsVl9wbUy5mf+WJrOYh7B3ZKutxDvCFNcXsKVe28gif8+DbGfAJBxlhchARuCToyitEd/DAMz
HM1XmpoIRK4tSWA8SvODNC+u8hPOXNvtGReCdAqP5Ns1ZLKEbfFd3FqzicVkN6jNUDhkNHIi4yC+
LxS6Ds6fbt22iwdOw78rvghpOQaga6z3Ac0n8MEZwD0hXMzThonXAWY8X2FrejSZ7zOOIX4M5s+c
+Bw/5ouBUBRIjhxLP9xFf1BPmSVA6TtVuXwb//HLbMKfxrZ6tXIfJYWrUe5DKi9NhvSpjFVz6lXx
O3Yiwzcc5yOd+oUROYGGUFaeTCKbs75TMBXwRD6XOjU5dWqGTICJqWSMD5Uovst7tqv0DmN53m5T
It1w9cGa1/AWGOzjl726Yuj7fFEA6POrbAcuUll3//k6IvUv0hwsL2TpcS5Z4cyaeC7y9ope6sGP
ql3OCzi+0FH7I5SaoBNFQHGb7vQ3KOyjMV1EU/v5glu6/u/ESXZ5mMe+gKayIZ6qqYhumYU0kboe
wbLyVfB6trSXfQ9Q8NYuaDOc5t2w3vhEbvS3LFbbMshv+GB7MNCJHOBd9RHIPb882+BS0EZPuyj8
ysx2VpHkPRxf8Ywxu1e23G2WWgOzpYFAV8NlRkQFCdajvOPnzfNA5RdELAe20r1HiF1BHgfz8WD9
oZX2A808jgfZllS8S6P7YbvM+ecR0SiVfkCV9tvDOlzz+XZVioAls+BDHUGxlwSFeml2FGXNVyfi
av0Z/Iw1BI7sezKUABNfDusquzAC953QfBIpXBKDgwu9Fv0VtTotFf+q74oSiQidqJwRUawgCA5h
QnyUjaNrC+m7EEv9K4RgxZLcf3DPn1E/w2urkflrNtIvxQj4InPwyrrmiybZP7DyaHbrTNo7BL29
9B+4jDleTMM2vFjkB7Y8tYz7KeqtTzw/6oqcTWk60bsIiUu166zsW42Fpm6ca0z6QNtJ7CzxYKck
JB15IWDdXfaoc5zCrGBG4XwVwtILZs8vbtzQaSvBEWbrg0wABblGQrpGEzivEUKA5+ZPGdQ2Mlcw
4oLU7JE8mRHm01JFLOuLoLKRkHZwvZWYJZ/4oHeXovKadqoNre8ddhAUKvqeYd79EBv8UhEzQZYW
I2b6kP1WbNB213j9YCeT+iPFc4zCLmHJ/HaEi8goopCOZc+njZNiOKdh5qjoDT+atFhbG5hJi7JV
v9OBsFu+7IjEJKG6n/XE/nPFoki1ayaSt4NVRaZHe6es5qnJ3kkcxB6vgmTPFXICB+1NFkVQK7bJ
veorcu2CmRCKLcxw20S4rj94VqDKLP5SvMj6H0ehJ8sjioHzQRwMtNMJhy0tP9vJjLIDNBGR7tff
oC9C2KPjp9nm0lpQA4tKN5vJzIk/3e2C810qjcixy661KbCyQWwX3ggxyp+yrii966rr+qoXU97+
xNw83YuuwgyoXw/wjHd38wF0lVoyNe+8xBE6BaemGndfw0rzgX6mkCXkCy2Od/zIRQK2J3OC5XgE
c+qcrvJOvM9/x2T9DdKOkMuLHMP48h3yueEsVMllBQS813gNWoFudTW+t5q7nIPJgExzAEtYuJVY
Rs7lSE5AuBWs9d4TiZKtgjMqiGV6nnNwo0rB+ZmYX4YJgMnHxj5kwc/FtwGQ4s2KqpPqMe8VX/W6
eLYQ6LBT9woKWpcWm+ySKEXUplX5ZqDBnMHpMJQLuS1N7VtkL4cuR0xz6pjJq8B3wkUbNrOwkYuu
cfdfgqbxdpD7kw5QYu9/YCroZwo7EIVzWWzyBS+Eqe45/SeqN0jQhmGr4y2B2HErRU5oaj5MYz3V
yqgvKSXiUkJ2ioSAVQhobJlbi45yda1rdYEnRn4bG66btXufS2ZzZ2TDVq6DIJgLlHcTXawwdPX1
f4K2vXS4MR2gXNjxyOIK/QTgw5OEWPhilyXmKHxqpkEfaQJm9lEJiRAY235Af7FDBMLc3+ieMNpg
Zq9zi0FwNxWOb0RFiV3/4nzaZdHQYZDRioTyqA8ZbAq4+6IcOvvaySku7oJ9X7NbKQKWK+vu9RoP
Sh0qW8e/5ycg2w657GFa0Q7DCTWJh/mgdnYE4Xo623z1yUgFNZMluQicEk38EDr+/oUwIbeWYPJF
ziBnDqRvVVr1vPUBjymaK7FBIuDkCSzTEmi2FQOG6XpjrrQDEPUorm2hYsY5C3/rsodjojgrIyIF
9vty1Ldnzk2ZqYOBTwsoptEozwHNFGNXi0rlGnQkR3QW2dxessH5SsJnMdaH+L4Ewyu0eOcgC3gB
+gBU3wZ51sms4EnsKqMRrREAQpaeAWXf4bFolmzP+hgNhZUUCTpYf9L/j96wjNt4B2hU6iRFXCyl
0h+u2MrlU7o1PhHpPisqUswD7tsjaq2p5cg37isxkr7W8QNtkZvYEe9MkFeHdO0sNfFmxSMlP/HC
qj2U3T+u9A82QVCsedV4BeT7HtARblRmbVoFZUH4CYq7Gnb8FA9/qzQy2pWn5md7CPN1fq/bM9z9
1R1AmxQmtGmsKEkT3tl2bQ32Sjoo/eumytYYM6PbJiDw122x1Sg5eLwQXAAm49FwIOqZVGX58WB6
IlaZa4ulOVCmY0Dmsr+DWXQssSZJ+16dASPx072vwOoxW5b384056R5Xa7g8Q5hNV0Oq34lCMyVk
FpsqELx7z35LNN9FLMa8K1KnyIZpM1AQHg1GkPoE53Vb/SuLYxRZl4KD2SmhtvdEKIgUCUhnKOSB
Tc9ULwm30r5uRX9oQNvf94C2IIj3l3pR9knU6/g+twRA0FFIPpTuI14/PPDr/wdy5yAgOyWeEObi
U2U9M1eC03YXCGTVw95swjGyKz4PHM+2+ErQ5AavprX5iIyMNTRSOSwYY++CJwRE1B17zYACHi8o
zf3CG6BTnDQc03hXx0HZXqgVsWUgPFVGanEI9EmHOoZMVAoT6gyIWAHszxCOPf7tn7/clp9WVIWd
PahY8KNxQWCSxKOyI08IdIWhmf7UTZndFOWFOnY8DFingpttPPJii9NU5Cv0ECzo8pfpzjYTEp/k
KFAUBJMG8mLIZn6hgCzy2wTErsnegDLaeWHaJuXMLg9OhYOgn5ZPptIM1qRW+aOgBbl8O9Jh+2h4
8iGDPmG5c5Fk3l7RClREQVzSolfP2qjuQiy1J4tEWw2Xw2TSM6yFmtJIUslee9V32DTW56xjJEYj
UVwSbJcQl5HBS+f7Kr7J6y9V8Nm31BuUVNnSLrlh1Wb1Z9OBFeVYYEtZ0jR8eypuUlXJNXctyYtx
JOtV0Skwmg8BwfNOgCZvAzVjQZKdXbftQFzl611rzZCJ1q062aCrJ0AFJuHr55AbyRgU7XaK7bis
xllo8FxxmdIfjI33XptSqSk8F1ZEGFy5mMrFo12HKcFCBIA7gdOC+Pc20r6tIrBtGem+lm/Z/z+s
JgTFSReUdCNp4G9rrs1ARIMcZ1J00Ebs6bE8h7ABrTuRYSFOl2kAQ3wuKPmTmM792+SXYMKzrBgE
0z6neR7HTnRFdmc14CEKv8REX6W6fRXkywf5Exi3jazrG8KGJgXJRiaOJsq5+303UL5ZFHqwTd+g
fNrywAn5eg2UDk1kWXypAoiMh8W7ZzdV2pAK6oo1lvMMIjHddmuqjbfFdLa/7hXCHuPm4Tcop5hF
eeaZfj3wXsbWafVEB7AmCeApEDeBukj0Z1h9ul+TaHVPAMxdJbwMTUSdSxIVLaB52fNkSt4L3qFJ
bc5eIg0ccjTSnSYbAYCyoBqRtadzLGjLefBgBjAAvvdZDuAAbu2blHXAI5NBvMmGDmqOBh0TLUJL
jN+ZA6bPWfRXl2hn0Coawt7AAflGR6OCAO7yKZd463BzAnuGDxgoHIKmljLVT3IYgnKgtA8sD57+
ejJ5NVrAHNvulS8a0PPmg/CtWgpsjy3nuY9iIfnp+z2UTRm1HGcFhbF0wDkTHvaV6X6d5B5ELWmy
WC5G+jdgo+/xTAGiP17a2ZumTwXCEGFAnPYpItZ0J5VECvevDpuiHbkj5i455CMomifCfcDxmVx4
Fbhz19fT7+8FJnfk0gRCMlpGdOfDfpFdEsvaUljJ9HAK55k/pbipiQlURUTV3VT3Sief4y/g/hef
XEvjfXUe+UgEEQLhrideAW1uPPYTLgPtfWZQRkTgM8g6b4+Pf1W0ELghX7gaZEoZnf/Z+JVZWXBI
WfkEtJu08OC12rIDM55CXRSUtaE4Xv95hVJgxF6wwXyHphnPrlwwHcXftMVMwhKDoJHTO5HjusAf
FQQU22O9bRZCDB3mAaQ4vTNTjUN5HFMb/JLX5h9VQHqImOHr9UOHYUnZkBqB5EpKG8aVyqoR0eMJ
triS2gOtL246X00wXpPOkGmD2Z+DhKVoAy1BjuGKuFGSk7PUV4uyBZ/4uPZkIclqQNt6EemX1v9Y
MOdnD//3D3ooyxb1NOcfAnfGUucIlGyutxdw2szs9AXC9CPBbHMNLMDJMves+YLjcVygNLmj+tc/
8JTxa+3LhwIlKmRZOJRJCdb3sgQxl5NIPaV1Tmyig40JMOnx73P5DoBq91lYA4fVW4Y26ByghqPJ
wMmMcZy33fGrrDCFfhJbvpqZykxbChlIzegv/G6hVHi+ZrQzNwnkMpmrohmLyzbaLANX91F2vsCb
BllnAgE4TG/ZZ/9UaPA6bUuRReF5gxVykESjGY2Fm+eryTpLHVKSB6Z0LP9GzYbFl3mg0sJsVH27
MgjuVwzJISVFlRAN163K057OuukFfX4VxnwhbeOiaur27iOkat6dSmqNF7a8ym079fzVr/kMhxno
Z90DUdFQrX7vVEpKDF1DzWMnBE1SyebKGx+7QLTDjV4VV5q0piLATldlEGIXC2UHgyVGpBXJdB4f
FHELiQssY55rZBsukxGUIvlW6GL64AfxmSkJY4FBquuNu457Hv7S+QSK9cvxNlHw6J8owNt3/k74
u5Be4Woefj6gLPgI38XZeLF4KBfimW936WqLQ5nGNCZFJxHa7MDWSVxvpGmOhDHnchJXqHngp/EA
WkVKs7ZeN2NY/VE7Lcl4qakmXmRHTgWi5VjkboKTHEkpHtN1FKL9UjK9WxmtAXAZTo2+bDx1tgiR
HrblTY/odSfmhFM7qkQdJVO7vtdHL4NFnGfo2zUMIl8BdsCY3mYAc5KsDIOwFbP5PuwJJxkuIugj
Kg2ldqRog9UESAx+VQu2HlslUa9nsZEw38NwuMD6NYcjd6NSC6cSQ1Sm7eG9Tq4HJfwjK2j3Cdvv
uwh2Woq0PEGguOH5pP+4U/r/XBctwv/ViNIwqHfLzTg1cDI5jzDlXkEbgbLiMU802ugSDV7uz3G8
aETmKrfWXWA9EMzzcG4/cATQINacAlNMMa+00uuTKsvUZCM/8sZXNyqg9drEE/PCBL+sZMSSZsjq
zHkRQ2+jvTBxN8Tu0ciYF8mllIK6r9mPQCqVXQ8p2hCF32X1uGzXeKtZvPNt+bVRlUwlurVaP7cC
8xOn8y8Gt3zFa9Azj1JC8hKjmvhycQwealuEJvKXCEKAyGDq25wxYxdsW9AaBxs+1zhGtH+8PwFU
nkmdWgPpGyNice1DvWErANfz4zIT9ELOdBE2YZ7nFvHEVZsfFGM/hrPEMCpFjOEphbCH5RrcSvmo
NDpm1cEx07onwXXdCJpdlzPXALr7I96j714lizH4O5QwL+BKG0Wvz4v4n8jg2FrCo89inFKtZ5AY
7bkvhdckzEEfFTvOoKbRvKAjRhl1NuuqZGJQ9HqBG+c11ZDj7e/9a5OPBW/ca2K55kpHWKObCdd/
2UG5w3/4Yp6kQ9iLyfTmboBS2VWIfk4fPzCdkeHS3A5XLPaP53VUhaUiAHAXYKFFhUUDSjLiMkWP
7b9uLV1PQaIGdZvvQvv14/ksDwmxvf/2XOOg/FmT91IctPJysXGZFH9jA9Y7NSVUD66dtP4BGTpx
yarD9aP1YYwCUYNgrk01B+buzV1Jx0YQDq1pJPuBJdVJ0DwvbJjJ/IxOkg15oHFe8/n+QjwgiZxo
R58A1poF+hj8nYjJWDd+dmkFuldoPWm1FNbXNl+1X6iz614PSmj+NYTt+gDSU9L0nb87XjnWYhmy
HzGRntnxVTfTNTyQkuz3naXuN9ch176z24o+MvTzguxPCTFWS1y7YEdj64r2TziddJtK//UGQ2g+
FmzsOZ9r8Y7+oAtBg7+hdtb49MiLI5yoInk6PJ4Xrt8ikN1AONx4KHgUOKAXqyOHJ3dD7FUFlBQ2
PcFXvC+IbaHIBHxKi87riv4gGiNZSoA8reRmpYOWgky4PMsZsnpcJ8ZVcF6ilTvLyFZOqO58xMLV
qMIKEy4QsKpNAqiXxQl0RwHvlss43tTHuy2kojekTIb0qPC3R1kksa3ZBTm5j0S+PHp9rs4lmlf2
T1aGaTAwUGuMcLW1JM6AG4oZsTZPoqW1IwH8tGWQLSK791fSKl2NFrqyZ+jr6E9QONW7cusE10dC
ppBgiZbKsJc/VAUL33F2mrQ3SQri9ELy5MqZbNcf8/nDiIQaw0E0zFQHuVKtOrPgQZ6xNtQfXAFX
rNN+gKNZ7dTXGC6J7U6AzdJAZvAvzidQ8BhjajTLXtSkiM7TN+ARKXLUxfjwM1XAPveyrwozkS79
Nzl3rvccXGyfHsfPOSg8e/F2Wyq0MPyBONGBBb/bsL+qUgiJJ4PdJTbN1EGc3YolUWWPwSrJG0Je
cpKiyQwVLa7M6kUeXA7NI6+rcbbn2+2mkMSUXP0EZgnATGzi4iqbw554awIcowlZTK7UxClTYInb
Q0mxNlWHBnqNrNubuMVIEoMpNY2HRs2eK2dII70AL5jZNWR10ZVk/UsDlbUfgG9ilxSSKZV9d5Ub
pt9drjRSDhD2Z4GudKsRm2xRRpsOmjwfYC4MNZ3m907DeQXAGimhzkC6+RgnRCi6znhx62FqpC8m
rZIaZNRI5liJhT8dgoWGK3VdD1eo/qWl4mLLye+ALiYe2laUViQk8LUGuf5ilFuKC/OMYyi1vAjb
pb4jnn2ZLmeD5udu7c0xluV5bOuu386242JGaD3UAoY/yhdNZeD5Pn6yPHQZ9n/NhcPqR2j6VWUq
XH08xEGUNAb+v40LTkP6FHMs6O2CFJxWlfis0VSnt3IdaB1kl1LUesrJIKWNJD2dMw52PBYWQ1rM
ltmcHej0LXFEackFT6EYB8dQ2WbvTYdandAbQ/bcSeAiNrhsYcpL55fVxd9sC+iPRG+hdukLFbWK
CEIILokAwTuAHY5V0UcsVMcHWWO6K5d0Bon2ltbBn1Yms7I0Jai9Fw5ge+Iwc3ig0JsqX0ALBvNs
ytlGV06RB+4zks1d2r7YLEIaRsIP2WhwdsWUs0XhFQLRg1cheDdJUxq38QEHg5cvOFUlvReMvMtZ
joOKIraySVSP8tgUsAUjKpjfJCUA/LpBkexVlPLIMtIyrqRPnn2FqYPDoiuq3EqE7gKwbFDAulEK
91LItceKojjrqQoKfp2WVOl1ZAQljmWssXKlcdtngb2QkPSo7EESkZFeqO+05QGqcRzHwOoNzBuF
dztqmdKUruoD6ONFuQneJJSxKT2Lfnpan2iAEq+5fGw5P94/50+KktKn6L1UUVAWxhzyQ+yWHFK1
udVKvwZp+FwjMHUbidVtqMDROdLQ/7g0yIY57Je5DZ8t4gSR/Vb6C9/XQXsHwiBloNsulIsTen2W
3jqeLHpqMF9Yl6tlwgirafrwssKeVan7/2AtH0efpknoGhbalBE61ND5kjPx/c8259plURTi9Q61
ovwdPnvnwfuD39jqqYzjpaH6cXsNIeYNnEM4VFmrYSHUDj+sLqgk2RHFL4MNC84qZ10p/1pfDsCq
hhdlF8RTBWTYgogTeGm/+T+fEVZ9UbHiF7k1RQmy1WPwImar34IAC0U2uOt5pwoHXjW+fB+jiWbs
X0GM42Y2b9T7f1vpEDj55/gJLwl+h3mce3UTytRnvgtFetqnqQWLyp+X31E518F2eZ7x+v/KlbN4
20Izl1+VrnLg3zqZvqUNOwwrCh+NZgQIwm04RN62kCtLQfOroYu3+0URRgtXyGx4kQ7Kj2ahONrx
WF3OzgsNABnrqyebGQi6VgUE3lEf/8/EqaeAvPIT96Q4QT0nf5RbQ1c11cyem4NW0c3vtw79S5E4
MU+V1SzU72liFip0a7t5TFEjsVlxZ8fHQrXkeRir3aZ+xW8zfsg4D6oTb2m8WaOQrt8Lqcq8MOFJ
kZaPu2C6qz4+z5mffdz8VSuUhwoIAPvAGzsXjA7vUXVcFON0nqxBasx4eGn+4bS5L8ls0cPQTbxn
7ld2orQDwsMobTJ0jQhVk5CHto8nnAkMSIxE5gBDOJVJwBsum4UQYn9VcZk/4rd2xHxHsc6sz9ti
HLFEXgDnoSh4zFonxP2F+cNBioZy2AcBbbR63828vyxHjQ/VSm63XRtmoqyPtT2Dg/WJ49rxbpUD
x4P4WHyEsgJEfEsBY0eRu0EbLjcPfJZeZGOLIgL0hvxkq4z/Oa9/fMuBt/s9k+JRFKo7xaPxU4bm
Phm6UzkYPvKg9kL6DzBYXidwOHV22yZ70xi7ITmt1TZtHEiDoanNjhQNXT/eAKcbWVy67fyXPZZT
KR/3yIkIt/ToBQDNWNqPl0vN93oJmgaf1j3cvYDO7+EAGYKIAkUXZ/tq9aUdKmbD6VvgFyKriJq3
MDQRwWQ94kvccelZ2OQTpmEU6BYiCq4TS+QhRP4z93OjtM7g4pOt8hbpfRao/wQEuuHKQlKrub4N
O7XbD2C+xyVsFfcXqR7d3X2Br+EZI1VBOhU360MeyXV4eDSeocKusIqXkDDiE070xZ5TqZCFh2wD
THq1/O4vJFpG5LjnDDQX6YrSRslQx3cqJsMQzu652u8zzTZ9GWqIHjVEJaGNu8k+I7eg0k703dIx
NotBhIGjYoq0dtwB1L3GOOpJd2D0H0CWH2HHxF7UQuSmxQRV2WQqSou7VGJVM9vGDJNjTpL/TXII
0rWDHctuDM+GE69bJfgL1cjg4rKWGzPVu7QkpjYn2BNb/s1MG+griI3lGZ9HJwLErVFVgFkgrrWp
u792vLYhK9vEo29hvd0V/NdwV5kfypSJeDK8Qv+NN8SVDy/jYPhyFox2CwCyWzgsJXFtx+vWgfYb
NqRK2JtYjlOXdBo2wrYauZiPqiPJjfu5RBW7C2gfeOHT/qdOuS3Pp4oWUU8b6O9QvzHxAo8UUb23
g2BCjPZB3YxUAdyzApWNyIrGm74ebdmTIhAF/LRvQfuIix1stX6xzhZy4WHS8ZsR7wySnQfzR3zE
yhs1Yh2CrDhMbe4vAcjdnhOxUPLwiW/hlQ7DVPXD0oI2snFjOS7ASiGjahPq8bp+hs57AxJLvQI4
qTt+6LwBnFeD57i0S7CPjA+TF/PBA0J/sGDZ7zf+p1txGg62G5FrwjwHg2KNczs8ZwkIELHBiDaH
jFVIoHnJajk4swJcit2GZD9njY++gnZMcKh6fp5VqhBUSl/EesLyeRU14HCQ3n1fzg9tJ2x89Yto
RmhTGQcuy8P8bb1YRvQVhbVFIo9XyuUh89tG0MXGrJx85vx6v2djDrEw46hrqAoENhfWToIvOZoQ
Vz80EPe6IL/vB7wT1x5y2PMBqAgWDEsdLZNB2Wik9XxTRXrzEWakYzBzqvowobgxHRpKOBid3x7/
cKCW7Y9yuxytf5rCzyS0xdMRKP9cdiCnEfw5RFvVYM0NoIZxHBbLZqMMv++V5m8wlKPfhzCsT9Za
8ZYUmnp+KHQ9CVOszteM/kH7mbUm6KBpLbKbGdAvT8JNXrMP1i+nh3XLGggwozNk2lL/dSUXhRz4
fcXzhbd+hR+NlKbw/BYXudqDP0weyGG9+JGF/FAE3gVkKAi+B+dI6rIsL0HtH6V8B/NAD3ik2Lba
XjTsrrnNjBpGJLd1QcOyvOq9VaIoxLmyRmXnfrsPLjiyLR3BoXIpqWWwZc109ArHULBBfSye6xXr
iC4454UqE7narjh1OtrbYoJZy7Pz+ZbaCzNFExBZKMVQ49zRa6HhA4mO4vI0oZB90CP0044UMdne
anwxh/7OZv2laV3wJc/WkCDWVjJckCW4JZXFd1bNTD8O4jxhAWLWfYFl3BC437Lzv6HvHqoJ+nLo
ioQj7oCzUahng+uZ59jKjgM9PcRf7pLIZTwgLWtVj5snHKyBGr56HSv9YES7/HND+Aol4JdxzFRu
ZGRA6H3F5+LpG5YS7+izYGz4ZhKNAAFwUkVxh4cU1idgfQFHhLWVys7fLzrMa2A//8ZX0iuPnhZb
aIyj8YpxXVfQSDSlFo0gVwFuV4x2Y/WSpoXLGvXSKB7CZuISSxyi2j+p39lsZpyBc+ioZS2+69zo
+YYGiqLUmhJUqyfIUFrvztux6s+iDSbPR/TTQElUudQGLQip/1r3cgy22x+nPDkNxXUJcwaZwzEq
wUatu3tkaHGCv6a8L9uO6ccrsdC/JubRgEqt/0G31a7BoOD1Vwqo1KBlKXBNvjcXthfzyig/UFdt
YM1TkvjgY93OdBryUeqLUh8MOwsXoLrFzTmluOZ9DbQyDvKUGkMGe47W8jaQbKW9S7rXk2+cjU3a
LAAEICCPZjDe6LlZzDENuKMQloZUeMz7jCBGsKNUR1ioEfaoYKfHNPh1mMPnbm61/VpCVdKL6Cim
o3/QZK7cHDYciK48FmzP2q2rE2chILm3W2yq1ciai25IG+FY+n/OQJxv5eiuHev4hqyyTHe8JjVf
sZiWEJK/5cObKhOoMOmmzA3OwLrjZMNsldb2gRzdkzYD/wdC7/zPnrbyZRkxqN3l9GH+34ci7ARU
0Ta7djdAXrwwaWNJIGblZ03U0qmWqnTfAyo8nsbqTuqjx/z0HDeujd9j9X8qpWFDvucy4pNwMJln
TPYh5mkMb+eoWPPL1NW3X7njB21B2tHUfcA+DHl+pqRHkAUj3kvUXm+8UHWEj/6N1wJkNbirDfgm
p3cAY+TB4k0Mm7LZBEPD1lKMMh1BcXvonHgHa52QfDa9u0Ylnt0DT0BdlXH6soscCtkNj4eKN4ql
Py7SkSUK7Xa72JmvbZJPVNWwZfSfKXEYxeXQQTM4NS+7uSpaylTlRrLh/1REvsFzt8CnE2hnaZyK
pE+7rh+U/G5oKL6RAg2Cg3NUST8W3VO3CJWxbuXjuHeAqIqkIvgvWkR0r6KYvsIypYJp8uoJ19Np
5szYeoRr+FFLyEZQnn2NYLZzsXKtmgwHOiw+ZTk7kEy0C1yKwGr4VXTmDpWOVdbb5c3nPKZvg1s2
RGQMzBc1ukUVKNV6FBjgk2F5Cl2zXs4JCCb/IaApSyhN/pO8uuLzp1iS0YOYohukNaK+Dq+o2no4
oTGN2BAVKoCkZn7wYDfuML3bwBBOnGrGX/b7UTjO0Cw0o8ADYmCfzs8GAO4xq0vNMmmbAnuoys4B
fQi/Goim5L+lJImyR8KBjFa1oIY0FaYyzUt2uf/4gxYW/j5c26ZUXwa99iOyJt2IVNVWxIYlt0BJ
0+M/iXjk9BwGlLUgPd9+2gleUn1VwwDk7RNZc/RZzUCLt2SFAx+Zy+tAdTWkPIV8VHFOB+PqCQaP
CCFsEFU49qO/zEakit0lT3oXwXhc4gm9kC1xuKC/BPbujdTKNz1/zzP844m5j3abw+IX2iUThp+L
pXub2lCQ9To5AEOaYkLFAaqnhgW0svRIxG5nnF+DspKrOtnr2Pcr45usv2rj+agtA8+Uqi5hi1a8
FhFueIUjsE/2OMJfvBfVqtXqRLfVQnEkWixEpxU79bMtMRFKT4p99Lm+AQ6DPG33Byy+sD4YKIzU
UWoeeEV56b19lb4ZAlABrwet1bC3VrxW/NCeJfgzV5NazbBTcttAM8kIKeucI1nqleCuJKz+xOIS
MSP1teMjKEdtjcm+mn2nY94migkCogGaN/u+GewZLm115ZSiAQUZXs9Y1XrRWhMMO0Qm/+wCV4uQ
7PQrD2wcVWK7aexfXsAromyCqUvfHb2FKUM+En2izcn5vkHU5aTdnoGhYWOXkELy0LezpGbUPyjd
A+cC4Bn3nACNLzAMQJQ2L4IbWxvz6W0/eJh7yIwKrKpE2IgrnzWxeKfJaWFLhv9xpCW45GQPj17o
Unn+XLx7bEtT5g3nyASGnSMntRaHEQMwvzizsEdpHazh8EUb+glZI4t+0heOoUgbZghziXqK/bu1
jDk6nFos4phyWsnXUXuCOxzi05tYm1eAQwQWG49DlArd3tcClsaC23QJqCmWDunO/VGpk+IVsTVC
P8nBRxDwNkj84ezNFEyZJ8BEGGaMXB6Bqhzdd2zKNhmQmGNy7uL+zefPi7jrezdSoSweY8A0LKEA
q+mabOPFsyZgauWeZ0zSq76aJ7CcjcZPEjg7+oJSF0P3NkJVJyg68Oby5VxuQRW24m7S9HeDho3y
iOaN0yD6rx/23GsBBtSdNPKEJ47uHL3gPUrnAjwyxlf5v+oeu+/4S3hLgTnhjLxi3WPoDUV36oZQ
hjs2rBnmri2hdU+EbuPgWNynqmzi+zBQSpdguECtHqgJbYlh1+U09YLtOEZckulqeCBleAffHzcL
Rf852SEWhDsodPN5Y49yV3t53a72m1iz+kW+RrhbXb7OFvRQHl+eZH80R7/W6yYfQ3kNqnaeyKnQ
hB7f2pvh/uQcKa3OJwocERsN2C35UpcbPEAj24Un7XipV8vdgfKF5w4X4G+kDCBY5Rgq9UGJ3IsV
lC5I3+MZow6Z5wWRa6mhyK7TB//jjYqWROev39PXZUsJjLhctaPN1VluHKgyIqjx7gJ5ZLqZhxS/
RwGRiR83JFO0zI0dRtKWVm/RMUz8X6RurK9nt5AgMju/GcpKUaGAqHPGJDN3lAPaCX5vBaR1ou7w
VEbL2TDS8NEwPYpOH8x2c/LmZlkkUPLqszIpyu9z8HYcSYRccj8YJNyaEbZhvNpD95Ed7aic+kKh
FzUovI0XRpJ5Hj8F+Ae8yOqSXCtgsh9/vshREhDKlQfh2aiuGkJ1qVG4bM5NF94R0FQ6mly6I3ZV
hWPtrfL7wYUqAE7B9OxPebKUWfaj0R1kT0WPAEbpXqc/ABNidHm2BToE6iSMDNRY9eDHPqAEJ/gm
eyOPwr8qEp4Pq64Oqid0n/HfPFHc34V4NxyY71Hir740/J0ObHA2J9W5JUlKa6EwOemXWVRjpCga
Z+N5AQl8Vz7XJaUlb4LZjKjc4E6MjFmL5goou5/73ZW7dXHDii29EXuiMuEKXDbiz/ur7r+ACrEX
obku8fVMhdRJ5SS2EspZwiEVeeL5CH6+cjh/ahAdPZklUDWsfOo/UceBXgeDTl+LXmmfK4cZD87b
DVIfPv5HTV67tnap347Ux74jNf/2vQZsBHikH2KbpuUb8OIwMsptxzLPRuI8PUD4Mw+NqsVh/QyA
qUgm6JoQunaGxworxZwDBGuWhpBcPxJxZCoRkZaUyki7Bkwdny87flCLByvMf8/NLtte18j1MJOm
5yTGQC2i3m7SstqiDbZ3/E4MIFa+eN7iIaLx8mlpG5X+EgEbPXLNG1FCOvciTjjdbBWu33bxD5IC
fcQvy6DUmynY35AOHhaplr5FV5aSIc2zyV2keHyq33pQS9L1A5wWVCnATZbXcFfw0JuBKu3f9fu+
wbHUlYHkCTl3SiQSu3Edt1d0xfndvkT0eMiwKU7ZVTmzz8LYSb/19ZxtupV0dg4+S1ocvy6ZB3zI
LES7BWq+f3zqHgowS7cyC5unVeyngkBZmw1ywkOlyH9nA8OExkY5ZKbgJWplLFyH9pVdZUKx3COK
WpPEPZzNKV09rCf0eepoEBDQJmv37c1LtoRF/f9Qrg2vP+AXe+AZJqIkakdkUgjuYtkA0N1ifbns
GoU/LA2FzyPcPwy8wa6GoRFo3yGIF6vBsD3LLFtewzTuePiYMrS7hvPiFPx68cTJAhkjN7o1FpdW
x4HyikkP/cwcte39XMVpd29FQKIBfhOKyS3+HxHXJ/MNrG0wUQ0bNVwhU4sCFx3KG/KKApfRnAuN
kNjvF+rIUo1MyoooaKqzRry/3q4TQGPDcePfVamno51JIsgFlH7gQrkr/8R6DmeEWuhXjh4FK+3o
gP9YMkKP/w/T/fDYvmxB2ZHJgANCxw22YiyuyNYo0LpAgo6OpV/BMMymYCYvWlkhdPRLs68MgEHP
unIHj7sebqXOZEVLY9dyCmBZ1+X+2mS1DUILJDP6RxGK9rV5YMdkgTNi9D36CRKorq7kiDyMtmhp
VKzauVvuWOMgvMFrGl33gdJyk/u9E8yUYIbHv9Xm04BeQK0TeubbzdPrmqjmD7nUgTwHB9r7nfNo
4ncnXvXEVx1rtWclWCRdxU5n1SB+pOW08uY7ykyxOlUEQ4gGRFgVZWN2O5xSa382VPJsGm6hhRke
rf4VR0C60nxGTiKfq27aocxbp6qiL2nxVgva0sSiFDAQ2SuweduoR/uPy1v1Q8btvdaLTOAC583t
+Ye7pt1XiZqOTdXmwhHZ6Rfx/fm1BfyESSH3FlgsMiojmM6h26bR4oRYRROjR+XNa8Dhmxhl5TWw
03o2IDmCrCcQORpAJwMzNFzIgjXn7EKoV2YOAL+xRpsQLtQgrc5NySKwgb4sg69p4DExgZHHKW3N
w2yLMUMWwhEoaGZ4XxRgwXQurchyMXlyzOZfxQPxpAuIUncIDvDEKODjK7L5tQNNN6QtNaMujuWX
WeFBCnNp56bUt/kLGI1fOtzxL8498pp/ewJvypyRSXwEiNHjiQklQsZwcUBmMQsnXuIEdrNnT+b+
UujOOdSb1CsVyHDvj5Z8QU5wENqRR/0C0lUdfCo54Vc2YLotPFEdJNSz460/VNDzO2m4LcyOOAU8
2T3G9zRz8dTRNIZPg7l+xMkiEHkrfaTCQ2Bq+6+knqFIhfmxhEejNxWM1NSk7V8pnGlZorPQli35
ryLeOkU/k+n/1WuCDy6l6tz9i56VCCdrEkFLeNbqXPIZ5JKDPdhSurIPP3AZiTRtKLalyeLPGU95
Ok5aU+iKPuDDMcMOcIE1+xGXpLtLI4he0DE8jNyWSpG8jsePzvBOef8ueXDqH4rYRDtAgf3Fb61C
kxq1ia5XPMnN/Dkp5taRk5XboVphud5X6W8Vw1QYCtoDWPvEo8l6qapQj+XYxc+DthMbRJIQ34uv
Mj+TVjcAvmrDa5YfLY89rg2dOTMXNSjaxxM5CzOGC+MQyT3yKfY8l2Y8U5/uAEpVaJS/JjYvI5O0
nA2eHW3vxa6QtFWX2PT3oI02NB+kGuYda9ayskTlj5YB58qS2X1ea2uXnCbyTmE/GwU+pIjsof5g
RYMv1a2ZCGMZeJC7QB0PbXMfCV6I18x/szJJu+VJoE8EAwiFHhAEb80pOhpHOe2i+eONMjJi2Ata
+lAEOwL6twQ4CbO0OE2YmuTAFPUrJqs29LE0q5UcX3J2byy4qKUFUI1hikESrEirfQcifDbG2zJb
G9BLVIt6e7Vk/eAoOXsSVoDk6wNfLr3qadyPWc7usy8hcMrLI++rsWIhYFWrnOVIKlG3zgmIHYtv
ftse2ASM/2ToNha9ZikS1v2t8U+FsvYwKowgWjfB3zlObfupZ6vPPyxu2SQQW++zVtghp8xY1dMf
O7VufZ0UEPzqkYYo5S9oCVr9r4+44v3sI4XTvvUehQ9a9q6Dx+/tW5kd68c3kIjV7H8+e/z/Bszr
AsuJ3+TS7Bq5VEzQ+FqHGOXgcTqfq5WE7XWDFXntWb+RRkUgLn9P6PimA3iTEbtN3aQLK2VNbybh
bNMFL7NuJvjalXrPD6LiOEM119/YdLu141p7HrFA6vMur+NAEMlDJUtL/br4W3/BpOTFQwRl+p9K
DqKGxVX/IX92fVqs6yd4+FO4LDGlPtChXKvWsALWAYjoKkVWLkdE4DmwAROzYU85x+6rLgV/vkZP
xwLxND6czrMZiXeM8RRPLliOmmUCvEYOgLQp3QVLqiBDQQH6lq/DCJXG/1nSulqF1pp98c/denEs
lKBAHOwR9zRqKNAppyWKLQRgf20vfetGN9b2aamJFv8XrO30LlqNtoEKfIsq0KG2/KcgsWO319q+
pwWNgsvJ2WGnUZ4gVZ+VUc85jRNZS0osstUNMrJR/GF1VNoQeLBDevBBuvLqvccYwB3wTD1frIgR
4Q+9hHu+uR2zG4tvBfAdeRsghQ1vrIYFyElWKAo+SxN1LMOYyT+G5bWl8uWIaBanveNVcIuLJw/a
IbKCDWbIsMhmbUSUHyIqQeBtM5BWzhGgmsIMNKodmC9t7rXKjNR/FSBuktSrmCC9WH592Ztk+9oN
HXIuKz9AYTo8MGCsN71dXyQU/zbZ53GIeKKp/DMAAJHhr+mAPsVq+TD1YwFD/BCp9JBK+QFo+bqW
bBPK5Pwqi96jZ2Z+i1+s+kheIvRBnNDt8UDOYLB57xrjWxR2fKjhk/Tl1ojArz5UJBZ0e9a7X6H8
dgGxKBMS4NlkQD9fm2mg4T3g9cg+N79jsiRaDuD4OI7TIHx+9N22TM/MC8m67mTmWWdcfgTGwGfY
nQ/2Z6Wa1FsS+quX0yBfZtCkgmdm4DkQOyO/OfMzjnclx39QJoaENqHR5mXgynjcuLL4f0qs6bMT
s5ACIAMKkcFW0L7DG4OLeuMUuL38No96aLig0Y7Hf74CkehfbVM/HKpdZtLoeo96sBCUkrScQpbO
aSeDOq2mzbf+hXJFLY1sCNRsdO6voE9rAruzY9i3FuFDeEwm3rtUKPSeBsb5/A8QwOUa2lL/+/jn
43YPhkfv3Diy/3aTN/5FSk68NTp3rvtD5HCHHqnkL9FvNsc1nryMGz276tp/ddpNMuwJ3n2588vn
ERZnKBe8l+QUkRMWJumN+xfae9XYHi1K/IOuceFw6kJ9WXIopZx/OmFm2NnRjUhl2j+3zRLOvHgj
SWoV2kTaGP8aBeQq4GG4xVhIMVEkD0fAg1whahNoAz1eRmhUBjRH7HkQfw8yJ5FemvUJSC/q2k62
g8JC6r8p2jF51+ZCTP97uwSIYdnd8pwF90sEUazppeQrWtvvwHj+kLCnarTfiKq0nJSPbj3srS3Y
IggC3FvH8tcLbFMmekm9tsIWV2cbBzbC+vLrK6h6RO5bwcDliXxJaNQ64TGYMz0zc4ItZVEFftl5
9Y6gtyll3UfLMx/bk6hEF71mIETcZkJ/OvJTAK0zQ6j5DQHlSPj501FJyNa+gPj3Fc33gOb2cnFm
rPKtfCbg5stuLm2Stn2+WljEwTLGEJizx57qHB690ojLVkh6Se5Zr4e4BXhJjIdk1/DujR47iAxN
/TXnkeb2EZHYMxC8bMibemDuvnpxd2ONR47GMOYAgIH8FYpncyLBF/5lAxTcH6ZmHjRQ63l/C01d
QiCLIPFeAQQ0twGRU/mp8A6hYie+FzeQMy8lvXR368aX5wV76VaeC4ANaFS4BUJtPfu6Jh7mO22d
pJ8L0guWFLFbJRW03Av9cPxxcPEQhRkQlCRxaqnWk05wT9udJuwUTr+SjgloW46wK0M5rmF//HPF
VIboooV+9sEHP2JBFpASTuWzn8KPvn1TZ7mG3oKssBffTev+qGlEFoq3mLLfYMIS63jYkij8mdjh
H+zy7JB7XNRxWie+K2+KHBgXMNHhOwQnS87A6ORGLkRWXPaMqWmYqwwvLmH6VhBXwRonp+JpkP5u
vLRGIZ2xuRJhY017xu5UXwF/xkokRpywPZJ9bj2tzxGyawjg40ekMKEDE+EmNlh2y+BFIrs4IoKX
vQtHTl7T1j81pRcKCzwjomoymItel45zdPFc3FhHA4qKgPjCQirPlfNDWpuyAF3TqsTkmXtNy4m8
XM/bzOuMQA9nRk8wEHx2WrcxCMQKGQMQlG0z4MyZ0CTOpvLcNWj/UAozEX5D+a44ZDXJBQopFF0/
+A337EQlSUoQ1AtOf/YSiSnifPCwkeHAFLYADV7IyKm/24ZtLcFUkNMUD+Wwd62gzN8aWGrTi2WX
2Rv6PQ5f6mU3uje9YUsrGTavQLEFAenok5Y3o1H/BzheXftOwLwStAzf9NDOf5TARXxDGeWJxzBY
DkCQvM97alqkltJDs2j2eXk/mhSP2OMp0HYkikv0hxG/McIYuk8udgI5bMaLJpa6sEWxboGwW4P6
j/eRAT11qZPduzGyaVlwU4lSGOM1m+T6/Q6jNunUu2cUdYNjjh9kPHUg3IfQKbwRvG8o+Z2FwJT5
FizNm7RMD7OHUiyxxmis8rpmXsKgY1WfN6Fr8dpKDJrxdJqpirLfBM+E0X5MJGFupJ0pMFE+F/zd
3Bev42F17H4UF7ndZ4c0uLgH2xikZyEiqo+/gmUYWq34SmpMQc8oBOFJWqjPEGmeA3LNRD/tDDXH
r0WO3dk4f6GEEhtRnPdzPhxjigSV1Ds9zdqUPQ6+Z/Qc5k/ntircVGc1OlTif5q+7FAXsWxSPYyO
x22/mQ2Ik4HtWq8lUrt7a+zQwWZcGlqwESRRuGjG0KTDKptWdJ3hmqXLhS0VdyjGcYNL47zDYJLi
mTz7J8UVeMKd4KK086rs3RUs1UVC0tH14xKFj/nsEhx4J1Hmh1iYTsEB05xWzjE0JSdB/NWtZFN8
hLocARnEmwxaJ7hBouzupXsvmWa6bIs/uLrWdF2QWGdR2lax2dCyVexujgGI05meN1h3CJx1ETmf
djZ3gru/SaCrVrtyEauLxImpOksOt4a43Fr2wH4yZmYNy9k+L4lUNSMQS001LBiNpIxHhvHEqIfc
zhWa16318jAJJlmSmtXQebsKqVhR/CW58fezeALAvCgqw0VtJtSz664ibeHUMwUBt0rlLN/EvBhh
TmJ//pVUiZoPTmBa/lVFGtmkn2/HcPVBZnnKVOTuuRL4eMglTfl3jiVygKhH87iIb7r9kI+FU76l
HfpC2w46BtT5BQR2wQwYtXvQ+uxiJ87nC/pKYdxptKGWtWgzGfxBoNQX//ZHzntsJaV5NFQBYoNK
cEkOdnXJ9WwaTFkZbJeTlCR0YK6HcDqGb3ENT06fy9j1wFrTbisVRevv75Rqk9Fzoj3Ce+a1cAW3
jENN3oV2WHfwHLC18A1hdu+jxKP97N3JGerrvymGdkBZbBbZ/ZnAIMKaTnIP0hsqH5gRBGQ2raiw
cUDoRDbM1kdaEe4ZR0mPuIt3+sbC+sid4jWCPKgZhY6LuoO4bUQ+CpXeAiQwsmAVUMsL0tymTnOx
VFTMXkHVkBd6bq7TGoGn10L7/A7H84jJDZYR8ZeCqpZa3OIwwyvehu/rhvazaLIFIuUxqraWq6/r
N9J6rPaUy4qGnQ+tiXTpuFtD/BUqCQ+wx1r43xvsSnxfFOIBx4iF8GD2v145+i0VgvD6hz37Jf0a
mxwFkPNUN0gHAlaEuOBlbroMAZfCERNfIw8kq5WvQLBGc4c3eTG30IYbIen6tUhQTJti9S0nOXpB
pO/jvYmyLiBKmGWWPMZJeKBkUjOOMOLbYrh1gbOEWkKk3jxAwHRTNmmhirTBlrzznm7ouh0eRoQd
aeMl6G3OB6D3AmrILmFnH45DU514xUyIArK0nocJSt84PEzw/aigYRalgBQxS7pGOlejLdjBtBCH
bie0Ul8lVdGMnrvlUQ1Izbk6qf/dV7RRMESVwDurNsGiT6NEndzHjDnJEUh/Eb/Ys4QfCjo+xIvg
+br85veSC7f2zTkcUalTQZ11J7irUsA2OqSn08xxDny26eQGDf1dz+xjIGEpISC5IBmv+QTiCPzN
u2+brC9DUlLO3tP6Z5jECFfz3RovCfR47Ju2s43V8oUGV7wmJAnEmJ7HeMmu+y922znjwk82973L
+fCe/fWpy/9q/CKgzgaV81Tv6QEXWZuBlOm1vWLw4O5XJUMx8Op4BdFwBqW5VEnYbRLfinMGWp0m
FVZtK2HZISsjs4SrRVvn/fWBDwNc/BLasA9NKtKDpAjnuMkHe7vh9YfyanqBaPGB+hrIjk967NSn
AFGWYOzyWem07gVEEeQJsyqWc4HxrT+IQLGQkGPA6zfjayCWlVWDfq2wt21G+bjP4UoDnl7QZcr/
XJ6k6rHFkCXcsmbpJr/IUGAQiFw4Vz07jKVMCqyfVbbhkTdJWbaQkmbpaD1cWWvAhTHxQKeWdb8k
Z9/Q2r8cZscoCgIQEEnE80jwje6yyyBr/D/8EZT5KJ/dE2i8yaOtLOjauLZzSjlt8kYWwK2ZbmvP
bS7HG8/SEu9kpy7fYJSY2568lCMELMVX6WxLN2dr2aXThYU6fRxskH22ycI2yqE22TAm+NGvQwLA
jPlp9l4si52Q2KL8jkqCOJzABtg5KI1S32JVumhfDsoUVmMHT4F52ImFN/vTKVxhfsVW1GoYvghC
qJeSnPamYEGLlX1eNoP2eQMsWOB0uvfDjQON6CaJUSXKeB3Sbgc1ZLy0o7aOXdEU648+uAeD/tJG
Gj+an0nGMZpcTmXEE8T1dl9MwXfI6snDKnacaMPrfiQt+AbEzoa57/5RZxuD+OM4OgVzJMz66jCy
HQIhoEEvm3laMer53NC5gaGK+31VYKgIYZar7gjzkFwS88cu6tc1bNnXd4guiorCborjKG+PbKvw
n388kFQWr3l1rO0v9Th9HYSnloXgnxtau8wJaeoSlbWt6Ako/WOIC3zQZ08bk4uuE5Yx48NPAx2i
iOrdsGRBzmpWfBAAsQb/7w9L2QU83rA0/HsTmBD7sL60TanN9BqPhizf65+7jF2AmIksJ1M/kJ7c
F0Ba+jb6DEzSVkXr27XEviRmfVxWYUsPYl0pj0DTP00Iz4DvHODH7w7LAzUMaXHuwbHtGF5Lif6Q
4ImblyESSC7vREyu8Okh8jnQSwmDMuRCKNr5ba/Qx/rMLrqE/thwR/g0NShjBKQEqTrVUkiMkmBJ
ACriSE0WFHRpcKMYBYuUnT+ly59qo328qBFP4oLakb7UW5B4sPX932OLp2rVZLOw3kHvD3CSwwsM
MTcanAjaLFlSwi9p/AWWzsClCfjOn5v5/lkmmrMnlV2YT6oDnJxJmEwLjA/skTGxzHgP2mnWWbDa
iqfae+9A0Et4Oxsfd0aBYsYnvDoyDAnTtm8PTFOrwFixhqnwY7sUfTrzmPtzgb3JM6ksOAckRmWK
JUWM6rLDjKRtNxVmgR0bir2fWqXC34YnebmivjJ5p51wgAju3s+qXWbAMPk5cdFa+VtJDpj2r86m
0+D8tV/E+mye3kqt67693z8knPg+TwGrPR9YnVyoe9PHFbLTly3G+B80tuYeUiEbpUZof+IrP5gP
nA5d4JfPqwkQeEdHIZeGOhERSWXIFTrbRdseLXVpCf4NVOamjKzoJPQuYNb8Eq7IqO6zs7vvHHF1
pVSIr1tzKa8aXqM2no2OdWrYy2KWgWV8bT6e4iaP5FM02FHigNO1zghWlKw65NJ/0funkyD/7+rv
gfmX9I7xGsbT+kCGJToenEnSR3LwbWQLvHcjpi619YH/rdzvsmR6anqsVKfJuxi0GU68cmNyV3J0
iWD7r6NAvAvlcvOkkBLqZrNc+UsfZ2+zQHWTLovT2gsIw/dOhbYNzmt+yNfNXyFo/BB/p6tCiM1R
ZrPTcf5uWN/gijBTSQnFxK3NtMzFxzy6vDhTgSruozm1FqTUC8ZgsMDNsg1nyax7/Vle+KRtQUG0
Nd7y3VuBLx9pTWRFDHhNbOgHQ9z44U6d5DdaM+S3UmL8NML/3UiqkoT6Vzr+5H8BAwF9qOi82qsR
GMlovi2geKQW8TCHwoxVsIc10DgDRma5f+QUfBfVMHxY2QWvlfbHLWYYy24axMTl/Do9PLsV/QZx
NI5Qot3XCuW1zU1GL4jSxHFwhHKBuD9fj3j+tnBe3zyaM54FGbcyrufSeBIt9Iyv2ykTzMDET6ex
/fNrCODF9NhCO9OVhARZQSVD6FKIqj715tkrAFb7ATYzihMn4slwWy9nhR5uG4NXz4yfWfT8tzep
BrFBI8zsiGXMnI7wV/YfRImIqH1Eomka/w4o9kTNPQT/p0Z96V9Fk7c5Q4nNdRPl2JSM2g9ghU7W
n6IIL5T+Ej8sQvtBHg08NK+EyBQ7JkC0C1hsRJfepQkOQnb3s2D0wZ3Uo5WS0YpT4AvT+XZrQvXT
+X5uyUfn1jbq9SeOX5mQrx65i6W9XeDC0omAk3iNJ/JLSXclt+ni2lxm/qvXlxiUcNUgCZJBXiHA
NzCyK5mwGtySaUnalOlFYqyAUum1uL/29SruTNDqt6bXRZOQNJLtUiP7LSHn0vyAZKQHaOJNeRNL
wxsf5vzLZdYMOb4PAHSBG48wYXj3Pk2tJVmG1U7rZQriON4rKsC9njx3Yrjt5TDTt/fKBfQdL/dx
g5WI2GifFny6m2lUzuX5ldOKVoFQtrsSgqOEasq5LVBw1xeESy+doXmJj/T6p77aEVgiRboXYqYK
467ViM1YTa6VVLlbIKV4Z3BrMfi+JAILTPJTy3Zp5GBxMtadLYZtn+UMVjFES9xp1I0us6We4NuU
hVqgmy5AXzOOU9bZ1NGoPksVAAKqkixgGRNATzdHjc4BGciEg6Yx4tXDqasywvDJer+onYDB2Fr1
9iD/R/Kg+/QYunavPvYaN8+44JmbdEhCuqgrQXkaCi2idc62Cm0I5ofGJs4/l6McTUunyiFnD25W
ZMNC008Q87VGQZkw2ZCtDxw7yb6yKrpWKMWgdkNoFhWMCnvUxBYh7ndCoSWDUSgnYNzjSosv05PG
G4OK18Rzbezjxat/PUrVW/JpIRxgsqQe53X63PXVYYkmOK7MKhPPLmhgSWfisWLb9y0A3heBosu3
Wh+HlWSrHo+fC5xd0gLrQZppBoPk/d73/9yzkKHzZ2mU798nfDLuiBPhipDXQjifCjoq1MuWhRUG
X/e65Sh+/HWInMkhkk7HdGuix+8xsEBV3hZDIhGFibc/AQuHE2CDCQwhzviRZBlvbaxi7oVyzkRZ
PPdv/rFUNu2teJaULuO0GxNFbhi9tN1BQCl/k4JvI6D8Dw9AKas6IsiehrtwlXbTjf2JlznRoL9x
ipm+Wnh6ckoX8uGu95nHSV6nXcGBBONJ0LOaJ+qLptcqibH+x6QjIkzYA+42CLv4ZbtBct6od+eQ
byNdC9L+90nnt461hCusAYjFGt2Xw9t4CPPo+QDvkpORBZ+MstY9qxmQEUHjQdA+/9Q3trWOVypn
0lxbBbqTW+dKJkBgNMLO0vCuSgQJLzun7s3yW6S74bOfKWamQGPum+Es0QP1rdJiB/cmQIhzyvmo
YY0J4r9kBDBUIbfN/Wa5kFSrVX9aUkpYta+Db0JAQp7sKb6EJBkqJ0315vkCqiVCl6Td6h7wF/sW
0+TDxY05wmqOuSDNHnz2HdXFrZrsAR0Bccnj8cwd0anIBKMfucOoj5L12tX7H8STIGR66wxS1FOy
NldltGN/HNfsPISIZfeanSVWdo4C/qg1XTVnbizI96Bc3JM2vd3mVw9GGYliBQ++Z5xOIGbqTi99
gKBRr1bDoxlDeDZmCeginshw4SrhrJz8mUzhN1VcUZMkhCC1+kUtiKSg0gp/BaLPKlBTUIXkriSu
O1uifPVeSoyaOhuz2lpiOFl8kJodpzuO7dojzEzsI2l2hQYyjRXaSlmBOTbDLyYT3tb4jlxc+FkB
QaYBbq/hmpx4F4TfEb3QyXj8/1jBhNLS2MTPzmLQIanTF6YYi0l7Xids0Hc4JNRzJZ3NUAzkgPHT
E0d6gbFPlAORnXucquvjeR3wYN0bvBvdoGEg+gmaAKib5ev4seztB+PmEvc5BO5E59kPPuzk/7B2
RIIxIDxewE//Pe9ABSo6Wl8Oe3Y3AawCJZdoL0ah9Dl3EuZXESvBcviX+lpo3qzPkW1PYP+FY28l
yB4qmBcgqFy8oON87gQlxOtcxX5c/jCtAQnFkJSNB6H2g3zZgBkAyKD6vvN0LWg1WWEY/lJpBGeA
Zb1W0LbIimqr3+UB3aXkjnsnOlHgp9W/zQf9clC9E4jJf2q5D4g9b0jISu0kyaUDYnTr+W+bEKS1
FLUmPhYK8baasctFVK2XaRSzG2HuaI8yO7Xc/ViyIFQgckFIzS8KaUu3GqCnbymLlo3HbQ/AwEUk
2WCLr/75I8uAEJ7/JV4gPgCYeJ0Id0/iUReEF/CnRFB7pUjrBkHofIGCJdTWi2rVVQYH7Kj97fMd
gB8ftmkBpgQGVE1A+3NN9tPXYI5bI1JOlfSzTalVoilegh1pnOQCB8bz0WOP5APP7/7bVcncG8qE
T/FiodRuS9XqeeMO77iM6fTaAqg/ZremgYOzOOLZbHlszWz5fTi6JuKdCnwSuXSWu66/kSpdXFw9
NmZrzl3KE01brHsZ6b8q0P6z/ug51t6S3sRxXn/zarB9bGlB3LXxUfcVo6S3rxd8Kvz9j2zeXO6l
IPv5WDov0WC3ARu+Aar+O4d/wROtOS0QfICybIJBVZ2N5Ltvmq57a7Zg/auPENYalSToALrIynW5
xa2CJoUU1VkX5Zio4T23YracS+8b1bd20miR4ql0y8ejW5+AHEviLrgYmn2GG1U6hoPbqFOojHXy
6IdP69ILEUV0pdhIAKaQSpF2K6gFOcWhK3viOpPqJGu4pm7S2s9sMnp7sTMrw6xCWxpYGLY4XzAG
/SaXjGC3GA1FwID0oM4IY/h3awGvYLMHO7G7T5SUOLap36Nh3Jh0g8YyY15Af1KJWtUgU3aWWAg6
Bt73FLJuP8WAzw72aIHhbxgWQkHeZ7n/re4nQQJDsvgqOeSJCmg6lAS44iZY1+0sJdNnCFKChJlY
lrlFUDW+I0JdX0w98aorcTkjsO1jbrNmEPjz2TRHTUEGX57diXuFcKa91e+E5UUY8g43MQ4nJkMb
EeMnPaK3l8KBfFusoKOZHVLm/F2Y9u6JvR/0e9J9YelniIfxTsGHDKXIF5MnIqC1f6/b2H8jyWBW
ksaP1dFLParymoin2bITZgILFoBAbgOr3ySV1aKynjFohwtcoog/p5foEoC+8HYrZn2QrvrJp7tG
w6i3NKhYWtcGozW1fpB7WkM1nVDLHpzj456lakrMI3L6Ok8ThwzlRuBE2WY4+jNTpbRGjYxJVxs9
dNM1iJhWqnb4eSCfU43GuMKXNxlx094mxp0fBz8YCOPiALPx6vrB1DF1ihYnD2jcw1FhYLdcGpQS
sfV1bKLc99L7MyM7eAiwvKCqHm5vPoGVvw2GZdKohxaSp2dMl++O+pY0yODjJO1mVuuhRZgk4zfX
E9/CtmRZ2GF6BakYGiPaGLlLdB1ONdtLMK3fEUgPowBt7ln8JVDrlPMrzCqYgpLsKG1eqkb/kV3o
3KSR+dFeGx5m5HkqN/xgUq9hkVTBt5pTaVpZqzYwUqYqwAXa30q/Ri06O1wkTHwO8nJJs4arC/YX
evkLD3UmYzPodOlBosJAPG/8IIS+fdeOBaVbWo0fvJeCtk+y4oC3PdOmFdJzav1nRMn/Gpfsffj/
0cxd0K/c8sGeorf6yQBG3XYlOb3b79gzPlgWsG+aA3a/w20NY2PHYZBc+f/SQtBy9x7WpaSN7Sdh
ycZM40PNbl3zr036jKRtxmC5C8yNmZFsF9kba5ptGwkjBT7GqYw2C51tyv+Nrhu4hedkRndqL9Er
jpW3IGTOHs8BXZzmtivCHdkFDT+j2ddJ5qxdNxI3SUrJhUh97mZpgOESgEgJhnqqx0NH0HB0LTE5
n8HdO2IYrcgbBysZZIu1VITcF+3UniyesZqCmqya1TglCPZ3W3WsV4oD9u9wT9BuJ+w34X/4myQP
sy5QGm9pIliD4OoAPoKyl/njwdKpi9wnbKHo0qYheVLqNWEpD9fvXpPMvECR1ntXG30/c2AEM5x7
z39nDClM9Jn20ggVPFpOIqDERrhjStJpmInzeneDUC+ZaFqiO5HzgBhf4EWYOZhhxVMKeZ9arFL2
bXYL1b1qZsDDrOZ8C2E44cxsVRpyTQxwUHwzCbd0iWz+joeQWTFxAtouyTc2WvIYCsYVxi9PD06o
I6LSZcDVJveScCtrDaGkVo+xGgkdyyuS/3KqtBJBm1poAH+NzX6L+udrYzpDMacKWoj+vdpfEZKD
Cawck2O7Wof+0tug4b6lYxBXmFgBgCHRA943Tz9Sz/wXiN8xolYcdFV521GrT/AR688IVz9wTiGY
tFNDa+BUER5UVC2m9m1mcLWYyEj/Xn6uoio6G37LDXF53yeNBgKVULeBaAihW3J+C57gsVzgU4Wr
0xwldNJMwBfHri14cQT+7Iq8tVS2ReH+B7ypuJeaEj/W5d2CWyr1UvVFmty1fTC81qrJBGGQUSH7
bdSUsBtelTZ2KgltRmnSJthua7os+0qfO4AgJ+RYZwlAVTMwk6qP5yozOTGf+qOuhFZLE9/Uwc7y
Gh+kPpwV9jbHlk6BWDOMplOH3J+3h7J/UqqEIhA1SFznKvpw3tzUrUHC1kPs58fWpHugnm+aatrv
8LRzQ53IBWj067HPpqmagIq3MkN20tCX57c+UYMeeoevKRIUI/h4GzHljBHlwIPq3kPE70XEyKte
UIdgVYaoR5wWhPG37tUNQbpmf+9QRsT5D7qOTjLfJX9SvOjLg9uI3JMIXiub40BUt5hM9lvcqFsQ
fK1wcZ6GxhFE/nQBREckM47U8YhK/Mh+sPxl2GZ53RVXflNFKvQZVK4WKD54aFdZ49X8EvZNgX80
8/Snk1TmyQoSopmmEXBKbr1vcFZNofM3V5j/+su7tFgmMHbJ22Pz5mvmIYKg6qZhilzUb/QvT1D3
qMXGaD+8AL+OeELl2Yh1IocGJri3LlcJjxkwEtfG9PlB80il3N4U7l5BdsjA7L+XBqRA2KrFzL4N
QXm43sbIjRJ5Yq9MGYKOmkoie/2NMnhSyvjuHu93g0vpO+F2+6epQeiCCxERHwR7E9XepTDkKkT2
RshEcel/Ge44GJ4CozPZyXC+zkFXfgo8bDe89uQGnSY6irXFfh2Zcbmxl7IN3zSyWZAQA/D2+fz+
IMjkPEIaxPuslKY2WjvaraLBzs3XDP+tpwB3fQ3P6pnwExjIA7K9fQ4lKqjeZuU8n7IMIFvX/++z
pDyGfhEud6wVmAIcK/mkLTA5BUQZpE1uhwwCGZ2KnlZ388Dm4vbFQTGf1M3Kjx/dx3AbOm+GLvzQ
gOpZHnUgcAD137vh3aQFNwV2LaoLyWVBVcZ3lOX2LLej0KMTXq7meMWIpANvW/46db/vHI6E+vgz
9jnT6grHOasvnvxCIV6J+FpIhhHdBres3b/QB2wmKJScpqQz475hXo91ia7vHKybGtkCWtbYKvd9
4ANNzgFNTcXR/IGOXo0+OtOIvyXBtH/MzY1Gy/PuQDsrt+fAtSpmFDDgfKlzyE4ohmPB/uA/MJMU
5Y2odb8cGV3XCDYCzNHQqlUWdKFjljoyRqGrghv86PerDUz4mkYZB9lsa6K4F1IS/llH1VbGBqmZ
98jR5U5lbRe2W3tlADbArH1hp5pW3p1GQctOSIdVn1PnIE5LTRWVU6QBBHzRMlgxSlsAC5sduHcP
FO3Lf7LUTS8qTJrCUenkkiQ/JlnGnuEA2Vep7v3YktDQFnZ/AY37MVWLz+14c0gsrXSnpVQaS4EU
2Fb2k1cNO9sOBXZVK+cgTn70E1/zMAkJHftVt7M3o0DIiKllwZJ77XkjX1G1zcoKebxGcW5JGEMC
3epLhS5iLWPdK5NzESGmSIO+Lf0zqF/aYeICA9h8QVLgtpSYLwA75gDS1Io/6oeeqJ6npvGfK97v
aBg1bzHVa9chuqvUYMIZfH0seQLECB+50dGTnCFvKpuOMjV2JiwwKwcih59dlO2e3peZ3S65+0OP
/7Bl7ualCLZXbvlGudIHFgL0g1g+84946KrJK3nq2zcsPiKPVcmI3QQXYzbLjrQ8ERXWBDrmmtF+
26xetfDMfinJ9ED6y29Ym/a9uBacJi7Q0iyJsKL8KaHvDS6iw71X33ZcoNdrN4/+nQVzzSXGoFLT
ka5zuDh3xpvsTd1bOy0awoMyIxNndkoQunKJHQrTuMhj2mnHqf10551pcIAy6TxLYsC6U4+fAQ3t
w1Jdkgp4vW5JrA4ymu1GSNb5nfRCkPeGVDE1ieaX/1ul8A+PGlk9yQ2/n8LySjYis+WnOXY2xSCZ
NaP8GZtOWaqY/KN46lQWWVPCNKmkOLDbx9INqAJ+Ne7az+yVo75O8Jk+f/T/H4g98CA4IM5N6P+w
t86+4CDnSQOXEl1Kx1GNIxFdFm6DiaAvEO4bSLEWd+sEKm+r24/dxX/DULdk5rwihHdjLeNhvn0k
Uc0wkOoovtInK6ZBHQYGfmMbWmgFNF5ih0Qoo1HkZooex+FCA8623YFQ3h9p6Wp9BjZniLLFpCjr
Fl/PY5HDLblQrhBCiGljStGT56gzj95s+G5sE+gdOKpPldp2ujLWrW/K3ek8UkESfRFLj/ovIJzZ
fySeDiGf7J0k5GEtjQVYTs/G58xsnEi8oFBYxjP6vESnJIPeo8l95rnoXKLYLMjUgcwHWDSXvbke
MPeuyVUosFLXog7QWTMnceF/ipUsK/ZzJbOAxwGcZLlIXmWq6SfDFvgLa/5ELFV0ZXs35t4J7xoP
lcMQbrfWbwRFrjp5UrBn/yMGCIy+TeraTljMo+eFq1RkChqQjc0OIyzxBRFKyrH+s9LZcU91W/XK
Bgz4QVmPTFh7q3D7zU+zAk4yCHBRwhLsI8dclQT5ZjWm/lpXuB3uZfmj2EVn2NO1NGRf+zZrVVP2
YTvziiyYXgRID8V7hzXwfAfSO1ozOFwhQyC063VmVRSeu016i3ogS02UogkigO4NBgpbfAp3aXNz
1SNkQF17dKI9PcO0pjrDCIZPCVag4yYWh7yO8LfXOA0u6s5ZupqWzJrkMVHyp/w6FhSIU5QDM+Vo
hZfgXyNmoKxxvWZFhFL7vuOx3SZLGe1flDMuiEkK7hvEL56rCUUDkksV30rbvwCNnOef4GHjZOoN
5yUjV9iRrirIcmuuojvIiB0BdiC4cKHtnBFdmXUE5x9XgoV1itJ2g+OtjJjG9kFRXPUm/OpiojuH
5wL/4VcE0UTswIbxCLWyQzRNhtDlzWKPFbjtXVpqeKBq+xUv0KCbi8IvozjJIirAhYherPtlHtlg
SnfLKFeLdqkdQxcaQJwAvxqlRkiIa+Zx+ZLoVetNcInnquQJo6a8C7O1oziLnWTgCNdE8G4bKIwo
1BhiK4PYXx3gsBC4r+Byv6VGAvYUWdM/ZGOBfSTTiIGVd3Ttr0M3UTmhEGHTnw22FUT1eAMas996
yXHvEw4Dubi16GVogV5bs26IfTF0m3j7JRPRlVJa7sMG7NVt7K7lO+lphpQxPnTm1H+ZF5QUQT0w
L0ImDi9jRtmmiF0hkS9Yj89+RrtnTUTWs8rEbIoTbKkyxPknfdq3o59WIl1b/p7puee1xxMMHpA8
YcC32E7rqmvebXJ4dfhEyxIEnVhj/RqzDvp4LM1K0jNYpQiG1xe1YsEMBJmpmSvWNFAf5/j6gGm2
VHg+YtuCPzkHXWq64hCoIkjimQQ7bTtbuVxIUmRjcaCP7T2BApESCi2KPvALXo7iIJfVcOw8DnH3
MmsfrSMn5DQhZwnoTc+y1FD9AVkf0tUiU99h3x7yK6vMz+RiWttLALY1TcNH3jr/opTwklvlSl1R
lROl5bhRlp3ht0ArofbTwWaTNGZRJRtR804lesIe8EFiiwI1BV/sJMOklYgyoLLjJJdt1OQEu4XX
Oqt5Z96B27moppAvdv7y3PWM1ek4tEdiDkCSGq3tElGZQyyQK6bkQgnPb5az6z+T9UcICeKpB2d2
jbkWmHQHCJfA2roW29fqe69oU98q5+hyoQ92+jmnnjWxUe5UsEQGTh8qjlNNzjk23ph0GNhxfQAB
zrGuaJhQnM5+CjabkeegcU54uUaWWHIF7hgriCG6mJzXq3ZHJlMphcZRYO5S0afHkM5J0ow7yzg0
+jtu3EM7S/f8Vf7K6ov42q17n/wtKwsRXpZQlzehkZTh9X+guiEP9t5dEkiyUlAN42bbsT9tgZIt
3kSrBuBb0fydNMbCYL77v8+oDQB1D/nz5eesir/64op9lDz60c0DG+R2zQMhbLeDxvxMIocGIQ+/
Ui9vDm7YEk1XaTpI1OhV0OPK3NztyxgipTBbbmnt4JcQ6KdnPdTNLHQPoJtdMju+Qp5GuOLrJ9tE
e3kgZFJ8nZai6YKTqvlIGyRHDKixdGtY85E9RqPe+rmYOuwEFO14X/1vruzJXVBvldEvj4QhxTCn
7DC8J68fSOHkKrPgq3U7dnPH4AZ0XuqQkoIolcNq4wKwQX3yKiSGrEMP4KijpLOTmQRiL7hl1h5F
M3RmaFaXgcQ4CmS+eG9HNhNYTl5+ZiOAsK8dtXbZUT++Dwd5whniQb+zC/7wHgnf3JYgDRqIdFAM
QhCV6qRy4Mz+YDvpNjXrNPBBjOW4F62nwull0KBReClarPZbW3sNrcR+4pfixxUt2r/Tjv2mOhiT
zNMQPeZGzzxhrK6zOllTO9zYP6tKbdWkF1JKdNWXAdnMnXjpPyC4F9PvlxKNKRUrtOF22m4oMFw4
cVYmYXeGZ1p50F43jL61noiwNTWLAAVNyLe+aH0SUd++ToxG4R/azaIARh2Wu1Dz1Om5V8gk4Jyy
tjSZTXRwdIJeEtazY96xnpFDE72Tlipm8gqIrHYFFJt07IHVE8h/DkEF/EPvmRQ6+X4Pzz1rW+DR
T4zg2GM8rJwwTxyBpWrZm4l/tB7Ou01NcuHlcXeYhC0qPM0DV0IYEgfHoouwznC0D4CeUzWUPigE
f+ZXpHBAz6Im/aFq/6Uhqg929gfHRzYZaLeNvYlVpTkNcHdsbYmrSmsIEB7Qod8G16YcG6BhzcRU
qLDTErDc/2+tS5O5VT8LlPCSxY0MVwPnMQSQ/3YhHB4mIQJhG63GGGhGw3a3GshxMQ8XEy6s5UMP
kfCXGawwx5cBi5lHPoEsV9GNbhuIacbxAGcw9+N2MsT1jqDIqtVrBA4thAis8Bh/7uaa30Njmxcy
dzXuqkwnFa4t34Hc8bhdcUnD/i9V+KXoJC5nT347jlY1BmRmu5MFwUQTLCbMFCv6vjfpu2nT6XBO
v3Yof/EB7dI5xlKuNi4vuUm6ykYASq942DJqX+6LFA9GrkJAk+C3fURgVOPykk8Z7lW5uQKlcUkl
yDYrrpUcH9+Mrq265GuFsRtW3H0xrNfRxd+mBmrj4It5Yhr6QX1o2ugBLP98IsmzIQxUwXauUGBN
lSUkcexcAnGTftMKJdNHmqD5bcZWEU2ERONhxBRUE7CALUqvD8xrLx+zfc/Zw7ed25KuWZuyuQgF
PaSeUPYmbZvgZmrxiib2PfKV0jf1mwFJITsR6/XQJDx1JCzfbrY8k4VOgD1llPitTwqh5/EQ1w2P
1pWg3Glv8mK3H8+hyqgR6QngUp7+oodr2lRthgSkagbVDthl/fFzliRHJVy6PLf6Sbqccd2sunMP
YILB6fVdu2Xev8eSdDq9C4DYDJB/F2aMIYp35UA780jsYIl8Igd0J1D1mAsbdygiuv0d9PC3QEzy
pjnWXpn6ygCXFp4BeMqEIWuqOFWzhhFoTUMZNADNKoailKjh6H2asMuH1jdJ6tYxEPH7ULTi1Myf
kxtkbGyTjxrCJrm/cd2c81+28JGkcpeOfJI9tNVLcJbUbxr9vXR1GXb9Ls9IjL4ZACcbaTBRTmGw
6XhVPHd4+mZBcPkvjjJ6M/W83BqdEyR8OfArEvRiQ0iF0IWmuSrJNDLWmMkmDqZtTESwGFgtMZdo
6ARUHvh9BccWJ+iHRcAN5BduKvchGNA+tLLDJ9Nz5x6244jHFlCBW1ZnOH4EgaNLjc1b3mYEI2yv
7FbWVvY4pxZHZ+/+vV2jd/Ry432TMQi71lzWrdFmzYIY5WyUDRg3wZ07rAnt2luvluSWfuz81hRs
cu9FcCs7xSajp0ebJHcvHAm8I707iF1C3/YDVevokrpByI52DbzEZ5Qt/bK9iN0IpLzCdHteeUsC
ooRxpOsk06T1G/5on+wgBYFt8JXpV46VrNhlFgBZOYLyS6RNQPXg4TaXQLNNJsDbV9bR9Sr+qtxU
ZHn/PRNNOpqMlSXYH+2GCCuivSZ2BTBL/8Flwoir/U2zC2LNaIi6osqSfHkia2O83XeMMSBq0ahs
QWxGVZjOAsYofW9E4yW9TE3mW2Neu3W+1FDlSnPQKEchKBQIZ6Fzc5KWX0JsyM6StuwZqUg170DB
Hr1Uz8ijPeeuZRxD8Pa7ZXRGNgq8SbUu6oyyfw2VAT2rRY6eJ2PIIu8K8RUAJzGHi9ZWnCa6hTpV
crc5+3PeOizp2GqBLl30GA8Zj9FdEd51TjGEi6SyAOTqCsaciYkeYBhALf1es3dDu8yZaK+zq4BC
iPFitHnWcfNfWZ0AjxTWlRLz123qx8+x4OnOneQQ71YeB6YN8LWvf+JpIBGbkPPCX7HEQfeAqCmv
mCdCdcaaB+Yon4zP0wi89dSFN0vVGdXpreooJ91qFjcNL5y/j3T9XqE0IvIYeHtiub2OsnW6nS8a
KirnmfQY6704ubFm0KluHNWmqcznIiqt5gMZL6UHtLbPRNkfVr6OUzxegfRfoInAQYDu3O4K/4rz
C2USrYy6WwLlrX610xniyXND9u7usQtLH4WWMM1XdgMJF1QRiyD3eBDezTe6TcYynVKIG49QPab1
amzkMlzOz8LZirQSfXpltHBZ94zYmSWbWVX+Ddop8FOeVYhazW+rRJlLuIXcW8EuCOzAA0UfFio+
nMBY84qq4G8Uy1RL2SMPT+qTzmlcRHWwQLzMZAI93jIHzev+cq7/qf1VQKLIvTx/UPSyFt0zT5Yb
ymjFA/Pl+Swpqvd2pfMOLZ2r0f6Mp3eskSTJ50ZF0/v7673SiT2ytfMVJVraQp0N4Ly/5OhMma+p
JuACxzsW/6G/BvlFuO+bQwDaKF90lIWDaigKLOSu6Kicp5zKCVjtU8lWCo0C5fkQH0IbrUu6/qI8
n+Hq8E4o0EE8Cef/yHRcbrRGgla57nU+xz3UGRhzgpgLfJswxR5U/qZdp6uktziUiemvbKq6hnFQ
LL/jr8MvSAG6Ij+lTmJ2bEgCsSiOzgCbh3zSuCNceNcJBDHJln1+rjVfRJ/oaHGt+zDfHt4xDFbv
WOMfE/Ew7+xBEiFvJSZ9gseAd20cDG4Y9aAv1CHHNFAJGdrlK2Mv0OCW0x8KqonhIelNigEb7qZG
IOFgkoad2VQHGS2R/Fu1zX2S9DXl7dZYmUM+aCNJujOxQ1tlL5Nz7DeYXMTls0Nk4xLnuu0hrJPu
ruI1iaeZy8tCU+/ril+v0DVFuTm8gjzOZuanzfkp5yS7WhEe1BYGOELNiuAIItZWSjng2QYC0RUs
HL2A9NJ1fFUPISwThwj3LCTgkcQ7frGhStdQ6Ou03BPnKJStPSpIYseg8g7v2gqZFeLSYdHN85I/
RRgl5hTL80GxmYsMNy4FAcimJrils/qWBj8YSmrH2fbh1uROdFYaVJHfb4yKYHQXuMipL3kBZnjQ
3IIQfV8goDvIyD2ZAd0qhP4pyuaMivysNKW4DO/XvtiHQF1j3wTOntKsl9PYThvZYWkSaeU1VOZ3
HrnWe2cvZERsFnZfMMvBBig+WE0ryThdAgcMZ93fNmEp4ttl/7zBFmcTdnoa1mfYqFeTcP9m0w+i
xoZ3UHc6/ukCcd7m/TViAAu5plek+J5x71OCDVD+BtL4qBhjhhZaMc5pn6i45kwwjJJ8XWBziwnq
PXuipVggQu1sxUezq02+5157NHjK8nd8JQ1MHyGTzkbNgO/FKmb8+UBpVGMgZf3M1nXvSriQRxLO
APTYYvaXHzGSIkZ6atQ6uc08aSHm+zNLPqENdn1nKHD+txQ8ohtpMXjc4TmRLd2WBk5EhftEJ+Wx
iud3jtNgOD6rAPnv5YzAxyZmgoqEoVYoTFuPjLyf8/2JIpctl7VNfvY6iXtAHxO8mqV14JFmPIMw
k/vebYpv0Jrem0wygGQngFB/xl+J58TsY0kDd8cx+PEFx64pL5Ib1c+wXyLI571zHVz4JF2lGcXU
5S2vhZ8JonBVpFgCYxjiIpXqzJ9QO5GC65iGkf7PVlHJ5QPV9nZC7sZGXUEsV3oMBCs8T5Sq3MVp
Sx84vl3Lq4UlnHijxboLsCPA+wc98PGoYzYEzk3+H8eLZrhOQJkWO/L6VRZycW5eyxX/xIOYsN+p
NOJfoBuGuth9WdfhkSDmpn0cVXZ+otETw6re/HsCSZP808wp8i7gwdLot9u+Ash5+XAVR8ciqCu1
oMwKxoKztYIg43S+AmJyZ6JaS39WangyLT/JYp/e7NmcNkGbncigAglovBpsBHuS5wAW6ZDnYiXJ
HfykHA8mf+Y7e/WeS+vngbdKApASHcJhmAOfibP8DAXopAxF/m7BOe8Yhx5fTij7FMDinLtXwkEB
TWkD2VDNeRmsipATdkJ6XthJG9nH0yuAnzTvjw6h70Qo1eUitT89czeDmJqZyvFPWf2/X7kGrvQY
nX3ic1IxK8QA/IAWdtvEAyEHtUI4dkis5f7MBZusrpMz2UL+TM+ZLOh7J0mQ6qs5OpJbUAyjOkRQ
ckwjK6ThyE07LELxfd9V3CPN+biadvJ8/FRFrgI/2O4zNosjiJrTaE4tS9IpclJ1AOifqR88SPTU
uC+aTw0HA31KdaDwJYnVlWTP5PSKnxY9t0LWDLkUHVJ3gapn2JrkRs4OFtRcnQnxRUYn7ViwqyAm
m+69j4kaldhVXaMyDPFm9xw11jTR7663LGTIXanBCMWGNehG8LB0kXCoFHq8m9aAVPNb1l7xAII5
KuhPEWn4QTc4sAHwcJ9Ye65uvViztxbkYb+1y0B/Ukfh8rRDEA9PQAOKfHLdPfmikxtBa+bJNj6d
6LSoh/d8d/4Oi7L84JrSIQn54U/+Jd+OqHpQx2NCUsx93UWFSrQeT9n/fW3wFtmoE2uSAldR+eqi
gJRjgA18Og3tmEYBqkjvjRiEvfGR6nEAbgmFD2yPuNTTqND/jg4NJRA3CA6aO+OlgpzUYHRRPi0J
+JpdQKLIX690sGu+fFo0T9UeugzDfRIBdwrWU0OxlLpY6spLIVYw8ip42kFz1jeMx7XAF7Sh9iuT
BD4cU1C3XHCxqcBVGiJ7ObH+7/nog9YESwYFFvYfo8VeoUyn2pYK3mhaW9S+9aYc0fCZRpmmQ5bk
Us3zvU4fXtFPDLjTmo4pvXl+D6+IdlV5gto4mXlO1qwHgbTzqQNXMi9B6efh1O2LD7NhPtVnykfS
hxzb8i7+F3ahjcmciXzwyRXroFWq54nZOBAF6egLQdHhiETp2EC+keZ7rSS1Lbid+Mn3P0s6n6rj
p1dYlWGrjkI2sHlB8/9qbhqYkIODGWHnKVULU+e8DYFQue69yvcyp/YWIBTpj2WXkap0G3Lgs6cP
vi9PqryCt39S8J7FzXNMCPhvAs2ZPuDleF+Pr8zDxTsFNzUTa2n+ZopRK3Ux2o/rfhU1KvYEnTOr
3U6DJPWRQt9FCZ/ACOSWBFTj6rmcMeMiHx3GHL2AwOOwa/GPvIKhSJz7ede4+kB71BWUGM3HE26S
UznrPjaI7J81t2vf78LTfVmJu6MF/KqTQv44PsP07+N8DE1nFjRzpFhEr+M4pcaT3jp1FF/t8yOJ
A6ELc7Z4USt7wTHjjy9dJ3pZVaurIyVj5Ql02McqUZwPf1N4nfSAcdSvSATYRFkb4y0KASPA3nmj
YA5CwJs4wcXhOdF9dFNrA5RwS8kDSj/Ll/z4kS55keJJilSAM75+82DfHdwVP4Lvqnhh/Qxnhk6v
sFWNX+t71AZrn7DSwYzxYDK0JbTY4BLDViGPwHYy3q/TjLYrRHloytQEiwuUMRHFeivkNZ3xeY5j
Npr86Kt0RQ8wdrcXaZorQx2CDaG6CLqRyDJIBrJvdgbIYEYgSvOfH8McGLc6e+bNb7o3433VTB0m
GhDLBFWR8Xz49DKtfg4HcKf0MwdL+1zozWL4bC/vV8MxVwb6s0AM3Kvevlk7ZeMIi14GruwaJK/B
bnGznrN/9//870K9Qeas7S3sVl013gPFkh5sVb6aT50IIGRgZYK4wdEAGBKCmEFtpY076Y8v2/gB
/cB6WHSHrXgfvWKpWCO48XBsMO3DPy1OmALiZvHRRS/XJK4cgfmZb2x17xqtCtZM4I1pIFUdi52a
PzH/o1bv8qPS7g5CzgYBfikzY7aNjstMk8h9Vdxr/124FifNgvVxAylwVnEZ4n5xlBB0L4gzzXqQ
LzZxVZ9442FaYxIDfjxU4amlEGDIicBpr1PK1t5KDkr9Xlt/Rh0lUkXuHqjBpPJb2Xom7pgC2NpH
QyHB8IKh5i9FxBWQOhTWiImiu+aG0DUTOT4pG+pmB95xrmqR5YwisFiRyjn4RlQfJh43s8aAKaV2
D5uG0LAddIr7iZNSryY4YkVo4jnZEF0m7DxwO2LRGZ6XFbyrEwBIXmv2oKeOfsOsuFZhSK36m7u6
cTx+KuLdD1jKc+tv5bgBn69wo0yfbYY41DtoalNH4iSHDku2z+US5P4f2+D9K8NnJ7YJxQazFrjY
gQ/nZu9NbCLHMb4mTfjiXmg/rvMDT97tg43RrfrykxwDdzPbTh9/kZs6sYc7pQnGyQx+TbZtqqQo
GsvhM/6pmRSQAIBiZk4GNCn0OhYjfP8NqK+f75DuDGmhqsrtG1UqG9ZQLUG+bAuimBmS0NMI9cAW
+e9PrstRhOtUBVLtSgdPEutO/gYn6JtHUVJXydwH0mu67bEtRJ9BViPN6JZqoZEcxdiSmWtaXy0F
wgU9iD0h2f1q+YVzr/nbtaJKRiaSctI8c4WI0wF0nwePs/m0SVvoJ9+B8sCQEYuxf6vScTT/xqzC
09TxVqCAu0S6JiISPzzAcuLQ9qpZaUycmkt9QxAqeCT8/wFuqS03u+gT9ZYs8MjSD5nO+CUdAWPw
Pdoldthfw9a3Tc7ReSKP9ZBcabx8MCOR+hNk+I95IjPU3kzqUfTUEKFC6eun6rG4X1SEOq6iQRza
UrejGzHEFE2mcxsIuQD4Ovh57Mk/Jry7hCLrc/rX9AWXKWpJIqSVOg83SpKHx11JyqbsLxnTwYYG
T3nXqNzir3dYLZKa45ZkU8PZpDJWe1QsOrGkJO2fp2avIHIISiUiIK9wv4EpyqyEvuLRmwpXDRUB
tIE3+kLqqIZxLpzlsfmbsXOhUqA7BAyxNa4UCT9WNmE5Mi7hbDNCtn9BQu6RGP8PwL6fPKXibbui
g0qBMRO/mVY9vBkhZk12PMVZ8GAZoU3DaczD/s8AkyR0KDXUI70AmubX/6rD9FSP6Ht+osgNjY4E
gcJnU21lCHAqxoQ40m+6EQafQH17r9cnMW5BdOld6CU0oa4ZZ9m27es3k97WDytYID2yhp2W1xUM
yQ/k5DqtGRf7e6URY8sDi11EL1gKyg4rr42YiqQ5iTbQkUneCGSqeSgX9JOFOxPRn++phn+jVtL0
kTqguYAd6eskjru2LCQBsPAfIDEoLyS3gMfBIeJthgyuLKYXuY2ChpTFKMDKbBQx/xJXfBgEt8EX
uNhIzE+blsVNEWsw2ySUTKcxgu9yFV4K/fsxbPEXQLZFE0i82xTxgfCFTtbZ8G34PW0ybpr1v9Oo
K5pwy+X1I4VyCq5PJkkv5TQSEnyJlHgxa6CxYPFd4x4Ylu3ccxhwKQPaRUvjrCGtEAOUCmBPprYu
d/8JL6+xoyhpuQnbWjPjPvZkV8VZKPNetsGRR392vmMsz2PNd40gTi1tfNcZb6AGaQUJ5LKeoqVZ
iEO/WoZ3LF7yrzv+GfGJOiIuzdKeF95Gtth6ih6fay01+qRZH3JKupuJJv6r4bSabmdMQNSZ3oLP
RqTV44szVZgQlQfpSnwdfk2In7hjgaXif0W/Doap9LuCaEUzbaBKRD2SC53wVjSxGRqsPHmldB/J
8ohCc0l5y2uWaI4RNJSB/AdHvLKCIQiapOqro1dlBJmD5YvIdU/5iXDLn41yukKWFghmI7d5Efv+
fA0IkYnp2BYWLBLIABYJuL8gx+mA3OYH/pkHdVK3HFlTwXo/jGF0byzWSpw/PQ+cAUeAR1fhjrQH
X0eLmdB3vsxEzZM4cfA3NvdF0ny24ufBAbb/OMVvTSXrk3AKqtiXYn83RdarZSxbgoSb7o8n/aC8
S7yC7Tvg66jaWSS7S2TnSLHCzF3Sn6n+YIkLicor/xAekpHPRZwd0071EkQAe/tu86DolqkPkory
xyNcDRgp0W9pofZ9NONwFg4xaoN9zEOkf1VGjXHGbZbbkt3i6JJas5ZF1OBa62o3EHiu4WPxwO9H
VfD9JX+qP+hxsEGs1I/7BWXdUTeHwSyCxoeqL7u1o7cfCRYxlGGBZvM1FazF7S3rsaAnzDi5et5q
Bu7nMhqh873R+kLRTSRRFUqC06RZ5Xc0MU72vxvKXdC09peVGiCdImm89yZ08D9EcYDNoXugn0Ym
O0MrMrZs7dGNgMWC4XdrfWKuTUkNG21F6OBpsc9pl+hQ0A1ixRqAbzXCqP6dXSpzLOTG896m3h8n
tHt3BvYnaCWRj06alG1uZW4d8S1WTJU0abLSOaXXbGXJYIPGdsDTJwnMFy3Bs/HHi0hnCm7eyF8f
Rs4Mf/7Bq1kgMzAHWyZLdutBLqPL2o479LqyiOYtaH8TCq5wQZ+N/Oug6EihfrHT7OesXwf1ZUe0
ZxyBhKJOiEwVFcw6F8BhbofW6kybPq9veawZEHQ2xtCVrqQltaESpnNetit4YqQZMHbvT8LtEabO
7P+TVGfd7rT6uYCqDzYguRDA+lxEohOFEnLrMLO3cytLpXRPNRRC7ESCpJHCYTkLZNWOKgzLbcQO
vP3m/YAl7n8O6WgALA/+5bjUqW+g7LSVwnvZmkhdeR9fFF4ux/86ZjxAts4V7ygBxHdSyFaqGG09
n4AD+zH+iBGWcojhwia59ky3M+fBsZbpyM8DE52pgnFH5nrH4nav5L6XcDH6xlRdSnowlzctnGqh
UO9gDfJdNkww6qsE1MvkgrDf4S8Dd+Jh0Nltd/tPL5/UMg+woEJ4rWE37COCi/VSrXGExv73F0ih
jcw+aMeO8zhgbPCdySi7KVYgum9pnezOWZYfOfVb4zltxB604L/v94zY37tW7RHNLnCaGOFE6tJ8
GZ+FvTbYsYFkchNjtlhB8IsypqvAx7NgxkVb4XXGtzgzP8qyfG/5wPvjBsDQtIH3Rz4O0Vlf8cTv
7ANiwyOG6+ynLeD1rzt5cYaW9x4FeUTWFee3dICh9VBrm0H+pe2YonWDq2P8tXwDxSbGUZ+lLt6c
ZB+17Nk8FH2o+35FI4N17/cHsale39s/H5a5sv+IMMWHChXkztyNj6nK1GKSNWMR2a+iEi8ub6yO
wsPnMzMTbMbADZxstqsnLc6vVNwOSO6zewO2lWp7qRvJg94/L4KidHpDm09e8893s8XPccJ8KxL7
JtcTGEbezehur9kA3kIM4nhtM+6cUwwz1+mAjP08jn1w256Y0QqtQVrK8FmSs1JSNfYdAZaqRYiA
mOIj1lQ9w0N+H4UPTgBBJU8NKK6oUJps4gIJ7qSiAAALRAb7Cx0SXp8n43QEUbDhqmItfTnpT6ZQ
g7lv9Wo84Hl58jPBHzkN3aOPzGo44QH07z5zUhI+JYGn06kIvFKbpnx4fWLwwDnUAeNFps1CdB29
FZspB+yOUsXnU/8mGv2VOTGKn1PzWlowETgwf2AX3FMYDhiaMc/SDZzrwfFYdWrJu9Ex1hP+iswV
YoobYxBWHkCC8Ht02i5rKut0a+T3vV2b9E5OnigRsZpgWfDD9ozFNJbyno9iSXVQOuqBKwlHj2F6
CpSWiT9J+MH1chJa1Z1QndUa8g3jC/zDACUDHt0Wh+qjkKydLRiPvP/SIybmiQwfVlFRdG5mUIlN
D1jBXRgTpo2wSXkuzIfSiIFB2O+U0NgthtGcjcorbzc9mzUdZKDLAbRnKSiYsz+frVoFUm+6B6t5
Nuot+BlYn732RdCTPS+TEKxaQQtpa94NwzwY94BXA1eyq+8oarb/70JneaICSGI9ssEgw6nbHAck
VBbhjUWZ9rxalsjnN/mAHX4fS6i0pnjFjwU/AHkpSgzEcvEr6PkF1EjR3cYwG/RSzE0wCXIjuwvA
LPQ5Qzt4lVwvCyWZKVrFFsv/sJfw8tG9qG+Maenc9SJCWJ3/ftRZ5eOx0bbpk3nDPIkuaw8HnAy3
pgbCguVe0cs+XUpBVqfrysNyv571EceWjVmFF2COmuvw4oL+9xUkQUgUZz3KXCYPsSgWUOGKUi3b
QMFTtcyypGN94YMdZ4MqbHeqX2RUonWQF40m82HgN4D8r5qEMzQr7HIwnJTb7YY6OQh4FXJW5fui
l7o/ovmbTj/vTvWNfmyDI0Wv5MLoKy/3134Q28SZ6bHrYgso1e/oXHZ3p+lRAzH1fTnEvq87eBn9
vedJBRicbtu7KiPS6UlzU6/z3ZK+Ebbmwrr6xMEOmIC0EbuAVB22FD/HUfcMaA0hw/fI+W31jYtf
MZUn7Vb81VsKWJke2F5Pg24lNYYLKKzib0DhoHnr8j+v1jWcVxJ0GT3hoqYtCv1M9Qrm5oLZTg0b
i1vjJCHzNGHhmjXOe7DcmqsL0XHclQGX5me4nHyzpGBol84lOpbYdjPpLbz/jpfqESn1MYHCtETQ
GsCsQq5Mo6fq+knjra4+Wq+H1AIndfBrqTmbFTxUHzLLbcV7bISjvtynTyfHCTuEFdnneSoYxRpv
Vo/jGitA12jqDZFxq0rTN6cMvJpR7xvjCYgm8WsYax5bgr0SUOeMIUJtT/8iW79ybq/voQMpssXG
dnk3DNWdS7nO41Q5rDZoPBjvIB338Rtg+R58LjCWczAX/zLM7+EA33b/ZN0/r7T5viiwjJ4+dXGs
lzLWAtAoqA8+kZaUdoUwFdcbRp6CgEshA++nJypvi8WwnLzsuR8Mq+vvCUTeX0HmcpMAIDW8HN3l
fDFdQTXtPra92ueu9CAhDjQu71fdHrgyZnns/5HtuzM1VH5kpaFYjG5/fipDv8XY7gGL8CagmSZh
Pjx5oxjj7hY8QUqQwL7vXtnfvYEPDjPJdGEcrKK+CgNFQLy1gUYyJCYYi2BufuvTbODSuGZQVzQP
F6dGgYTKXT8rRmP0Lq1paul+ijFVqaK/+p9XautJ6JR2XXV/YkT9oS6/sL0xlDPqm7nEgOxHkYRk
O+O4kWPfMXiCkmtW8ApdrJnpzqTa3WAtyV/yKnHpT5ZA7EFUFTahX9/pqN7v2g/lcp8vA7MEM7m5
AhSanqs5nH7QKbkRyKMdRC2hjx41SgK8F0rdpob8U3wl71ksUuSrTgGHuGc0j2XfgE5cVkQRV1EF
1LRkJDZtrBEECghcWj2/+Dwc3P5LE00ZY91+elYMMHT/CECV92WJdwqDgwQYMe/1L7oXNYiFmtkS
wvQ3f0LqryIlEa+2gS+y2/WxJdMqU0a6BAa6QDu7KJmskwiOYvcMrBfz+FzFP3O40BMFOmxu20Al
51gaiBeKUq5Q4J4aMKknjKOQ9H9OL7jiBvXu426wyIOEwJJDFuhXPq45/vtp/6+jwITDOoj8aFst
53rAvMFdXKZ+A/TX8xEtAZZns/4ATOcuLsM+WMVgI6ek45FbCFXvd3RhkCWtnsibbsZxH7ZAZL5K
ttcjWw6i+nrY1atKDXDkRbpiXbU4kFhmXTQl1rknNIn4JaobbNi+mYSHcqcQpVruT3e8NW3xCuHq
PIDpKa5gIN95/frGsrtBu9EpIf545UMYSqnDL1+dBPi+MMcLlIPJkXXqwRDVyYbBhglhWTTWWKAx
HvW2svRGFUsw2L3ezeIWzsMa8OLxEkjmDFfdgFIzzvNArc/dQvCTSIexbJsK3t+L4uq9CpTFRHIC
6wyo5B6fgdWsUwJKJeB2GrMp2xMiH4nYmTXvsnBg0xBt051s3Ng4FL2vrTboziRrt06kFxYFl+ac
JPiD2/AcbmpEy2c82bavUX4wVlypHrbFQDapEtx394iMFZfDxrQWZmAPjSWs8UJGOsxrMS7nmzXc
dr0k7jWn4iD4x/lf/kIuODiuFyRaCOaNvVPaZS1l6bIH15ITyH9aI8NVvHPAzHpyoxSKdGFfTYNr
ZD/tmaffU80Rbm7qltcA8l5TwPfFgb9wCzvB0M2XxgrBx55BdqFjhdXuSDlEIl5V8GxDL8Ok05sI
hLfTTdnfoZT0T6A7M45hijGuJ6EPYVKEAp/bMOgrbfwSKD2KOY7gJzE2KG9vRjsfQUkIE65rkmi2
2r1THnj+2vnRVl3RtHPc12wvnys3whk0B6z9f8UFAij5kPcgn4L9ykdUwOIJIhLBU1h5krTodGV6
qkMWXUpw55PnxMzE5GTUgSIPdPKfsCBZHwofLQZS+1JtM2z8NidvV2LAxIV6TdHXj/9PEiQ3/Lup
JQQQyrHyfS1oJ1ZuMgaI9o4CQwqJvjXxGRgtWYMEc2/PApvSaAoKh6qSCPZb1L/+QkU8W7xEzhk6
4/fqwPUxFWTGfeVqIxC21R921gt+4ut8HVA2XvmmEoTEpVobMvq4GijOJih+Dthz4qw5DETohzfy
cFxGGrV1LMeKGTgJ2evTQIkfaXhDkTohnyoAguRZg1DEHBthigHFThCXR2pCiXXpkuzr9v7SUCG4
Dso+7bO00Hd/Kp2XhuWE7FEqI61Pf2MV50XimAunO9bpoDlI3Hh2F0pMHZ+A5HfOiSdCD0HxEmer
thAK2EqJ42YD+ZPPhUsfNGFKWf9hjjj8djMdR2mHp6Mg42nLFJDZPsxLblNLwOLk4FOdt2MqO3ix
AGosZ27TBVOR6nFMfCJKVz3kbzrp4I3WaF6MHL/P01wLXGsW+U7qM4ZxFVw4Pfoa+7e0iTrq0yVy
baYgh+Ok96hkza4bO5qkVvQd1vpNdzlQdN5utQSPu/XaqYtE/6B+S1+c/IOt15rSrkRG36KwHw1V
LyDf+FmcqAePPNLkc+32w80YTvAgUFJpmoZiL3A65QA33RLAvCAC9VS840l6J27wR++CqoSQXzpj
2akh0gR59UnuT3OWvnawiVgwPFrxZOdalvGrTf+zzO1OqsiExxuI0q+vpZNbdz1NQ5be4/Vdiec5
iymXanX9nzVmw+rcF9BIxO3iyR28A6xxiyBkZIOTVYeyZ8bS/QK7IPiAAPEVkF7THGOgcpmLalw4
ZzxoHm+oqlC8VUCXsEjnK2VKfNWJu/gQyXDND6y/cbi564ORwsjbz8SJ5OM9cgTFGTuiETTLrGla
xWfXcscA9dfp4e3Tftibccb0dXkllEXcVrXcpzajA98/vYqJViLvxzfjV5Cub/YbIgtw76dQRjh0
5Q4VkD/zMyzvVqFBB8Mw7xUuNg7uoxl+x+Nqnds3SUWIRE4T4i6asI+IryWQpm6QT1WARc2Y4f3w
B+etb2ahwlxfOpOVVWWg7RAnWeMhyCnxxwrImyDtslkyzz5extbpVVKklca7KfAhBeK83kZ3ho1n
maboqZQgODtvf65KMJsEPkwIkAyCWPekQUbkcnT1kxiX83u5w4Zg66tv0Fc0tI8ryS3t3dmIMztP
K6OL9i0cMpuPOP7h4QAqhkx2y7vT23YDZRUDu5a9wKUat/owU5uWVAe0UoYT67MC9M0RxrgiSbia
xmjjumGX+kWrbGBhjEG7kexzdKxUpGBDN8dAd1qpIieI6BScymWLekCgtpFXm7p0yHrGS0aUKfZZ
qLN5KN75/6C0/mgNrYgXahyVndPyFvCNqO3nL/zrNMANBbqDgjOlLowRD6ACcRS15cCrEyhkjljt
UBjDY/qi9LfcG4ej7sxjis7ej64XUb3vAjRDyvZakcOsM/qPTB/Xf6AmXLVBp1/6Pm340ResSxtN
OXlCjK/tEASnXwuJHszkblt6G3HQ8WpK/f5eesr6kckVd4sPySAIQnmIVepu7zbEHE2nwoHwFCk+
lJSrmXjmd/0Fmx/qdOyIY4mYxkPpd1AM16Ifr5AXnsvGyRmN3bzGBiOG/VlSPxRCJBL/E1xSQUvP
Zt0q5gEra9YLVkCClenM6jbx7oFDAPL9lLQ6U9smUlhSiBXrhGwqXWpkYamQ/hXTeyxkDFPqRhww
rCLukPJeSq7khl5Q9+v25MhIZkpOrBiNfyvFLVDsaxsyuB1e6vkPjxkrj9XmKzSNCLmiQkkyl6sV
YFg01GQRztIDTY2HWRHiPVnBkKEtZ47BZDnCX+hpRQ43YLrgBT8G4EKoQ2ZChhxTpEMzrZox2Fmq
sW8Ez1TQxoBWJCDFKrGdkQcUIqVryX1ecAFcVoJN15rgyc8EUuS/au9ui4qUw7IEKc6ARXF3S0Ny
7tQwLTpgG06M3y0gIzDeoyIXNeC9AtbYC/c7kcUgmgoLT7iL4hOKRIi3BrLDEv407SPHTWU4Nswy
Pxqqim43A+MRH0nuusnhP4OIIYR9cwV35VX/xX2dmAHfh/fOfhyAox295UsBNS9fZd/4Sd6CbkxR
/0th2EN8DDdDKV3dPSzWnerzOh8UTzMCPoVmmI/1HiY1aAXW+d3bBIcmi7zctJxD+F9vmQxM5anK
7LAqBXAdto0miHvsGMaqI0CSvL2HzVr4RV8QIwXs0jEE/Xn5ogXoP5rQ/XiOiDJCr6JlodEHCTij
qNyuJqvq8xLxBCrcqvuycvQ70yR8us2rbXZ5aQHkFO5zIMP9BFshcJuHIZQDMKSN2x7GtRHpadPp
keq7gGh7LyEeLqAttF8sLpw0UAQsPF/0ObA0JuFeV5G6naSWDeyJyYrEk2JYqp2hV+UtSslytA2v
2s44jLj3cwzxBE8qDZJjN/PuKIQI0QJ2cB3Ymk00KKCOjj4kiz2EtmRPeGnPH00hzK4zT0cesOMN
J2t/RPc9oa2E5pIxrnfSn8Pv0gkTONWm4hIGU69t7FSuaxn/Cv+WmImX9P7tjkFKPQdOtvbMy7We
wTI6M5QUayj4TkjeFW7q9eH6BWg1Y/njX3K2JXijXGmGjm7WS/tT1DFiYVCgMeLafq3qCo1QwMwv
GcS8jOUjo5zD+Z5+pxwglgiom5BAD1s6sWwEHBFdnaJ0gVPsR931BFLlzQOo6fbKsLFOwq5dPeFQ
w/Oz3ycT+y7jhnsZ0jNUN/2OTWM25TuEmYiWzySlXuXv7f6tubszBExxHQdI0bGfJb5XbdxQ3oMT
58/P1PQY2dqETOuxODRhpzfrz6LfM4V/7iTu3MwPzt6ysfO2EaJIVtyse7+Nwl5ckpM6Z3OkK0qo
fNIosuyHwDr82ch+ynysL0caE/UED2agrY/tCDkzGMeo7CdPMT5vBAZ8u+WCRP+wH+/5AQpbwoS8
ZBsV7qXdtNSaE4SRExSItceH1VhE2oKP8ZU32QzzNRhLCls9aWdH5QCGcpyeQ2ACZCdh2CHX+qlv
3rcx4QwIUZcSY/cMQikBdTmpF2fzcPI8Gg5bPn+4f+EY3Qdt4hyFidfv+7P6HA+WpM1uD7xwWfaa
c0Feo9eDpqAuz4S+p59NrjWi0GQOkDzXymWSkNb1pa6ezxcw7FMX98iztEd3vBdmJUpi711kWEiS
EWGGVFLqHv5RA6OPduT5jfdyPzqp+zDAKQwFAkWtCM7pIce9+KzspgEEFYBp9rudsx2YaqKtLUNQ
ZYsESutz41dXEtFH9OGC5r0NxEaRUXiiRHP8Uj7ZCR7l1qa1Cueoyo3BIPQ3KdN0KqNI92SA9N8M
J4IqxxWtzOp1O7vRMeFWgFFux5zPLbmA0OP7pAzSFkgrwliMGSeorH0r1Xoo6XdrrS5mG5E4qk32
amKP2iwSVyj4WykcJkpLWHMjb2w2pDpydnsV9Gycy1xY5vtqUgBlhgcSmbDhhS/tR7JGZz35ddLl
UI9xuo9/hOiJ31opZkRk5oI9VlkMxFo+SwfTFRl/3GvaWrOH0MKZJ6Nghz+aG7x9ra/wefhSUTNq
vfMRV2yB2Tyqwh4I1KotcFUVZfKFZltM+N8TvNY+qIbfGgPoM8TBvf5COwsB9iF4D5nED2DB/P82
FxK1D3UOyPb2I9TaARpCJu9azBgvPynJQbirANWV8Fyr31dRXGD4oZ6JwOmBclQxRWs7kNk8BM2t
21VIooxz3x345N+pJpIutyaGdhmdKl8I6n8t+yDFQ5p8/gRLwqxKzoL4h4Abf7y/KSsS2ZDGOEvw
e7QtqDRJb9hQNDvb42000PqDkYnVoJOWyXpGbIp+YqWoOTZ0aTZ+OyG1/hVjFSvQQAeAjrdF+MDT
1V/y9RoFv+6uMjwZykkQTYfOiQvMkPg3Q35UZEcFMnaWiDiMe3s3xO9MDwcGGSqLdaamXKysqKoa
lLd1NhpEg/T5P/aerJ+tbzYSPsGiOkD9MmKcpNVS4OCUBMDfMaVJy3sOgfCTSLoE9Jyo+MlWZwQb
pBRj+GajxkDiZMSpmNrJMC4uAIEJeMoszcn83CGZIL/rIkKbZmd+0F2yyzH7Olatp5KNqc8RpNiX
/kDpaBusw1Onz4mmXO6TXM//FYqvBH+jtqbJ/eyOhFZuJsZD+/2PuvAPTXo3QeQGuDXIvOO9un96
0zGWv78rr3G8Rdqi1iTnAYaUULG5x1lbA+CzZWUEC2HhXcP5Lk0hFomsLllN+t+W8O5d2u7TcFh8
42HcN0lVbeMuOsiTfmitr1sqJgz+IcdTJLy4nz/MDQQW2Lj3UQ0UqekPIPT/GnnRJGoTKZKKIBhp
Pzcayzh2NPLpvQ2Rhrw/hueeDOt3BYQI3y0+LJqG9EFFUMveRwMqQirky7yabf0vy3oG4QKZ/t9T
VTquP50Xjqd4PLNRSBqwHQexSox9qF82Z6uBuyTcFrhGiSv19XRwvEMm7mfehG6wOun2BUzRXaYv
DrUeTVQSXnuoUNjNuBxMRUuroFlRHMrY9afAx77FX55okSHWPKvmY8way+K1WKz0LvBc5ylSqbtA
VJAtseEilR6VRF9qieyYlMYliVp03arU9o/AAIhG88oDoqiLZ4mtWuCGfTtbfqtDu59inbS1nBTA
PgKn55ht7QtoiDce+XJQMCybrcBj1TrJ1Vo99rgByHwoWmqXTuE2gmixwBb/X2wBScq9XMznCsHl
FbKj/t7P1EquDfCuzghtfrd56vRfjxVi3tcknr8c9wN+lmJpfkhZjk662ZssQ+6T3gvmXQSa/+RL
9RlKAhMpmXVLgX3MgkxB1nuo6Vl1olO7OZrPyhXn2i7EtETE0rnkC4pCz7znOi1M0vEjZY0IKgoR
t4w5lFxjHQbZbBXnDqytMKD5OHr86Uvp65TDmu12WhQPzgGzAy2SbT/Ol0TBIoRj8CAS0bP82kUF
kRQxnrfIabjFU446upoz1qGw45QmfIWr10hZDWAFc9BblggnkFjO291g5digaOp6dBr9bqyXfxF3
x/7E3rn/1k8cKktx2A5IZrTWZoq2dbpbcSQHkWdUbInBPLmX7Z5OeuUlMETQnT9WAb8VTXn2Q2+f
S8xp0ju1tgUEolaZeMDTWNsRXSAMSUqQsHU366QyY8snQZP12b6tJ3hChk1rK0e2E6LrQxUBHrWK
mFpLy5L4dPPSclEAyK6i5Yf194BvjpHl41Q5LXwrsDw7F/gJEhw8JNnu3VvnpvJ6FWgT+byD+Gxr
FcgJfOMo/YW9j1r2BDz99dit5C78c8zph9ylT8Qq53pc60wQPtr3BEkHtu4C9zycLDU8+04mE/KF
HjWt9EBFMaqofRyAIBHHbG3WdQfnpkl8ntKnOjTEmca21aSRUIXiCPgepHbEE+k2rde5qQAdAKd5
J3W2Co2eJZJUG1PGMrOze4VxECEDjUnFRZIlF9JyhfRGjMu4jh7MmN0h4ngQ2ctD7AA5JjRiOYRG
D5+uh6UPTn9hZbDjfKHWB5oT9iV7J9jENcp7P8BS2OETQdM60W5rE3iFt/6dlyElH47mW9WC/B3A
j5dk2Gwpbgyu6oN7IVaSXD0bpaDM5ZZM6JJGH4BePkV0RpFOkTfOFsC6p8DtMCKf8MB9v7uPb7Nm
Uwlk/WNm2VywT1qbIwE0PoBzjHNbPijGMsnTAtnQ81+uVkFFFznFfL4eRWEoi0HTTk7HcElyjSYa
k4m7tLfYGpp/fj8Udu5q76XGXLgf3bO5ElQGNTC1IJaErZF4lmodwuBTY9xp3a957mLG4iX0K/GB
LE/T7xAqirHFN3dO1r18MspMnEJTuoii/FNxYYVoAAecU9c5MCSKpU4W10G0hRITzibm3zvo73qp
r2r/kcMZTTnh4TuAv00OEmzKFyvXk5S1HC5Z7VkLNXG7QKNvsbsVZY1Ubzi/f0TmHcsE/R9CZ0t1
MWBKZ+26wvPaHsWw7I+WLd8AxEqH9wFARpK5ExAzv0Y+UX9TAoLlVreEj1n9mouTRAZJ5NyJehV3
wIhmeAje3W3sRJTfW08N6gAIBXQPE9ZdixE5Phh11JFwwX+no0ebkWQNLbdetpeF6tOjnJzYOifW
+CBVDo9Bt3tEWuRWr2XNtLMBviLTS2jvzkdCBEXiHUnjMFCGIRBT5CZIQwkwsc2uKOrc0IzOcAzV
mHCX6/AliGRwCGZgdh3pUfo41ibeXJdKzUfRs9Fkz9Qdw363OvkljMZv93ShVJLh16kKO0jvRjdJ
yE4yR4wUz17BYXYuwGUk3K174z8hOgiSwxDv8q9So/VmgwYu8jLJTgu7YUaT0IKYD5U/EX4g5Z7o
hbnXHnoKagB87mxpDlPYlFnABVtgA4oVK/FSyC/nB/UuKiJ5dp2c4itu6uHg0PFjr+ksZlWmZuJj
mzSYoXEom+jV1bQei8kb22kfs9ncRZplWU5fcHVh04NVrpj7gPzaokn6XD41enCP/iHaXXnxxtqZ
udOWe0rX/rw4ad3gFTJ9imIfxcXNKBLOr1SHt5T+xE2IHzCTNOuxFecT1BGG32a6wFE7W/eovzHj
X/Zo14148rpxlKq6nxz7BTCRukCv2oQYwQB4+15sB4psQUYMXvlJsuIIAcqW0Ma7F9aGwm29gSvn
8qXVSJi+zV7FkSAlBwT2yLcgBNCCovtwGWp0qiOsdPJ2uqM0ZRhqHQg6/EWh5wcraB6SJq6Dgxuu
q9UFHD7Inxse257Yrgw+JkYb4srUJlVz+Y3DH++lkUF1F8Kk8T92bQgcPQrb4iQqWY+223CnTkMX
M6Ux06/Hka3OcKam1qXAghrOKhBosSwvEaOifUk/JXlB9h36BumfpfwKi+xVwmpIHYT+2o0vaKpr
j00wnBQT69AgoiqqYsCz2/V3sZ6Y+ucLZ2G3FnuPBWnU7ngp9bWAtjd84BcYDD1Vq+7WjTjng8af
1XldH1PYE7JcKqA2Mlj7Fo7apSLTAEy9199PR9opOedroXtJFskbF+rTYw20UpNx2zb74h7QSf5t
JIYYpURo2wdACBxxxWvMaYNpdaKuZ0kyXn/Jom2vbNDRYMYtWNkNh8OVhnyxddzji/KIkG1xD6wH
0UqjjaSZYzWsmT/nLRgbepuo3LeUzHRxsdTv6JW/FIm+qyJjy6lRXSgThQ9feqHAPnIQlWuArCSc
bSN/2FmcaMZGLgwQ98Imu9kLwMNk+ieKQfNho5dIh1aMlWqal1bFWHnY/K4VQSFiaJ2oIfxVDZDt
Fan4WJVZ3arzFpEtoG5p2+bxstyioBDsg/iQoedgqXa42iWqs9Tb1lhxeKmZTlwKLpaK5Vz711xR
AGhksbxWz1ytqul/W1qIEPRQp6bVuSJqkAUmvgZt5jkvuS+LQkVghCiAF9aL290LIILrd8jcrDMo
hhMyzndHPKRJ6s/jDoQ77PAmdW8CciDjGY3s/aTWMokB9ME44TeldJia0pYn+J9VFbFZ27oC4Ar8
5QLT21LR+Vb/raAFbCTq5EvMwxDhyNfLZIc7i6vPJSi7U48mot522FviDOUB8kmA9Zr1W1+coM2V
Xh3yK88w9OcqyJbByS25yTdr6b10upRxhQE8j+IIMr2GLq1v9YN1/wxS93Bn9ecPDBne1XhbVbCI
lZEsrmx9Z4WRGGFEcm8Oz+/D0o0jaNinfq1lJQjUn6xAdb8949gu+lzWp6kEN7wqg3VBYAmOTavg
+uVuzBsDm/KO56XA4mhsGxtou2r+1UXsQPS02zTwPJrbkIO5XnqwE6XyjjqkzvfP0U81pYAg+G9x
SuAR6Vx1qBpJYnchKpyEr8JuUoBc86X3By2d+yCwb3CnbL8nwIsiJtSNrX7mYr37f4qf78TDHTkq
zqoxhAojmPkkF7aQVjCN4g4fqZQaqssKhGW6DgegBP5w9o1iHmVZGQjSceobf0wnyOtIBlaqFOAS
oGkt+WDu0eEk67sjR+UuDv339MlZ/sfVyU4tUboyd6UXecjpsLoU5PKcPYL3daTaabB4fiUqteuJ
t6XWMvCQIuZeOuYdBKljzdMqHSWP34v5rbgOFpDIg8oQySzkw/v+ijQRXjonHH1E2tkBleIKOchm
lgCVcAHe9TupvKm1i/+aZYN/UoJopwAFluDrQMmz35sG/rxon2VpyxDAcF7lMekhK+hySanlCryT
7jinFMI5GrU8TGsU3btZDE85jX/yXMo5FdddlszK8zWRTDVZbrOcPjTT3v4a+fDWvUVA8G+7qzLi
KldEDC7kkm5+oeczZSk9DZegDSa2AEFO0VwbmEVeqmXavJZKsKCf7bZPg8ai1bPfxt4KldOZhhnh
tgN2G02tLzroOJU5Rn0mw4blzKS3Pk4taY085MRt9qxQJOClTkLEg+YzgC6KcuzcsShl7m21aaWM
he1ni7PFW/USKFkBOfG/p4CA46ZmT6hJ3KSmcNZMcr+QxmJgsoSJsyUQF89mxGSynSqnq1nVsCUx
x8pLpxvaPphoRlbgfmzkc50j48sRmeIcsV5xB9/Je+d4t5jFzlOqJEME1EG9oww5KTdbdHOozpbm
8mhg0wATXFax+s7IHm24sFZLxFTaRAu5U5Gt3YBPBnz9WeKlTKzTElscJhQje+PoS3aQ5gHWqhci
xeKBverg0QuGG1VeSOeacdy2mgXhly4Io5Gmv4ajr1qv9lIl5Q2iET918UZm740WZ1X57w9Gk6YD
YVSFR9NR7BD/Ln2/BVbLd7hURpE7YP+I9ooD1cLo5xHr7dw8kJVrYSGIeEWVwe4RoXULOfdNBpbW
Y5eUO8WlU4Tlqbo9uoQ3laAn4pBcX9RL8dipw9skBOxqjk8ZLH54XmUiIAob8AwOzfzpHN40/1xv
2tSnHQ0HHuoo/GjZiUOTRjuq7GuQuPpWH9K2LYwMWVL260Y92wO1vB55V/weKSWnCNQxF4/BqtyT
abJsC49oJaXYCxMBna8QbDw0RxYWl5bDj2eeI9x7clz2hlCA/uSZAUXZAsMhvC7fCaMADQnJJMQF
Txdd1rWoJ3GzvShQ2OlC0ORF4iKNp5H+PJ6RjTKfiVYdWduD02hItacpRjuAD/Q3ewDAkfbUtva0
5W3An/EWEhiUgfihsJ/0d1XYXigzsKQ0E19xEC5W5kVoE3fjz1po5AiweN+QOanvCNqMsmfzNASn
mD/YVJPqyjdZiZlMlpVf82HilQbzlIqFctdCCoQe34/Uw20FEau1VNXebUUQs2u9xAYF3meCSHSl
rUtTpN6834aJBhMncpIQAl9/LhmhQV3yWWxvod5knp1Vyn7j0D6NfOWuOCLNDJRQdN+Y+l1N/hsU
BFh1MMkrBZ5VNP7JgdAlrSvXzpd1OxQRZgx574S8UqAgpbyNjXj4Np1g1Bt+WqEjSIi0s5a0PgiB
/ocDPSWmOzU8TtUatR3EWl5++6ZK9/DH96JZMgbKq1EzgmtHwOYzKZ+yFYKJST0Ev382gym+UFeN
W7PNO28/uBBNWLq1vI7uQmHezBcDQtqCj3+2xregKV9Hllo43r4zpkqSaC0oczv3MAxV20bOr3bd
calnlgeYcnmgYAZsBI+t1e5ai+u0OmvJ2rYv+sSZen30RF1MlVnHwXnoncfrA+fWIG2f+d3gBIow
dL0+iZTfxm50/VU9tRHswqlPMflug9Vc4f+TTrcodF6sWRIdyNjp+eEvwDIAomfrqepSdcYKT6Qu
GDnUYbzGOJTBcZoHLQITE4bvUj/kgfiFrvqZjTdclqD6HjVbmdFXjGi017NoJqhBXzQhsDFEwsFL
7UlIsFKXnpv4a/hyzuR0+0LLToSsnfpxvQbQxuken85cPC6WQd1vxVLQIniv0+u6aal/9wI2GCK7
awF0KHPT5VNRU9QcY/ausCWngDPwZEOikpDAyInUZtTKy3VqWpxCx6GENgaN+PaTKYudQ6ugGipA
yFH4klYEZILF/XXdl3H4e5DiI//V78d25mkxsoqTI9RCGdnrk4QVQfivCcwVgKKbnLHB8RAOX8BM
w1PpYE0T32cWWO1ueipfq8KETpRT4HrMnO0ClNwcXHsCwvxwX/zjf/QuZ3k/8E1grrIKa+xTguG5
e2205rQNiNSXc33vNMwkgTJ+5L3rRO5yozJLMVpCJ83KtsyJcrIw2/4DBmSB5DfZZKoa6lf7xIn5
1TtqpJtO+jN7uf0yNppEuyfF/8IpvVCsFnkXM7VsEZzFbr4e0ra+li5pmAr39BnNDUCFVC0agYa8
fcqg/jBatwc2sPP98+fo9P7HpyzdFx41vZD9PU41mIs9B+/BzVdlPMPbRJp9Fhkk3WbKGyqW7ebZ
Fv00TbMt0/cTNVmm+qwRmpDPxBtrX9yyP59MQYhOBGSmNIcVdbAMZmWd/+b2AsNix4Zceat/EmHs
o4/cR/A9fBJc3t4zR5y4tg8FyL7KtXM4eUdZhq9HtPfyvWv4QDlCcC4BS2UalFI4zhhSREt5vssm
s3GHv5upHNEOKWSEsrhTO0o03fK9MiIEBqa5QKiSGNVzPpvKKRtE+Xo7Z5zvEH15wj1cbDyuteTj
aVMT02jo7X/Wdf08Bl3aWnyTffy+CRRKtNbYcA/JHAqLGYbWFfMVl1zaZCBmG+c+hAs1idOihDbk
BVNchw9qR8YhrEMiDl2KQ7RooEcYUY8ZMnZnGhFjCOsHkgjMcCccK3TG+BU1dK8vERnFJO8iPDae
4eSmb4YgmgZBkgRBOCE1g7h4+kkp9byEX0vtxGFitx4AXAaAKrxnTaMFrKGhNiRBUH0YtVgg4ooZ
+MsAQ8NbJwALy4cfkS5WtwAcNBTpP5nL16UaxlgzL6McDO8bepJVnFgdRIz5v1q67JZXNyzH7tpt
GO3ImeG0wRHM4NbNBoMWEgjDnXtN/gZQo4Mpkfmr7QJtq9vCPUFEMpCRucCzJMLDL+onwYLDjiv4
uzNT64d8RgIDS/E9O3FFo1eI+Gt8dxkZyrWSoT/sxfdd1q0WSNDlD7OJCzqziX7Bu29EWWWaKXhl
Fh1gpheUHmR3E7oRnhIvlnz+cmGjDFuuT6rzVf2onHuV13S064J/kZrrl9TueaeaK6gSqJrgohpr
CgfoL7m2SCUcJihLVjBopjt4a4DIWOVDzHGo3GC93/9agUrTrkQHdtzupz8D6xozbXBWDcrRZCfE
YyHHfn2nuueBFdC0MSdzHtZ7UXEbMCDGFn0M7k+7hEFw+RmAS2Y2Q6qBXim+CxJIW+bc+Et55b5f
gxLCJm61Png+bUw0L52YSJZq+dZUcggnr681KiFsZ+sBEiv5WpLpHXQHgc2hKWVNkqSm9kEnTvet
V4v5bgnPfnCyUNX6wYiwUNKUEoe+pgmoaFcxpiQCqSA90l09+d4dwqKcfovCr31U/ZZLuA6GC9xn
sd1viIKWZFloUYjWQbwbbwMwczG5yq7WTq+7DUxwjDP70CRrhPOfq2xpfmrkx7y0KVsWgOeRDj52
YYr/HnDb278EmSCYBZ+QehJV+ahoKF/YtPLmRPAFc0xEsKW9fHMw1Sm8n5tYz9ovcSFWuY+PtJNj
9f2Xua7n/0FatsSoHQxf53vISYP/U+y9U48NEPZ2UlZJsgOLTuJcP55hp+n4d/+1LqpxuAjQArku
gYt5TCegslqOHGTHFdCb3m7++ksJoXAIqH9dJgdMmWVORd1kbelqzUL4/ETuU3sAaZgGIcgIonTz
eHr+UlHTDX0KsC0DfMvqVRXMJBIXq5FLMqjRU492y9CaekzhFsi0WdR56zMSepZUaZUgjH2U7dOK
kPbYBCP9/spqrizZneA8WmjJBUKP49+5/P/A0hWz7ViIJq1chB3QquuAyR6t6F70ofofjzqkYXG/
+sb6JIWcU83x+Gs4mLiTdKjZ4wIzkiyM7Euit3VVXWSF0CK4bf70h4TNja7xULSsXee0NlAQok+4
pt+7uB6Gi3YgoBZ9f2z4fzBMXmBxh9J0MJVoMtl5whpuy0jztAiORw0BFfaiDdsVY1UVxzaBjpYf
eizCsC2jXdJxV6csz5QZx2K7SKoSMLXy4xmHh+1kSPKrkYUPtUojZRhukkrvOxq44lZARgAmwfdk
4EDoHR3mcdiKJLyGg03L0uwXv+6VaMlA3jdKQ36tAxb49aSPIitQhEEUwHuum9wSkjHwX0l6f1lB
L/QOF2mCHNbjnyzaLI7hn6GAPK60JAD0/EbU50UGfy/0VhXOn0lmwaefMKtzrTusbgHpJUIhHQ0T
BgyFofZY/NxgN7USLEdMyRMYjSI1wCGD4VaDC8kuwAhg+wr8RsgxzjJQ3PJvW/6DyCBROZiQYzm4
f8ZwEt4P6tsO3qK7+WgUCjcl9rBRSQP+jX3iLTUsuktHz681s+2EuNm2a98TdBi0X/5eHpals6Kk
0rcNrPsSrNyBwhUVWy04kQHYQ56rgOcpUno5ZdDHnDsAcW+1QM2ugZ1oJNXreIAVFvTA9c8HmpyA
+Xuz7Rvu7ckH3hVbyaL/NUGoB770/WR00SgoYJA0E9cmrEu4gFlitZrf8auE/teRc1sLtbgIaC2a
Fh9U2VN02N3YYdlSu309+ii7pZK5K2kEKKRZ+2OO8jIB7m/JQcfYXUoNBN4Nkpt9xPaIrMwPgVE9
cKFxwNQzQTeKuxDw5hIbZUHDAp2fYez14ZJ10jL1AtHXykHjsRCD6lYIQwuxaHbK7sf6d/KP7K65
9/xVQURtMBUU/hPGGvj/yLWvzfswt4m0W41XUDxy1vUGOd75gV3zAjIhenKb0YaCHSUql/018S2R
xGEQCInZdYBlPyEo0jmlqF4h4ybaliyTqxV8bWj2Sw8C/3r/SIQesp7ARjz0R7D6VMjGis8/1ZaN
aakQoFiSi8LCDE+UYgwhh6arbKbr+YZ5eI4i6DFZgj6u9bTPMARaUhbsPh/cbyL6/tQaXcPGoV+a
zHiZ4YOs3B/7Bb56W3jz0beijgHehScl7xd+ky+jUKtb1DA8m6xCFzGMuBfNCKtoqDYDwG3CWMiE
5nj/zXzj6LqAHgkLm8CrZPKgigqcj3Dn8o2eIHeD/oArRcXzXhY5SC/U/oT7Th3vjYScN8AEAzxv
UjhsLSHAULt2glYnxx0CvN9Q/kOD4bpYvhG4qGAmvHqJ3jHnDOr/BNF5KE6nij4pOtxkOe/h/IUg
WuSBG0aNPMDEH+R3iodU+O9357riUeJ79VzK6WG2CCPKWHQibOi2JNBHvwWkGFu1klqW/tPlMoaf
rH849J5DQaN+z/bnmAPuEE8XxKSYD2/zVISkWF2haDuCOOB8uK65NZV/U7FIaKeT/I0NwAkWrGzF
3dPUHnUF6RLCgqTNGpe7UycV4dzDFL2afUbh/jptifOildmarhtYNufH8nP6Bi+LEacs1J2qTzz4
DoDzQhWQJtwHTchqGeoNoWMGEQB19nW7kuppFD0POJN/GnBcFcKxI/7Pyeercw0QVHuVEJTnw3o2
Fnee+7/kPrqy/bvkg5wFIJs04CmlfDHpXgpBgmSDrRQBhd1BEUzaxfVDfnM/kOv9v7SThjpWw6b8
eoLzxjjbx1FOOqYgBLCezLdrTQEi9YUzkhcHGcfyZVoDyR8MtQH2nRDox9jju9hzvu8l+aSeciv2
rUW8QanuT2t5TF74EsAjVzHTOM3qlmbFPqEZ8wsiV9Gp3jfvXyieg1MLiUtjc6oD0C+lgL+0G32Z
K2L6D8S2vHDClL/oDprIJ56ZddYA4zR26amwAIqRnsCjqphjU9UtXM3weuzua8vIuWkKtIv7Mgz1
ZGEpF5wrNLH7HK61kff67Yd6haj4cna8jVHgvE5o3uNhcTHgdfrfhoZmJaSl7g4Tcaj3j+xVlB1Y
5fChfZxpSt3SD5MqFs1S/olwXJZuOjH+ZAl182gZ0It9XxNfUUxnpXOhWqlFEhbILszPayrTES0r
p/b7V7mFrjID/gcYyR4upQoK4pCVMTwq390Bg0+2hilr3ANsI7MpMcd9Eg1bS3Kx4iDRpb1hEFji
sik/6YEZWGRWkq/4OOlTm/V8FIRm8xwEcWgyyymillhMQGtjbTc2lGdrvvrGuhP+3BbMi+PcUs+H
udtvSoSCWEIu8E45Y5pxyvyWR/hJwWq/5+uC0nlkZ8m9ea5V5CxouifOeQu2kqBYVhfS4NKz6Rpt
uhmQwjU+pciwdU9+eNGG+opWkijfrdRiiVVIebEuFcHlO+KraFPwl33deqVrcWf6aAsXBPKwI0vv
5PnpJO7/uCPzn93ZpzTNLb9DYc0/RezGv6L2BWlHSqcU9POnwBlWpO9eZ36WkXFWDKsHumzDNj2N
nOPhX7VSwxl75QHNWsA4YGL+2zrMta7pVTYK3AmUBPajcx452qIblxEIYPgHKWDrh+a95LVH9W1Z
I4AVH9/jPQVKHegmz2H+ZQ4bTEekIlyqHxyjHuKqf7JxmFLGNWOcFKztSHsyMml2hbxr3+G9cFkI
Y4VIa2USLkA4KBWQpe+yBII87Fr38PRh8a0fawz44r5RhZUhM8s+hP17zheZoYp9d8yDaEVNuheR
tTVTgrpEQ1vD+gVBCvTyTzP1rgWh1vNAriRMz1RSEx0D+SsKguT0S4qJCQhlYK4XRmtbnQqC1LoX
UnuCygrZW4gcz+fEh++Gp/LniGCRGI7FSRDQvzC7fGDW/qpzPHWCOnAg80pt9exWBLQM9ad6CzGs
TaDVkT+fp47aKeQS8g2oII6wZPjcu49Gy8KW3fZ+jU9ndPjhZ8sqaPFd9LNNcV1o/4uUrS/ZMupC
gmbifvXr1bcLUEQrgC9jODZJlN3zh/GKIyFaLrm54qICceanQgowF8S3BYnO6FadpBuTTYa3N3B0
cFWs0rAfzsvX6psc/dEUv7iemSMHK82EUpmDnXBkGqGod5NCaYKBkQt5ltMRNQ+hhL8kmBqhTYc9
E1F5q7hWdYE/ODEs/0YePWMrU6mQJEV5CyMMDxLTcJhf75Sv7UtH7BI12fWGb1itE4ZQKgQnGXpR
RxpU2s5VXx+SQkVDKVud5Wl1X5xbWezWnB/FA5kaGjeIL8UZG27u1m+WiE8mSlkEi6lb6ZcbT25z
p/i3H7XIE5XQGXVYSrLVzYKyMWL5hU8ZcHSs9TelPcOhc9wT9qWWLC+SL5ZNPIkyC5EwzaMECfQC
m+WjYZvGXJoGiVSPJVx4gQ57f7EgyhZnuZdL4HtXuFrFz0BRtro2X75Ei5YTNgfyqWm42kKdPcGA
M/orvYIud+6qzVMoVj6U6wHEexb4K8mnb0L6rHyHBEwE4uDMuU89bHKSFv0cdz68c2oDnuae1U0n
8aj8BYGjCE0u9/8FGqEupVyE0XZpB9bSbH9FeSsHVO+e9RESA0wUcSd2ZJ2YitEDG1CwrGQh8TQ6
K+wJozWod3UZSRhmtt39lCSlS0DXgr1L/+4qcVF8RtVaOo87tqueOPLGL2uRlrBgVu9XkNWSOaFI
XjVY11QK3XBm64qipXHK2VnIhILyWXmLuTmGo9aK4wHLP2SG/dzUPlYOWVquCsurkkNl6u6gvPb9
njvF4mTaBCDcIbo7SsJylLvLB4+KEo2D7Ap9AWQtn/lZt2JB4AIoXvfKuVmibZDorv7iwBFCAEoA
5HKpioizqgZqzqsOlHGqokfogDrwrk1L6c/yjq0o+fhWbjheowfUPagvv/eEG2j0fsq38TPR9vrm
HEa3GAK8sv42G80sOlDLPEo5KrghEXekdBi2+9/91z2VsbVjIw5BI0PWtCZJhlFOqaZCgax0XYj/
xz0B4fQokeCF1UjxlFWpUCMlrszV3Fr3Oy1PRfRe0840Wxs1mz1ZYjgV3xjxbdX8bM2eh26vuNyC
5OLlr8MOy8d02YO6xJyZpWk2qmaGtI0LC4DJKyeBwdjdbHV8FgYRm55yYhyhfN8zWJVGLH9A0+Iz
9zafOaxSOHrFdX9i/QfDS9ua21YCBj5v0TCoqWzHp2zVjISvPnDiQRMLYs9uwl2Z7sng22NciO9g
FfpUlybb9uR0/1CfldwVj3+4GlueLYDrFfqRzjDmlba1l8xp8VugbYTa9nexoAod7DSzJQ2MM8ky
wZzsVbcBe9GEZ7UBQSq/X/cI/OlyNg8GTP2cHJ2MuuGiCJ7JpFJyv9HSr0SgTsToc8U3SzvvflYK
mx6Yg1GqgZCQqOYroJnM39oW4saZgGgYTadPwiC72c6SFfceQV4dI6fsuO8etNwa/VmEppzDiLd4
42apvmKHsssyiWFrF6cXVWROxq3vysggBFOhfc3F72dQIM0OyfC7YIOxj9Dv8CqZ6xugl3FVkcqH
VoCehnbqYhhbhF1WJ0eJdG4u8udlVBm68RvGrhGTfcxtvzzRYojZshhpK9g90e5AX4wmvyzfhyy8
EcFjY5VmrpPuSaDI7IJ7xgM25hfOgmfaul3grozVp87QB+kgbeveuqczg5nqaZbMCeGEG12M6QI3
YwXgPF7Flb3I1ELP+YTaaVFJ7sR0vFIJHCUTk14eaHrIawI1x2bBDp1h1DNXIftXTF8OQdJ23W0l
MwWHnc4E86f86OzQnaG53qhrNXYUPJ7PDmhK5QQN/qPsilIEOPGsOCNsyg2WfEJPSEp0yWXnm8qI
8r7Apat2sqitdEAOkxlVIrthE4cvbMI0iCT3t6aoHylY5nYs1PyAU6h5UvTT2U5YvyciMqzk6SI3
cGrQSeMqpKWDvSzsTEDyuNckdoVT3S3OUH4v8+kV+WO9Z37tOZpLi2gvnn/hTvHyV6Vys4HlAeVX
2PL5zWz6MEaFqwJHjALokGMRbwjojTPl5VWpBdoR+x2yKbEiG99jIS7IVLe9NyoKK4FDQPra44kv
lTCAvjb5NoXQkcLa2/IOJEwpmjKyewiJzvwT0W3zgbo9S4B6u/zoTX03K6DA8fnXpEYIbZ0M6G8b
xXvzDrbNlV9covJJ52jqJaAozPY4qc3WhX4sBOz4ezkkdViVLBl9tfOmR/S+EvmWa5jnPhRllFgl
PzNJzW6vZVBDryT7U+PGnFo+pOy5K6b8meQSBmy4LrGkM2w8PZJIy3ltFe2Y5S110K1v3POEPaeX
98zqsTNWPQ9vV/0caZ+iFg8ToS6cgz0yK4wUtye5jlBrKqPZVbEoEE2oox5ek8yjuGWylYi1FB15
K9nByJTrgD7K5/N2Y8ajhGNgN+gYWRpkDMHcFGOrfYu9vhB6RfG8O9qpWoEM116pcrXHXV6g9T/q
AwwO6gBXqCGMI1ZHeuNNWrycHilKQvxzCbvHCZe3xkwffghsKsuOhjbWi00YC2J6QU6ygOdfyRCJ
2aSViN80FzjR+qGLtJFaCeKJlTQvwThralQIET1BzUZZj/Vd+BiVuQUGtxeOA8G8d+O74jKa4u9g
wT+jSMd309E6w6xp9uv6LCEp+tN1fJrzktF9L88vK5i3VEs7JAp5i28LlQnLnaS2xR6xsQ+p2EHh
IUjtoSEX20hFGwkMEg0lP8WolsJZq/ObT5+Z52OHkzUKT39Z5SMs7vEtFAuzv6tOJIHc8LtriVt2
Dc6mSU/H0D5FEYAYnkKuFWuW47dKUz5IZRfGUUwThFvfgD058n/bRLhoR1/0J8nkT7St+vDrC1TP
EqZOsuL9LTNYSBUWAUbC42rq2DEAaRhfUSchEuTD60/YVnCBCNQaYvz6N4VEWZ/py1SmHI4KYxpH
Mbm4eQU9KfHQDWWnTYpUoUfreW2I61C0wf12O3devPb7T4Ra7DVstVKlLua3s6rIub+fKVTAvdVF
HdasxEhHDuoKsCFN/6/NYApzgOvOa8bEpzpEcjqJRyrofysCu1XCr5BLknG7YGhKEE5x4AquvVkj
TXpQSTSj8qAYIdS9aIgYMvMBSaF1YWr2Jq7zP+6P9lwajZa5CGf6wLV4Vndk+yTNdL5EXh5uWpRt
iplP9lu9MM5mOeXhXdQWOAEgntRw9tdnxAxdGsRRoqLuQgHJ13YWTCi0jOKTTi4tNoGvukxi9Oa5
+ljh6b7v55ZXH9sUS27T/k4zvKjxCXXoFtXg7WmCQ/+II4PEgGU2Pw7+6f7HAtOqkryjpVvnsOvG
oksjZLMkxED63TJ1boq6s2eqjwsPkqswtQ5L+6i9oYGnezZyjS1O1eq+EcFadYpNFd5AzKRhizcv
DUSVycZbPnbA9m/twyLwsxKUpeBOyysS2koTy8xTdXiSLC6GS2VRjBrC9aw/B9U/ixI7GG/66E3g
VA4h7qTQM6qbACbjlo0KpNI/ttI8otnJKDHDyT30fuSEacLiB/nypYKKQRdgS8MIMzjumr9d2nBt
ulFLltTDNzyKHgRL/IHnJ5IEEkDewzXEC1oME5dBkdVz+mwSBrcz6Esq5XTFeSkt+KnTf1Y5jw61
PkjvYceVo0kDk5LxW+sBbpxZPlXbu5mME5Ub/82+C4Lh0Zto6GTFvVA0JUSBVBAU2qw+EkQ5sgKN
PCLNSU3g8d/qp84uynGzIY9Uj1yYihmrnoHrdv2JC01oYTOrrqnFtPpq93kRmBaeA4DIJD75XvJE
8E2Dz6+oXZv+AvJ592t5b+Xnzgp0jylxNQZNTX0/CnzKx5wpM1EPEfcjJmwadVv09Bg10IhbAN7+
Tt9Pw2i9ALReYyjOKPfvessFao45Qri2RRx7DB0YhXRl1clekgTg/m2yHEAUyWnUrDe1kWMYsRb0
TN5CZVB6dAS7BUnOfWJG/cnr6t3qY5s8H4uJWvxxcAgw64+Ak4A5rJ8Z/T6IShc9eUbavj1gbXTm
5pD6gbXV/+dHskQs+1/YS0lEF088qiAK2vLaG1EKU8FAfGdL5Lbur6i7bElE0GvkRvZeLCJzX0X0
7epdrSnSi/CxRvDaiaM4UHmuXeAb8NthmPlMX09aWIapGWLpHIwi2BJb3u5kyjixIeMMXXHXi3Mx
A+y6cFhQBhvquoDasXBhDGzNBI3c4iZwZkyv/+mS02VnISZGmo4dPGINJgBLqmhEp/qa3LUrjoim
oDm8YTyqZdkMGEt76CxnNrpYseMBS0MOKgv8fz0Iobmi+ubslK7NgVc5Uai7Eml+c1nsI8KzSFfR
um2LQ2mWalqN5jR6EE4ZTE2y9YFRTNNLKGwz/YD+0wxrkWiBvq7CED58vJCggwHAk6wzEV9l9JgZ
ppBffzcauZ0/ZJR9VFKBnuv1X3d7nejRezOc5dJKC43Axz4/jOBdOYVLi46J1eoyuHcButTtaZdj
JyQat06G+oRgfRhkKuof7/O4VTou0ge9zHDLw80tfWJrKIVwA/m7EiFmEjQH11AuUxZhsQsvdrm1
zmpPtpTgOGDSw4WEoZKUnLP/6dGuqk6gcB88DKrXN4WaXDPVN83QBJ9AeMKP0tzAdQNls6jwfJ87
Mio/1I70cfb2G0sRhOX4TZ3DZ8Alypo6UdoDdrmkV8vpxB0MMRSEL+lp1tKegPF0tKB2mmdWHIDK
8od0R6EO2jyoQlAF2FdLPK/A7zcCRBpBFfc5t5+9lyBLQat1NRIqS0fAvlbW8Sm/BRo+t/W6Ztmc
q0xodV54dxMlwyySJpmsG+NHjdhPZomLv/ialv4wtaaaf+wNAt7NGlbOk59mZsImRnTG7g7rZAja
uCoiC4BMMsizuacxU7vOrlEgxE7H5xERBPPfwtTzyIK9j8fMZ6Dv6RlTPljFCEUHUz5pO5XlNUZ9
OjinBnkMeHwUK8ocE1/sNieMxCxymlMbei01bhJXzMGkypV/rIWJF69EffMRAD/zthMWHnwdFStu
1+tbuiigTdIkP/J280MhExeXrcrpNUbSAoqnvznUrqbnzXC42hoHyuwGD9bFfEKDcBj/xZmZLDLg
42Cxmk4+bcPNKNK5NkicM32wH6tIzw/Uo9JZPPg0Ml+TUHfVRQJO6lqI6+fo5Y0EyB7f2W6ZpXix
Pu8y0m53+uRwWgeRaTKdnIenZx6OhG0iil7+2aS77IM9RAflqDulAnPJuBVZ9gvVQ+CmODu1J9nY
dSLfJSwITKlcAWKX6gorH090DhfMlmfRBElU8hZSDj4pgQ64IG/2JGNL4D5844olPeDL1yeIIDm/
0YkX1zQu9koERT3R5f0gyVJtRSTy9iMi/i4FDdn+k5e4FROGTMNyibVrSquCEMBlhAeeALSAbIg2
vyNy7anqkx3X076zksbVTmQkcxJQ30H5S01pPpZEVU3fd35bn+WolqmYaj1sIPtkijdYdeSj4JsU
AYKoEdoI6oRq8ETN9WeNMhuo3KpX521PKLVabvFigjQvE+dc7GaZQWWeyh4fDsTiAroei9Gt4l3L
1DJUg9s85DE5VgrocDlTJN+sN3yCPponXiMU7p2Isq/1kQGzxYNr563S61aH5HTh+nGhY8qS0ukw
96HzvqpFnYjiSF1KdvwCjY99N/RQBV5gCC2KLx15/AAXdyteq6ROZzkxi97sv6sbX0cK3WV6c3lX
SjN3iZE8OcZQw+mXFtgnzTnxWVl+Z9kOteDeksqi6DezdpqokO/DF0SogTD0qIoVG2DUHRe/Fqex
LXUxagymGbMgRjBpOQCYtE27NWQ4JWFewtYOJFS1dOicKAXWqABPJTBhPE6AdFQQ63GKSNkXjEby
nHsiMQJVoypn/GZg6GWgbjXhqbS4a9J2n2lnFNCIDj2Dw4RbEcG+i122GvDl334htMjU0cDpvAa9
F8DAG44D+inqlY4iMnuWpqq9enfRU17gHY2QXrK7HysVAQttA1xjlXrtR1gpYaAgk4LhsTiEjVbU
ZqSywkeb+VhuvXIESgZo5TIcXskT+Lg+yIP5RozgNhatFHMW4v8HeyVMaM/ZDwpj763Z133c1OiQ
BzojrDVhm1I6SlMaFObgVXzjLPr8D5FonTIX8NxNjvQdlG3KzmvXrbgF0qvPkgqYjq4pebatAPOa
dUsKASCP92ING5mCxc0Du7KQ0Q8E0A5Nqs+EZdQ4CYoLv2cgbafEvDArr7dIe1nmZ8G/Hfp2xuyt
NfMSLSoKnnQcM4YjUwkaQrP3/I4XBjQzVUNoaEv3NqCNnuJHwx2f0YTBFTRer/4ToI2m4R6dF2bm
QqwECcfJ66eUgp1Rw5Q7xrBzY2HCyLN/FhdbgD9QrTg1f4b2cUNzAeGfHjV3WuFbeJRp/V2UG4U8
7IR5XoR0gCpx/Qi4d6ewm3p/wS8TvzewXjMpGwZ96zdlAqI/R6ADRto6NmMvSgW7F7Ce3gsu/eYZ
RhjpTBVHdsOhVg8LJUWlPYlXb2/dv/Qyv2CwRM5C1ZU4cvpuhVVbirt+VWe/PGBd1Jdxq03hDLnA
P2paL21IM8+MHwplFkpmrr3sEboE/bIMPFz4VbvvknSR1Foi88eQIqH1cYPwudSsIiDtZKiramFp
YzizKoygjJz6pLr0zJIIOvIGotnv+gkpqPwjoXVXhHkoDuA5ZpzOwq1WcherUSaA7ompC7Rv0ijm
0oLLTTkUcKQ6zmy/BPRd/O5R7j37WIMwfVwYjpbA5TJLZOpuTsuaDDXvILJVQOoQd5CE6X+g8Nwl
UN8086TTLntn6IIVV1lxWuKTjjZlv4620jtHI5czklUf1g4vI93H7vEhOjkVop13WQWKvUeT6b59
KNMa4Jb0dZSzHO4N+Jsd4NN3CmjHPawSsAAbCjJqOczPtLanK8cnxFFq9wUE7n48FOsuum0aSJ/v
WFTrgg22+aNmFH3mFOAJMrhaYVIpowXHXd0Rh1ewgb/hnNODfK/Uruod4Gn9fJrdTIfYz9bStUdi
qKB1PQ/TYqHqri3jQgnP+n4CuPWyKoaVMXrv6alFaAfec3dTDi0NGLMQBP8TiSHQwPxndBeAWpmm
581VhsE+X12wTdqazlcPfL4F1kbi3rEHQItBcFyt91EcMLkIMaC0SG5+GeJ8700E0ZMKa2PAQdZG
BG2BANjDmWDtDjTYQZF+8iJmB1L5YoiFgkx9Vzp71ECCBxoDydLQSKSmzmg+xYlPYGqYPXt+rr3E
cIIF3eya5AZGL0THCn5L8msTqGG5666VffkSa/HUoOvtak6WSpyDrfVr1i3nKz1S4xs78DLg12El
aNdfAqAJx7ABjcnVzPrKaoievG5o+Ta4gNzYHBq0P+wcuiWlV5nWGupAwUIlg3Af1wcTW8hd1uV/
O1i3VWhWD7wuElF7fPLe0AB1oq+X9prgydfTkHBxTiIBbrwlXfNoFlIKNbgvxkNO6Cc8TzLpb5D+
eCcOYDon2kcNhzUaoBW1VrQxibIj0LWzCK7/4aswD2wnfT+x7P9hPp/L+lBwgCee9u4xw6O5FYug
1OoNfNu/S6Fkdr959enUyFRtyc+95P1vQxfUXp1MUvfvGdUY6OP4B6qNgdJ8ha9GHhJYOi1hbviy
iIrJ8PS9ptTqLnMtAmsmRuSNhYSqohHMbYwxfwXsGWJzf1bQQ+yyzWy4yaR+3cy+zkkNvqwNCB3w
xGV4akl6M9ZcRRPOzozF/toRoKRDrYAs8bZ3DXrPV8LmFP2cUInpbg8fMB0XDkSiiLt/LML+zsns
PBq3TXNPAFTeoyWR71Rw5o0J9MTZNOTDUqHpLt2r1mBROWQSP8nif0mjVgKuFWiL2MoxUnoD19vC
vQRfImduaj/lRJsVScJUpLe9997iFNIEZ+prIurHLJDI2KoG5AZoTq86Os9HtJn27U+v3A0NTlNA
0k9mZrAPQFS4yThTb96FR7MZSTNaalHZ7Q6L1BzvcbaW5urjSd/opqwKshmM3cV5Tq753Nj11X4V
OGBaL1M54QGx5u2J0qFHGEciQZeW+WKSwD414xVs8tJ3KM0Og/y7ca4H+DPcYN56EtmrjEQJITQx
Pv2QA1gpF5TvqGRFJt0ffwU8F4Z52YT6NBryEgYYPTmhthMt9jD9m8R5plTxPQ/WPH9ncu/kliPM
sZrVksPq9gaXW9SHEMXNsKX7HhHUi5uWgjXFxmgOzQdi53cDCnuY95fa16sG1PjMlILWHkgpfK71
Z5Gx4O1wC4fNptPFSdECi1wQxw8cMEZ1mhojGqGn3t8lxVzLSuhqTiCdRm8T1BrGduKPitA04aOW
i/OV1kU2zi8XGEwG82QX4Q0qM+hIeeTgLkDZQ/TNiIoquhbIXIiVehVaK3k60uY7YKBLJJAxErlh
/sMxGcwrQ+Jb4HiZjvMBRLmUzxLXqfQmDm0mkKqdTTCkPL1WqnJxJ9bawDzn6dhHr67sMLvxWNkM
YRExagQGseTO1XNu/Sg3kZ/wKnQIjVlXuq3yXqYz16fpUUcYU0IUijKhl9WN4hbGsXb+9rzWKn/D
sBNdCy5wl+gAJHi8OBYPPXftwlbkaZio6YaJNlzEcDkN+j5hQhjKP3brqWL2L1XImEFHPES35G0F
7pxlliaK+on+EUi+4KfFwFMx2GVIBl6dlZtiF+GInZbN31aMwQZ3adDzFVeAQAn/2qhNn9cM/2FI
mntCixfgL8IC0hhwO5+o5ndTM8vJeibzdUr+y/B1pzVsXnUteoe7KOzA1oCSFLLpfLfWmX2ndvD6
KyzacNEuy4WFD2FDKuNn3RPuhMnDAAe05gARFAyA3YVY+sPfnNFYsOUar6kd7hYwzK2G1l21kd90
RdRBa7gBiXJwfA9I0ARvnwvsiYJz6QOMQg97djObtOl2H38Kw4HzQEUKaeXTpVoKclBp13EQKbfi
E9ne4F5AQHdkKfcoQvYM1eD/MOT4qyzU3lKaib+SJCdwlMSVVnXJ4ePo9rjLTo8tYHYxBGsnJAfp
CPJsAbSbYOQl+e5lovuD4Kp1BZuu91J0Y+M3xmyFDkzmVZeb/AsSntvnoFvdwX4GDRMuN6Hch8nV
lNtZMIRXA6lFKWSiSlF1wJV+s4zuM7KZLj2JWysBBEzBLBgVyl0a0kgWcrsJ6p1V0hKBLQki19+x
WTJlmL/uHAA2xpsjFkiTCECT+kV0UmaAT1PPPMZrK54I3yaIoZ5eLF8j6j16B3s8EjU1fTMO8Ahf
FAsRaKC2ioSA0fwXdkHdrTtXDMuTWgcrS8wYIu4ujz35cdYq2R07PTa5+M+/thMiaF55+luMk5uE
zQ1U1p3048FVe7bJHgGynkOcpPwyrPP7tYWaqVLTBlrT6o1jTQlD4UOS8wGfIS35n7jwHjnoFZyf
04AebxdWQOTS3IqnZTBeXopjxHImoKD/zXJX08Wt4OfMSr7O9T78Bd2WhzM8JbkMhK/G6gU4dgKK
3nBgMqZnUvYTkEy61pzeGdax8JxU+6QLp6WRf9H0dUA0K1Wasj4Pnks1NVnIsqwqH1L3C7+oxQd1
Z8AQtFbmAInSarkVeFOxj0NsJJLNkx8UxFRmrJzqnp9R/rXOTBGf0IbZOzbkSvhs1OHKdEbmIV/L
AVQL9nvr+OhVCjTTVBb3kI4Vd8wbP7PCOLMWVog8+RSreZPaoiYGsoapWUWJEZ08vtBxPfrrR6Va
wNv+ttBOOST3E1DSIBaVAnyP0zdYTpolpL4gpfrQ7UfeUNkxD/Mshl5YLxOwNgmsFx0l3VglcxpC
YJdGs5AlljwaxxDjQChYCt4ATBZTprpBVhQ9cbMLjOVWq1+ZY2nt2zQI9ITZMSL4WHJC0lwIIWnq
Pn6gELnzWbneWL8FxPim43cqdWxFUPD3pDxhHAJSqLtbmUHhgGhx8MHJYfXS27BGfK5glGwM0PRZ
0Hc7MQ+A0ve0TpX8FcD2J0XLm5OJkIhmFjYUoboSN+K6R0n9rhf57J4PZ6zPY2F6wOxGlZnNHHF1
n3SHMM5qUSrLPuF3PVSJWJPyHUSnEI2tr1LPPAJ8swjFiVcSdt1RybaRs6Nm6PC58dndGAKGPuLz
zO8mm71mZWnlll3k+Dqh5IJKFXkCPB0hkijP6hrLVdH4xG9m7KHEBYhesfmDFeKat5B9cCy2z3aR
voIdn9z7hgnlENoEdDCGB+MXIvxItbM1AbRNImXJcWSJ8eWjm2+9HvHdViYWPVnQStk457KMkayr
u7JYDLjnE/X02y3siDlhLiixIhBUwPP6/Hq5sNn1T+sZbarEpKIuQV1ITW9L9jCZiWrbctu71RvG
LSWEYLwlEyFYQvB82xM3Zr4VronlCaEMYSrfjURsl7P0lmk45+QWJI7r9FyI3Obl13b2MNUGJY6P
ee/+mpBWBVATMbKdVnfAA9GScQQxSluLULQzMu6ja7HaDAU7FmtpfSPirc3MFcrAC8EbQRmPl8A1
B8lMNXi9Yfn0hx+XLNNiYXGR2OmM6kQ9ph5SAFzHIXeZEYZYQoMUK/ye9RDTmZkolY+XPBzGWjle
C9sv9ZpJj3VJNvShnEtEgq2NdopjZ8Oe6/W/FIWa8MUGlSHgAMqzrpFwPqvt7Q3IgTdt6Od/65Kf
Xlb3eioOrrodnp8p1qAwvybAHIwF5mXZDI+gDVXZpvTtN0wfhQeHJ4i1k/opQ0in49JPMtzkenK+
vDAYgtaepw0LXhd0X9EivkXnqWQwBUzK7t/hfU5N3IPLIjDCnFDloorD/S6YEUjDdTLZYksyLIpS
xuOVPNPJB1ZGsvxmC5QQ7QmDHSR2OFehL38FZSSnF/pPiPgmz6DNNDat8cpFVMm1dgTe5K1Xg0Rm
6f0lye3Ru7u/eQYScQobR20NmM8WPOfYKTBy+8IQ07KaQ2v2ijvwsoPu7prgiyssIfICRPrt/zXf
IjV82AKN8poQMLdjG3hurxpwljU6ZvxQ59gAjmcj+biuhfxHSJLriHPFgsvoe0oCs+tvhyD+SWd8
JtbKmsybxOzngD5TghYc8KLUs93HjhYF7GGNuRJZ8FGLOB04SRsAy5yiflrytyf9FvKxpK1XVxxB
MtT5AgbFefxX2HBJrtiUGHA7G5Ku956BlNSWcyM+pcKhTHOgn/6q9PU3vKsKYUiqe1tkPJWNP+H0
HouqT8so8OBpknMrGg1ybRo8cLLG5Xch5Xl2Fa8JZJAQY9CNmb5Px4UhWF7vacQXhiqfNPu+rxnQ
jBTSw4VaIPCiqhPd8dE1R3Tw2oju24c1hFOfLqG90MOFfcan0vA+Pj7/dvAPGmZ1DLQ0xJRKz4LM
VURrMx+0RN7MtgTrgDSKZmG5w9BpF2LuLVjcESRiXsIc88/6Y9GuoBB7MgYojHzjiGshs5mwo+c6
VGK1guRKa2gy42KgACqcWQpaSKRvSB6zkTQyyH0mo4DcCZJ2on/QcxELTVw4M2uTegbs3etQ66Tf
kuAxyBBIn1ByHQLXVp7co48dB/s0YyD3p7NdEaCiEkbvxno4zcrF/Ldf+egC1SqqK6IjLudVzhQm
ZVQ48+DTpXZ0MulWQKq487n4C8PZhzIKgMxgmqBvcpuJYa9E2BUiV872fFxn4YaesaQV46PqKGGt
ncQmvdMLPxqKB3+6Ps3YspLPeCDcHjyI54qqiBhiKOTg7cJHS23Qnd6ja0eH9Xf3Yrk33vSem6f6
3Nto34Z0WcMojCuCSn9Y075R9Yz7MwxN0YgrkRjrngKrpp8xuc9DE7O49UvAGxZl1c/POAWI48cD
Ri5FgCe4oqiEKQ5jowRhI1ZnGWetJvq26cPaxO9J0O7HP8ApBhy4P5V/iFmSGC3MlPEZStQvMYmB
NobXhKDy8uA78q++kPp2VYwBldkSH+usByIsMBkmHAIr5RfDSHVA4NdrQhxFu9jQF+Qj5jqFIxre
04miWXax3mEHTr2r+gn7NvHmKVaVXNm7iOLWpB1yuhGF/n+QdUdk8NK/z/u3prAiBWSTRCGBcoou
LkDmwYb7Fc9zcbN8bk0BwYEpJfy9+k4+2HoawDy613uUxCz8aKR8RhLdImENByvJ2iwrjAW8ZhzE
IHsmT4NJrmCwvxg63jS692N8AXlwNHXoeRS7I37bv9IcOjes/s/61xKrgfvHv25wLODfKYDO48jt
9wWBjrlN7Crnm3ifPH9CPsax9/6esGuORi4px06mKKcr3QBgziipxMqa5UDkBKxJhYpjAWEYlVRZ
5k8/1nJR0EtmjcvVF+dH7mP4roqodPK7SwrB+vUQRH3TkN1MWpvY4ERXhBRdgk52H9YqyJMe2u7C
/jFAYqm53M93mD6QUeaqcCm7nZWKXJEdogn6D5Aj7CEWGoFJhSdCjVeiKTMfp7l2RixMQXfzd8Kf
5R2Tnb1zi4TMwiPYSc/kHiSLTx0IxuCwl7xaGjrbYEnMcXOnSPVPp7UKbssMvIV/yZzwyqaz/S0T
LzbkNVfk7chD+9AeSt0MD8MKIK+vo6E6aXHYPMwF+otwlau85eCkUkyZuom2ljrHmc5DA0ice9Ww
0vopyipYesSXzmt3oeErxpdZ3fVGw+eGcFVJXvyDrcsP8YT2OLObc5m076o3BN+OhyE81iCVT/Rc
djHtwbDC8l4jRFVRA55CV2yCcTxogAiz2lucqoeWHkYf/MJT0xjtGPAwB+M3zWzhQ1X6wA2zk+y/
12iRyR6IfNafBJuTpuT8Trj06C0cN8QxFVQx3Lad5zwrRu0yDNYRoKULliA5ZuG+0dwRDP/LaOAc
s0uTRcfU6BsSNZRD0+wRhPEo37FRqeUvF6Ov3CsQSRAmWqvzak8Z+A6bgmMNgpLbt8cjlfCfPHZR
b1mia1wIBvNck+985nju+4H5/NLleKF7HlYTeTZTVkm0nu91ZnQG6jOon6cXbYe3/Tn1Kwx3Bm79
LdeW1c2hhfFspuT1enRiZcf8EHTJpXnMok46HM/b8gkwg6rBC0Fbl76TxQ9IiXaxOOvV2NPJn4B1
WDXKdluwC26+iVXIo/Jxz0DRoeMwI+vBeXdnm8ad3X3RoNnzJI74jdkZ8xp9ALF1krBtp7UC9hQc
US9bdYBw9JnCb1iHYeEdOn9j8f/gvLD6YNgkhgNgt0St4Gl01rEk1zbKtU/kBETM/tXhQq2P9QZs
cadE0rw/mRumsQglg+900blOYa6eBoDMWf6stEKNNOght4KYGJaFpzoRBNQqIAZC2gcSpZ6KVjiG
b0YEFjmwvGnU5yFrEQbpj4uIU/kdSOXqkzlAmebvzTn0elWjVQzsWozmDzNsDqCKqIntc/7FUAhG
5hbkDkdM1mHpFMVq4A9iqOlcNmP74SmZ4fzHvn2RVmlXMp2ALofZtPVGDk17cKQxdz/KFvW1NuVc
JFnfhsDaxk/zcp/kFbVUUSqTRGJh6WxUsDu9tKOTnjs2wv+7sS6mU5/tJ4DEhm0tX1nc7TlCAiSV
eoeF5EC0cqyGSnLa1bD8fmlApyIFGWwzG7A0MLehbHv25S+O1+/tglTlKyo0EwVrENGoM6K1XjKr
zIzF8FKakoM7WO1XRcSDhaof7BNPBLaxCRKP+uP1hcqH5Q57eO2lUlEKUYU6ejGizCmPY7EXVwsd
i3dPq5gz+IGlWhGD1l5g2AfF8hSyVQkOC5oP2SAS+Xh/k9LJ2XxxF5lWZiVx8HV3YSgRKVBWRfz1
gd/WtymMiEopvf/2FV7+/O7vMdawFjH2vHtXxK//PV/xp6/o5tntDDJb1ZVRqakNpW8ndWT0EnNm
UhtSnn/waucz2vlt5lFzyTnZOkXdwz+v8p+IOcKvCZy3v3cWQeRZiuvU5HcMYdaAyM8v+i7154Uz
JfzxIgTZ5t3S299VJPYTvB7xAxyi8ln1OG+DWzuTYuwXBBi80EVq6jXZor336tY7P4/9gWGGVagC
8k0BjHMDhwSSIVzcUXr6IhtLeQqaeVlew49DPbFdXmOf9W/yIbPJPFUmS5/KrdImJCfP7DM1gi5v
SykLdUEKEQEk4E34ySJScWOhHDJGPq+QtitrxwMrG9YO1ETHegJ1Gjm82oDqcVNBVu2Zc6qJ3NTu
4ux+uVRYoaYAa+GaatMmMw1WKqGQxctngwr/sWR78+hNVTLwxfLdT2oU6VskK8lxkfG79jkOFUZj
6s0jTNCX0styqBUZ6B2Q3ydmPxhIId0LMtbMF4JY3lT1Ds9ClgPKzRzqr1y9FiAjVbnwIcza33gg
mlodoilp1v5JMSkYnOocblXDP0FJSx9JcEbc8vOND4x4mzGX2Vl5182WQm2hPEPI/haKwaaq+n02
lDypMxxtLJ6AYt9klc8HwxL7t+/YIP7Sy1dQjaBm3lbXOXlLpiJVm0IOySvZrUcKjeBRluzLpnbT
WW0u9N9OlydwYeIPviUjVjx/zIYeIoAFPFYRalbSb3750h6jHbvreJTBLyOXWaIB/Bd6NJprtrFl
Dcccm89yqWMVErdnz3eZE4zS/cwyIWG78mCynEO8rIDKGUhG4aKQ4MIuWBsz394dMfkdXlzuhzSH
RzvPwjdqMAeooeMINot8HwU0JAspar6xjE2Inraiw2Msldx0PrBZQpU5bv78009wTwkqR8Hufd4w
COH+k23IvqyLtEx0h6Hx4TZ9z7kCt//f+rm2S0zLgo0of0kvNlhxDiSeZBevWdOxKVEF+xliT7Dy
ItWGPF2LdLusryy2S5quO5xDFPKZoQqwb89ZxaegDBizjp6g+TsA+dgMcFGM6ZNbi35FuPc/yLTi
JZoNJ/FpKEnuSvLwtulUuNDI37IvS8m2VSDhhENXB/H7qmD4Ey4UitEDtO0kbbKkkEVPxvSS7xPd
JxfsG9jlKtnSg2np7X+7VL61iFoAIQmgTR50t3/8zXyfijSLEoa8nBIyUiX2GqLLgLa1QZFbMw6F
9ip+k4OIwwJUulumDy9SgdrI6DW23nDdfYxltN0y8DZ8ozVEk/mLIPa1xNzzT1xMyb3XE2OTSMdY
YYYsmeOfrSOgcHAJj/y1Xf2rhVLlJSmNF7SpGNotg+SEv584JCnTAZpq+fn1kABr4d2rfg8QpMbg
sTOeEnNcAcuNM8EqfWJbrN+R702/y/BVeMB0iLS+nZOG9wootK2b0L94ZHE7cK3EC8z9+STRrwNy
BUDCl/hL/FFQVBBzinP0Zc/nYDEH88c+0O/2UWLSjRDV0bHTXkxPHfxmOrQoaZluIUMl85m9eTgs
ctm/DjGM4OLoA4vfFd71sGo6AQH8cn+z8jrlYlb8Z9CeI+SbV5vLf6qofS+DCpc0/w3fFdz5VbLy
mjcgVj66ZNBvOI/maEHPvYVii347vEEcKSpgj3Uv7UAVBgbNmDkJr5MXtTsH2jB50fAdskEujD0b
HcIE+TwbxXAXNC/nnOW/o869kr2bo07OTOyLfhBwwf/w7mYj3UxrC/CnG0+eOkqoeJemNAyj5tvS
Ce1UtVT3Eaq1m+EktPBeJTSKpj/BAxKpHSOddvKpbScGrlF9AgRFzc/YtVb14np5VFiHfSsoA+wt
IqOnRoFf36VGaCzQi6sIczyxvsJ9wDhQwMSkTEcIi6g0ptWzai4SG0OlL9uwlNKnDwXJeoV6TDvJ
K4lWaDZ6mvOpu71uMoBmNAFYwk4nibFE2MVWFrahS+ui9TqQD4EHUMCUZ6GUqYuj1GV1v/30e7Ih
MfPltI5QkdtNfIHdhpu435Qcc/hVCAJ61276/7ejI/PKe3SQunHac+C7nShIxxBWlwscc4NavfrW
HY6Gxa2Ud9qyox2xWtdSHrCMfTTMlTt02lKat9Ho7bdfeHT6GC/doyqq7cLBP/c+Dus4IpUQCJkJ
lqBC29dS3mnenp/mwOx7NxCxTT4AGhuFNPqh9nOFsdIUJoNmJJk6mEUYET60VNq3u1BDhwu2ikNe
dq1fc2DJn/oAwCNcBm2mjHCwaOTDiN+m5kyd2o8n7nkGG+jeajOI8QC6flA6JG8+na/S6uArDx8N
VoDrXEgkf9YOe4MBGEyMMLKO7YNkHpw6pJPe6WDCihClyy5E9LGnr9loMMY7NXvbYf90oROEyT4m
MglPmupqTWKt131YJvT5r6NXsoYwNatv9KcjGRYI8ipw+ZC9WKspicV0i+aFuq9PyrJHnpHNjcNu
ZnIf6Y0T90McBqDnV1EeVlWlkf/R1UILR5aypWXdlSTSNqLS25jMTOwZ5ETGiM4a6HEwfhn6EUXR
0NgT3XpTwro20l1JZ1FbBqpo4HXHsTHsuiR+gaeCHjBPqd6W5na79K5zCfGI49m0BAR488D2ac05
iMaUYJv5pwxmkFqPiV5vkBAOszeQNLxDys57qK0j4jt5bctaP5zVRbPnXGDe6uMVV7Hm7pHhWN/p
PibO40yNUreSspWcVa/v1nAQV8Dc41etc/7ym0HXYFXhCjx9QTUDrxYaFw8QFyhD1U3qg17z2SJW
RLNiclDsL0FVOYa6p+0DP9Z0Tcdb2GEM/URDx3/eYsMPN/fYDJKvzlZvC3xk/kn6NwU1l5A+lLQZ
8ITizdE2ZMOYBEPFvJRUmiB9HSpbk1oGQHPg1gOlMsYj4ZL24WkS9OV19FCIOeybCEbeyxQwcdRK
iUoEhhCB/NzYG7jW4ZvI374jDJJLuMnLTpEKqBf2PPi4v5eZwxIP/DnbsepFf+bqKz73zupAXi+u
nl96qi5clZ9gVgbPuDFN7ujrg6MAf9iDSl1+sbCD+izNDZrOVOrlJtzay1DuLZJmnW9PcYRTNbyG
bYAL9Czm2BTrHQOy7uXKa6HxQ6SYYsNeSoZAvOIBjtzbGz+njj91CeXdCMghxHr4916pT5YBKI0J
13biYLwr8j3OnIKCf/xDcn8fT17WLhA3AUFmkZqFqa6yjfMObgvVmtbL06LELQ901bq+hSEZPqvz
iQ+vpklZc+WYm1tjqaSnUk6YWGrJEssQYUIhX7WM6oBq00Ff/fxbp7lJ3y4IBZpXR5aTDbl5jsL9
ASVtN2FDHm6HzuuJeNDkCA9tAwkTg1IieON2ZayN9AMgsv0rt3jXSAhe7Es46bH+9RTnp6+tsl7X
HGSTtZsDMvr5Ys7kGl5DEAhL7iWaenobgVdVJ9oSnfIrFVM8dAmRFfGVa07maNnWNb11ZldaXcdk
wqluoQ3L4f2OpX4N2uC629yVrJ3zQQeByxpWh1lzOOZ7PbxyuyPKoTGFvQfc/vq/kvr4JbHq3Byj
VJjzFy+phXibRjsGDiYoajJOSyN9OzHrpPsfM+xNYPMHptrFDA55uIsz/0xYEYjCfMR+5qPWWk67
SZOXrHEJroD794/IX0DVks9VkVWLN4I6s43+T8vfdA/Z1VXqS5l2En7L2CT4Hw9WxUxSAsjcWBDp
a0d9HKUWQqDBtYu44R1B4e7alrfdcVs4reH1Fi4K9PP4HQuIviIfgkRg7kCRtkX6G1rom4ywSo3f
dqzdp0XpJnQ69mZI5sMh2rYQ01Yp8nH+d+sC53z5WOQ1WQiINGs/htyz0DLx00v2qRxZk7LnHTA9
XMD3ANHUMPGUDqdsTiVQzlLB/MTTgjzBFzVLzer0YaCRBJRlqgANRfp89gEQh7YnlMf5ZTP+UHLx
MBDr3DOQRb7Knjz0cbarQRJwMb0Qc8DSsPZQmsH2RRgOeSVOLyfNKYPPI+nUxBABYmar1NpVc+2b
el8DYTaj0MUlM8by0W7JuoPScoldFSnIbJpG3Zx/33cXCC9Pj0qkrigaC868EH0arLGP25k2mYvM
b+FsBb0SDdLW52LZ59ADUAAwoTFg/JXtLBBd6Dpr9M67VGet53oLclz3hNNRO1Gc6eiHko/gbFBZ
o+SaoC9r4VoL+uL7ZKeczY84Vf13ZfZEVnWZHd5NwYmY+1zwzViLM+VA0jAbajnou/hdyunweiWJ
4tEXbnGiGaRYbzEcNAvYTJlaeY3yQ+IlTS5lyAEDbxGJAV13ec9rFJe/U0Wx2uA0nXrOZmRu1A9S
1PwJIoBIpgorBe/TuInebUyo7Yxq33CrWTO5E7+1HwJP88xwd8/0uhhuNWw2z975ByM8tVhFLsU7
7A+Ghk3B0Qr/2t6FWcCsR4AqlR8BvylqSkZeR/EtNBhiBtRnjmMByME9fnMAFLfbrMcJ2ezo433c
yTIJBiOas+MdOB+qylulI1dNOLfRgm9X6NoCDtXysJawMVtJowKsCU91HEnI3tESyIOy1LV7R0aS
+eIWfNgn0FXJBBP8r6lrOS6eYKiiavXCMASoeToGt4J1/sJKIBDMZ1Qt6M29eoOyHXwjk5KT3jJk
ferFMBHlyH5Qpy/Gbtz4F/5tclqf8QcKvEnyvrOF3WxqU2zaWyU5J5/vgKtqiaHzHtA5bnNnbEns
9O+kdDoCkvCWTsAVZpAnSOHpa5H2gjTsJR5Jg8jAIQlb6zSP7/oMpA1vjsZpkn1uqrbaqC4LSN/Q
FjMMalCFw0ZsH0vQaD32Bu+s3RH8UTgv7BolxMWOx0FnEPb+eUJmnx/KsltPPAvX51/C2AlfGYCn
/kxRoIPRRidT9CSCDka3/a7Bj3M6VuNVXmMC5poGHGAFRXPsm4NoZolzRtUap+4Tr+moxd0+hCTM
xm1KWsPlyxnCivQJkE4SM48udkshrCOA+vO2xOmyp3SjKI2hpHzQqsMMBJH+qxzCPVi/jj1RWYF+
XxkTB5CqkKKT6Lo7zEZBnv1ChbS5ulz1b0iBLWOV84nz7Zu2d6KQrQt9vIWAA38jluwJh8x73E+j
Yyhu6dL1Td8mjHfn24jcSjoY6YGwhRPv61WCxI5kugu8JwUChvXa9Ft4A6Xo+k9Tq/Pq+Paz6GSj
bVMH4JpNbShdHXMFbwIoRA1UVdoAeGdKZIS2hRw+N2x2MRqRwBdOb48SrfkDHr9/bjWF3Z82+VKt
515oo02u5DzlNBJ/C3ED5H19PsRv0t4H3oOoAxarRgAo/VjA+fP109agDm0pYVAdO5WB9kOTvCEz
Pxq7d901xIYlRarAp6hqVDGaAGE/2HqlSBk92s4u6Uih4g4pjpARnvndEU+7/TyJRrtamASy6GAh
BJQPuOW5mKJUqcdRsB58/QP6fnEsdPnkumIRqjzO9brZ2O89UELyfeXKGhnJA6oThI6k49vhqU0l
yNBOWW0ub7d6BOZDMUk01SB78WvRVYLbcJXCKUBaJAVdDx2a+X9D6vwtkS6nRCiurvfxwtjFxDAT
5PaY+f7m4wgq+ecuHeaweiUhzokHrn6q/jSPJosZ0mWSErdzNzMp0vWM4LUhF8A46+lxq2Mg68Lj
nMw5vJbEosnggQy1+qI35lgCGw6ZuKfX3z7zh5tQfTCxywA+Tk8JVbefwU2MBTq0C+c6x4F+Y5zd
C7WcXHvpnLztyQ51OjShtUqwtYIKEXhi7b3VRNnkqDUuTdkTwiB6FdHqVZX4wzoEfKPlhCrWSAMF
vgSyD9/ZXzwyP9GD7Uj4C3K1Sk/6/rxZdOze4OSB6r70rkTWtY9aN2dYcdarSew9s0jvMiV2W/mG
XQqbNM+offx9GaGmMXnz11dwOVmyLO1IV7OBbKUQcVPeurz3f1BWzfUgKKI0lzQmV2RhKX8sGJb7
jkb75/jpADO8KEybrtMVlRBH8MfRHMGkevTi9q5CAPdYPH64xpuq4RyupSQkjoS/lrntpSTcpL4K
Hoad+UYQZIUtMZbriFZoOI/Ejp6YfJogimq2lVtgiiG1AsPGhlA1fgORAYg+ELVKYRhwZlCVwKDj
xcLT5LwFTTv8VXEJJ5yxzA8tj7D8YcB3kfaNBP5Yp+tQ4ZpE5e0wf0jnb4tAymQQKpAmmKAbTCAh
Y5imYx3oL9iqFn50aGI2Sp8GMzzQAw6GV6L8cbTW2z2Vya8wk265qH7Fq7U07fRfaH+TV7zUUvoI
pRMCyp9r0Wga3omGm0V0YjlKFL0WbnMCVVfVeybJF+80xwou2bg7euaKotTAKfa8E8s+I4rfMIVW
uVoOewLsRvoTLOmhO46jkgOoun6YybISdmysBhHAwLLuDxRdrBlJyFkeRQoR2jjKjJ1n5JmgC/0F
oHdszOh/FA3M+pBr3QJNs+duAqLLzvIr7pXI5Kl6fwaN8/HK9dz6zJVadKf7/66Za76uRFml80vh
vPTjo8y1haeQSQVEiu2SWts4vlY6+a/FNVmHJ+JSp+zIGKSBLo0RDTJUBtJUZyY2MLX3aepbxG0k
yqyZtNeSo+VtAI9iqhGvu/p7MNyxteVu83Xf6Xqb5+B186bfJule/y3HB2W29dRdkv8G46H0GxzH
jjfcEWNFSEBHot+fRUScg9UZ7IfPerC8Cd/1dEgQq7e6L/450ISicqr4sNpvpQdeHw/1Pj4uit5f
uGG9Lxfj/ADl/H0Sp+Fazo4fLX5DttKXFykbcxLl7N2jVgsXl4M+cuGHtK9IE5YkxsTtygyLqWz3
ZtfYnq82TKzZXxJKNK/Xv8moKriATBG1GJXdCdDA/L+svji4dJp5zLfrarRefMevVKw4wdbj80md
YoRF8FKtATV4bqFOHf4wvRTnnG46bW2uAbrv8OiYzn3xQqGn48plMsbEqRb0qzjpjQP18vU3dybu
/lGzSsvnhnM2xg+DM5KxUoveg67rOfAyXx7RHNr/Rqi9XcOtRBGLOq0DWeWmdhJzyAIgCq4OL2Qp
Myyy7o7k+9YYETFvY+AYUteOalgXz9okn1aDZeS7Ax2gwsxpG6JXlJ586KaK/0n9QTuHFLMzmG9b
BgmOHFois5sgokMOmhgpXe4TylzfogphBm8MwilXGiUOmErRLKdyGkf5YzqoBQ46LjxUYLrjYimj
km5CkmBlxuFk+bAi1Y6oQMLVqMg076fSW4DF8u/x2owxeHqChez+/M2xJpDEMUYikS56DQIxTYl2
t+7sYlkGOTyomDXlb9SIjDb9DPNc1mgnD+AN3Mvn2lMBpONQOlZfZoQGpMWd/3iPNyr84JAtHTsL
GxueSiYf6t4MDFyIQjoxEnzmvzJtQkGY5PgIPv2BKeo8utQRk0fvgSwb6NJFMX6m3yTFQr33jr/F
voBrpFS5j9yZE7KC68DrJZB4GgrH2QJLEwBHAweP+e7V3k3vL4Si6lz96VCiRNou3DO/kVSod7DM
eVMxayA2hRyBIptg+TYiprk48cMVfM4E+APkg61PLDprJwuqliELE0WY3g4nA2bYB716ji+5HC5n
0Tf5lfXW59drgo4E4ZKWR6KsyuYB9Q1vNWrSLLW5u080eud9B7uQhdtfp+0JYno85etcdDN2dxj5
k7sLdFJqyXdMsy6QQn+eKkC+FkCF+/X4SzylRKb41bJfKEKVHjYDq0fv07LYESo341hN7Lws/g5L
/i8Ye4RtcYr9IUI3cKoDbuUECI+y/NUuUiuO4FvR+XBK1ANsZlaVZ0Au15JkgF0Sqcy5gPa8wUkr
M6Nc9xbE6YCRzoOxjfDD/IKZUbBYsmO6VYUz3jYzj9G4QTCfygthK7IMtROkzFquTEauF8ynIa2h
GjVKrkD+UvpZ50VoO0F8LJS0hc6esPp39F80EWhfIb2SyrwEtrCt+lM3WyNBoBL62F+olo61+m0b
+lZq/RehcFonR8PUeI1Eas8e4X5Iw8mhri85flmqnuT+69xtJjIq8srRNmJaTeebbRShXwgmueSF
FpqazUocJmqwUJ7HEILBNR+6V332WRPfP5t7IOffS568cd9EcqAiUhWCvjfoGBEbQZF+iTyRO/HO
q3jWc4ZGXuo/315vnqQslC7GYEJYOUsh+cJeijr6u5XhvKHfcNDdbMYi3Yv8vvlvWo6HM50sIA+7
Ipry7mQRNWWM7lAZcZ28GR9IeTGV7Npikze+sieWBW5JfJ1KsQuhsUqPNXMYzL9vEOo17JHGdJIn
exzRfmxQJPJlydRBhaeDuw0ChrjkaWqxxTWuvf0Idcd0c7HUxDt+azFMqHCpizi0wnxqsCRROn3Q
AFjXz3uox2WuKDcV6+qjkl+JZ04xUSJp+Ss+jvfBWf45clTrwvZDNpXPu6GSy/iQdJkQ2Ky1a3Gq
Q8nmNMJVo0RDf1zpHI7IdqNOY/WjX1r9RoU6eN2VL1mkV0TTAyx5ygi3mtKXy6KBX02UkAqdZFHL
Tp0kaPOBvNSbfSS+WX7VnPbtYTshAdvuXTQYdu9QToMJfUDkRlBcxaFoI12eiEqRpSRi3LQTRuUd
xHNZS8XLpTfqfKybX+lCtBB5P2LvYqyXNsdl2EV46a4LERKDnvodUx7jz1GDLqoXlraHt63z2D5f
NPH54SGBP4U4ZM7ilUWLZM9FN+MkwMmdIfiqdHcVbqXcQPg6Nf0H+iFGVVdTkvj+pWMuI/OKldlP
dCutdhuvHhqR+K42Huc6MFl3H8Ju5Y6WnmSkLzS25Tvu/N9lJW6wRPxvSUg5dtp5LDBpWDJ+Kx1Q
4h3epbWjAQdUYAB+UzgoBbW/nuw9VomGaYheybXj7pR7J0cE0fB6FsvWX4xk11jajL6p70FGyHUU
/4Vs8tHNUqOzHZ8mV4Dc+5vuLD0zkCkNIJnnRXyx3Jq2UBfsx0WL2jLTBHtHbjkaw8I41PCkSzSx
IJSEC672q2x+HXZP1WBull9o+w4RDh6sGXDivq/GMrWEqRvKQvwz+ma/xmyjWzkh/RVVcky68sll
dQVzVPe0lbnuSpb3XGF912bx9CYXGwGYttzReNXGIppZDEoz6G8hqcoiQbfkH+nP/tOrCzL9vxq1
iaZPVXXDk0Iu+DbWC5Gs66ItSi49lJhNR7DdCDK0ox28T3Ugvr/Ei5pnfAFzt6lZ+QUzZkBTB8AM
OmlLey3PUlXuzu9bI5s5OPqsV8v1BdZtVw7+b2iDfYXIE81m/PuyaBmS8WXVjn51c+e8hLohGeMg
U0RY0j9oNYJWu0QNbohi7FjOqylqaWUeGXpR+jD0FSkZeOeHqnawm2Ahm5pprb7JryWDKbq2C751
turgFk/8IHn8hOJ6nd54eLFkESfV8mwfwDLCzX9hL4Igg1Txgbra+KBYX8dbfOewJb9gD6dDd+NF
QOJa9Acoc8u1daFblAdLgtDgddkxWrGEumFJdqBSsbqJAeT0GFiEz643Q/cc8BTwE1fx+y0R0tJl
qfvk83sOKYgusBo7O1wOLzRAjTNY3NK7urxjGpU/Zozs44161ljXhmk47v/j7/JQq2SZFxx/dQeb
nVhtpR0sS7GbLOocbNaxuMdun/LzufF98cBsPaLsk4fwQFvykq/jSTxH1Fr2wwVfOx4tgikXXlYE
QQHexxx9psMtJ1kA7rsnOEq/0l06LLRG+lwQWFbSOgZJfVjcTTOkH7uVZvAVFqZA7oIIaalBh5rO
qYjIOdwhO4EqcmHQJfavwKckxq0Rw5iYPr6ZECitnT+OkuiHD6Pp/n+PJut/f0cV39nGgUsu5tmz
nofsxv+G9cPJmbQMUEUyA2Y+4ENXGYkl60SRGRC5FWmNLYaZe07pjvWtHGsamA7D7uIgqz6DyCPF
llwbt9aFKoJpswwwbBa65U3eaF7a9YBdvO7Lvh8pZ3FAZGSqtYINDH58oz+5MzqYCYZOPj2EreVQ
XvqvASBbGzw1jC1PFtFB0fEMvVyeh30pdUPwKpZQp6UxWqFZeJhluOLMaZm4huRFasaq/TSI/yxI
CbDe2lQ7xYW4H1iJnx9RpjuMb2XFRwpa9YWxDIjAeuQlZ7aN9AqwEmKSVdWksBdwnaUOg5SAzk0i
2Vqofynw8oYhhE5fcwUx5xcCAEtwgBmXyEkCU7tYBDaG7oTNvBEx3hqMuuCUK3u4WQgXwyUF5El6
kj+eyOjxOi9ZWnkw0HCa4/tuxgsKAhmHEdiMrC+Ef96NFro5Jq/BKYTNZI/W5broEIquNEJ+oDp2
xxTmmT4CMJaRWAplSSvgNASz8zdaIops20Yvo9wbv37s6vw0XGS0pj4f2izCDFFXqy1X5gtDNaOn
lezY3XqRZz0WFU2V7RMducVcuoHyI7wCzTpa4vz6v/NitSw5PN2k0A/+5UVZ0b6TtaHDXtU8eXM4
o8UTzEmMBz2cOO55PM6eHEFrTxvweR8JTxhhJetv5pUS//myiJm0pM0sgivHLlwrlQ4AKAjJQ25b
WyGL59vu+DcVEZxPJjODsFGRGUof6FyWXRFl2qe1I0APIru7J5HXS3N0rqFIeZsbo+zEexpRJWb6
K1TG11jRDbE8bA0dJgV2Ec9cncwRCvdNVkG4pn/Or1xG0zTi8p0Dr7AnSweU4cy+Y/TqIABct3fq
2plN5JbUDPpjutfUdJoGhvLCDkoFtK3dSt56gSrwZA6Q/IMwHnYS07EkiDRN0dduIP6YnimFPKF/
QRmGHJJzXSsEFySvFplFPy4w88lBoZ2OzEB825QaA3Qnedy7AVnm8oJLfRBI59t+CuKrob/p3CUT
/Cnqv7hwYfHC0UP8zRNlJTlyHqMHeEl0jFFDsQ/GDurYEEhtgZ1El93nf/HptoqDVlVAnstXo0X4
UzgFWW8sBHdLQbeknJi0jgjGB5pOQtbsDZlcrEbffFtYmuuCnB7+Ej4FW71JfA/GRAW5Cr2gewE1
5xmp6qTW+3XRvG+PwzvRnH9Udp8P9bm/7N0jnSpW93ZGXx1jXOIbuSF5s2Ky6JKBO1pzj7RP03NN
zICajI0nHR4YMLWFI93xLPZvz5M3T5UxQ/SFjtzwfXf3ICefeyay0A4jxmIPJYDWY0QBHLVPHG0G
hIbtEYsBeizuhAE2ht3oSehXDmNa2FFaorjTpA5B+qrZsYYhLQ2FjAa/8TEY9LtNlcss3uM55+pc
rI7KpCMMB5MRxNjUWePeJAiwgdkjm4M6ErB9f05hXTv9X2UW2U0dajSRAPGUsSU+OLegtRAsa8Ez
18/KDASusOUDT7ly84p9bOijfr/gwRlfmwOQSSoCbkCPWN0dvnnVCwrciU1RPbGJ7O61HU/veOCW
CVnpU7fNjPFYMyKeCHwbDwjxt/6/f/WFW1wT/b7kF5kFgF9ZSCf8hT3sprSMwFymJzAflGJmhaGt
3tEsyziMlsLd5lyyQBVQudgSNvLAOjWjd4l5uRFx5lpj2LJRSr431HuGv4N3k+eJeExkwvY9gFez
MspauBmFSWrN0WuqyEGL6DZX9EQRk+E72+MbaImKjXLexJhNcuL6s2nPWeEks6MthmCsPplM8IhB
tBf5SLI4XBj6U/jseOEpaxz7Q/+ZNfh2Gpzis7reC21LNjiMMbP+6LfZIpD38akOuweZopvQdQcs
7hWaYBGSAW43Bz3TO9saPQSuG6jLxa6QfaqL/b9MGzldW0FinRLYavlKru/VvGWsj/pm94gtL+0g
p8X8PUxlkryJCghj1dyJ+P7Qf1fmtxqB9g59RxWhOsnoHCTjr4JldAfvUHWO1yYgF2ue3+b5fdMS
EwbeL6j6kMwd5hXm4JIa1pSvknHfNCXtIh1ua1BEX/jNDiA2TSvpSWsqRf1cugZp/3xk+uDjZdr1
Yn9Zg8gaHN08uMk+SFeFzUGmszbt+ZOyIOB0fOQqfO+55hZ1CSuZFgyJj/95yQpb//MDFnB9jpzI
7fmjhimdeVb/CDesseZcPPDxP7LY5cw6fEZIeL9r3vSF/MIR4YotkUKhEPpB419AN40ElfFfiWXW
VWC2vJFsPYVnije61kVmcVfEC/3w2V0O9bJX9OE24KdZusGyQK9BPxXy3UqTY/EMmJtLpcnf2Y/P
BMO/kLSTb6lK4Vw3SVIYPIAPslHyZSvzfuZZGbJppPl7l2+btCEOY+1+RBsP8lgfcR/BZQQ4c85Z
mU79OuWgT2YX9a5aq8kmbUl6f5I/yPJx+q55Pg25WvRC07uLB22l82G5mXtXNBVuMz9L6/+R+hcg
YTR5BZw7Wm/QIgJEBVRubdhNZs5tss/a0PCK1gPgwH3PhGDEb4qSYp0ltaNOoIN6yu9RdyrrdADs
ovFgb/g4ve0wvcQ7QQs09rYCCOhC3Hv3kr6W84GFQ1oaamhyBQukDizW1MOWOdw4KxA9OvQyKz+j
iNOc1GUgwCNdJqadQoQ+f6kqGqkd3hiiGEZznafL7Wgw/TQWMdWhrDMHFjAhNIB3/t70eqdVDqfg
uRFZfu2ogCkv7HBQ7et98BI13LLXlKHjG2tbm18+xff9AGn8Lkbbs6AzcFmX7Oi5+k06QdY015CR
OE+/aOoryMy4lsXFAjLkjvlGkRlDma77a3ZllpU+85/t7tcB4y9/oMAWeSHy7vIKJLWuPV4q2eQ+
F/y9AyONSY6oUe47PtOnmc/FcEHF3j91NYFAcvlaqWKGwldCYcWg0hJRXxxjnbo9uF+QuYH/RTfP
jcprxNfjnxm9zpbP41OE2k7+5z5ZcoNFsGVq+lHyCmGd27w+jt5ViTM9fmPzw57PRHXmYfDmsTxv
sARfaB2Gt9iLs/ZHUT9yPfmTAZepHCBTj2kuAeSBV0zfoxg/QtqA4Rpvl05VtuafBxTYxu1Wpq4k
D+gBviiGSI16CFvc7Kr8ELe4868ozskkVe2e0AGF33hZezVL6XrqnQ66XkBsnby2tYCgVjUXHTx1
BvISQaiIkYy1M7k4WGe9a0HpCOALolZf7e1klZLxQuqG6IedP5bOBvO3dR+t9Caz5PZe+6JITJZX
LDHQGCWa7XZQU3/fSdE/0p57Qteexo0UP7EJluRkRSGEEwScnV8MdbUGo1oE5gZxBAFpbS0dhttV
dYOa2EP93HFXN+zfSeLJ8KOs02Q8SSF/JIKzkpbW/cSrRrjfIOQyOkNhfmy/NXvwlSs0f7gCVMQo
t2/sYzp/NG8vLil13ltebBmLWWjOGBddBuqDBDgMEoxHqOl6AP0+vFrpsqGtx8kyu1twPezRql1e
uJgGC/fPJJ05R93mOf+H+UNpLVawQFgwvZizIacqrFJF84LjdUEuX/S8vNL5fStyWmcG+hhkOGC/
2GQXALGAutmxT8voqvzMv+9wmHL+1S0hFpv0fUHmlxHTZ6TXdu7E2nNIxShoXaiXb7+YE5TiO6va
qqhg54cCRKyI/5csKP41jGpv+PiDqvE2rgi9EcHvruNSO6D6X+QBZOumGpg5rKfZezXKgnsVDdfj
P6R0ZYnhBVTjwDqKWSfuvKMMIZrsipB/WN5cWyv2MN7U+N/zcSkzW7FSF3JkDbVtqs6BJQw/Ohp0
MvOJJ75TYy9sqkLKMw5j9MMam5wpIh3dzHW7CcGFikqof6+s026UJq2UdwcDpV4rP8qWjkimobpH
k/5rczfHM3krIgRyw44W7zyDZZwl+89wJR+RQuy7EtbRnM2+PPfT0kgFqAvAPhfwCmRtOCFmVmop
mgeJTRCNoYFkfZshNanF89Rmr/lRO72z3hCzgRDEtE33vCxgd4dB4MVk+cp6U6kP2GZCwIsfevvN
q5O4ReAloPCz1JayOnqUrGE6BK4LwC5ePZMVZYUsvgM320vlwyhw0YSXXe4gET9DJnjHrC6MZ1Of
2t76w0PpqHp7AIsRL7pbXMDWoC/4sTbTq9bHzAKXyGhzIo0a/RY21pL9Y6gr1j9fTKrWvlzPFA7a
DKxLwMGBSJj6JFmJV35WQyXbgj2kld7icw0zChjHF9Ra2jZoDOIQyyprycAp9c2EIRGGIyiPFyBo
i3pDjvmsbiKwSNg8mMvCe4KyKtcju4wvp/1glEFNYgmCXeklumyZM9gG/NjWPhpFvNkcP2HMWuYe
9hnYzO7fGAunw9lOBdu+ScL7s2GTr51mwJshdX1rjHewyeWAuqenOGYYc6rRdKnrEBskgNG9i66m
I2xuqOfkwvOSU9BmZqA3CebNGBcoq6RCiPeFNDFVqIK/DHyBJGLyDQ0+UTQp7Vkm9YfZYcE/KH8U
KAxnI7ROLFQe0X2Y6rIjhkrHhCWSIdTDyLQF4c/nX8DiFcWvQ4nQKO8ZHmGigy0I3km2f8E3fQku
lJE+uHlTDzS9btOE/ZBlL1N4jFf2igGHGKoT6s8v7mzdTfbAHEltpxjI4arta6pTZJOgO9GNhb6b
exNXYLabZDD47wXyOfHeac6RPm5H2K92MaXOYaK0ALYjrV3CBYRipUuCsJy65/bgNm/LDhQ4LSei
u7pUIp3vf0wMmXsWYAR6UopUq2NB2jkt/C/LfhmevklTeI+5vnA+Q3oHtaCktovgqAZeUjhWh8Nu
fsP748Q7XNBIDAX28/FBpRgmuERePf1NlGC5gMCEGKsDSQApBFLs+nAWZfA1JvvON1LLS2QNDAoW
AKpckvmyZOQUT1VX9qHU8T5g6VhnFHrvnH31gS+I9pmT6CLbty7DlomACxUX+VcZrKPvExEZNU0Z
iKMTB67MsMJekH8OIY3kRMfO+VgOEnXNrT9zQdsq0u3NsVUz96lwTtU3AClWw/i7/f4df3aEsqct
QbAyFN/fT01hlCWXCT37a4L4YXOrxiqOCXdWOZvZodcGn4697+/A1alU0/Z2wLSL6TGU6wnn371a
Po4TAs2wv1NHIkz/p3qQvCWbZFcnYhqlar2BQvVrikSZONNS6HkIjGfTwdLjMV7Iz325/fvtFSwI
CyRcthM5f6PTw2oHXnGojPbllvqkb0qs5/dg6Fr5cGy+WN/2YZ9UqEU29QS3dPIwpppUJFtKOq/d
YJlKevNC9ZyBgNgfd47+C6JakCSDChlKvjLo9KSsv3DBy7TfGylMbvPer5JYBSiEZFmaZy2GkkMD
WUO8VGpchDzTHaVRBU8eppc0C7Hb2RQi0cwWWFE4X9s2zguxq9YaSyo5RQMxEi9b3ZvNHEaMmsZW
kyF1GLXPdyH+r9EbR1uWWeygeM+yGh/gu3bEcn9o9DwugLb0UWwzTdYhRazYR1zTOFPCg2mM2Ycm
93fiTioWEoJR3yeMzRb3AgaCb3bROXivwJxWiJtrM3x4Q7yDHhoW/EIq9CFX8t7dJj3nO2sL3jNC
TS8fYd92EE6HczaCAz6cmg6KySOf56FEhBY+tr/g27IBtTdUQsfV72moq3/99q6k1hHGZkTZzgUv
9i8+qmeVG/ZntbYNBlk3IMLsB1cDDU8798NFBbdwPwPnPrD5AiNP0k0RzWtCc73VJhNkOBQJyHex
OxJFlvEyen7cCyT6zRHupSoocegbvhp7HnWMwOEn3WDx8H+vfk34HFsmZ/wUtGWiqn0cwNGmdxVu
6oTysc8d06UrtkH0UtFaQYffAdw2ut2XWSvEyCSqWmdQLxp5q9VbpjOE4jAY5coeZEhYE1BFGKGi
k68MgviWfgW3LSt6unm4LA2d9wGNjh86vwk+U3rcoq38A3kMfp1wm23HBFeRnjcC7Y0hXscvLF4R
dZ2S0LmSsC+8RtTB31ITkaSEQWXwOuHwOJ3M5X0yFL3dJiKyurMnxfACN8oj5mr+P0zG57UrUXMx
EJYD2pQdzzhxAw048tEfLiTDrDx0bs1iOvjxhSDgLLqGx2LyuSQFtl4qnDk762aFPyG8nhU2TbeM
qAmEd43tH0S2B0GTvZhc4ICzSO9p7BLYQiZ++WqUQkpoFK1xywMDwBFC3uecQYbzCme50tOrC8C3
GfDUCCN6vul+Jn/kECOeesh0a02I67pTFRl0MkZgGqiqqynNtHgHu2qHEx1ktpmBRceWUhvHvlLo
f9le7p+lKVqvO2Q1HKqWSH5KT7iQAX9wwUeK8LUaUnCMysbEWQtEwTRuyQt5wfuGytetvN17EqsT
7rx+Im2KSLvy2c4mX7M3w7Bq3HZeXakSbqIFjaXnOsMG0VirAVGrHL9Bdthr/EzuUYR/5LQ34QVW
uUbvrD4Y5ygooIJtpv3XCUwRw2BYaWIgMDq2cemIRUQzeOjHyTbiBYT4uQmDjZ3XDvqYLlxOtJA7
wuOGjkJUKc9hyuEVsNDjosa5RlSqb7HnFc9eg1iJgxDQ8N0KNj8PHUo6bGP2Q/1z/TlELjiplGno
YEG9ZFxqKYEfxF78zAwfpRY7EmlUMOICTfvn+IB4rvypUA6AJpGyl7j4u+G9WvdojvNJeelA1hRA
5jSzGNOvUkm4XW4D4zELmSWQzoUBZskk974VhyEmUi0eJaUsooZ2VrDHEs0MNLnLmQqHXGsz6sr8
XkJVyhmI67dEnPhBxL8ZLvbDImsYbpzaJucc3Y+VMjBn5aMMyhnSpEFiI2fYQg3HMQdZ4J6zmcww
v8o16gcrVsJHP2X3YgniRdGYTtEY6Fh63WihMoPp97lfNBpxk4wHHalh54xAxuH9iSOVdmWRps9n
FjTuouw6V01whxxTfOyux8xSFMhhQxu4rwloiKwud+pSexEGMWV5J4f9a1B+klys/xVif1Gon+3y
2uKFkWykoFK9/p+QuHCDLRC8h5dHCCOU7SYJvglSNlRcCnjEOa6zzonIqvq9KSlQqd7U4LswSAuL
dW70PH5tNki/O6jpiyFW8LFOEyzoAOLR6riD9zg0dj3NS6C00dG7AkECSmPVOkCdSZR7mY21a6fO
5h3lCxtWsFz/HjihVchPseyECaJXYmxSWkZBxGgrYBQ80lShRx2npRsBfefl3YIMJUjMx5drgLV0
qfwvszW+8J9hpDWy7WnEpRufZaNNgz8OsDKRTGcf2CSlGCRZAr7DgZQFNerZOu4mADx8AxfY93Jy
hnEpSKj59aIAbvxcu+q8d2suKC1+Mcn360gkaSFgaYpmFBuYIHK2XyuGc10Rs92/fTbkK9oIP+dI
vHcxIsk3TAFL1P9jI9kassENnuMdCkj9kU1BQiuCXIJjYkyjD7WgLBbhpOMw2JOP8Qzsk9igF7HJ
hk0gzTHqWFdc8ow3lQssEL9Fc2feeWdRVRLlFN6BgKsFuWqJr9/pgREsh72N4Os1NiQcqFvdnNa5
i9l8VGObUcyZ0UYUOm5N2qpbPSpU5QmhCapLEoRWP/K+vv1MCpg4VlbGMNQ9sTszd+5zNmgvITzm
TG2CAKn6j6FIUMpnDlKJLYwM9a5f2867W6hE9L9cteVxCtYpPP1Sug2Gcb3cfgEfA2dKkQYc4CFx
PTu48j/1nPTtzWO3dczjh3jgSJtLNkrrmkvuoCBFCFA8cf7N5DBkqxa1JtRwqqgJS7Bq64T9L/uQ
q5sh6tNu3kEgABKNO3UzP12j/UyR+QgOIKpLY5QIzJcnYnrVBxIq4wqNTaK3xxySb3woddFysP8I
npnULJGYGwdCixFeulaw+13Kioz1Gnkh7q4dk7uCsTaQPYoMkUDQOjbN4Kp9m+f64sDZCW2P+jyU
WdhuDkfgr/grnpl9wN9RP94mgZYc7qt2ZUDP1xgYb4PbNbshozRJsr2Rq2uFi0/MRxjzqE53vQ4d
mvgeKUVxuB4jCQtfUgSKC/frrqAv/mMO2tfZzYojQHbMs/oF1lZdDx03sSkMKX8CYP0B7TWshAGy
RAhraysjHJN+QTA9cgxR9KDglV27pf/p1PRBIVLOvDElIUge9ns3xZ2HB3niC8SqJTfi8RLDMZwX
H4jRZyd+otng68jKzHNM9psp7dSaU9a/sm3St1VLLJ3RFc82ECMqngOcNuzHzsDgVtFu3ZDL4MVf
Fr1MiD5/ewq+ATJRysKeOAfvPAV+U5L+BAxpexhkZlFG/wlQFoeaZquvKv/UMPBDJr1It6ixSNCF
iEcXdwZ4xfmM7llq7nhqGTNS42jisFbQ9aGnggvIvU8D0eOqiejJk/fUZLWoy6v46a1PxnwwM/So
XuEDYaRkdDMc5zDoZHshgILUKTBZZtpNoXujQjwMW+VRapHPdL95yU/88nk5A9gxmjy6g6EmBIVC
xc3xUO2IzinHl8ftO4XB6qgQjgy9roNYjan0e/OUehEuQO1vQ0NIpeOG8mWQpi42a+lHetBKWQb7
SK61iZn0lfvh1GfXWwAUxtcM+ofLZEWWNf7rwczsznZ9jQ1M/DHpshAi2K0lJwvNKVyeJ1fTEOL1
KSzTXCp9gWoTkYqQZCnv4f07GQ6x/erD9DrgxcQ1XjcWlP2w8n5xG2wRZe5hhKG0T1Nx0iW30B8D
vwXNuVE4Yr9NlqfPp6ZQcdQWS9M7wy/K8z1F+EYd6UrbQd/VBET/dJMQTfrxdXuUNYJ2msTbpeeK
I5/yHkQmJquq8viDkuLMAVuA3U4R3yLBu4nHcxzq4lBhX3MyAjL5v2suhcrULCdFZv3ZLVIg+ABl
d+pGfG+1WYhhpqaCW9B/4uMJDpjC0pPzbRa9Yv1np192FHvapCHOC/XNEpFRUe/LrqDS4hvbrgf+
kCRNvMzEElOdyIT5s/Px7C88RAPfS6dA2iCEYtpiQkKARNUV1kQc8xfXzI3k83g2e5aTfes3M/e8
WS2OQMg1PKwFsjKOzyfk5/VYNzcPcmxBr+U956BE7pIqvtA41yoBK1JviBTdFAIwPMAIdRd0mNfO
pW7z2L3Kms6aZY8E9THnbJ7dYfGWvkChotzoVnUdnQL5gzU2/f0OS2cZ1JKmKH7cIkC/B4ZOemwS
XBypA3Ayfo8QsnfOTv3VRSj/S/BHGQvKYR8TiYBadyiK9EpnQImDhkAOnic7ASfdXqh1W3pWtqWg
3YRolkGkugdr8YD7zOMd0SGBp50zMp4/Ray6lmbuhPm9Bk4kNsRrcmBx/GZFGrlcwGf7cpRj+D22
QGtYTrXZnS5ypRbpi1WyViwKy760Ttdoqt0mXjkOpQ2pM5BukbTj4DuxCOcll+oIbylVNVzwQAaD
6zkqq3W7GZ1EHld8pm1Zt50tXzAvuM9zCiYZqTja/3F2oEuA1ghK95qW5yifxYIuIwEuFlKw+EGv
Bha/83aG6J3mUuIAN/oDwi9GBAj+NSEps3fagr9dyTuLQneRBO+nIio9uSOup4hD+FNV0o32cv6M
pmKRXpYTAIvrxz7uxNZ14RRngXqo6GOSD90Q2pSvpH+tLfSHy4J5ZGk5TchFgJ6ixGD0aHM1PR5O
7XQdAau4739K6HWCW3FXBBem7NPJWWzCxUkxt/8AQWOwu6MaySr4aFydTTVjMdYfkLIIu3a1Xc9L
DXv0r7a1IQL8+Dn0r1C9Xv1o0KULCRl+MGkc8tNbex8Shfm2DOU5bN9XP+WsGFYrT0dwajbeuCO5
LNFa0Gf+pPlvNogqZ/cm0F+kxq8NsKWTB0r39rF1RqReHo9/Jhyzu6xjOLguR8WprjDpYci0Sgdo
Cqq7mVaCVbCR6F3wXFqJATIszjVCgGk81NwHpDF5RuSwbMNGSBkiS4eILCuToBHBQpZDZP/KkoMH
phUgliF3oeIbm4O/KZvEVG2rrwOQkke/TdJGUbFlUuQFgZVoeUpC0xniRzlXq0i95l9G4tkIjhth
PhEZe2UpRBe3w6n3BHRW3jE1GTKtmFn1Trl5uTrm7JvyTz++ZmKALeCy/+WUcS6OfwBeqpXX71Wn
fD69IzqNfG+GO9o0Xhw+R7frE6sDWYe40lrtjY+Ew0IceNlJJRcacnJ106G22wAoE25XkqdvXwEz
3qtIZyRHlj0f7SZ4uxsmyk80PY757ESGEO2KvjGamESyQopHbKZ1OiL+56R1CllYPduSm5U23GDL
4UTaopdmKqvT07ChUtc+52CcPocITyfdLkYahg4QPtfmlS48d8SNCgKvIb8hTa3ctZWclWU+cH/c
y6gjzAaul7+1QJWtyhHBMM1ZOPW4Gpn3Cq3HOAhfZq3gXQ0DE2+UezkBUq1tz7aegm2/VqJBstzj
nnKHx4dDDq5Fbkmpx/PS7pjhgXKmMWoMooSc6ictCQEEQjOtbuDADD0VYVARjGYf9pj97DZCAgYm
NMBNwxaz9xvbA5dE69BEEG6i8NXSkbsH9YxXGRIkJHvEPQIqpxvxYCEDaqBEHhu4MKYvjfqMVmU2
rI3xfw8rjhqLPW6Miawu0G+1UUwNoby/KI27AkmUdaOgsCOajleb+KI6+xvhA37jQUl9dk8qhLnG
DizR9AuT6e0wWU4O0i+Xz+bQiNkZKkQmydLJKG7bmI6b4gKjT+rY15u+dLnd0N0fVMxL/ke5SaHX
FmOwXJxGrRr27ev1RWxDdAtIQDsrR5RBeH4XObftKBPISSgFCkgve2DP3QoUZD1j5+eAfBPynOia
ovbvn/XyziQdTJqZq7Z+QB4d+Ei1SJZ9+6b3oMMLeiNu/zgP6ikUpnQxQamufX67z9Hw6B2hSbMx
LXeiHzdPh4p/SRLdF1G5EBkhztNwd9/2bsxGQm7FAdkG7Puke+FTDPW8dBCZme2nrEQ/jJhKTRwB
MGrgC10Xvz4tIpY0Amw3i40GT757VSVeN7ucQsI46hlRh8eibiYCmJSYWhZV/uYmj43/2UIwNEAH
pGY//e8cnyIHhKGhCcg5aSmuwPnkyaMWHtvMyQak5WQ+UUcFKfozlMJpGLAnV4yCAWCOhoLAPsDf
+AdfSGSG7zJTiZ2f+LxWryf2PIzvEBRbw/65obsB8i3+iVS67+vfOVvOE0sES161g6H1ED3uiuZk
c0C5Q4Ruqo9JHuxd4NBlLbU1eFHRFKQR9DbNruo79/ydR5Ytn3lbjVY+XCu7Sdu2oRa2g3BEWP0q
xBRNb+daYUQY3i/M3vKqo3MJwMftdZH1roN1X+GCeK6tjcC7cN8xTjMHIZH7YtFgmAyaBO8PdwF5
QacwekIt28fS83iOvcsjsurKzk9LLAMnYLv1DobXifLBwSlxDfT/b6r8RkOvnrxE6We6+fMrEuSr
w0ntkkRhAGTU+TITvoozlnda4wv3/f3ggy0Zk8KCapxnezhT1bAqE8BFMMet1cykze/9XvGJP5GU
yXdMoy+dfFn8DBb2wep2aRXrZGfh61sJQeAZ4FEojLfS8FtQ0xa61HJsJvLoaeqHRzruEh79GVc+
OpfMCb7xlhVvKYAfZbGVTp33CrMrDZGc0/jsJnJU8Dqc42wFTPa33Z70Rewa8XLWffW3UlDO+9Xl
/+weC2dg398nf2Wmw6tU+3Fec5wrTLs4BJQYlPhZPhe2lPZmah8bgbl3tC+03E96Fb5+RjO5zq5X
eOvM9ztI94GfceY8juJ1qMYu0EVQ38gAhfwr9ejpRTdeRq+K8ojt3Wxk6I6J6ONf88uk41p1V8RB
EePTcMai+Nd1l4nU1j/C1gR+yV9G2uFv4rslMBeP0USSS0EBNrIT1HymPToJYL3o+QsNFx2JvVlG
XOE7Cat3Vxvd+yMHjP2ShVtNZ7Q7S5lOSUDj2bN7miEEOD+WfOr8kgQW5I40iMf5PNqi5fSeLRB8
SqQhEy7i4pfLnZIlz9mJJfI3EfudRTu3LJoGNigU5O3t7dfbd0vtdV+PBdVUXUQ3+mR1k249RR0V
cfaZvE8NLfhInL/lBE5yC9OFcG6jufY/NABpSThLmASc61A5lO/wTlq9OxVbGLoLWa7EWBch6cFf
jdVyGHURN5rAHBLQB3pKEXJBeQOGLr2Z2FidHFswfbS5bN3cVF5VTmV9wNrS/RKBH8Jg6G0G+Po/
T/qrJGF60usAV5lZCFe3/Vadimri65PYdkDaffqUN43nkC4U29PCkHaSr+LlRk7QfwFlVlq5XEMv
4JLmuxgWkGvJRYqoijd4N7cYJEg1SFpIAncxo/gr0wGlN0yjTNdU6r3FT1jfPIycyt0z6SfwXppS
jOjx6Rrvyfm1yjr1Zg6JCdLMS2LmV7Fvij4JSS/VtQ3ZbmFxq/ZhpQy8edECzJJBctUb8MUgJ4Zx
sz8PqZyK4WlrMVeJJoyeFFGaXL9CRPMC3VAOLlKUe6itwKeF/v5m40tvRTxUEVcI0OZd+R35jP1F
6Xs4YDQteuBbo7xeKhotuan4i3tVIWwT1in2ndVz83g+pWNqI5VKJjLHrNT35wqqcrZKVzczRuZ1
23XU7EA3y+QV59/BM2G1fh5009jsXdHdA8NEWy95/CcqAXB5t7I1AFuv/7BeOQQ7lD2OklT2ei/e
04iFldS7TB7bcExk9px1tW24GIMms0L2zb+E++u00dqp5p96KSTKyr07uMYA5fHw+HLWcmMg22Di
lL8M++xOYq+ub/94q6BHbxoIp4om1t91ISy52RihQzxJkJuYtiGzYuUtJGmogKGfs6bDOuWFKW+P
6NisVfMgHsZ5kKR6a1TZCizeHSConFV1i8+70Qi0azywjFxZBZi7GMr/IR8H/wp5WbAnhGHPgmSx
Ru4JZ8xiciKvDNdJKCyX9Vbq5esW+IJSohbfRZnh61IGyq6/0Z0L7/q46MMZAf4V5SBqenBvyKLB
UoTSgbCrx6Y8PDJ3UWz8GJ3Vbrm6mpCrjjJx0F9yf306uf0F7+laEaFLSjhKABjz8XFMSXYNOsQy
yABJGexa1Bd7nr11qrTXyEB48PPl16c9AKDd85kMAoV8n1EMW0UuVAMKQU89mqQnv16cL4DNKdvD
yzD9oHEMHTVzVmN5V6yCSZdCrGjEN1DcZNia4vMzSUh9nF1yDms2SlTddbFR6g9Vhv+Bs8SPdv4u
UIGm6F5Z2sNAYOkrVw6HOO/s4HVNa3hHJFWUEKaT5KThvrIi3uG1yh+jpeWmg0LNbDPNyJqaWAsD
5qxVq0aUbB1S7cEHcY3Sy84GwlegbkZlF7Wng+4O0mo9f6yFngBvc/+/rRsW3i1/4aI13e6xniPO
4XQTwQLNAyRquBsmB4XSSrghJ3OAHkhmN+VUZZan1a+baiZJK/q9SlHbn8ObZnSXUGgKrEkVJ1qs
xnyFwP+V1tuvHqgcpst9+30xUZkbT77mjunFFyRwKO8KI3M2iK5k3IShgvpyzDTjLFxkVGB7tw+Q
z2bWnMPB3d3z0b8/rVWxd97UCj62f3ORSPigTs9HICmhSMFDeQNno9Fsl0/goP2taGQT5FQ8V2Ec
4rXYGRBliGnewgFffOlsSvB8JTQuMIMUUjOhCcUYwaBzo83jyDpiuIgPmVw7A0b8PQ2esGLsAylJ
1cfsZ5C5eAEiCNdPSqG/VYbwLYoPAI1o7fFyPN4sxlRlkIdRlz1biJwEigebDdBXcVhX0sXfBnAP
6yRt3iytVxzHjHyaia1iDjFB3+zVAOOXbMqea+YQBilFeWScBoECsC2W4zpPGRPu+ThJnlTUWxN1
GQ10hkvK83Tx4r+7fiQN2F4tNambW3RBfK5KRl1kpPJ4aWuyHGluYiLjxOMV9XKgAV1LsQt2C812
OCduRRG3RH7LYauDlYTzROjIX1LPpVKIrXQhkR2oaT1idWsMx90OvWfB7i9U2FpDePcio0Aw9hdI
oDkEK+N3D0UIY2GuVT3Mbd48jNvvdtM/l/oJifaeQgQp2+SaTv0uECuTOvQjYU2V3HkVdEx77rQL
7auqVMSa9+Jbn3mPegFRpHuSl8CeUldDO+YVHF52yOPTw8FcOcjqsKjeDgNo/1E0SUl88U4z+NFv
0HBahCRFbN7EA/jDS6rhCOfR8sR4wV79O0d8YhZu3a78b7OKc2+wks2MTySm3r7q0KgLWvWCkzzR
Juaz4jpFXsmSdkhzg/3sDV0jmmuCbI7zio6Om82cUm5Qg9kc3S4G5C1w8vjw/ItOLgWr+qHA1wSv
yUpAzlmD0IrHTh/vPJCxe7dNXF15LyrnLEaqOUJJwfVy0aRVw82V0Wvc9RrNENRXMn+CAL9byd4R
RiYegXEH+cbfYEZnCZkhIDMPrhBZVXXjZd9kBvcsMyxnHc2rhJagbCzBcs4BgIbDKmvkbvUTbrjU
E/lzEXstEszQ7tnzdbUdFK1K/13nF07IPyzP5IBMJjr5umCpxUbLyugb8hM4jgs+eneNAQlFRk8r
IWJfYXm5FZauvcbbN10Rc1pjIs4e5vL8PKXPEtJPXEK1nCR3hVgx4db1Yn7cHbSVefA6WZqqF2u3
uDIMV02j4Kc7ugWZnWPTHrxc4WRwCsmGAqOGmsYZjJQFutR1Az/lwUyrc7Q2TE6cCw0B6PfZIzpR
dB2e2WYuacVzKMDj1wNtslQuo2CrfzNOgaHmq/axBdlLYEZn+m5+eIfd9YZaRQG0wEv4cWBXtLBb
nxqyxpzO9LN5Z64HZtkuCLtaOuT++t2P+W04Ngb0VHlm9th65nuuZisBmfXZQ/VmfusYXyDhyGfu
CS+I6ZyNrtnSKMEOrWh6TP23q9JaxTzbpcsyVcmka7Fp6SWxDpSuPXT7Ip7yN4PtqSGbh+pQSFmr
cibmBJri7b3Uul4JAWYMD5HNfkD8alanFj20OmcsmAmvlVi0Bu30rB9bkl1mESIM0/kFpcs6kGzc
uyp4r0jaG1neylWh4YYfMyHQXUNrhJ1FENZpePJ6JwuZ+1JE6ofvD4fq75Lt0jj591hA68cfyuKe
4COpRYqVt0LTNrqbcghsPz3gc28dTEW6YqLnoCzLS000e0/uMDcRtd7ngo5i6fFy4ALPZK2nijr2
r+hSR17gPuPX2mt4kZBkTQ7B8jg4tJuJjZ2MsoTs0JVaHKKaMDBAClTnLMXraYVeLMkKPSWxJfYT
LLJuWImbIhVaVCJNrbMTm5N8xgvfPGfOm6I32JVFIhZeRAtBLPOc33vMMasHcDqUA+gqhLlFx9qE
jX3qWdWltZ+JCmepPC5j00v4uJeJZDCKuK3S6iM33LSyEDQoVanH+U4kLHinfxKSnyYUXD/sDyQU
IxDCGCw46l+LWNh1bV4zPDrlXO2ta3FLZOU/c2bwfJZ2RAeI8PpniB3kcujrXi/XxttAxmVVLebz
1wPjOAJbbDylhjde9yQbD+4XjrL5oNCGFwl+iMX8ktsjWY/ipZQL6c/F2ffzLiASwUmTMXXD6WaU
3C8FE3Xcj4WnOScaQLxmtcH8juF6CAr7DwtkO/F7MeLMIXqJ3VcQC3DbWo4v5vsyEY5KlsBOqVsB
mWiQS4F0Ni1agkpt234R2uY3ziqUyWAx1czgQj/bKVcMXMWCs2ym7AsmNPoDWDH68qgFfOXDwUpU
/U1P/8N2H0P9ztFbHpIFEArJmJTmmb5INgt9g/BGCROO9FR3soPQv6bXV2TSM166RSL6Tn8ErKti
50QYRS+FctGT//uBaglA7/EqFKj/BIO59eJVpcYmQjBxbv8KNSf8uHWkh+/6teeT7YBxQJ6r0QQQ
tynCal8iorb3+1Ez724lOTNoqDAzAsEbm8SeBr/RzLx0FB1g1U+amdrW7Rl6rdY49yvGTyz1Pz3I
0ambIB6qD6MG3EfIRZ545ytD87CcIjOe1FIdfi6BdtmwE+bTuZzB33qeb1J5SvkGIyedyb/BlFPy
up3mSQoQ+SbFMj4UdgSCgI9NaSR5svoCPWyzn9fn8yZUw0R3eCeWYJYHQ+EJBhx2CtxXKeCMqIWz
FQa9vuPb7NoSnR6LXMs1db7fMNazjh9tR70togulA7DHHK3qLhJyVbQJJ2e+4EOUH3FzuZ2mvbyW
m5E1rUg44uMGyQAodAV8+ssM2ssXV4BfCBJeBeozE31PWtoEAZ0IxudMclYW9Mi0/7qyzOMzTCb3
P/fo3XKcZDhXPE2+UGgjOfOHiXmRNG1PBaX4RJRiQH/Dc+bhpI/3cR3orY08Z8K0OpmgS5npc0TG
gmJtTgn7XW8wM2OpsWgSuErBd/EvxHFIY6Xu0vsPKXGmpJn8i0q81xR1dXLIWl6QyCq5c+xBkvzu
vhSL3BzULDqpckBL66gXoGvzXr7XdcuB4O5k8epnn1EuNsfK3kaxEQWT3/llnerJU5MRRXpU7kcQ
SkcwhTfESXdeLAZCZLWOIGzGnv9HNdMjeBWa+52hSj/+lVfR4ksC0QSBCnN9TTkFLbshI9yDxrpF
nrRBJa8HOewmKIVJ5sHPAKV6GeJB4qvoIohdIQ8kSsTeTEaWHU9FIeAgvzxzDGntvTEseuSAlP2D
vjPA3zM7K99ch6k5bRAWtZavOexidtpZjGrjV47lPTocUpp9PMah+E3I6KzoJri9TA3jEU/g9z23
50yB6zQgkb0E0rPM7gpRwFZYmyaM7iP5/LHoCvgiq/oCcbENmXw7vFPfR6tYCaq75VV41k68gpPs
YC3ykSUEuWxgwJxTNrQuAct0RYDvCJ2CiGxMCCvm2J3SdJ+UaWlsny9R5Szf4hviEsBvcAssTyJ4
vHfS0NiiJI0cml/SyR0ZlvFxddrUU6S8ZYXhCgdAj/ZeoP6bUKsK0ZLEYckv6VoLVWIlHcc6fIFu
HN40iZljqP2tcjhaJdZCAj6B/vo0PxswFIn3QCWn8D62/Nc9Hvh2idAs2NsJodXJ1DpP0Z4HYlPy
LVvAIvKT0VHZFCyydaEkv68F5DD7D3cYcCY4PzmemAWzbu6cht/d2BHTBI+jJ/WZ5cs5VwwAkoXr
JnjEEIrWnY8d/pI5K6w1p/L67qWAKrlvqI75x2Sw3Ob+KcjqwJXBrhA9fGbgX2nXYjOmNM4daT6F
ctHf0hmu4unsx2tngMNab0cWbW8Gq0HudJSOv13gLrLCt16n+apF1P8Alejm+YR+u62a/QuC+wZX
R/uBLWv0R31Tieq9hDNpju7CbEIZe9pLrlJXworGidGQ5yHyS8+N6t8gs7bJbRwIiTILhlttAFzg
wU6SR0eVxovPqJ5+jqGjcqbVBVmfsOV5oTpcfjz9nBJ7uz1qKComom9PPYzdoAN5vH8kwYp2GV+K
wsNrXCyp0rt7Jw7qjVw1KK/pFpuVNcEcgoGg0zoE1hr4SscnQ8KTuil3G20ZqlW5QaonQkmhzx72
eFQJIzwDiZg3pzgj3OW0wD5NqYZbJXf3MNDPHwDMcVCjT8kDjUX2pmexB+c9cta1aE1ChWIABU2n
eh3/3vIlYQfw78mf9Aa6mfEXmQ98fYoEPWkhhe6HtDqFJtW+0By8WB3uCx7LKtypWEH/NSHGy7NN
9KsdslkmWUgKIci9ytiRbW+OQLuqZFJve44tNVRm3C/lW03GAEWk1RZU/c60j3Nri0VhGmdCnN8O
DfhLVyVEcNPt+41Kwf1Qk9QjKzeMPzvxTawRLBx46lHD+ULBlQabvrmmmoKcrA+Fcb6yEEl5xph1
DILrpOAD80sc41EZv+G2qsjna6FfuGFrCyVkTdhAiiLMFtnCtttuUeuOmOrEvLw04bS+bRKQlXpS
Gxk451+Ew1Xve35HWJNlRDWYqIax8NAh59R8OqFdfZXFK7kWmI9FXPjr+QxD/3Cb/Un4MGvuTNx4
s95Jt68OZvEhbR1dMCLpDyI0ICxS+naz0BIWcvLxkwgiwZoYwmmMcgdgS42eL1rEdO6QhnNI9yyL
gimdmgu+MxxTurZE2NWyFCpVm45IJP8Cl6QrS89h+zUHEV8VC4wXpzfa4F6sWxDq5+qe0kcRVTqW
3SQZDpbevaQ3J9wnlNJdvynysYlJ9ss7haoAQ1O5HYmI82L+EjmcBm2ejma72AiDipCvJgvPpIHq
ldaWGTQ1JnUthH84oD5Fp7XhclFpc85IG4iqWIue2Z5qfnmenckIVnGoFEqIvgZsHm1ZFmQ2wCU5
+SMSAFaZ6l7xvD/V4L2OBreWcFzSAx42WUIHw+Lz7DZqKWtDRMsh7ew9GNeWky2b3Jw/YRJdFDYs
E6cCGrVNBH7CBfhpELiVivDQTt2jc0EcCJD9WVeYRn5U2nJRApYmtD1xpqBJ+C+daLM37P4LdGJZ
/sL6TL1r3VJOrU4DF4EgWjvq2CTdyko4hltkctyVOdfsxiQuktFPMlWFrpQ7zc7PaVuCQkkdqFSN
LNNfHW4wNTUQPYUfquIru/Q+JgbecJ65QpQ1uHK9abDVblk0Y+ZOve+qvsC4AnJ/o9qGuNwc71VQ
VLRXvknL2FY4Fx6z0OtrW+ZxmkjWcUAUHBwbQCwXHGMxB0iFwStPO0d+hURjSrK+U4MkhIfPqxnj
ScDBb3u/AKU1tMFPdSoFyNPKcG0JTfeLg2XxHOCINOeMeTqPrlMT1IoIt5TyNDeBG4myE8UEOLz0
OcaNebZCozgXZjhaAW5VOeiKF69ggYvjXo3SiNSroa7Kik62PLPf8CtOcEmeahd/IGQT36gl9jQt
ebdiXCfAGZrxFrhWqyNMUyzi5aY0GJzBwXTc9VD7N5STaObb2KFQTJt74zFAORHwUqFbdTvU5ad0
dMKOlmg+Lywh6vdh4n8XpNYP9JkxHvLRCBZT1oYCN9O0+GSuwkeh67u1nEPYUIBYFiINACxPfURR
rpTJf/l3RgknjcgeWGD9T4mMdJKS+1IqOxzRJjEaqLVGhKSSiDf2pWppCzMALtBuGfOetk7jN1TK
VK3AIwtI9+M8+I5BVLmTi4jAJ8Rf8usOCN9jsj2ZMJ/QAG8rwzROgX3ZUVf5ZtangS21jyhVlD74
CW/TS32M+/hhZPa9WGOATcqY1bxknPwxJ9q4ex+czuncI7UBjNU029xCxjKAxC7tV1iGsnbt2fT/
zWTlMWQUmxDDCWixgv4+HGdSIsJO/GUmhUl5msavrq3jlIvIo4HXS7jSqqB33wEz+q2q7aZXvAwx
V4fvUrL1vUqNefvz39voqNwT+7X2OJjIAGu0u9apfhl0aiLpmHSBTrl/cp3dwmjxvYvskCX4ucwc
NQ5EhU7NZz9O6CdiVdai/6vszMFhQdAgx5AyIdQTjslUYavD8+8b84m3wm5wsCFuhQ/P+KLTHdvD
RG0wyqE4aPCE0d8CQkFvHpNLddH5b3cM5BjPg1w+x+dLCA9KWYjwqkkmJCnnbt2FY+2PqalKFM//
8xvmB7X5qdeXbqAEMjTLMe0TkRcVs0nlCUuqsvkdoWihkRGJEYszOw7btbcHBYaPC29m0E3/429/
yAbcUw9JYDzrrDthy90Y52xzpnvw+iC3Sck7xieQgPYPHh/BbkXmUy4ZnHIYg8KJfCsJp/wIXVg4
hPU1cAeIUhzdAjZF1qaGxmsVZfDHPKeVcMCBMOF8BUQLrszTrg6D32Q+81z2WRV1U4q9BlPYCkWA
H2FgmZoKPWJcKDwh1KHMIgIp9KC3ehXye8lx1c+3Z+q8+XVi0EAZjY0CTP5csG0T8GLkatZgJzN2
nX2QN4e4GPW/7g9kGkJOsGIc6CwxTaMOw3mQt8BFOmwSXJoSEFF7acg8pVNmWXdnkClPtGsuQY5n
sYV5TEd1eDXcpYBogfC/ESaR928nDNFXU07eU/Ws6aaOh2+Rh/P6FTdI44tIz9hC6Fpb7/oUs1Fl
++c8tZyIOA+CwYTYNyM33tqBOAmDxjChETWRzqYzRkdyUO8xpGEvnJRUxxEoVwDhQo2hnJXussxp
8z1hihEK1zLjte5msm+XhYTLXB/T4O+6z8JiYpcR36tHWUtRF0IT4lIJDkjppLmhqh8BQkSE0tGp
QmXKaWb6SJ8lBZx+pXbFNhNjRa3ooWsJ0A+eRZ8TRl48NEF5bkRLciPR6c5hLl76z66sMbWTer4b
rIWTadPgj7o2UnmRnMgprFAn45ggO9/aNRjynrcCm8ZjB1QCofHK5ywth5mOZmV3dhCFCestPkd/
X3pYCBLW/u2xhvnoylgGoIRqNoXkkyy81ZkgOwE3SnqjJIxOtlJ7rjVPD3FUguTIZhBXACbIlTe4
MXl8adiRq/Y6VxPzKAiEhABDtb9xIiv4yAMYbmG3G6CoyLw7IGEsEMsJeUrr2othOfWtAFWhUDDP
I4JLgfVh+ssQVG/EpKulRS60ZI8/tpv4B4pzgFI+b5IxINT12j9GLvVByp5z5fysx/J/viH+Pv7j
417AVDegaHGUcrpun8XOZiKvtZY/bS+JEAIrFZhUpZXeKcBRa2xWc4weBsUf2MtmAIkj+Ag+bkGv
CzaENYBp/OU288Cx1fmg/Xso8rlzQf4FRESi9VIY2uo13d4sJsbRWyvRwDfPjlFqTXJANlNdj22J
cyQ3pcKPg5HVAqroUCgZgDQsCGcFHbuxFBeFt0G/SMCqvQyDZ4jtbh3wBTZ9j964vw4pizDoGIV2
TCNyDWAtw37AwktsVIDkAPk/qhgf6aDYgl/W+atijVuz47sOsVgPgQ2M30OPAyx6F5G6d4aFI2N8
cujl6K/mrezPkk8artky9wk0ONbOhjFkVjHt8W/3olaCmqDheJpkikZoNCSX6+1dHZ/ay0JNbFO1
se/8lyyutYmsB/P1YzdKELIJVP99pDzIUH0GAimXYhi5TWQw0DYrTZHqyfe4SB2UoTHQlJeTklVo
xIrjD/40BFEVv2y+DGz54o1ZkQFDu8Bhl10UXIOhnWcEuEgo+/RLl0D8OL/A5/ksiDdvzce3o4pM
HMC0MH+ef6R8/EE2DBuvGTu1F+ToPzjyTWiQAzttvcD4XfqE9OOzvkAq97pBaDvVJlXLp1jOcOrs
bXCEmwJiFpot85Uk8xs7UicwCvk3MjvSGHcmPorImjBwEoSa/yyCLgnpyTZxp/4OuSeuPCFEJkJC
XIJqew4FjQXsB709dTfqM9j1GWY+CtKMrjzn2FThqXX0HicT/tzD6TJu/QsPirX/g9PeXJg1KeY3
EYA3rw0/y7iVzTpMtzwLLHrIqEQsD7AY9DcJn7nCakZPQzkkjtNjvvY9m9bwgms4p40nZGmh83mI
r0k4D/Eq0+mL99hyqQ4JFMz6zCO8bBcln3wqr8JsRaaq7an8layxPBAWy2/7SISakvvk7NE/W8bM
k8ulwy8S3B9rlPBFxGRKeIk3AF28RrMXzRzXX2SRzlA/lSdZZEs+ONFrqd4/3qRQkrqkZzknQJjO
/zQufCGASaNN7wFjSwBadxwOZH7IVJLXkj2jxFtKAdVo14iC4jbSlThdkhvsMgDur0T97uM7P0Aw
cySFVFQOTx4NMZFFliZY8RrRwdG7suXG6Nferj1XeNkPhq6PYCvULXEOTiIa475K6c82Y+Zcqdbu
MkcZm8t9OdyFGXsSXQ8rWO1YoMd4j027aC5HJCXjHD8AZ5uvMLNxEiVYPNTrrL/bDuLWswr0RYYZ
ot3QthUE7wu98uE60LaXvbyL7LBJbono1peFMVrfMebMxQbpsU2TBzbkLK84MDdDtcoNJXosNCKT
yqkFSDb/IcEk5rqejOnZI6ZWPXiGqA4JRtZfUO6qTMapZkGKosKhXPc7SWWW+fyO3a9slNORPvQt
5PaRdAah+t70mY13aSCZNgMoAkp0nd1HIGHyTfVF2ifHb2LIAU79JBtlZpFZzUjlPcqzq5nu9Uk1
1KWNAma5sHu2AU7sEDoYdCZ4wsi02YzOI0NtHZPfJineUu+qdY+UHCL3W7AjsxVqIDcU247J/gzX
m/vz8kb7G6Dd+HowDDBfbG3sj/9CRC7z6yj47Lyr8pFdclyUqZaOYWZtV+sTSKQ8WRMZjAXFPKM5
ue/7qlxSUHrM9A765ANXQHRdBVBwf753t3hq580p+k2jst4lVD82vb7rqYYSme3jiLYoYod1GfRp
+ZP9eKXviWEfhOHjTNNqLfeoHrujAN+v+VffwAukrocrFyp0n0jkK2zhe1n5jmFm4NR3rbaZkfGL
CvWoUU9xwpfeBqUAvZkFt45pFlIwcI3hSUlF5S/sOaJ/mPJL9/8IfuxcXRNj30RD4PE8Bu/Oj0ef
ILZSmBeGgtaWQHlje+vWA3j8It/GOyYks5nZ3UIaI/sHWpRDrnivJgc/t+lVn8ZLmLEY+lhjYpoG
Y9ecx0Sp7Ut1Xr08984qRjHkewmrWcEMAKCReyfx9500n4udtF9lkTAGtw+0NghBwK2+40zyigAR
BD4UcgrN57nsvunIo+p7LIDgFkaY9ySsRqHC1CL4x6uF5aoC9n1Y0j8Jwx/fOE4/FHe2ikavy17d
8ug/PNRtaZ7tMjfTKmTd4B72+BugEOJIsfikh1n9XhS7fh8BDSxDorRb/2Tyn6gYAkl8bZsVCwi/
Xx36RHhcGuSOGnIGiYTjkDchRoMYZrO7k1tT/ihjpWbWrtlzHl02HxZEOb4Bu8xDUl3uZyiZtOew
WfKxvSEnjKO4nqLMLyvt56wgfb6d6tR+ay0VjrhJr/9FN4Z6En4s8zAtPS7H/wunIdIjXIMf2mX2
xp6GX6KFuFZAOy/ulcqVW+HQYSilffqye8dJBQ9QvWooXxsY4qBSNCfayBhvmqS7tYamcQjekezX
LkdcSa6fZsYnEfAk1ryv3JxYtYPKB8oqSeOQsS1YHUANUeh8QcW/Nh3LOGhxcTInnD1y9BxYNjfn
r02y4Ztjy6GpmNjBuhmhDZUK/7NY08oEZnTy9hGliWZPhos66GfpwWqIYEZA9ceko0tF994LeFd8
y6N9OCOCopMM6oMI8o2bTIVoJU12izFr+JREwbgCKMbLYrpRmrY6lOVcMHiqcInEwTb7i00ieiOA
kR3VA3BQ77G//LwZeGt4zKBj5VQJ+7jMzKM0LOvcodIC1U22eh433q6xDUKSOOSwk+XcpXvkVzzX
3WIVlD5Z/T+77aqgW/pbK3lLkV7oO0sm3bCm7PinKdOy5oFL5sAAiGr4NbjJ0GP5a4a8aOkWGgHz
AdeAFVB67KET2oS1BcnMw3BMLKF3eADUkF838S8cv3dyKG79AXlSb3R+LhBOxTEHPbAjT4s+NuHK
ZIW/5Q/Z6aKVpKrSr5LxewhugBE7gXingB/1/VRdpShn4aMiULvh6/3kGEoF1OM7oCKy4C7VHFM3
GNGQOX5RXtCVs1tYFqvp2xNxRRTwx0P8Dkkw5QmvQ0avsB5OTyq6vHe/x277+pUoEC5p3MEtOVGc
K4Nk0bWscd4N7T03B2xQuYSGwQMTPMB4VwGBKl36gNZQF61NFGbA+bDe4vRUFSux8I5JPOAiclQv
p9aplkwfGfVFjOIZm8XaE7B2+2/ZnExH40WiNi6A+ro/ewcI1o7/ZlvzWezV8R7Fab6pebTR54UY
hnqlJ2HpKMOPgV1u7bodwjecvgpl+n9frJcLKYY4Zgx05+YVVfXv1dj8AV04MEZ17YO9Mpmff7Ly
6WQDr4rJENT/K4eRhnSRrBrCNoF+zlrM310s4zEqDG+vbBw5OHLQFQ32sG6+E+DuwOVDRcNzw+ry
H5pbaz8wt9nt8LAbRrRhvm27PCPTWYeB7KDP6NRslrJ9zv8bYHDafHbtSVZSF7EgxeFcMz3OcBwm
eh9wY5JI/XYOPuDNQKztsb6cDiT+GLDbcMC1rgDbXvCrCh61EejnJdfuqWw0PIx+pnG0yEeoit/2
7qpgDIhq2wGrXybw4hE+DcYIaU0EeebpTIlsyqBFaU2Hfzi1HUOClBcHN0W4SS645kx6TUEpXH7C
YOFPNA27dmppsX1908HVlbGPBKVTD7IpuT9ynZeEyzR3jfnM7bzp78EdDINsi3pc2AEHqAXeyTrb
jl4u+txJDBa8wJ/V9vMrrEOK006ZNpv+MDXlOot3ZA0NuIFNcTUjvgtuLGQ2W3kU32XK0xFfDolf
MjJjKUm6QtQcfqmT/q6IpAvC5NdqLc2EiYbt/0K6ON6jHAgHPgiM0zojC5VUd1mKrKLSBnB21Yp+
43t/ek5IwcK5e2aD40VTbNx4pjyKAHmkZnBypcg3jtOn1k16yqNrOnQNLIf5SwGPFHVUqWYxESHR
aB6cgjrnHRVRBbkdN8GNNYJ/cNL6EsVD+WiaI2G0krHObRP/V5jTnVPm35fJV6ed6m921W0jDJwC
hQjU4Li0mp5IQl7n+IrqWkQLdObiEP6Sr/uv4Uxrc86N7q0cc++mbOiWzyj2RqEJ90f1PUZMGOoQ
MGMPoPwo66I6GoIzwMtf2QQxV4aQglta8qAfTiWfsSxi5V7OZt6GRIqgnFFNms4MVTd604KmnoYJ
3FKw4FHzowk9HjH/xB8I+ThN09sjMt7dF9xu4/urndtTSzpXF6hfHPoryMqVfhOCIe8edmhuUO6K
vQG9tv5xie9Efm47ddUWjzYCjiVf+DasgLSs4cNCkb/6tL8HLlTzjTxiIp2IMsviDw2P1mCK+X8D
kJrA3qzvezKVWThgacOb2/bd4joWass+m7NdWoSSDhRDMWmBk9YasNudbadM4CAz2xwpLliLHxCZ
gXLKLO27yi3Ejb5qIbPs9qxSi71t21EuG09pXWhhAGWPrkxLf3gSPksdZ7Sd5Fmth+t3XXe8DzED
RRboVs0bY5vL1SNEIzl0MoR14JTh1zoZ/yCamdLmA7OIaxICRPXy/oLJdxmFwZl6a7BTpmlQyKUP
lqtlXSzbtu/o7YgaQpB0iuRuowYln5TRcnEAgjDZ8xZmjTjx3S2EBY8iubnhKHIqPiS8yk1iLcOd
7vTdkpnublUAoDzQttePIpBulg4F6dUnhPERDdXzzu914gZl8hMf33vhD8i8JZnkTKEOf/Bfs74x
GBjs0HG9wHa9ePW4ZpBozHB8qP3ChHEuRuoBdXOnSLt/jQqzwpDIJp+lkmb9k5UI8ryyCxGuY8l9
+aDldLbfzWtpu/+lLetv0j6iqhd0emcOqimWrG2yHlr9SHAHUXrefKhm+N0ff6ogu96NK+s650cL
dPQrTvewBFanGbBBNvfDe1LCYICWudKTNlCWuioGqohwQBlh4z1OvMNPmJbkzNgumu7zbzW1ImwB
T+cOfsHcCV2ROHcXXKovN1thU1sx/yOYKEX3fTm6Kg552j7grAUMuFfQThcJC0rNIBrIeJUrGjrb
qYPr8OyGajZFlPk8kin1XGgZHi5eHaXolmpmX7B751RPS9+K3r0fQlIRF5skP0I8PG/nTOasNW5u
FtuYjUDNfMJcIsyFhm7WlUT0pYeYUmwRU4MloCHWbfswGGwEUscR007OKGdP+i1mOs4YyLwBD6n2
sJh4NXrVWwDtJsuItjtQM+gXLpWPNdP0xj8VSeBvYWVgpqbHHAf2726rLB/TO1AYrNlDNCgTQ33O
WOHoAMsc20VAZ0hn/Gg/9o2BvckJYvKCjqKBOOp9VMdwQnTr0PKQr8HUypqHzGFBQ3xIIURnQ8Y3
xo3rt2sxIWLncMvdFfxK5o9YP20xApVtqjEk6VrNCc0pPyyOAwNXhxdJsgRRLZjge+GpGfEyQhb+
PyA7DpYS7CDZ3BNHsDux5ze1txsHyrONm0oud0cukMw0ytjXHqRFGRCSCTOebpFE1xBT4EQ80l2n
sI8YhvVGg17OJ6eGIWv06ELr8S4odPcTFFga1wJ/R9DIFhip8vZjw7qzvOAdaQyZczZEUGh/uSFy
FwXgw51aEDjaVj7TriThLwpRfn3h38e8c8lcgo/LXbyIFm3OxxcJ3Vmt8tqKgwqjIzsyhN8RvibO
Y+Eyd/1RYdIHaV8i5j0qNw/lAJhpYt+ArOuY/qHNJIInJd4E+TRQ2s2czxxRG98EtTmHPcCVbybA
mtapxVJMGc31LOhd0TOmuWS5VzFGquF5bsaBu8g6ThpRDTG+3zAteiDlmQNelu/fbIYdv7oweaBY
VjiIrKXF0oifg/mmlvnw9+E42Hd0obhw6+eDsJ1HNivv3XwNUlX8mouE3T7UaevvA31tmF442kGL
q6uY/zQmpSl9Vx3UPO/bqq1x37aU6CRinhUXuGhrrxlbsQDRhEGab/U7XvSCFAtt65UwaL2WzWbA
jVK+HLr15IdLDpO+DRTWZE8Bvly7lNYZTN4Qtf+ed+SYgElN9N+wIGe1D+NgPSRkYHuLOgWt/Hxb
R/UJy4Su7X1iK4JEvdZRtOUyAysqiiuqNnSHgcP+9kQahv8l+sFtVXFmaCQSeX2T+qYTQy1D+4bJ
a5M0+tzHzgjVPGGWvtTZ7Mf0W6sc1ZbfBT7gr1KGicVijiXL8pY2DsjvfuEVY1NwdIGHz42/kQtr
e7IFzdzs1EI0GUlyAifioZCu9gKaM+Sx5Rc0NZ1QuclvVB01KMrncv4gc7g6u3ImvI6/CoBECtmP
/xAtkuswO7cpDa1ZV/+e7yvJOQpHomewv52qoxfsZAspHUyAQ1NXvj0n9H3E3EWudXNASZnStHbf
AT/NbpvGaDRKV/cTqn5YKCXLVa5KSCnHODTBfGia/6irdHVef1EtPFwbukw41e8z7FQhrWta4BNe
A9vNHg1ypduUtgUDIJy+9p4/o8wiQEqri1XImEwI7dY3Z2inEynmtgPSWgZsq79BbUTMifr4Y+c9
GkVjnlHmmvJRA9smb17+/p1whZtFlG33hCtVVqlCqa5Vft18DMmyi5F84f1E99GKaOK2dK+BOg8o
/YjGNG0CUbvt36XVzw4CLlX5jjB5MlKu7CTV2PpWAwojbI9bVOZ2IrdIx7W/dMKW0Jq1kiJS5Gg8
Tu6MjZ8m2S9lUYQ1bFJnwIRf8SsXyrG32CCCKK4LAC/YZDO8p6lBq/CAX9/TJ2xeBD737bYC1sO7
J3hI2wyIPYYe/syxY7OT/CGQjiF3yAnGcJBUWNInffFdccHqWTEvijbJdKZqlP8Qhvwn/uWD2QzR
ZBesETKj+bTMYXwAIayxvY3e1fqwBDArO5BUBHcuG3sGR+VO48cUlGOjBjua17lyeW3yuznAzGJy
MnoT58bAsS1VXr4O4JdoZkySaN66qscSjhidGS3/YwOXBn4y5IzuLfgzb4+C2cKQjk53inv6qbU0
ff0r1PEMFDWW90P+qKOuWh4/1J3JLEB52K1zLELqakmK6BA6EVb9h3GtbDC7Jx67y25NIUY9jwKa
gzEi5Y3tH55azI9ZscAjtIrunw4JQi+FFkeQjUj0VNyxY07XIyVSP2bjyxlePCglFILMQEjOkRbb
LpfKzWZs5MYuNL28elUf7k+UMHIacnBEbJaNvoI/LeHon6DOiDwj9MTcGWofAd9nYuJkBbEIBDtI
sYiv6dytxOm2rn/UcUyo94vyIj1NTNLQx6+JG2cPWGkJ31T00FRVQ6PTnu9DUn9VAVWGol2/4u7I
iavpLU5p9C7sivrkG+A/0ddQyg+o+KT+rAFb9VE9m/KgXhjpWbG7KmXOQIt4CaSmp24Pke+8ZvI4
CQiz+SLdZi452YQqoJEK9exqGyvkn/SP0caM9htMGlDpIo8WCX4BlkbDbO6DPcjWgUx67xCElehG
DVBjlEXRMD/J9Hy3dznCY6iZMm4etkQWymwkv46mmVr6ElAIxwGAqIHjLLY0peyrfEMaF+SDqLI9
Vx0EorkuiYgGKG7IDiEX97N812En0T/THkKJa1PcbVr1y1/Ii3wtOXu55FCb0TSvcTCeCytYo9tw
24V0ryhxSZAcAfgBIfT6g3Z5y0T7Rb0cqfRW7iVCR0p8oOoEPHSYs4a2A5nKexUMgbiHcDZH7Lbc
zeqeaREhCHME9MkYZ8VsKwfcWFt7OuPmAS+SUG1/FtFBpkRDvTN7vav8uHdFMV2vcb4EIUdrw63P
Jsp+WcGOaxhM0TD4Dl/1gf5iOpcWJl1ZInMguuKU4VZ9gHQ8HhWifRMgFeSp30CxwpBEZurE8xJY
KJh9OvGCWKCkJGtYytp0ntv9/Y2itfptdfjUVjVlD7CZ6bGc9CvNMxfVjMcihvfuNkAsgb+K8ELo
BBVLYrWZzguASs5G5V9Zga6UzrqLi+i/6XMHV1MSCb78i/BMUid0T6gBEpvQHwmHS0EJ1brk0bOl
YSjP7j8YQY5Tmc6bapd53PQboAFYXCl+4XqM9s7F+F0CoHbMiGzGPMJdvyW8775H4QPMwWhRkrXI
P3tOLL+m8retcBUJE94oCNUK+xUoGC5j6GiOUShyZi9RIBXHe7jW5ESPx6vTJkuJPd1IP9uTKo15
26y1++WOa/ZJaGFaWeGqyBuxe5zED431u7YMiPovlsA641JcGvfOtkiASsqeE+pURIbm/M6glWZW
GvMgmIyB0eC5ale36CcqKfusMkR8tPMwMoyAwLYvSP6SdgBDiwCAOL5jZn3zFC61ST1ay7KfIqFi
tCH4vckqVzYzjJVHhdBZ2LpmCshE5fnWVyzBdGskKj9X0nXKQpmbYkl+NcCnFLnNiCRUm+kPj4JZ
yZRAp8f4oaXekRQ01Mo+0ErNnCX79JwK3Fwqex/tSNpEhd6bsJyJ8zHj36d7icBykawfCMC+Hf1D
D4SuNy0+AiuxdyxktYNyiO2Uaet+wdqcIwizpTs7LZCZ9Ivxr4UiJI9OCgRQZ6zkSBGsBJ+S6BO2
SVdZWb12fMaTaBS5udlosfVvXPhA4foaAEYKyfXVzUP92jEEvmqldlHDSgZSz5Y/2jXvMhaIx4cn
GEot4abPpAOj2/Q0IeRCvrbf2EAaVpx4GCTHkQX2rRQ2GzencU/VCF6bm3KQfFdI3erDm2mtWAe1
9Vk1IXdjwkCR2rxlxGq+R+B16dbKOHrzLNr45m7/LMYM45++KhW3UynjqvUwz9IDyujdmMyjKFLE
vBsX56LzkpaRTD5U9JwL3becCBaUmj/e74Q/XwvalRSaeRkNWlGWGvjSvNtBliXAwypt9NN6iMhm
oTeEm82L3x6DlgQMxq1sFdHQuGy/6NHzuxQRAh6nlJfzUHc1+IgvhbOcw0FM4jAbkRWARZbNYT4O
yv2PumLCJsj3ow5g+fVU73naMOs9wdiJyMgtsx+ve3sc5iC0lCEENoYGyILwTkvYIPqY1Duh6mlc
vMCbpr1JtK9IFTdEllgLuAbdLLBPCb/a5WMN3pOBG8w+fWDWUWlDmzlHOAbwBpHlxfQ6zwvT/G2s
EEqApQf639KQC7NIdvrCJLyKCQabBDL1TopPH18nACBr59wnBUzdhqfFW8E/uQy/QWRs2Qg0YyLh
lxGeBeZtxHm+226uVWUIfLHWVNR1hb4Ev+aKh0dhaG6nxPFVxFsFmM28HpnL9apIjsdT2BZJfwjL
obAp5QyNKZGd2h27zEPPX9sgL2sz3+XRh8z0IlA9NkhtiSgSpMsHmfrdHsXq3QBddSBdHFScnj1s
p1Ct1YPTXmvtVQniifYMAM9vaGDfDIgSv3JiAjYPXosFpqlsCVvNzm79oecAYxo2i6YANJXLX//n
GmiqUcZRVqiI565t0TFAVxV3Y0AzxSDdBUK/i+W2YfvcZ4zz8c6KZd38wF48v/m2HnUHGykxZpl1
lKSm4R4J7Ep5HhZg9/cMF0Ye43LhY5R6ZiuTJkYtqL67Ay2jwa07GFgIQyuH1s3fxXltZIktz6Uc
mJCuM5eXj4mChAY3jenEUOPz12BftR1pTa6//wgwetdCrGSywgMHae3D+din9T/4imhxku+w8fJZ
M5WBksD/6PwYBn0QXgl0uu6wJVQq047cSISAn6Mv5Qscb9PK1/2hXnyW7Ayt9JbFsCv4vz61EX9k
SDf+m4i/DMYZ3Newl+IgaZgGrtRSsuAQUcc3HcE0YZpfK4l7tORkY/G3EgLPGqpqWyBo4s9A0q2t
DL5pz3o8WvVR6HbHo/dPc8tdUBZ1g0vrx9YairY7InqsXnx1dFCKrnVQPU583wZjDw+KcFOtBsP/
V++G1lPnNAokkR6686ezv/nF6P0Ecpw4fTHEHLnfXQyxAt1lrxX31/oYsIcf41ps/Dhy8OF6yLoO
8EZhk5bCOvQavdg5zuXUs/BBuM5kz1ZF44sQxbISnqvTcP4vTdLFM9yqjwoZGEEwFLGG8k8lbZqM
bmUiWjlE6e8kQj1Tk1PjVm7D+HNPrPWr82wYBkhcd4moe9eo7wdX5QQa31frla53R4L1r6hcnZDG
Av772vNHfA0StPwWffP2xXDwT9aM+71rB5uvr2K8OR6vo3bKoW3bLszmYo+1UcNYaT2Y80IA5fcB
LnUWxdxjvA4Ckbcd99rYtCNafmy6hty0Y7vUbBUrnTg+IvO4Lde19qomlZuGt7tRov41/IiH3LDN
48lqRVJRTnaUCuCO/efBE9Fge20hCeDyhp4yCpNEfEPeucslootXrFQ+Yzd/uuNZuzxuA56fKyQl
LkZBOjgdwMmZiUMzE/sY+drlhK1xJfG81cGFfyb5VGB9IbuU3WWhiiTVXKD4e31n8UPlAi/RMKNq
wuDUDJPyHdbM/UF0OwQ9iWfUNwiJv3s9ypTrELGFGQPM/HNahznDSLniiNBxDJkwHAJTIvdRAWPn
v/0BuG5DPsfI6+mncDQdxRubLBzdOoubFGC9hq2zRpJEezz8fZ0ckHOk87tgDVJR2fulWBCPEcHS
AAivajCDOCBV4op2n5EI7ehqh4QQDqPjko1ETLdZTfYFFdCqNn9m+hP4WCaCwPmm60HjaVXspX/1
6qNOn782ajItQM7zhDr5bq93vzHDCOuNcGqjvt/QaK0BW5DTl49o4UrfPzqYoPiO3kXOXsE/J4wK
fQRnvFCrd8vecgahai0s++RBkoryOgONVxGIZt+nHsEPHCK2xyWtMBPzIIDT0BkHi7xwEUwbKTJx
jKcDsocprcodIA/vdAl9vg4fI2i9W0oknkMtD2/5QlvyceqU8ZfScUneH7cEmdPgKCPsgY/Ffi28
ukzFOB9Wep0I2p+n32RgUM/HRRYBbjphgWoyfWAbrSysR/aMBoh3yVE3Q/8d4RF1J2XJGWN2lfh2
VS5bvdpKo1rYaIMgBrnHThPtWSKNj0bxjOCzSXofTh44SRA4PCsv9QFnisgL3KFk2i/l1r3k7TDp
AQwLFXxaTBCD75uG4rb1tMqCJm3kcyFLNrufMxEMAPWThXh1HwX+0K74sVXcQkzjPKagLbskktUo
8AtZfvDEqNFirRY8iL3MpVV9eYgNT1/eoSxIbbcJK6HuvmeMdUnQTHhKKDtXU8xVIUuVPVT/VBiG
1WnnmE/jL6rWEJBQDcfDmM1sA4eUBI7aikxWz1jGng6bJX7nQKq4RDrandvJ4QBIJj8+qnW93MLU
ODLzjBEj2d86HdBIbmFqj0Cnb0PvRCluMFiiOnXATeLNbgggTSsQLgEwm6GjIKpf6dLKgXQlr/7h
ojTtoisE/poOJu62OoZkWZ3VGb1or5bUXtThGBvDF3WpKj6LsIT6RH45tM3VCNdHIBzhqR28ppvl
hYl1NhSBVvQ0GedVaJfrka30ud+ZEL8JM2+aDN6lPYCZMvniM1Do2yGYK7Z8QPjDORRiKy2Qq7mE
Klqm+pcrRidPn+jRjgMdpEDSnPhI2fM/LzLFcg5lpTbxNKLBqKzDfu9RjDB2X0E2gauujRO9F0nu
mMF9dBTRvZ+pvx/hAiFjBSZycvREdfCvt3HA/vX8VKjHozSTJiWIBo/l0K5PYiaE0S/Ki2cnWTry
CcgMxa0ERdfyBp4ZeTb+tgmEyCt4c3rcfDo4E+ezHYeUaFBDZAQc2AVN/IXqqs5+ZKgsL+4Hj/lg
8dDMUKS/6MH+zhZa05z9VOu1kLMk75vq9MS7VAZSCuxNjqhxCD+DU29pSJVjwz6s4FoAfnoCK3Nm
tCR+x9w5yoKgXF2AbMCHIcqNQQ2nwULvSEJBjjWN3/ZFgB1MRL76O/BzkM03uF1TMNL/bIX02QzI
QKhQE39b5ZnQ3dIVp4Nz//Iq/sv5ghdWAyvd6VcHGsmQk6iYTGQBV4jAOY6X1tv36Xim+W6yiF1H
C49OPdxob7IQHsnIHElHMWJ4apwuZjWyxwsf9Zs9kJQsA55gMdynPtnVXpmBBPAhVOud4VVl+Zc5
WClYRlsUP1mbBgqobom0WIMAThxFeX5LMKeT6kxH5bPQ+DdTmxx/g22bXdvOUyL3QhAg9l9C7fNM
/8HuIdacFL4cvTdTjOMk79BrU3qauvsYvNkoZEmU/qQc3IhZ9FWGitaG7b68QJdqUTo6dsc0l/in
L9L9HIOeJPjCsW98bMvA/6sEKO62fT1GXvgHlLnF8//c65WD5dtnbBnqzCJbmpQIVIt/ufXsIKnU
x2Xh7LBz689ExgnCKotYcQdL/rSyI5qKIcPiyJLx5qCwnMCsU6gWvyNBC6rwDq4JHSQxJdSFAeoS
IwsTZQDf0cZ4t2HSKAzdZu/xoGkbPPCcbail1rBt69kpFGH3y46/JXB/+zfPHQoCb0ciholV8KD5
JBL8JwnVa883W8pPJixz+hmLdcZFNWiV5uG/n5Ma8jVW4S1rnaeyMqCwvQ/8P2VFMhGmukkmpnnD
rKw2S4XAguTk4yut6g8te6Zpoo9570SEGocyqs8S7tPuILExFfHo7uha7gcVvir/cdUaiRKPMpz7
02HeCd91HDreGsiaqMmXocg4d0zQdujSx1osbclieToi78y7P5LjgRYUzhH/gzKYSkMgsjZHSRtH
2ZH4gJb1Btq9PECj7aDT1p6H9agRjq/5I49Bf2DIno8FiNVffvL2Gd1pkCbAWCsSQfBPEyFCEX18
WfsGHolBrtTjSRj6bMoLQSccvYegIPj5bNCCWdel/eZVZ5ccN2s4SzCUhu1kSAPi0IfSKB7gHDEl
lpRPzeitaylVEr7lRNh/PsBgnlWMxps0DqYricjsJpAQAFH/8wrYNQ33kI3OQeD9nSHBoPCbvITj
8wrN6el42v6DyrCeuphF7LbHPGvub+FzlNEKilD7I7jyuwC5X/wwDpsiqfGtdS47VrCgTkVKHnkR
o1Jko2Zo8ncVfFIAj4YC7vu+Q52HxPpULhakg04ymjSEsw8hi5TipIYAg6ikLPB32BVOdRGTl7sl
eGoG4pkYmuuQbAKUhYSgzqNjhtngiswlxzu03eqEFkoVbVtxvF0szxBQuh3iRE82weneFs19WuON
RuOS6A2tkLx173AlWIgK9n4c1oyNck9gxrHeh+RNR0iVtjNkVLo7scyA2GQ/mNMEP/QHpdNktKQh
2ILPuNn4Fn7vrV7AI0xTQ2qDbneGd1qBekTTKHBc99tcfh6p2ccdsa3logzFKBBM5lPAR8txNrXx
o7FnsIcaDgpOoSNndLHwegK0MsBtU0q+c6iBBEnjrnGoyoH4YNPJh3a6+DcqFuv5N2crvxxsqWYy
kGNpmtqJSxzrA8hIOse81qrEJHF6+A7VsmdGinjoMsZYtupSDaqVaH0HFgFy3CpSmY4UQH3rt/4n
ZBBvYiEOEhP7nk/LznjQE7JtvQ3W/6gkLRDPz7DjHpY4wmXO70xor9eKkLzolWYxodZIs/9v5F9t
kzlwa/VsEEI6FbioQDoPyYn0muCjxiBzlV9uC8v6ZYhN08/xUW5Pb6PSCeawxb9xQrJCchg2JzuE
Hv6tJg1mdobNn15feWU837UPSArDLXSwm1IBLUfMhB2AxvWzftWRdW3fkIsPhspjCOo/CkHswg5Y
U+sAkNup5RVbP4WbetvkZeWmAmmwElY2eciTaoOHtRZX9x3KR2CrsXTDE+rKrI2ol/23CMWOJ1r7
3MOJavPdCxJct2f0/uFvPGEtczp5QAECxRgxzMZ+uBVe9P8sHlWmD1g+mvzlXgeGiTHI8Cxlk3Zs
ByDxuQmBV53kXl78JO8d/O4Vy7hA0f329h7ElU6tqgz6l5jW+K2vZsktk9Lm+JlJfz29+QR72TbS
ci5dL23dfXaFkLfIfqeTnVgxW/X2YBwMYvran4EVVQIObqLU8XFTQAS5uk8A8AKcoGQQsfWpqvgq
ydwYFMzQLkDR/md1shVny3fa4HzUz1/2E8aIwZ28NcmL6Hd5v0ZaYWoQ57eMyExB9AeOs+TbeHCT
WH7R0jZ1fdscreq+8K0lHHXd+Ix2evt4KLa21F/aQUjLM5oZX7e7SmamVx9kUk2/pbPX7kDBMZZt
EOvgFCXVwQCzXdGtVbkS9TMKZla6Qh6xEyuDG9s/AqDdISuDlKCncyBPaWhxXy+LLxJ61/7wuEtj
g+JY3+LLY6xQWFoQB0ULkBJVBi37yuJeMqwFYjvIpi0Uc+tCBM6dwXav2XsIOCoRWXzTDgvIqY0o
X36Elhh3e49KyHqgzcdurMXCKrDdGzMKQ02SdPM2W9ZTL1fnzMd5o0MBXCv796ijdnoq3pabF4gy
WMIlaoSDPcpaY/wVsBEKINpbSwjVUNO9UTnqhd0bTizOICs/NVRa/cMDjVOctXWyxfu7czg464Ek
xF06EDG2Z/VizGAPTxbOXXg0U+mwxOguB3W7bMYKTGM8KEo0J7tzBf3vvV/O2sLkBdnEyWOUORnL
tmEiXXvGYm1c3MUh5f0UOCOKFKOhDJyaMoupM8qu6Uho8T9wXeYfEL3QXNXoyjbhGgELklOvr+ry
dCFZXG95rM/mh499qFBObMIbJuLp/Yq5RqY3eBpAmIQ9X8E8DUDJVHn3OwUZQ1P6tIE9/N/uizrN
scc3SkKzNAqLqoNbXwE1KgLulQ7Xws2TqGku+aHqJ0H/yn8VW4ROiBUYEymxn3c4bVkDPOWGR5aq
/YjHV0TahxuZfT0FFikPk5Boxoie4tqg+3+kPr2q0M6tvR7Sa9SM9uwyxRxtfpdAcYFncUOUyr6c
POa+MTR70p80kjjYtdPofB96hrZQOL4X74T5y0VqShP+75gtx+BtWNLko5Q+p8nrh880KDfwToIo
WYeZeCatEJgJ3FC0F960sssgdUVZoTwesOvyrCwphlb5cGlcLQmlyK+4rT1NnSjwqnz9WSdkwdvT
M0GyWvDBwamn+WyCvRakiNRaq97JTbB8pRfY8tsGQK71YPHZd59eN8/UJvsuO+flIWki4UC3Y7XG
HIypkW9KwGBhDP6fBaXbzFywQdbN8PP3QNkYa8iYZb5DfF9m9Zvcg19sNiBbths87/tC+lkSrVIN
/NmeLjzRru96aC48PMTB6Nvu8xkLKaSzsOgSCxL+/v8fMOTSYeVe6r4DKkZFwKrK3mGo9qBvRZHg
fA5EJ12SdfvCKzlOdch0s6zeM1p7+FHqllHAepF2z5iQciepnUBz4VT7Bgjnk1WVlH6FEcZWNlqn
Sz/qnuvgooXPpCGZWBxJ/qJAjJ5sRo01e1Xb2G7OvtskxEqBQP01RLauvhNJlYxVgkuInuauVorB
LhLY1s5FyDxCXmSFOeMuOfejLIKMbUCO5BZcCSZcEiNMTrwrQya00ZXz35UhzQwPIyfXFCnnmFzl
YzFQuCQjxgcZIe5o7raWW3J8aE1T7cgVDXNNzkSQgufjug2D3uXE9twjs/fzbzBD5fT81FqBtq/G
zHWehyd0ve2ZydQ4pxIpGabO647yZckAm6QiJFP20pHa28ehMPzzse5vMUvFD42Go8AsNgBmrmA6
hsgU0bMTGyGTCRhKr0RN9TY37Y0ZMEspho+FkwgG5a9SQlk4TxAur8g9/F+pgUaatBLh1KLCP3Gk
MW6qiBDmMu3/SfEJvchfJCf5HMgE9gW5+iJzAEKyQAcZgYs8+xQLPPP2tQiMV2jgN69Cc6xTR1Ae
N9z2WegCUTQqlwLTF52DhYKbuEN+5hzXZ6s0Aqn1R0DFMFt9sVEYGVy3zWAPpiJBXVUvyjOj0rgQ
ur3T91IRlLsslM5ImDG0GlQCsBy1DTrD3nh1Gw3kg6Hn9O6DPIpRuk16I4Mk7M+OmWSzUdK1e0iB
d2SyffEBkYwgrWCEyWc2SWu8slFR6qj6HWUqNJQRW/tyi1JHSnc8kycsfuu00rJPKc+Q7hiZX/Ue
fv65b8yH0HVo54WNyCTqQvIgp0odxiyLf6PZm+LLahD5uzCeGKdfODPshNik3Bp/yZsJSPefza5d
ShJGxnVFReJsBb894psnas5sm2EjO1aL/lpic0Zs761l3XSoo8RyqV67BVh7UiUsPCd5o1HQrKFc
YqvNQGBYRGtY2u3sHO8MmlpX+CWAIlObdY/rukGHUIlLmKVs/2KW/N4LuefoOVvwPO1Z+QN5MiIO
YbxUCdtioSuCPeEfvWiY93lElBVoW5ch4W976v8xJJklms8LqdZIA60//WTSayLBdj9e1RwXTT6s
/XkV7actnVEvwZQHHAy+G3orpY6Ha4+IeMcrOdZPOianNNt6TK5kbHOs+xdHrwt96T8nlsSfOVow
GaYBxim46QidAOuxEY5J7OCR75QiwQtVvls8jixQAv+Xww+l+V4Nv55Jb4KQHgtikp3ABqGRAi+Q
YDqvmrNeI5vEkFmy16CG1hyoc7k2mSt/DR5R7nuTwHwyaVkEBGmRB8rp8UVEprG5DVwCaq0poHTC
VsmL92o/F8a9mVlKKq6tK45xve2pWbRdlqHuFgYsM6w4DX2BoHlbYQHw0Qi6czVMIlOg9EFEk6oY
SfGFmSffQXDCMJXUusIeSZVRbpxaQeMCIlIbBP6k4//LcXy3jH9Y2JhE3Tx6CNW6jPjrtxpe6y9b
HYKl+mhRI2JNoRF5no5b6ZkiUmXY2+KsoIVF/Gq/pQsTrsFMYRav+YpFvR682IUkhcUKkWSBJeL7
7PlaAUc/rQVoB/+1Fvr6NLJeSTchAItLWhspjOSno9xcZd4r8w+tJlzsL7VM1KQ5iHxNLfojkpq4
K6od5J64PGBbwv1MNvRkCSz4PsjHfwNEFV4lTZbQmVG5gphKddyziUlgttpcbuA4Xk/jpqEolQg+
NMyDwZT1cRjE+m0aOlhEWSHQVmw9g9RZwL2/d2V+v+8c1gvKaTT83g5CnfrRvlfensRrM3AN1z4H
vgEZWCCrjPlEpuoGM3iXkGyco0+SvWb9Zr17i8WC7Ol4GBx4PZZsVxdavBeBJgH9Z9GzLpksDQY0
/YF/oFHKgUEIx+ZTSp6ovDfNWaGNUD+OdLyV5YUT9DpcS/MLHrlKlggmIuI8sdW5mHEa2hgAUrQ0
Jho6GG98ZueAvXXEm22KN4lqRhKyo1mGU8TfwixvdTC3UtYY5KPV19WzMWJyf0Pz/SySOf/y/xnH
MCuJDlm1Y2R/c1U3J9zzakBodqCKII2Dgi0YjaqgKTs9YJCN0BI0OTsTFa4ZNG/HmyX/9OGD8HfN
3krD3aukpWVq8L3S6ziDO76ZIKC23J0UzzoG+pBxAMmv8xOAWcevNd4AahmlPaEh1IcAKNcnmTeu
6N9TXwkc6YnOS4fae7H74tPOX/pOXNKV0p/6jrTVDFuaoQ9iHuzJ28QzgtOCwrNsRyFkxbg7zpXF
IUZiAGkYUyPvNbokcv7OY+BmlTN2JcDxgchIk/HmH9IRJZy4HlQMl6f/Jn2FgdFAfybODQrdeksa
zh1whmMw0HrniozxOuov7jk+xqwYVP+FhExEpUyK6D5Pd0+gsKKCdgPZWI3bffv1vjlqs711YQhs
l12QyZFMhM+GyeluoMWvszd3Es4WjFySNd4UVp1WTIipsAOljSlx/kFZlTlIwt0iwt7u5zHNOWeV
NDtZig3JiGOrZwp0Kk8W41RT1c1klUNw7ZfyhqidYs2jFhCjN3oSdWt0AM4PkicCGOfSbC2A2qts
N0Y4+pyDHAojsj+IK/4HGEc3LCF/Hegi1FiAnqu0NH6gOT5R22iViG6IWA2ZVLqPafmnKthk0e1n
2kfXNv9afRp2U5z1umZ4lkipss1vI9ENUKu/WZVRptIWtjeULeiUSqV950azo2i0wCKCQIQNi5SW
11CVC6pm/VRR48GquBhwESL66/2NpDubo6bJDiotLIzuQoKXL12g6tsBSKhRr4O5VZoMWffQtjfa
1Uxd3bnZt0WSr4i6aBAKiZoUfyIOaL00euh2jtY6BLscBAowcjH2hW8wb4YpNAml4LXa2cOhTZIa
jcAr6BN78oCs4VOSj30jp+IuCgdPQpfwg9d82ftS0fsvv/PCShaKtqDUMAz4ph6dIGl0BEvC3oSp
oWynor5prBEHIS8SUu6aJujq7hx7waC/cTxbC3I9VBaoRi9VQ44OOCuw2R0YgE7eIfaitHlfDULU
7d7KsztT5ax/9vCBGNckOsY2ulYlcMrOK9H6teKoZy4LnY1/l9SVyyx5ZAuuz+rg/qRfIN9YTzwR
1V7S7WbqFs+TbQ8SrEw+Sd1WBcYbktQ3fg540NPmZfScKgeFE9HVhOh3TXHnVWe/WPAz4Rh/D00g
6LGAoUhtd7ERLYnpaJZ4+8bBBFy84nJaFUxKecGhcEId5x+t6w3zrJhf8dW1ydBtOF6gYlOA5D02
yNHL+6D2nUc2qnEEegBk8uQ4Tli/GBv3M5vdQFAfel27JbfoJueSiWxBe8OoVz6MuwDDtrKfDirW
ZIRo4BRajuVJShtHJhAO8OPsRL6ttMvE9JPz1KeHc7dXFHYLIBRUgX1EkpLrgl4B9pU44+EzW/Ya
zW+RwFtxnCuDV95MDeN90g0VmFLY2v5BlCczQa3xJZmWoI9A6yLjrN+Rx5+gxuWz6qSnQdOsB3Eb
mOwtVMUEhDBYpwZn7Cj7Wyawlc6OR02jHt2lUGF5NHKnR0iAW6kf2ByToGNTmXft63S5PCJAeaGT
OxEYAxumiq606NU7b7dKYejUKvl26utuPNJRM906qpOmeu3ZcNLyXSpMRS5E04RoMIyFUDHkIgBw
I5roLRqBpG6qvGAFqwykhwJw3Eh5wZSHwIGdU8UpKHlF1z2Y3Q4N0AsApj/ha/0WEBcIeDBjz+Wp
tvVG4zDmT2cSr8vT6X8pqaYXgyq3ENy7YCqjK37rXbDy0V0h9g0D9K++GAbQ2ev4qfl5Pbfs0b9c
gUA8X1z7VXHipCTH1gTfo4fjGAR7lzJ/7lavyUQSTM8hLK2LXQSYY/LrlzxJVYf50KMZZR8rxxdM
8yPHeC6iXOQCV+Yh6A0F5cseHpkhDEt4HzwiOPB9x76DuN1N7ehzbWbjlBEIOMIYn8hMHgY7W8i5
pIBlnR6Mvbrvx2tqWNjFMM2t1TcKoUkFWuusvF7MbIiT8hnZGGpkPYTNJNEzXHIaeKoVsnuveOvk
8E5k4hmnRNKHcQcDbeh8bQ9/Jesihnpmpb/3hbvIZ+T4wJFcdyI29xvUHBis3G00W6hDpLFNaMch
aFvVUU1HACkcpat1p4Gc98+CdYAuqp6N7i/0F92inKlQDhHnK9yr6oeatZAjfEbwZtqMHIkUD625
/S4AvUbRM+QeXbfmG+MPPcu4cBeHdngCMyOpPB7b2BUaEISWSmm1Dum+z9dS75kFE1erAaR2gDoH
ByrOobx03Qm/PMrAJ087VddQa+zTnKDaAI7Q6eCfwvEdHogvJ8NDVYWaBI4yDkKGMDO7gopnH0Oz
bzD2HP/wHd2VL4Xr+Cj1fOeEV+oCM4nICjaGG26uHLQiLXezX0kmNYeaXh8xxcjOuI+eSljkTpTm
67VfbakaXc3PBsXKSJoV4QRG2vZayfCTayN2MgTJMe32hydM9Cyk8u4dExqkYDWJH0VWDc/Q7sfz
9trbSypfrzLUnUrd22pxhkJBwnrcUvPn08RFGJF1fMeqDPMogyCu4pPs5vgHYT0JTebw9z7exaqz
/XHIytWac4PfpO8ScHuGhLzFPhiE7TCw6LRwa8zlbMrlRUDUdky32U1KRfDYK1nQ9964ju30aBmL
QRBTyjDkFKIdtNssMhTtVICwx6UsoQP5hbkEubHqkaJbJwuj+5iVZ6o9PT6zjslRwbOkvEVMLAoc
O8ipm9s1Yuf36FpcAMIJInfTTWyrLC7PWuhGIztZwdT5swkf6zpxG0342nwWjcB6e+5HfSvs5DvN
iTpdukhD5Ju8PZ3eysdzPQbI01no/ikCnPCFvvzdmdUAa+RHPtXPjR2vzTl3L2YHs0P0DeQXwyxZ
qBHo0Xb+1zZ0s2hcsfHf3ibr3dF73npP6ky9AzwYuWqhYKWF6IFjAXrr4/WoiZfogTj6uNYqpam2
sSByq6xrQkOMOd1JkuAkMehn4/3WxaI+W+4e2388cuIAZz8cY9CrVkCTYGmmqILBkcGC+puxszgL
5gbzEiNZZnuqZj8DsRdfTUxwZtK93MbXJP0fYKiphXcamloEouXrtt+UxlLq36tND96WCLBiKWif
7mqTb7AfRERW9fC/dVTDFqPsToWmMa/yW/hV/ZaM+zAUkSqLcLVG2mDyGI/00B7k0aYoImVkiae8
xOxre3DvRaR+OU5NN5+5PWQmENxhMoPS2ecgTZtFGS4aP43z5NnwvzljMWlRkIFE2exphylf5sO4
fEE/2yxTAhVhyZeJRMigAPTNTMCEpQdsDjV2OOjDA7gf+59Bq8plEvtHG2/xBnKMaT66PmgLYp1+
3F85AMA/qDbSlGaEwZ4mXr+QNsXeRLOIWHAnPZ946dk36sQ8XmqrU0Yvus440EdSiWx7gQCYaMt2
asolkkiVdFkGfeT3O+ufbykeTxsSfI0fxTf/lwTAqlgpaRI6/7840NxgU3Twx+MmIWTVKHzZWyE0
hsVRJwjsAq1ubcH6Hnwv0Yki1LPUv8d6pR/YrbSirCU1wlnsIEGK8l05Tns6vcVpraew5jRmsd59
9b8zLbP3cphjEx2PXrzIDIu7tQ1dkQNm36v38jDzhoz5im5FKBC8l7ICvhg1jKambdWJojkSv9Qf
92P+/MtyvuSEh6vZeKztmMDtSsaLRDhv6gXRLnBCEBl7N/W4Yb7rvdKfn5tjaiUc8vZweQDiQN/N
5zI4GBT6OdadywSpVcND5UrjdYUMfQcs3O83/W/zgexFVksWMJHPkXJKKajAzZrZzN+rJeevFUg+
VLSJgIQPpglse0VOOBQW7cWgfdmZb35Q09vq54mRDLwKCKaWXFRC6blHZe+Aq6hwvrg6z8107wvM
cAZanEVLOCdVO9yxdlMX1Tc3A+qIHMMsqjUwt0t/n458UmFWjCF75PMcRsrqhdg3hc/tqcPuKxGk
2g0veEcRAw94ez7Djh/AYkp//VysdcA2JkUqknwHTzk8s1CEgGBMZXEqoepVuqs6wg068BKt5Z4A
F1HQltWqf0GqhlKgKSuOA3z8AlH9VZQ2tcOrovP2cDJYn3End4ferByTe+icxf1msSouRTQYKpBw
7fMUOR7xaAOV8DK52qglL8jzTew/XEjRSojSSKqcvqk+UiffirG2HhSzWSP1MOzuHg12lh3WmE3Z
B3yJyqBnDnf0mvgb1pH9AI1bHEJiBZOO5Frf15DetAcU1+ReLOXcTgTwc36oyLRAFNBcSyswLJ+x
x1zDu84806iEwzFHHPoSX2zod8vu7zs8krhWTKcyxOgEvqzqguBT77ePNuMC+8D+dNrWB7U4QT/T
05dhvBBukMR53QNTC4aWNvkC4nT2uLtz1yqpEuv2Z3TD5W31IrlHeWqbVuT/gME3jfU9JH6/sfZk
QBc5w89P3NRfiR006ygZ20lx6ISsUvFQkDUGS2FPGDdvyebqLVMu1zbMf4W2EIrvUrLZt+LbFle6
8jVPV19rXrWZBkrw6IEV7gJfGgRi3E0D22P9XGVstWPWfqix60e77C+Rim5Qm2gF/zBamAyQq7GA
pYmwlbArpiyD0upcwnJ7+UQ5NKG8htnS/ek5pJXwYVNkCFDbDtuOKgCFl2d270yTHrhZF8l5AR2Z
6v8duWqGZyYonnQSBs8x7M4V6Loa/uZlYLi44m0P5JT35evKWIv8ssjCmq+/y+p+7U3o43qghn8x
4R/60TNtimNwskq587P18joRKbQHXSVLYQTlCnGJKEI6YpvT6s9Mn4K1l0DxnbcWnkkjL4GQ0UFt
L+pAKS3uK5poFBt/pzZQTx+CM0eIrjSApmtCM/64pmXI+yyvqYpT4oUBffoPB8/9AuLC4yYVbM5f
amrYRo5M8DC2iij7P6NlA2YYkHh/oiZ/Vc0LfAm3M+XeDJZJq0GaiwD2Un9cIuhhAP4gtrTzKdeY
Qs4IzTIaOyEREYgNWx9HiM69SE5RUsJW/0qXqqSIoFkGMXT6iZ1mI+ldY9OQ9TK2cex6rhio1vIj
W9dN1QDyg3CDBKvYeTFhaljSbAJCy/s3mRhT/OTWhGCPfiLMZlx1uqC0VFDHNY7XUrQ0+KXImK8y
uQmQSpspSYqxEhazOQpRjdMhvxPaO3IAqcVgZnByPiJP3H4iFoGe4b3XKkfijSvLxqR8iCzsGe9G
+EbnV1Zoe/Kq1E1tRcasn+aShhWP5NWNn7phkyIUX0G+pwpCWYk2H6kUwUNCPJumW6BCUFMmu+it
hLh1OBiTYj2JNsH31N1CMEc3oY9aw25YLQwJjn1JkC8uAY2Fp5N/8vD6/WlAAFmzkM+eCHz5/GeY
2n8klFN95kY6nNjyMS7EArcnnnSOS076ljPFoSmtnQboBG8nL9pERlXfWesL/kW3pCsS8dgKNvp+
qbilM2s6dHgXIaJge6S8hfKnk2AC04H78eSuy5FdisU5sW9pln7Hh/2yH7VucFdby0rjvWw1g5TU
8mixYn3EVk2hwPuuvT/ZZCfZ0DHYPIF7tx4B7VN2pVr1WtT3zs5OUxuZQOy2BNowbLZWW67yYMrZ
d0dPglRpJUK8mFmBpwsBf763l0wKx9KaqfwG+t+Z+9tsExbMNjUsnF47MX5LUQPkrzIXk7nuzDJi
+pvzKaI7hohbFW9mYRQ4M20l4xWbFF8+CBbMUQZs6uWCjzS1dJGZyqbe8DX0GmaiMK7m2oBs5nSO
9/4TRbmmCSMxJxxyBfILW52mnQElSrBJlllNMmoqnwbBjMmrUE2fuJuyVhGCiT6FIIsmgw46vTYF
AZDxSYdGbdQaqvgFOrcYQdSukT+aIvym3oaefKMJyGEk9BxESK0Hq8ICqduB1bZm/4zF1ZZXGcqX
Fe1I10eV9GXw6iGgP+OuJ5e9aPkmqpmr+IuF/Hu5zT9rFAcgn+y+Co8cEFKE4O2YFfi7mUfEgLoy
89TIBz1ksClY9dOmOePZ28ozIz7hLyj2gWWgXt4nigw3zvAw+O0u8KWVz1f1gll7aUF1ALCBFCPH
o5SIipwbQ9j/nR32p9xGPYaiAB6MitCVVmERJCHdcNxGFZ+aNvlJmbTTzdKB6eLqmoBhkUmyTIBn
tCVpA2mLlBgNquEZXbVeexejlQzsnm4p7xm+BLvfphgqLezIGJHKd6Pcg4WROkcpnDBzBsApQvev
5l/HZiPn5qsdI5Hp52XEeuW1c01AVOIJ9mxpL81qu7Uzteakp4BUsIVFl6d3MnG1NAwrNhKbxGIN
8qnhiNR9q4IR6MwataEk13CAxfOAxNJfiAz9mUtcbbbMu/KEUphT5fLdyP+omDVZGGL/Caz9tY2L
Xh+AHld+ACzwcPl/skgKMQrH9oYDp3n+7lTf9cU2rYCr++JdHM0aHPaVxtg3/w6g2omYEE69RiVF
pdwVyQtRpuaJJmaa3A6NyBE+2+wS/Edwo2w4jgPSxdiZR5c5a1AP+aAAn9DRy/QnLCeR72kImqok
41AgsVu8L0qm2ynsbeSnvOHvHbGk4CyZfUhGlyHQML2X1PbXVUVE6YJg/shevxGmbvGdQiwMq6UC
sTW+mByQiktI8OAvEjuz7YDRWrEjordYbLQV+6cIMHNmkWXcSxsdosF3RbKEmQZ853lJdE2C90xy
8LZNySZ5VG6NdSwHsrs8FQmr3fixgKut2We+2ELU+HUFnLGlOA4hKI0ENxfXm9jXKL8gu+b0ChNx
E5X/Gty/RXlHtEvQVXqkYTlvAygtqSv8FEGJaThOwhFQ3W9xhv+WvnGhHmqo29SKYnkLfMSau4q4
hN7SPw8A4aoN2IWgerqDItJNUSJb70i9K8obIItmgQy6JJrCk23G6ZF+i9pIQGm/kIE79tL5ga72
7itD6r3yfaQ/I3JvyBXPvt4bKwbX/z2o4JAO4foa37xtiCOVHzv0rdyaQW963B9ohJCD3ccopzxv
F2FDWR3wAj8KJWyigS9jXUxasE8+sYOeigdllAg4e6HVNGoHmZlOeWH0yS/hk6qjGFq2UaRHmOWp
xAWeOS5AsuZTCoM7MzRahqSWFVqGV11BATCqd+0sTaJLvIy4WZtdBR5vhCsEN+qJok/hMlu6KvzX
SIWL1ZnI1tS/U1DB6JM5n36I2rSbGv2qXq7sVNuKxaETWmfyvr/WRs7E+0BIXX+UL/AM87i8j+FZ
+4O2I8W/2dbbD9Ob7UTg+FseFLPabDoaua4+qaNZL79UiMreemqWpKgm52h08Raceal05raMggvM
BjIH59phLWgwqz+dUEZ3PCx4ypOQgUqq139MFBcJYtqWVm6g2ieJoQ/W/hQ1QmcxWAhicYof/bbN
zZmx403HkH4p7dZ+rygeEoh7pgHyrGNqI3oyyRlscb+RN8UQNVwDN+YhS9/TekM07LP1cr9EAiYR
UOTeadf22v3/iyVeaWJEdZ1ptgXDwBTdx6MGgkvXXAsY8egBgtGx96WK4rTiTLFBjmBgGY6fyOTi
r8GrPEXIosr9MTlzbsxzY6YSqskyOhEEY+jqbMZjiYBrxNRNsHN1mITuW5zIeMLwhs6yj195KkPf
hpmKkSWXAYtBsMaAth0i+dqdmcz/trL5fOxqO+nzskR7RiQt354ywE9Z6bBqLjZXV/fv5jrfH81I
PLI/jc3YeTIvz+09zhYDMf9/WrR9rFUgP+RyrvAs1Ct7azXaLnj6Pv+LeQo1nwDMjLPaRky5cBwD
rZJezka3yb2HP5XNpBgq4Lit8x16SSHKvnjH+htxp2UwnZfRUdfLdWaFcVYEHAqhbAsSgGHw61Cr
cEWRX0Z+4xOcWPMp9xHev+H4zo0MIuDWQYY40srZqTpPcBFsejm6OdphzA1nMJFl5Ru2zMSviXOy
r1F1Q2YIT9o4zjb3X08c3lvz+W6kzBdMH8JKNIne4L7YD102bDuHADv8qia9/VJuUm8nNlJIFTGA
TAkdFwn6AaQqdlaRJOrh+LuZISLhVOzIWYH6/qNm0EcAEnxwW/ZCLx12Pq7iz7fxcRfTY0DPpGiz
qog7EgERNiSBhFa9vgxxwuuUMIojHleNMnMc8herWLUFMZzdnNIvZnDvSRtVcpTN/NRxK5Or2+0X
UhwRaka7yVHJdYLLDj/HLyzym9nxHGY/5nP+2e4eJvEQv9IEAu4b/HgVLN2MOD8vvljeDhhYFroR
wnWRMoSQPVf7djj6oQdUAMruHUaC/QszU8q/EDyxuw1EpH5kW/+I5np2fvum1OXlcin9Eo8n+dXN
jvd/rA76nYlDt3A2FE5mRkDNNDrKrxoDgGQoBtIc3v2Dz/S+3BVMS9tq+2jmEVN5yorUPa+8lPhC
hYeGO5JErG60+HXhUSfIrvCwYBfG34lj+9kfb4OieF8YXu+McSrWPCmMglyRoCyMw0OMDzFVEUPC
f0qgSE3tNP6e7KFcXtMWSyFogMvNtiWavo7oAFgWl3SfXCg6Ks5WSqseM6D31NnkS6JcX7uopM/Y
HPhDJIWlIhx9u7Dieh+c7W0/hMFN+je0owFMIJHZWpfB+xOE2Q5kVy+GhLkWniPK5IDFs7HmZW4A
PlRnQk0ix8p3qY1QtIggaGYNWmlQW5dMc2AgD55ftD3KbKGx/Xq+ZmmTn//cJ7CefYV0E4RCH6Cv
Duts+vco2UzWp1Ne855IzNrmmomriMRQrJSAIiSmbA+L7LfvVuwKDXw124TfbXQwmgfAkXFGZ4l3
N6gAfLA2RRf0jaXS3p+ZmVkI4iLxeKMrIaftBAqlxUmqkz5JerlSMaZm5EYCAcfvvkyA/Dd5ND2W
8gPSh9eMdYPdGgOlg0QjQDCwyZMmvy17YYTF1ZI6LaLxpSNgzKl5YgHW0YG3KWF42vv8mRd6gGyW
B0rtYLBM1wRxIEdvnWDrACZhgnmwhDlDO0ExRuktfKb5hGdysxaSpVDcSNvLjxWV0hqNx8k4VrD0
7M8dFmPBr2QEPVhzPDcZ2Se7gGvoZ0ckXbQag40z64jdnUlsN4RBP1hlPOIBTZUyUSpbMorANgPe
1zUTQTJTINiEVkhrJ6szCmGjz6z4kaRwTcYJi4jtCCaBge+KWAsxf9ZLY/OO6+4qMVoCL61LmsHp
JiF7Ezlhz2jREmekcUlFexaXGqoDX4Ag06HCiPh5dlXE9u5othOn/Hj57J6q8XCc/482ifTjKJEN
In3UqnkfKywmrIiprJKsYvusL7yIYQHyOuKxZ6HRDiGN+L0V2jpbT4B5xIPu7umcQAnS44gFZ+Vz
gOl2B0XyRPin6Qdsw7hTOdJF/uX8WtQSZ2uD0/AHfHlL+K7PirhngLwWI4jsZE+1ZzoEQVzSbbQX
PWWk9ToVFUdcvFxSySqGAhR3xp6Pgqt+ounQnWh2G1oVGsAWW8LGUIGzvwh1+FkHsWf6KXXiL3UW
ozVEJ6cjU+TzpkONvBYt8VXYZbHaZ3ZZShepy0unXxVSZHOG9Vh9EJzywRenQjB/6hU14W941u1I
VxdW1wZlXUO46Y6CEX9ZEREvnlgua4EFlFG8OiBFgWQSapEQ6KlEFFZ/d6q4s69hbn4PJzw2+uzt
y9AI/m8OdMl5EgRbFFNQPO34H38xzgNtA9uUZnJeqgmeeg8cMur2GJwoea0WGPNVQCFKSqVxF8ms
qO5W61v0CYs76wh2096lofGZh/VaZ+4khMv+XHfvyW5+LmudgASghVfzNrgZ5z6fy5mocR2gXu8/
MhvMi6TiXJliMsNtBLUQRH9YS+6cShku7ANRU0VKMrlEkeq6YKZHYBhbDgFfcD1XI6sE2X0IamBq
F6mDjiouGQNIwIMYt/tOX0/ag4yLeTk6mqrNcTxPP5vAz87eLnBi4GIrY5hceeZusxpJc4WoUDaQ
VZz+UzY5ZsLPq3WzpZaPZBbUyGGVfIBvUcWJ/bDdaTJVVdl0t7+j6WtiKTEIyr1InYFMdmrA8yqB
ccK+47gpNYYdQD2bdtxXacdWZeiOwOs+dn1uxAY4t7VnLjs1ti0LXu0TwfeZDCpw9OBwb9NmJ2cM
vl+G55icaxOCrzGLMWgZ6oQ5KRfDv9SlkB0AWJwi89p6idW3knVaqLmLtTx9dSpz0cL2tC25ISXx
s/uRzdkDa4TMp8PBLVc6az1EfUOQVgG3OB3cTrH0Xug04gYdwOWh/CRDdaZacyyZJnzsJzyFztJL
5VNxkTAewLE+k01bqBqbZMR3mTRqBRuXN3nBi87UnVf4tdyQiCZM76U6abtXvjkoCM/ENF5Spv1F
cAGoKKGqaocb31jXdrZtVUzUvOztZoCQqQReKz5UFys/CEDOqvf4PXnt8JNoisjSBMxBCGDcl6d1
Jti1YD4wRJAWH5lI3kPXYl7xwmuwaS9JvpvZ4j1JMGP7VbQF4Qrgvob+wUitHUVqADV/rWPdW1La
7YCC3ChwrHOXOFA2Sc/kwav1Ap96DfyNGlp8IJuGt0U8h1J/Wws09ZGr4flm9GdE/7Z//E7447OK
ZsDD2wKLMQOGjAxXKfP3GcOjV2G7NCRZ0pT7d1moZL6g2W+PYrNjnH/UkKoTVUocqU4eH3ugLHLX
xTy0cwxEGwbsdnpkszGcm1RiwZKFvUvBCg4Eh6nDY7LyUQTBYTSmP9udiym0wk37MLbnuSQXQO1N
T0ExOAIuUVDuEfln3SHh22PYnHMs6TbWQeEqbdMlIIlu9xKlzKSzbbnW7X2gBwR4g/6ZQHzPCJop
vljQhKPzzN7x2Vcr9ra0XiX5gJd8vZsR/VbJRykAmaSWePh4+48/KYJtr9lBo+2t1rDV3U/81axc
cFHXJ2sXYHg+EJcuS1K38BdLRCSz01GCVnfGovJ9lg5ZS/6+dH+oatmDKTZNecwxTvV5nnON6d7+
VkbYMUBJEeuvAh3h4u2rxBhwUWDHKdzeLSO+5BlXoPJf1Rv3N7CMTct1klNYIdX6wAZ2W7YB4Hj7
sYC7DL5vUYW/IOJyb/tlyl0Am0PtE2SrEOs6jFjhpwLM7Gvm6gBM1jy89YCrflKckeDiXwpT6mkZ
N60DTg+Lso8MDbjnCmdkVt9CLvtCNYKNOLcsI8wJ0iHa7b+L4GbHFX2juaohJvRq0qmLOnV2ynl/
+m57G9NJVwds28C2h6vrGBX+WAQNN//zxx9HVRwOg/Yj4A+TEC8CDea13jXmIdjit5rmBbP2vfjG
C+2QMRuLKEAsHfx3BGNvB6iCu/UlNbreK/jVwcGKpghrJ2mT+uZV2osrTmeVaVqioMdwObDp+C6F
lZjrXkPo6qKSJEpGIhJG+LtnNZVcubIrWrdv7sxrHvOrWml1PIcI/g8jPwu07dgrTX7ykdFk1VMc
zy2CKMDwDK1YTV0QJ6m7II8jbZ9CVHQlf6uioYt+BbjSE/j2LKf5wWocCr+/L+ujZaenmyf1IKH3
4MRMmsIgRAbucreSmEFeIGUxmvojkt5hOg6T1TSi1R2OHch062BgkIVXGIxvi3IRhXqTYcEo0tc6
z3w6U2p0mPdD3V7McPchvidKGuLzy934+J4fN+NtNXzqj7WV8mMFYSJMnwkFLKD6Vzp4yDrSpUON
ou0Eb3tWEvqao/PhtV0Ev8bWpKLTRCD7KKIuhCepH5XeH6FxcnqK+tyQ87GSvKOhfFVNCOd9n2KD
doFGfQDoTo9bmjQBiNQQOxIALkFc41eM5PcFXALqMhndIhvBYkFgEUzpXRUAIq9JUg+LKD7NerWh
o9E4sc0HE43vWc7Es92nl9JOy2cJmfi03SKhIjC08mE1UAVUcnQtyojhLUDYB7q4uv2A6zJI+h3K
VlbreqlWWemAbfDJJOxsgHz7/fAjKrXwNlVYWYzr6r7dAzjVO+i+SzFqGLMuKUAgnr542YQEjs4v
kvHVuhmyX6ucyd/VeHV1ZDMd6MnlA9hMHYLP7aj0kmCMYmMq/2IElP6PcsLAlMurJfDj9A99Pi8F
JIBRrHocXKtYesqtyRntgaYeGdVO0TjibEt2Sn/NzR8rkmrnJ0TsQh4XvASSh2meSrK0xKp7NxK0
7rTAR84i7Svj2vCaVGszNmip1LxINW/Td4HJRDcsCCV6bDTmo0glsisSuytVyhMygJfEuYghje2F
ZfVmIWtLCIs+36/QMhwWlAH04zGUneFCB9cA+uWHXc4/9AsEmpZbMfRHQhbuP0pdAyNyT6Agnd5s
yR/PSa+Wp07d5XFG2ocZsUmUAT0EDJMNg0e0KOrDhxRe4O+7y2wId1DCfNh3/eOuTz5oyivqSgZK
bLYuhb2ks01LymBdTHB3IKG0zADy+DiSSWMsTO1yWgPkwpdmXvNjKz29I+/AZ2mK0NS49m3mWHKS
2mrTfn5L5MDGKykkwCfgF1sU4w3rgPnjFKjwcB0WjkkbbDF5CUUbzeAT3sU7Neq/II05oKjwMGUY
gxSbGNV1+mQUcobtqzxQtyGDspbo4UqAQ9RmGQpCJjeSfzm9pn8lZVX9Ef7FEMNBq2JzzB3DQJWI
S3tcKwMQLMJ1vOygu6ydKDdfprXEUgAhCQXQoCLdgSs/Z4J1b+qr9RQ8XSA6n+8zW9dyIWid47+h
xmxWHncC8kfnK9FpwASMBs12c7Y5fIe7C+wvNjY6j0GS3Kl7GhWy4dBj9n5P1Jc7PCbohuBzpOW+
cOF/eIG8SXQpXfA314URxKK/wdaDA//GH268IWdzJPPRTS253st1NHYDvOGj/iSXuCOiFqLQ4yNO
/cHRbHVMkY4+zlPQtEilYqZlLFMiHO+qJ8VqcD73o2JZWmrr6pDMdABxhPjaqkb14zzvnT5gDDlY
40ICkk1XVcNcXjnZYqwgVSjxJ7w9+dXTVQ/jk3+r8d4BLELuR6wA7bvmM7zxtDSTF92cCLnu2fix
G6QNUt+KSRgtDbKbDJ16diUF9eA1Egqh4lGGyLAuMpaMNkaza4pxZZMMzYr54Elb6CwLOMJL+oOA
/zAEI9qgcH/aYCaN0yKdRvaCemstPAupwhnpzo2yWyOwHu2u3HOZRJK2S1OGlz+EBvQtcLp3VWEr
kOCCLtVrXYRrEuPayQ7AH8pJOd6qJlTzLIOEwpIOpyKKZnx8XiZII/TdZqCTv/vjwrl0MxTAXShW
D0GfvyDrarQJLzVafnFbbbKlXWtrqWr/OoDavzoxJZcpKhOxcv2IYb6GkdFTpMdTEbBxEptyZZum
oqH+Obe8X2ZYHu/LzrYc6VYGdBBjVFZkh0A/naf0pveACvg/Pn554VYiUDMsx4l8U6pGyLlFd8Ls
IVTpR3YjKZV+tajZmFqGL142lGG8B6hbOPsCTNbzk4eiNaGIQxCPAq23d+IAc7UBYTSuJ5ovLKr4
uBTZGRiS7h0tPcJsMh9y36Aqke4Lvew+XIzjIhNfzgDQviEy4//IVFfgFhs/IRPRyGzbsp4SWwG1
kDZKyvXlgqHn8c1kzxh+1tuTko9laIqLbujF4CAIk974QP9D3gpW/+aXd6NVbB51YT2UhXbGcPby
3NFIbl0ZheSWN52Ez46TqVw2Tt5usrfbQ0M3+6AIx8TPdFXJAQFtYklBfiKfSxUQ2Rn8phKfhf2G
4QGu7YdYd7kD3Quqs0rCRrHyBAFCBuvLP2yRUGu4To0qO/AMp8ASfKn2eG5K3pNPfOdK+qu1Poug
meSseH3Gh4YM+EOLbjTd4gh8SDhGFo07ylK945bfPvncmKw13YxeWiBB9DrxYk/g7ebkdqH9I5Wl
5ZJZx+z3l5uvcdn7EmK0oq52cNPvKXMmJrGt9gXG6ofEkSQT/SI8BSpy99hUDFbh/lUTnZRp4aDE
Dch55J0+0Wkt2aspkhrLvPYCoxLB9vyBuBd0E+na1rm99seUHxhGNuFJKwZiZLOOlqa3N5BUNdMR
AmkJvSGEJ8fusEbP6uVEXPMnT6tMU85NTd+Xyb1SxmbV6JnHt/7bbet8HspybkJC4LLBftPnHI5k
INBMmESssFY1Qh8t92SzTwhbrYZEn8R6rWXs527wn0oBYlEkAKciebDJJgcWXQ81/ymPsH12vdFu
vfzkaMCSUvlDSewLlWynkJwQJgOJPgGau5QKFwSFA5AE9ncCs4wY4eBHns2if5UK9t5f2lIKZIQw
9i88v7eIePrQApnbdrnIgcCw0LMxCUEmiGoGeJj3tEJdMZLM7X6ZvlJxUwB1DZ9x/lHtuagXBWU+
9sJWnDPKZ8Tr4b03OfphN/rMsV4kWb2J9vZ7Nc+CxRzD5GGiHhcq1u2AXaaXl8sXpRRJpeu5Srx8
pIIBcJSB2BrBUOiO9PIekX6qBJ3Omdcu1+yUHmhD9+kCX8PyPQs0IPIO5Ks28Y5/0os1Crfcw2Me
lQEtSyNiehQ5m93FJSSRC/qjNur5GEPLteAtlYkxQpDTYoqyPL0MXLhXDyK5it4dRtSLAFG9uHSU
96+q46r1PPprDnO2A99tWemBYNQ0kuZzmWTV86SdqYfLATqDhHg6C3bntXt0c2EaOhLo85Eh92c8
HT85PuuXJgaE5K30l0hiH+/tQu6wGfaagQhDBdP/f5Urnc7lWZDOi1v5N9kswj10fGM4ajjujqa8
b6JwHX7Vv4/TVMc2jVdaP71juyfZ5fqN2Q/p0561jzQbXWtXp3pWp88uoRXBGzqoXnVWlhV4MrRJ
ShBWZz1aHLlswd1VKuQYiwOjS8NvkSYz6E5qvUs/A0VYJ9VRdyyv2fk5hQMJbQo1T980TUmB9MQX
J5HLu0+O1s6X8SltDKDMD3Rn89f4bx2bsRjhmdbu4e2BdKwpoOR1Z4RX0gWUEgacKiJ+7HRMIHac
le2njrhrTKoyKcEIInBsvl/vH5U77ODcFMu1znhuO4E6kbZKBUSbFzsR2f2YNn478iN9jXYa3EIp
Rk/pJOSKlDOO5zMI66sHlVhvwm6NAs9XUvScUwVKF49fgyVLWVu6T91PTvYL4G/kxdy+b+lGmhwh
KJ1AnWi1rus3xc0p3uZxSRrD3dVBWzdFNHHsGOaOPMQWftg3mdCW29IqoQLknO4bbzKLljUvXbds
B+MMwkvWSSOCtR+hDLl94EaKxlP0e8T6Wz/nZ5CWTesEedc6h3WU+hkCRTia/9xeTkHnM/EMz92H
6iXuuGqzDo6x11913bJHPsagh90KXmD+flPs/K941OaLYThW626SBxD7dULbWq1x32q+bzGTbRFE
h7zrfSo1NwdfClCTcBeBytWVqcX9uXWHvM66ULDEmUzdZMp0ZmF4E/1nmt+lFCjIDNKJHvOZnzIL
ps7YeUMoyjsMMy7pXgRbv+Ozz+SyRqW0lfdbwvib0EcUDIroXgU3IECKvoZhU3OJJJ1OzLyKm/yQ
EWVUJnL4uMFpT87QyyEGmkvDYJ+Hlm8jPv6uxe3vUqVrYtyPEM6JZlJSMLQhR64dSWNB+EJgsvwL
+tBTw0Juha69G0WbYG9K63vdjsRhXufa/labUOBZaNYUdXersN+oBXUFUbOWl9gbO7OU4GxjERJ6
Sf3hmWdiJ0SxtX8nCQXgUXnVfyxT7hLcoRJF03d2nb/ocYDJEN+LYaPNu44FjEDKRUWkgurRj192
VwjFhCehEY8wM4ZMWSUyt2H7BB3znNMaRShLdrc6IaplvhJHp9KgUfumtrAzEze3DYY8fx1LBiC1
zsoVw66WfG6edh/ILioOl6RlGN5m8cvmX4lH/W3rvYKTSPBlfFsh/rPCevlq7WTDr4s0npBtjdV2
nNJwJ+GZlt8aviJaIfJtTBoZ3MnvYw0/AqDsbRlmIxsrucpM91mqPE6nKg7tvk2JW0rKsB0yHIoV
wd0/u9WBPNumduYwsGcNdD/NjgkSL5RZ8wA2FQqYG1wx+om06zjn2hc+OYKNDN9K7reOfOIfKE3A
K/nyNsqj9eKNSTru4PnRadPDEsJpbhSpWI6VJnfQEo1/jpIuoVMj8ke21Kfs+3sjKl7aZPHh3C/j
ykkddj6KKyimPKkvsxiuQXilCIQOMe4LaVp0zsjVstC4T6qow4AMLp+66LAkrOApLcUJkOJRcMpg
grRjOZ8Lgh0YBOh+E9rlkxeH2ZW+llRDWtN2MmmNOeYt5p4PTMNVB2m2z2LyZwYGitE6xlSdSwqW
Bs2k/LdCin7EwmfjgiuFAoZ+CunZRVskdHDZtoW5EphbVKm5F3Rswvletk1PMHQV9dNykzZIjSHm
5UO++o1zWJmRdiuq8X1xSohcTQhItpKgXeKJ79meOEHohjxVSbnfj5/grqGml28TT7QeaoE0p5Xm
gqPhq1ERknKcd6k1LDMOiS4jNkyYuQX0aSvKj1DvWhb7H8EiESK5kS2Wd5loZLKL4P86KFz4utsP
UE3V2fuDaJ2IL7RptqCRqN4Bn+kVcDnxZx2fLtDPzn0ah2pebed7xGs+1D3mL/82Y2UpqA49QBlI
ULoJKMrafd1J5VzYdPylhY7W2uxfus3qaCKptK26klHMa93H7xJaY6nUAPliYun8VV63ByvAFgH5
QA59aEdGDvTV1GfGMyy1s9UZp2fgG3WozlopZNZT/gssa9e1LHRxnneYNTt3rgq1XUbTN09H9Fue
2KNZl/X4aY/vv6ic1E78qiFV5wop2ZhtekULR7g7mM3NpUNDylyImfw05wYMsuI6CblHCbTY1fNJ
MY473K2cLURMhXN5FzZjqkdYbN2Biscjrbp9qoOn2/xGmQUj3Rmqx96Rw03UWhMC61YC8SDIskFY
qmj+lHZfsyQ3+gGXzcrwbuJXY+sqpEc9fCvhqGQy2nhnYfMUsQeqABtHHQ6YdrmtyJCh7WjgeZyX
fmlQZjrgGaOAciQMeoKWOqxqS6BZmBvAWIL5l+OVzh30e7+73UWKjHLz7bu3bcTf4/XLPTYKE8uJ
a9dAvRzyUrcNQes+y65eZNliR/D0ZY6NfDSATRLs6zq6qdW0h/bqXvuDoZeX3dtxI6f7Ufmfd6vb
tEf2SSBg1hbn0RFEhD+CCXZzhLjPRUH7/N/WFvJdvL4jRkgd5p+wXSegUlIwvqmkMBUaYokMzvCg
UsusPKqcz11EjncYAOIfT+7Ql/ig+fG73HwRKpoTRJF2f6Z2IK1h93sLIcYeqLqn339pjbPFIfXq
p9oHDhYpecvw2webbxhrIlYAFTs9hedvPoaPWxvBhZjMFJfeo+ZH8dV49Q9CL2pQF2ThuhW3RORT
LQfDGcpICm3oAfYkl8l0Si6QL2CHwcF8yXWOGXEyN31DDj62eyXfRV48RNLb343VxA8oTKTOhFgw
eGxRnGhkh2oqF2BH/ldi+kM0CMQco5ssTI+QWows+FVJVj/ns9LS2tgmemP2/ZNihNZGZGbszemS
ID5VSjxQiaYuai5LFi/Nn55eKdkm5U+rgwvDRm1/HL2OBZ1GalaD5VeZAEW/mXNevUEmdCUCqPAb
Bh9UmImV6IYfo4GUjHZMhJUuNgJQ6w9lK31COQ1oy5Yk7IP6qWYc21NZXmmdvZpbVbLZRWv9B4ur
zZTaYYIjjrJlvin79778Qlb9XbHeXc9fk1qQfSippUerdrOTsN4oggObFtTlTpb3eBkG8UG15+cx
QZQNMgmTnXhvuZGMRj2hjrRyJAGkF3dTx8gjVndNtYmPxZgT4nq9Kxujr9hHHV4nyJ2Zfx/3yoeM
jVGh6q28a/ptfSnqLFRE1wmH2ebfSaxDPOu9ezpsOywMrWsf+IfNTfsi94dw7g+jnbgRBSQ4c6s6
Xwrl4qNmUxENQPAv4fmyybeLc69vdNRuy+Jh5oSeDPcnePQkPfxGbmgXaiMeymgbTt4ZQDHHyP3l
hwx5X45tH7z67NykNJFRgCE5yw96zl7T49f6LzNW8kHINWIjQ4sB3yeZ91eA3aH2AjwwecxTje5u
8kG9Y2QCMMwoQf0ZI8gno+WlT/Ninxzu67pcJ5t8aokKGTM8yuHDhnTH6JszwdJKmv+oJBl/fGEE
/PafyKTG37scxED9nD/KSDpXouEY+wUtZH1GOoRDozGo6RZJQ0gpDNuCVf2oyiWD2t7y6M0NW89A
3Ky5W1VCHnGzjuJKVmJjOgirIoMDrOCqmSQDfeEUfWgyzddpmoL3+sZkT3WsBCQkGm+iFDvk2w0L
exVa27rBsEjUKe2cOmoyLjOlFCzqXMuGDesk2eDh8dETOJXGcTXQj6owrpa30+JGogZC+1yVk9Bg
zbSrMslFDIA6Fudfrt83Y1sHd1cQ2hs9LfjOaA5w6T2NR86yRzli2sZnrDD2v27QTHLWTLmcAY5d
1nITLJ2cumVv+7CMTn8deArdVawXk5ccasCQGYfEp4HHAxJAEgX26XFo0rosVcNVTGwENlLOJ88+
CfCltVCuiv/u10Gt8LOo81LE5wuUcpQk9CPNPKPaK4aqWW9HAPAkF9ewvJBl3JzIrpPycyeD0GB8
Tgyw/U+n7vbOimeoFLQnWdxnG274R/5e9R0jhhfE9YhfvUVAsT5Xfyzt81NvQL9aeqHR1C76gaYg
LpeUo3nknVWIo3cWwgflmb79inUjZsMs2CM3PM8jS/SfvpRGfiXCXIPJlpleYyiKpmxfs34D9UTX
42xaEouS0vViiutnFI1rA9ZW6r3JYbdQMSyfiA9nv/QlAMrBu89TbAGX0M6TYABX19clf2rJVjbh
QnBZ307qQ3mgkEPKthjNwGBTcqx5v6b2onnlvxCAFnAtuJRMBSTVgZ2JA1FPRhUj5/MjkjSHekQr
kSfP7xShNnUhI3V2m10dl+4FGMPf6Ptuw0oyOsQEWkNftlAQs4ezAAYn68weMCHvnB9LEZBKzY/R
VxdiNcApAC8XQz4S89CKbrk5SJfjEfA5Fr3PLdHRtgFg/2CU0yO6yxFjk4MJae1uEX9Ln8XhXOi4
OPtxgyHiQ83pALzXLyhlGzgJ7hra/BmyFMxl9Jm2ZH1tnQ+6Y1l7+Z1jmzGRlAsYNr1hWPLpYHGi
Y36C5MoAvCDso17qW7aciizsQKJS6K8slczfm1M8AFIuabuOCh1CnqxI1W6A4MQgCB1gX1VOeNgJ
a7bQwI2y+mpGO77+6iU8d9pxjfNFwiz5+lM4dD4+lF+kURCveOvBE1BcdKXjDaiXpU5gQYbZrRA6
r+50bZ7s06bBfoIB8WbTA+CeQ7PwrC4HNT9Ma0z+crgGIpDvaYaGla8gO9UiYtrjOjdmxjfYp70M
UjpjhN4l4xbPoLXHbwg+vQENVJIcwwOyvMOpaUTwuxrRQ4vP+775JW/Pimufd49jdiWb1/5NKwW3
xcnBJLuXKRwNEBtLOnD8X+8AbROUrX1YYUcrF4G2K32TExzYrklS2KTMzoXbNiQ9rIs2glRzue+N
a41BD2CfY2b6jSGrEuTKtN6E5sMYWEH5J2/dyOh/CGROZvjbKKscGE1vLPYsGgJXCuN6u1+gzXDe
f9tS6yJIsgedBhXUlvPNE7wsbpSfyqJbUZ1V74gyYCuD63uWk9d8iCz1r3nZZVHjH2QOaaA0GFK0
iEtmQFfKvfvVH6YThjihMWJNwqMgbktdDaTAdBlCE3m4UpHJGDl4nN3bQb4q+SD0uesxMAK/2eYh
lHNs7CzxZlKUyT3AnolRZVQvMKdKFTEtWBKDOhzhRAjJGcf064ysDe5g1nJY4nEEdrkIi3LoKthj
C4TjIhmKXDw38cLCSn5gCjeVOYJGiqjAZe2qPZh8AMbe8kQLY/OHuf4n+tmlqnshdApJPfl5TY/L
dC2aou0p7Q94wvNzaM1YI824qwCjfGH23eCGmNX2vDyKt/U8/8HLTaTIIMudcmPXPfkKk7ucQvQu
SfOugkpct42ciFC8/CL2+ieh5wBiShm2MFkmEFy9FLNnwoYIqbQJd3P0nX05+D/lcxxTeYUfbDIk
/mbfeiZkDjsB98ucxwEQDM5h5028PNs/2NWyMynLNhc12R+V6jtIBZdlW2YquDue9tKYTOtNomli
Y0TSqsO/j+KTi3e/mTWogB6uEe1UYa+L1l2l+MDteX5tTDgEtxeGttkBjYMX9J8d2sRyL1bkJEEy
lmu1fBGkoBiOYeZ+eqfnN9dQJq0rQKGJFeCrsS4Ap3QxknJ/sIrBlf0ZIMJtWPtxP5Iab8IcVT40
FUp+O8H1TOtUyF4hJmRkjYQnSGoxIfWofkEyWGiC7k7b90h/TUi/k+VvAT0eKuYv4O6y0Q+APOgW
WE+y1t811LVUIyG7dRiHeieyWwgDe2foRUwj65BgDdKFmbTyPt3hPQjyqJvaRS4qJxuFeoF67W72
SLT5FsLmXeVSDvRX4g2LzYUFQAk5a2q6Gi6tlza6y5IbZumEavUFFO3nPGYAmARy18EIf6EzS0xt
WJJlYo9P7OPIpTDBLE4517Fl6hzJxL6TekQUkPlf0xAUzG5+whBlbTZI94xKgDxPtCidqQgCqSqe
FdPY4Er9fQzAECoPPtJJG8/cVW6HWLqaLuCDdd4c0vmgGGwu3wjCyhQgpfmiScYqNClGS2v2Tvvx
Sjf97dTrUNIQ1z6Y+eOAooZ9v0T6ihrcOOO7xi58xmW5LEUOJcrEy+5C83w9ae2RSJGNWVtTzUbk
IhkTyX7pF2pZF2s8/jzAXf9cLkB96rxmX7XAtkOY9GJGxWrt1fvXbtr7HnCPppOYEewsRFT8MJGC
rNurxwRN4Mn0jOdqwuiXOXyAUdeHCl0hhRjse0KJ4f1DdViaVklAttiypkdT9kvL4YB1BpfBumBZ
jTjYDrucPwNgsNWQEoatugYw2jp3kFffXqoDUsoVDOqB7VB2tMFL2xbfCmRCYy6FEt8NpgfH/+1d
Ir6U0UkGiSmFFm6mkaPuOQnOpRRrHBu5CJz5tzODxlwwSstByXJjX4Ubd3MTB++5+c7h3ik+5Ept
ydZockQQp7RCkjA2WHa8AR9SPhUIxt8QbsSMyPnnax63mMd0sP/NBTodtUadSWcUNTf+xPSLaxYM
Cr7teGkbbcV3qZrK+Ny4nsYcXqX2URS4LPOh8HctN+kHJvGOfQ6xZIn3sS4JLLwuZs66PFyU4yq4
ia7VBeFC5UyrvWX/flGf5S8RC6heFTdlIGdfBXe9IVEASbB31RZJQww1oWDpzJ7uw22pJXg31qCy
wqjo02itYG4nsrcLYtjvt6jzAWnN8UMY1F59sMjZgMZ+biJ6MfznnD97brEpceIuwNeY2zbU+IHi
Njsvc6LFvxMxkLAyqHAP2MqcDqjwjifynKMUEGwrkLq3bIXyGOsIcvmOzIo1gTIf7y0gcxsw5AQl
upZYIDVmI4J6x+15nmQQC/MK6p0n4heimsv3O73oWELwoUvcS0t47CrJaS5+pptUbTX1vsjK3USG
Ta4K/Ta1ZxDy2L804XqiDXMF3a6+ZzZju1xVoRhUOF3Cgu5YzIaYtyLjlz9aamqjlI3zmkCW/isD
yoH5soJP5n9KyfW/Fu+yayLZk3g75vjo1OlZhphJrxY2zbYBB2FAOeGilTO3EdfjjWzsVwbx5iuy
RKNivPtoSMITGK+6h43iixXImIC0dqygclYsgHKkZjhSZoWirDT+jh6t38WyUfBIOp0eDKED0oyu
5b71gP8ce/1ZvMnrll4+SJq0YxcaGw/jVGbwobaIv3q9f4K0qsORnvJ2wvZDHlD8z0068N+lTGdQ
uY/Wiqt0GzEjWer8taSMQSOMPqnuTmnIO/s1mqF0QKZcTiB2lOReD6h8aObHinXvNEQCM8ZjeC5M
ElnUuCM5/k92hb68PGsUM21kAxxDFFJBriOFjCuCmUyOVmqZynmR98g+u+R1rEDQIxccXwRka/1j
XCxuMVrzqWvuAKMUjbSto8YrV6qRzcyiaRSEeGnB9Ry6qKBvxjuXCdCroMxruj+r3ESeAORRuBEJ
+ntn6+TW+fONeZ2TC1Wk01dHE2yHiOT6gj+WJ2nqHCzHgBmO1wd8UF/mgp9F9uHciIw79S2pvUTu
i1aZhYbKfCjkis7yum5eNwrbWxZEAH71FkLXRHj21bypVqdj/6PCkJj/FOLbgP7SOG2w/Z9+5ZiJ
XfK3i7EYKj3Gx/gayFQ9BIMLO58X2Uqf0PyY/oZ9HSO0xIaWLg8Q/89ko/dQgfNVhMGjcN63nl2u
mWewqwqgzroCrUmH6AImK+kj8/w9EE3Wy3HCuwPemARsM95cjF7/BByUpz/UCE6FKIYykvho+0xw
mKMqPysjM2WRINIa5u89hYaESD3ZIu0mI7+CcabE4oCoDdYXG71+uE6oszrTyWWTGdK1bo0S+FA6
cXJKRgeFUhznmpTMQCOCiKi0a35e6/YGRT6MibrFI+ySC2ASVF0NrgbldxykAzSg7v1yB+ypsSee
MsPmL+0PBQ4orhCZhGlHa50kt0tgPPhrtN9DsSFCJIcZnpaThLdCZszK24U2rLNsbZ6W1czAWUGO
cM5UZ1ebkLxA+pGtYjnEeT5ILiBhumbTLMsZR+7c4o8BErYriKSyIgVpdrItnEi6v/ZOs5AJXTnN
+h/3jljRpielIFkeVASKAnwPYz6IlV9aQIg77eXoV7+iFa2A9xS+4LfOacGDHLqDjTKIAJeO5BSu
WSIqYYuSaLy4Kp6/W8iohatCwYjg1av2K1r1/LBCFgVpAX5PTdXc0Xa1puPbthThVdxsrjO6p0a0
bGJsyA5TQNaqtOLPhfMxCifhCqYf9eM5phVDghZfJjBmA9DFRar4dA4CpS3KP63CrVpyPuK6hkco
IO28MacjODrVmffaKtXGs2M2gVDlt6Yi0CkC7MLaFIUmKjNrbdXOmhy2hHnt67vkvcdjyqpjiM3C
4tEtnZMfw2nsXdMYUKyaaWDS/fVGIR7uMuxZFyFGj+s6x6AYFg+r2OKbVvyKPikP+RMD2AKQ6sff
l/RezkvPbhenozMRcnAeABYOqJwleZa02MUTdnjjWjs6R6kHpVN3ZRBKmLcGW1/IERN3J3sWkiC7
eiCsexQrAzuDKjr4AWHtIz0YNEDdOOfHRMKCuIVCC4T9Zn95sov/NGZlB+X9OsqQbP+KpmGEPXyu
j2cWwNJZ0lstugSyK59rddleduiA7/SdI/yQ7M+WP2irYpT9S9DAvHX7H/AeE3xmkBDzDr8fl/rV
cSzdni7nXlrPIbcJO6i2Tg2H0mxWze3+2p+D/wrnThayfGYDr5lU/+Wp5SbUXnfaM8NbXYFE9pbd
MJINHTIghLJ+dfdYuTCsamWmCy2l5Kzl5/Kh3scqMcJmQClQ0q/ry2dUjPSnCc0UdEk28nEBPz82
ir2d1TU1fD7RqFVPGdVtxAW03HpY9wBIE34j3vr2TP8sB5+r+Tn88dfmScMpslrmXE55KZ/xSa/V
DOrRY7MvfluD5F8HetAkzcjqtkaUXUtCLXVz956UwPX42gfQZrBuoa0a8bb3s6zLK6czJYnU4FEB
Gm7fRk/3e+tqM62SqwgHrdNm0BMMCxjqvukwkzBwyZ87Zw3gYcMuHyaAVNaardbSNybWPlJZPeRU
8zb4xUMO9x+yShnT/3fgF7KQsXgJD9/FDgYbParwnXAOo4JLHB6Svgf5FnUpnev0mqowqMXyvBBk
SNj6/o53CDUlm5mBEcaCQqS0T5mEKr9M7lpjo+NExFb+w8fzULggJJ/kPSngZdeMkbA5NhdY9ApZ
5f6W7sbxprlJpDaNcKc+mnHOqQORhU+rHFOZhiOyevvt2/Yn2mSqX/4tvqlrGrEGdLCnCDQKKJkI
7M1vaAMrYPBB1V6e/0f2PRxd3iXNkF5u+KRMig1zofB6aGWAHRNkIEL+a3AWWCVUJ+XBHelWUzcY
JuDR56Gqzqx9QABsDlXkHlCEALSEKtErYihnsKbCDZmVzupH6PMETy2Cux2IiYXkG5sjcIS3D75A
heo/04kKtdrdssyUTA7vO9ny7MMXpKq/WHly1q3L31AMVQMzyXt109BQNauHasoY/988uSdh7ZAO
w/zwLSC8MY3NuS0V8zoVHFtbAFvzLyZjiV4uVfsUlqjZeoWAfj1uLthabj2R4rKqEKC+//w0Y4UY
vxOE7ghGYcBqaH1fu2ieRda1EQ0SouHg4RgCpIIDWKe8Aik3p0pkcIJLhlePIY0cM27pXjIIOqjq
6xE+j2hrJoYcx1K7NtaYXq/NoIKms+lZN7hbCaqM12Dqg0gNVhhSQck8LDopfCUckenjNwzNFWs+
Pt7ZFDnboM/MFYgdvXq84kY5jhyUzt+8FOzTVjmqxz6NtbTpl5oBKb4Y4OOJBp22aBuiRxIyBfVK
tq55iNvwkG8I7WIHzOq4OHEmd4BGf9B08wGe4AVICOJSTIK8bxEeFXumKE3FdWnKgokjvisKpg3U
vXB/mkaB0X0mw4ySSeCfBR2ZmHeYMig4nU3IjRNeZtmsXrvThuSLJYdB9ztF9249g4LyfTR89dwU
B3BJaIJi2qaWXYa1+dVyl7c996g8htjmEnAsCx60iybWqoVeyclh9EmlkQZqLETSGadz7Vqqud3y
NH+ke76tguySxUrwG9quYXF2Xp+Dn8EFYpUh/DBZI/2GzNAjvMAPtKD90yN1vIs7vQdjOB7yMbnF
pI+LQ+Up9aDpk4WiMFeLuwKuSvuFbnBxfFsv8+3vNzLzK/uGpmemr1mhtk0272i0RL0kNeytmcwY
TOMAiUdR125GtbmS1eOeHkt4XygC66jbikL2cFxcFqfj0lDiAhODZUtkHhdpwBL9CqM9JOA2K/fw
L/uzx7ZchvzAslXA+nxQO0hPJ9upnTQvtSt8ZpvY9x07czfmvxxtrt23oDeYIEkpm91rL0nf6qbE
UjHyfuulOp33NJmTnZabGEjjenaWEchDloxtoOtmBeAznvVpFyJAOe78//8xYDvftdXSvovDh/mM
0RbCRMy4UTRbjFkX0D/8QZb9iKZMreK3VhYIcZF6rqcm6JUtWPRUJ7tP4ztf8rCyssoEh+zQlc7m
Gqytqn8HigQQ58SbPwxWPPMiMAzqV1gKWEwOegEypq15ByL8Y1wOpmNxadyYYnpfF+k6erZye73Z
8XGMI/hkfL1LHxuXmPItd6kQNlHcGor+Sr9zJhMq8HGmKDcfuK+25rOgtsXw7Cji7yJCAvsr7wk4
5EN25zFlUCfs/xRKHoMylFqnBFiAUnllTIXYTSw0mf2kGfj1Kyrt+G5GOEQzet5r9Chzq0TiW93B
A7Kfkusgx+Y3jGxrFGFms9OIsdN86l3eJz0W1eMdtEFmvwPUXoqJI13WPdzwGdkjUmMDqHa4vUSO
/NDTmLDtmsA4qpu4j4nJG75yqBp0eRfiYzhPDPIALqo329jAD05V07Y3KysRXMfEm7miQpm4atEa
lT9pBrsca4x8BGPKukuUrqyu0NC5LxMaL9rOfq5ThDZ5Kmzy31BKYgfiFHXGUzISt6Lg88911kaf
jbNST8T4azDS9e0yxojVyjsRsYWCo59NuwX8GJ88sZacziCNiPEXCTm8HvRQdo7uyKQMgg1k8GuK
B/RiyS/r+23X4lvVmPAL9U6KW1kzb88DBrsawiwbYcbc1CT1NNbIDU+4rkC+klxoKzhoxpvU0cZ2
eOHHEaAu3MAMZsghO6M0MWVCvD/KrkJwR0YllmhZyTOvE89FHSnY3zZqOSv9DmP+LU1lu7yg0iWg
VeVOBbp+47NPp7mPqCDWQpZ8ajZEZRXNGJDfZiBvprSK/vmfQajWRYbYAqsuJZkWUZuflBMcoY7C
/mUnLr+ul5HPFn/G6i+BdBbEjyU4qMcOpfGLlXqz1OR8pmyGdZPEAE+o04vvR+XuHq0qvaRfH5H6
QuGXPrOM3Lx9YbOkoAE/Xi1F7/GxaOpMRg81XdRaVdfMDmhZ0V6Kf23+eP4sLhcKEm81S3b/onQt
HpSnlDqcazU+SY9XyfnA7tWylcKGvU0qk+RR69yHGaG7y1kZqrrVNu5WnZsxvrjcIHd+8wa7EWlN
ZrHxCgfD/+0reqAiA4kpGXRw8dYlw3791F6iFClkOK7hMLLTacEk29ZOfAk2GIgYT+30VehR8709
sFPmonFNJUyL/zLCDumNvjrSALOfgrjahk+5DH9yHAyVQZtkUf8SVjl3yuztl2PgG5+3ExWDDhB8
icPP0BxTN7IyfoPQJNc2RrfaZU1jYbj6ZhdA48lcFKUuHy55C8YuDBC6bfFYw6qUkDhTPfGSRMvD
vdclwyBJNrImzlL44nuzeBlBBlOeL2iksJoWYKivBNi3tkkvUBLX/YAtkadBjC4GYCpRjZa6CucN
LmsUOPP8fU5rZOU6jE6pOn6UnGL5f8YtJUtjkaEaTEBPVcnbzH3wWoCFuEIe8HeUtQ3mn909FyLL
ZEmXkH4chv9DaegyPMWNuNiucPG/A9SHOaDnqgP66do20+dVrNlGREnnylya+68Y9EMNpYmVKVZB
rxuvfuPA5REnielc7/h5B61EwnP/r2Q0+A8wxC7QJ/pm5zkAbSlXO74HOpH7TUlGa0j6vhJDqYAm
qEJlYEcktlzIoI6JjIdtO8gId/QemwenwgocqBN3udugo/51T9YPiYfpXbN8nF/QMrPtCsHCs/WI
2RWjWvtoNPwjQwGL9K4iomrpI4EYJD3uA6KImmOquPvAbi4Bg6O1YP7vpKppDAVxqvoEg/qz2W1a
H5R/zAKJ6XAjnF7fNQwVvbz847kJhsS8961Zobx5njCdZEXv0jIBDWZhcBw71SUSklMBdU69VBnr
Tyrb64K8QWctCAXqf6SjZtvY2TfquwlnvuUGu+0fqbeG+MTH5215K+dsLwLatwRtlj4xS9qrAMtj
JyFj7AM9bCbDzevAevsRf2ZsyV2+6Rd6jy5Z/i1m8HHsVpKHkxL/nRlKTb04Vhp0EAh3iOXxMvWO
tmsByHBtBFh2IVPTr+DUrenW5MZw0BXJ9vBL2wATl/2Ajmhoc/SFFMId2mXAYsH8DA/xEHyneZuQ
JxnmhHYDpgM3oK5poNTxZ6toM7IbGCli5oVO8Ovv4kM7psi0eANqZugjOVchfx0F08N51E5GpVsG
uzgKp92jJETjTbAv5/SGeCCjHpHShF5Ifr1wvUeiHRxCqAQ7te6TowpT2H5pbiGXIoC0TG5yP2sR
gSvAP9T7QjR51emzMrb32ZwP6xH0pgrenyZCbXnCLbeczNYUIdJzEMLoAHk+XqlXeg6PapF/uFxU
1egh6IjKTrtaKqFzjradAAmbXPZU6e+NzcMSAr+1rBAoNhG4A+OlDsxgqOiUDxdPLuXIECrqw76Q
CNLxltTiSbJiWwUc7TJoH3ZoqW2JQpLinu2bOjGwG+hYyHajlQKVr++qiZYIczFsW5/OS/Co7eat
+rlIKVLDPrrl+21mqFa3M9XXiYIg9/LqCD7OV2/t9ipIxomcgd5sdGpaLHSXAODd6Xq2WOiUP6MP
58sGIu5qbCzB1Dfq/9h4uOBkkwJ/rxIhu1IpJD+YzVjS5j2/BykQtn01s0wTR2gg3EbqJ4Tcg2Ef
BiL8FBYfUfQ1+A6PtSEEJRryLnUhrGlD252R3vzh2bA364KExARDYk2q9oX0yJ+1pZfcODaIiMGZ
zz3K6B6+rTkoU6MyJymp8Qe7zoxmq1dAZjuMOHymcnXji5feAkZKNTXNKbET746DA0n/z8WqlCJ+
uwNTAybriygJWsQb0BaFq2RMBE9TAd70aUpmvc7kbmrw07aOpAWgoi8RAS/EGXQSYVZt5aEvqH5V
Kvrh7WQtio8KfBsOSxgyl/CUxLf5TWrctsihff4uZqDIYXN7JBCnJvKz6F5Zy4lOv2+SRRQLKEaa
CvvwzBFyCqsx4zY4D4rSX0BXMy2LYO1waQOLE8akmaUV06tj2FteHTFSxDnH7bc4CZZ2p7m3f7ig
ckRCtG0aOToQFPwvrU5t7VevqvH0mNMMk/BwthyhWIo+4+BpQkVRJ0l7iCaz93hqNAAXMsKYwb8L
Ml1+YN2ZwNaxQ5vaYUaB6qnWVjd80EI/1vdIwMwSbm5Dy3gpGObk7sfaRHZwClVRuEqOgqvT8W26
hGdJ4zlbyZgODK0bWouh68m4nnTiGiZmxGxa28J8Daav6Z0vLci9WnN8Yxq3D1YMnBLl+qxrGX+j
KPYnvxt/WmJmJEdRarEemIdrAFmXzDSeqcRTO0fiRlACm5Bc6lESRPJ9xpoBkZMZOpW+GNt0hlBv
GZv2YaSguGlV4ptUpJchZfF4lfQN9AhYfms697KnLb9aXdGRdPGadY3eJGvmZSG79jmsNul8ROLT
iei6NJWr1x3I2QeQ3nwDTTCFzKnpsRJg1t/XK1e/iAVMFJbHgBmnVT3iXwg9phw/zDLN0SZDCsSI
2h46esKL9E9TovYK5XPy1SCtXgjrixMEb8OCVk0q06PIu6Gn4Y1f7IvKROlj9lBqSHWImXdqrpN4
mCilWJjpERj3RiBe/KSIdmB122ZG/uY144aDsPfAvxItkDJI2XMifWVRaoT46cUdfqNG+3w2NFUe
P3nzK/4oXYIFhP4lNRz4vm7L4QdPvOlNjNVnlIdTYHxx32g1BZyMVicdge2BNLJq5Mq2w94ctyBD
SxNYSE9L1mgHFJJ3iZZY11l+6BFVAnlW6EIszGtjGMjadqO8SelG5Zq6jDHH6IomeZeq9hw/aUVe
VrH3wLdQ1XH3yte0GN/iEeHRdxqp6OFsi1J6WCChkhc6KYARLTI1MctAV3PiWpV69meWFWXlwrzA
4fs+w1MEzBzqGOant0fsoX0JBUxfY4MMayzCpqYI1ahEx6b9yd1cbHRs0y9Rd7MYkie1SwbxQPjR
pX+0E4ysjNao03z7nhrODycMINMRO+WQWQviD2kTO4uyr/TmcyOsr4G0QNVrbO4NsyTNkfhcHHUM
1kEBtpmXHZWKRmaBy+RJRHIzqz0iZ9y3/7PVwjMN/4Fw/r2gi17vyyy8Yewh7lYBpDegA9iRVxcb
lPk29GhU/i8UkoDCr+dz9dRxwdkpv63H2zfboMxugCHUc0TjHeCUYSiDVz387UPOukUBxfULJ/kS
hYAwUBjwK5OI0pSb0NA5qKPGUmp+4r8xfv71VauVNfMNz2R6+YKU4cUNV5VZStAHHDY2uvJqXJ6L
3SlGByYvkA/6nQ+90cE8OvSfEFjGk/U7X68EZnkcu37SbfJnNZAs+J1HP+H/ssgVKgY1DblHIlkH
WMm3LPLgWECCTql/M2rjcecVVFLzXr7xPYDVQMVZA+0QZtvT2a95UlVN7oUGaDDfJfQAsFI6JvHk
7ZirMpiX7xGU7Ge1Ydkntbn3j3yLSQzjPT8zAqCqbE6jWoWZHSD+QxDyyRZQbaOpXp/RgQtxmdDJ
d3SwA106BO4sH+Qz1TmKCxk6ZRD7M/1CCWgpLqetTy+RWtYsf4iBANiqcvHELISAUO/hc6CSp42T
VD2+kQPpVeb+O5CkLuuEBPqjtpCjrwnpQ+7HabDIMwl6N76pM/aSnaVhzlvWeu207DtBJoGCALe5
qNZbF27qJonwL2uIt8NqoIFUGjrVV4+dqP14QEx0QQfrx8hrqTWbVVk4v2RZuYXTP2T2c0t4VGvu
luVTbbol7lY7zys/+rXrMBrtW441Fj+BLKvZkMYsXU0/2yzdMfw1PxIDHic7qreo3DVA0HQAlztv
uGimyE5Uu9UcDuGBkdSOROY+1aOwI83s+AharGnJ6t8UPJjF/7UpOt6MZDcXml4njXPJDVsOtkR3
9FueeEa+3soi60EieSGrZ8+10Pc3pGk/3PHLMIEbYuLVatS9ZdB0327cEDZaGt+2iR8ko08U2XB5
VbbWHG666FZhGNf1kN8h7u2nZANa80EOJeYhdYfvXIyq9EAsdtZuacVWM5IrvR5EljBe+y0OpWpT
32zN1/6jlh05xMxq8XI2OX7mPRZtlhuhK8yY7Xvm08UzW+9AxqnB/77srJXluZfYL5Gw8/rARxOK
/WZcV8KNX4SseFP05bnfeCgHbMy6eoIonnlCLwfFGna70sHfapdlYJHlyjjAuXSqrjc9lY85pE38
lzm2gCQUZTBrRnKQeXDEQaY7VI9wk2ctyM1GqA6Iilb73Qt6c4Xr7Od/jQobkjCNCgGu9wgxsOtl
opW1kqJ3WYUXnTMCsXDX0p+twOQwxfnuyz8eti/ftR8qgKK8eNlab50TxpnqXb+48cL3ELle/y2K
c1TtdF3D/1ItUaY2gxS+mvE1FgZDxsdME9cneGo7lNb9gSIF3XXcYM9AfpYh4uhcaZv46mwK3LSe
rcXE8BTQO/hBisQdit0n4nk3mT3se+v6ACD7RIy4qySYlCNhk5Pn/8i/8o/RK4ZqFK9GzcWqawiy
aoY7yjMEFXLyXWVwige/SV0bkOynst2h6SdupEZMCziNTqyk6fKqh0f/aTbI5mZdhDh5XxK5fSy2
PtvarAnVw3SiIf2+sWklLtlelwfvGUj84bCqFMA9tcerPLkip1kM8aG4mcvn5nZDW2OUhvca3JdD
+80Zjva0UyQio9I0jSpXiTvXVgWDRuVKHSnikg4XNdAsWv3GGAlpTVw9BLP7QVDtXfdpH/9lacH5
1146NHwvA0401ftVahZBte5BoEusn/HDyfYax1sp4nJifi860OOPlqmlyBCR1eVXc8BdxWFxJMLA
+HwurYRcUoFziZy7QotoNy3qfJgBgKQmpv5ETSfdeEWkwkfksSbqiRRJBYaH5ZFno4kLWD0eZp6f
A7qghbhNtuYNyi2qsTyw5ED+B/Mzo1795SCAKAIGGoRD7W5MvWNzDXMBGzbz2grqCzpNX6o2+9/F
6KxjZb1NyDnO9o8CKsXGWAvbED2EXi/CyLWEJ7MQwRSc6uVTTCkiOAEbHqOHnIQDCdVzuAsmewcf
zCFUyRzPGSStKaP+KtFGu2dcSC1pR3jkbYTzKd7CsHQOWA83fxYA6nJHvEfBHUrorQTzatdxEBMA
+l3xpelTLE2ep6A2jxuMB/3Cd6lzl2ajF3IeLGZhG4/+UqOyU/0SsbWO1l5TdROy+FJgtzS5cNhG
ESibJEsanasmbsNKDge0keV2q2oXjVl6nw3AYsKIFMkLLyS3P0k9KCaTXxQCs/hcfTvaAPDzGTo1
PUhymFqghbm6wd2GI4FchbvMJIdoHBHDUy0OapbsAJNxH0NuVBPr4VMaFmAHjwzJDB1ACxgLVdtj
w3s079T+IciyJ3YSEweHhz/rbHZ2WOA1clRbNQXRCH8aimxD2rquN3Wa7aemBzJGK2swpTSuHqJr
rYrKwJfttPd1E7N6XFWJ0vHHRtCSjyh5kZiqgT7B9GjNnTnIpATN78EEEmzlJGr4fMkwApjZtDfg
8uU+jlPizB+WVcBclFdmYWqPkBCJCuPqxlIF2gzmt3l28k8rJ4HPWqpiv9B5M9clOsfQOc4g0L9k
I+1RXx1zbcUWfWRtcm6R3sVuG+3ZkXDjHayqLJqp6CWnrJPifxzhGKAbDEv+hZztpfGAiCOhCauS
cKp25QPqgfxp7H2RDzMrO07Am/z7qkmXgY/0Y3VK/hZ/o/otjnYRpt0S1PlZPrOZO+fXGnopZKtS
I/tfNRwqAivz4lye6u/aCL2JEwhtLSMX0R3YzzQH35lkEQR9v3yqsTbP9P68nRy9fP5g/1kqt5Ya
LSFsZ5jNqWJq2lbQHem0ZVe2tIhpXPQdrgMjAkLyIdFdR/jet1XlR1E6ZxX1LiX1eroFXcXZ28HU
b923D7EwUl7IVMf5skocZMCYmmhin6Dm3D8g57y16JZWAXVGzTb8Ur8uoss20xtxgr9mvEI0w7le
lEB5eRp2UtdSPLnnceS46pfxPsRAlEG7mkl8n+1O62cblK+xZFPS0QoX9/twCwZ9wXatphqe8Vxl
Dp/HGi1+QPMzsoJjP9GsaOa+AfLuAJ5BXuYrdpDKa1xllN2amkhX2hK0m1DY3+p68Ii0WEaxp5JY
+x7W7jXoxdUP8PXABojyFbiB/0ppLcIkHIQQ5aJXZDiOo5xX5IdQVlNO/kdDB1SP412cFCIO6Dmh
OD09AnLovo+l0jidmqpQu2GZHCi107Is/Q+l6Y1f3jzWlmx4gIPf9+CINSa3S5FKVMy9FWU9RzdI
AzC6Kqcxfil4ofNWlSpEEHtVah6/UYqSRhoav3whMrgz/44O5N+DUEGnIafN7ma0YsLnlzIdXsbI
Od2ahgaKhJSa0a6enlsLdUQJsR/2XDjrI7d2jMWKK0LrtCdyzACT5ZKNWrhIJhkG1RnPUYIDit3J
aVIl1QXLAw6j41TGuwYvkndjBkC176nEEf1NSUmDyI9Kc9b9vJSX98z+TxhSr2wpel8iOBb8Phig
lU/8oa88UBeXXu0hF5PtecznN9vZSu7+JrWuvac+mgH5D8QT45ji279PM+f8zfcA3O6lWeyKl/6T
N91DYy7vhr7Xsv7Naoe4yoHpYarwYlfDnZdQ28VX+nbqxnk/uMZuU+9jsyoAAXqFLoDeaaPLqnTG
yE/51nl1+N6JeA+b162mi/1yzpy3KGV4//1ObN6R6BWGgZTaKluG+PgGkD8UEIeln9I4LTgG9hhK
bfrGBasFlQ+ow9+CwbyGzGEGc2EObc+G5u/G48ckz6DfsUm0I0GMWikC+HSe+zfjMDQiLanKZVcx
8DihAhcDzwmqQ36fCHpY23lTdkFICevsA95C3kJAQSw6v9zoN1Y88UKEYw9M9SgNMKbPLAT8+7BF
BpZwKGKO0o5OdGtiCBMhq14MPfv/IY/rEARUqXJBqxdqYQEVxuIgal7kf3QnQQCvSKpvw1sEcp/2
ED+7HTu0yuEstOfaPJ51g2hMoJab5x3ZkWrz4OhoqPd68iA1020QdcuqZLzM7ZJD/UyiDKVri0Dh
S6I6WKVhP8s+oJT4nakCWrMF0Se9I6KqnJurWPO6Z05b+pe7/9qrBawU/rWHkKRrkT0MHW3UiKCS
c36XqkX6oWaqughGxggbGRzIBp+gbI0gmli5vxl0uoiXcJD1Nlz4mdvxgHZeRkU7HUcxmwY3LPkF
3dN8djkzAMu6M6Y5tQxd7R2Y2nj7XsaOy4yCc3q2rcj7dEjLTt0z11NWAxFS0aFoyQzU6AE37wl2
kjDc446Bic3HTi5gnY5MpZrM8lV5yAXryFoOiG5AD5xiasabFgjfhWVS8zvCYhUo5XmvG2d5iizs
DUnWq9jyEhdSEynZnfAATUo9Bf6lZ/31TCAy9Ngnshmb3X16tvfNZA4FaYoPfr+qUjN+E50Z33eQ
LuP0NDXHOu6k+UqHrna9gZeXfJ1RHlTtRBNdVm3dq2NpOhj7eqOoSykU8JJBw1IAJ58lz+G27io+
97ztOCMjI0Ip2uJyGekgSR333DYg4Imf44qSG9j84S4+RZ9lxq5a0C34TJJxdIWQPp73TEBWSRKM
wtFtfWRVdK2QFQu/kGK2JTawx4yKm9WSTC6qnA/URCgvBlf3WD5BKk2UrvdVQUCCla1Aiv9fM/et
EWdi+G4bWClFrd1AKX6he4SIjQBhxSAtCxTRR3EiVY7ErBhk2LExLI8AC85zCWETxFdw1Vx62di4
yNWm+jkgK19PoJRVBRT3zVS/1W1JAuAY2rSvymahwiWlVDZI++GfrjD8o6sHEX8J7Qt0BqHdbcS9
BloBOtc2y/SoiOlau52N9VOpFDah6Q5/rWZkgt41A+abfgp5drUhwsMQtGGFoVfPstmKRfPM+Fz4
iSLAbAxfhpzBxSgBDd+daKhHtOkqWkQIp+oZ3ApXiJ40RqMYbe/vYCYnLVyvIO81SmB6sHWtwqQc
p0oouUYQGQFddVNS4jpgEHVB1ReYJLeQgSLfXAEpniWHy8s1NrCsb4QOm+HLOGlHdULfeLvAkTBi
RERsE30M0PKGky0/ALowDJt8xQXiWi2dGr6bhKg813XJQAvtfiMC89M+FfIWHUd+ZhVau5qhP8LP
kawdABk0PvRcKdIXwNz39DmXBPQf5C/l5VaoWwJmyKtAShsJgiYamcTtlWGpvyOUoi2oftSygpn5
8/yEePch0RgLPGrhaXALewN/liMSHEr3gkkB8m5Sk3NVtnziFTihqRk8VS1JacvkmEHtsVwRoCgf
ggmL4ScmIH1WQ0g+rH0DSVI2s135gW21wLk6YIgDysfhbLf0dcdrFCeOarRFhwpN3Nb7OFK4GHH4
NHmPzmVX8cAHAf8BbMM+9rwoP9PSs6qwNB6ubr9DMhwWMDfi9kPB3Lc4+9csZX2702ei1oyEH3AF
iP2SwBaGpJO0kLWW7jYnjiQu1T46kmDtAEjjOIygmPzuEpxDJYHeHXfcNbBNoilve+5xFHhPb+jT
v2GRlOxPnsi8dqU0fv15dNpW/XbINvrHbu+gNknoSfm2FxUJ4zZkQuPgXIqMhlX0Lqf79Ugb6NLU
LCQ2GlvQ9hpXY76d+9iGGXDds5xySlgPoVL/nFjwnceTCSHc0DpZon4oKm4mqiTzLcxOMIMfO3N8
NUD8kxRotwhdGxlOATxi0QNP3tcq3hfIUiMha4z7bMaBO4S96LAP5Ei/wd5NzDPrZsszAgKKpUnZ
psfxyCoFmqycWxTQ10TrOQG1jocIWKtGJdQTVMorg6VCR7DDs9bR6K4mFsuIfOIfKQu9YGy8ubGZ
axUx0DKBoFm+B/8Cc4KqB7Yedv4vqFdy16u/ZrL1tSnAtWKiQ4rYJAIqKVST3xvWDMDrurEJJuyC
V0Uro9v3D7Vj4lQGhLyOIpOnvbYsfZ963U9nBTU6nozaJAhNrjkegQnukbiBkS7jDtdT282mKyEX
lggcBtbQ3X92BgLI/+y2M7vDlCRrq+d/8f16QjRBkiEpz20H2Iv9CXGikgyLm4uuvKqVXloiHcc9
u2uEe91fJKXD+slx4Eg7wQ9btixq+M8MT39T2v2Id9yqCFD6QJb3I3mEjKlDbp0bb91AQNmkjpfN
eINIjIYaG0In7Og8y5cBGAWgHnhhr8En5CR25eoGoF2VQm/+e32bbd7xsQfpmf+CzP3f5nEYKHxQ
AET49HXx8CCwptFMTbZRGpXCX3Zu6Iomc3DLQLKwy4rPhU/g6n1qVQrjBhHUuh/jsBZfoNmyFX0i
78Yvwp9ypSjjobkwLJ4CBVzT5RE14XMPiEXEPWFON6ohmw1AfBZwC7gM4QhFHNKidsM9LK538EZ3
sFx0zi7weMvZ3et/oV20U/wx52Dg5/165goDXBC3bEZ72w0cFF058Gtb1AQkFTBRVLgGKQmp9y/t
xK6P0EBxlqtPeBJVcmOuMeMLYDcJoCQAbbDV09EdaEFuftS8s7AEjJ21C1kdgXL05pt9avMif6p1
hKGi3ch/yPbzbjSJKy8HRqYP6K41iQNUhnupwWLq5PYA7sXPANo86my2Y1+mQEV8zBbFiOp5LgWN
SZApaguH7OIWdlsRXNuIPa4QiFSnUUpX5L7oqTd7yckjl5dS3QQXo0qPx6WgW3be55focZs0dfh/
JgiFYdo7pyO1ZSp1RCGsjCxYi9AUaNQKLDVmblybsXtwhQO1g+/lGAwyeRouPoZJJUPvh5zZUOUx
3XU3/MAwzJjILqVQR79Ig3yahkLn1clcV9JaO9q/kMRsBG8uDnTrJVPCn1hz8ZOk9zKfruSHRcBy
+hMAONZM9IF6urdSPgowvwfBnNCqiB/OTmpCwVeMpmFsetQDAXHrhrIdZZ+xEpI9vabKe41CDSGJ
3CNbdch06z3IOPkq5C/B6yieXZaY+Fco7awYYTYHBA264wNN5UxVZx0fvqGd69FS75a2vby1gTTq
16VODDMfeQeIK5sLhM4u6MVM7+l2BfvpXW8IC03VoBRiRmhDcB+Gd/nUmV0ZCMZTddDDLbHxhe0M
5ztMEhFJ32tp83QDMuLovG7wSweuFE+H3BNKRmocpuu531dGxonHH/jVkgIeAdHop/Y2VAF+JHp1
w+KzW1usQc8OOVkxSCWyz9TGv66X3pOfKolc4m9InyOYMDT3kRA8USui6ztaAMJVijnGIVS5wQ+e
wvLsx1foqu4hDAQyF8yvQfDwQQbXnv0B2Ya0l2tkTc/NAoMrzWBDMeI+oY+lKr5r59VUWJEN++rl
2Tv6NXQJjsWUVO32BzSdz7+dsqCrCFiT+1L6UGIw0BEDxePBT2M/muTRQlJPCFAoZdmSFQOXFgA5
QPbjfN47dBxXN6w90g5P4KPV3RBEKZnLvqhy/dfsrA8/jqco8d9f4d4b4TzXRq1j8IdoTyj7P427
S/gCLqq9rxcA94AtNmM+5JqrMPybQyr28u1+8G7vAJidF4FujQcGiS12ha6U4yLxo+I1wgator0x
JNTxucOIdvhnmivZZfCPhiLC7AxZ5QAitJSpU4Gra4xtpyeZll8mDrID9wlVmOUjm3UHAYCDph6G
7MxUHU33lsyQu0uiEk/13LkWgL27uEGQRcmL7cAc6+9DmGXW3zTWXX9pY8RSXQXI2Rep98VLKryg
+bbLM/hjp3mGM7fZjw2Lf2atspawNQqzMA1aaavIUhOz50f8n97PCWpVmQxvbuw8z1oI/4UrSoUM
pceIEyOvCjXQSHSWGZBllM9Osce2CHdjlafdp+TGRw9PXo3aRtR+hvj+UTpJB2nLlunrSY9BgrCH
HQBLpX/y41Xvbmp9crv+rudntdvukB+kJ7reMOCPcub6ZMaHYF9XYvUOfrniOnYkCVPWcBULokbT
ABaMtS+dDpxT4+HjOCsrFFwKAihU/ryC584ZQbk3T0HinyKVUK33mHC2dsc46y6dnX8MYX0YCqqZ
q26f5h9FpyJpiXy3w092aLkRREvjMlu0XDvp1BPBmtZJ/8J7Z2lRsBlrz4xhs6LcWoJX4S2HTQpd
Jvt5+G1aG5L2wXUFWNvQHQUDKOoE6HE+wVcuS5fIgBd9XQMEClTAXtmKBIy8I2FBFKj2sAU0oX7w
S51sBLRWMFjO0PWmOvBqblWfmJKZVX7Wg8i/0CMZEC0fKHmYpn+xofT+xVGXmLOpQH3ptq5iwLEp
2AJr0lrEchJHdu82xKIPypaZZVf0Mf2oLIEv8AUC87lQw8FFF8eg/8y80v/+csOlYpFmIhrmIARz
riuk4ygpW0qQ/aAf93P1+TP8p5YXPBe6jDkvuzjswgaURcWAuu0C7lGGZ6VKczPB0kS3feWVBV4Y
nWi+9bt+KXIg+d5A3LSEI3VaysT79Hs7yktyteNUiRs3FONcc/IF7WOYuX+GQI/MGdJCmE/XULY+
ewi+HI6lSWnvadcNWfJtyfTZN0woQl/HJzibctEpuAia9EmHETu9DiiZTAyawYFxEg9zMDJM7K74
3pvAzvx8pyjEfBNo3mkK4JC+pEs12WqC4G7Y9kG1QF47YXmgCDCtp358FnWdGhn+Kz57Xw/dODAG
8FlnngHUlJPRrLvqmRWDScgYk5iE9hhkU5L4lXyb4awwkRwpgvyn26axnrqOnd5ynQZlFFACgqTr
B92PNREJQZSbt1xaY5ftwxh4gEBj4OG6duFuhZNofMSJu5Zeu65OC+EuftyTOLy1LUz4lgnEQmOw
cuFv/fL/DTZohDNhlSsKNos8D5Y3mKYRPTwxPV+80gQUmab0CKYAZw0Jti6JAbrl25Mm0H8WR9Ev
pZnUhuIwXppxYfgPDYHBsbCodBoEfrEfm0ZTkLNDHFdxqpYjZOhJQfcYHInXmlMuub3fjZnKKlVV
RstWXTJYyTiJzXfd10bzXMPaISB0ZMKVJPgsHFHY5VTREoqAhFnaWv3jVpL05DkdGZ7aFlqbUmVH
kSdPN5YzLAMWHRdboGVVbawTwSrlEneQ9CgKLRKSWoq+PBNrLX70MoZCbGmlElgD/AbYD7qmJ6w6
hL9TvBhWhMAJJEmpp9IWXV9Mc5q4wOO9Fag8uPbn/UWzaxs+BaQ+N9F6NU8oP0+QsAA6/fmRgy8m
V4Xv9Rag5NjRd7FQSG17JhZGyLIrrH5Hci8UxOeWiS3hCt6dDYI07i0RAcwfM7KVvz2SIIy+pkQ3
UDQWRg2Q+e4O23QgenDtwsYvjg+ZJTkcUefZjpKGBXXDLnsby9IcfHXLl8oAZhFVEUTeTffmstGk
SpGt5yyTQQgmnzsUtXSNFsaLVUqBpQ+a9sEQq0bSBUwGXhnmrTLNBVwg3Iy5zxsqiEJROHAYkV9n
FmeEkux8m0CLs2NrUu3dTYqa7hz3AdV3w/owHyGUGiPrYqWFUMQt2zyWjyXEj8FNaffYCZOfPWvs
uK9kBBhonzpGCSYG8B4pxRNIOq1/qaeT8F7dQ7HDjrla4wjOpBVUGuad/k2mxOsAUBwusYZeRjPg
7ZJRymkE5ADiGB85QMFasE8v0G0YZI822BkCm56IP6uF2FqNBNjBGO+UIKc1rBu2pLPjHnLusVTE
U/if52D7gojWbMrekukA1Xm1qLFHhRLA2mgdPzkGYy2+mwY24fp+g7AmTUL8IZCJDm3JXnAZ9Osm
HM0+URzwKu7FvNlxcRtLW4jeeoYay+uu2tCYL2X0k+sTLIMfqwWw5FunRUK1+lD89BgfuhZe+k/U
zbMQX5XbkLuma4MR7YY7e0j7wfJK+O65UbI+JMbojrIhHp9zuRE7vnJECVBVQmt1nk9fJQmKgf+l
4Qvehmtn3om1cTRyXQvkBvXwsl04eHIC3w6WWxRFOW/YfDPUnT6ORschJRjNH539smSVQC7njjcP
Frb9w/REucDWsAkVUcSkLwezqs7LSSv08UQvd0puRxIv841rjsyfm5U3NrQ+hZh9rLBQu+KBvfq9
NUShwdfONreLgDRm/Zvx2RLSDACpMWnI7/DXxFOJFdpuZ3/YvokS41mRwkvMvaEZEW6cdwsUcy2i
61qjjq8D5Q6VCcuuZJ2alTzMMJaVAp/Ic5L5G8hG1C4r1WX4gLtoW0DrbNSTQBNThCy1jld9NjVF
K4cqVY6C8f0GfaD7hJskGSh5QwdeNs/vdxtDjXkxaokG7Azqub78wiPUdhVkrV0+c0xyiizY7hEn
+UPk3zep+MopCVlReJt4Zhlothl3ZuJL52o6Z+5T5/q9MPBjtYyOF1kjKgcTvlY5ppU0b/Wuw9v5
xZq97wYG1MccPfbTuIsvvLYM4atDFVAw/E+t9urfooTD/0eDE72fiDoJ7MkjZ7X5NUh07Y1BJEoa
xI72Z25EgxEltYaIdLEdScZTvU+j+xr8wq5tje7D8kYjYuRigqyqlY80Lta7abRyY585HX0SyEU7
Zqw/xZ7V0yVib4zgHZbvDpoRu355UpDs2UV5s9TBGwH3TCkvEK+TTHKCcuMR+C9iedpfW1XajvGC
2XLLEcwAiSe9hbP8UogHI/m7z+D0irTWfwchMXu2UsIFjqgkx+4qvgORSOZCcjIuHAPRSPtq4h5y
5DTlpf52ucB5iQPqZ7TKAyxM3tSmV9WP8SfVxhZBrl+T6k/7PWtQdwmBfzLQwxNSBrceX6s2JRQj
AXfm0Q6vDG4IGsIZGw6xJGL7u+qGYhGI8Ol8CNZAfzBA4cQ0JgEULaV6WJMs4thTZZDYHDHdt2YJ
g8yAEilypyQ1gscwV00c6zOgrn6RsC0fYQUKcQW5Bmzpj06N88vmFhLJnJBAFvwnsmsY5tcJWH7A
MgvGfOLWeAlYsvUDSU+NejPKR2NcJw6V9u57f1Z+ccl0MB/p4EMs4llIhpR5r3fKuVgV1qTHn8FT
I+oRkG8ljbXwZuuOgRvt+0LJuMtDYbqwmX485Xd7pJOwkl0WDtHEieomN5R/S0PJbhhWT/jvfh11
Pc87d6LLobmKm1PINak1dKKTfu9xFHNNwuWSHtmKZiTbS8G00FBC97DADRtM80g6Lhs4y8eOV1PB
7amB53bg2QmOJIRHHQ4xrAKtfVIJD2GuQaawGkiFh0v9UNu95Ea0xGyxuGAjk25Vip603rV956Rz
2M7gu3wEyhz8GYWKYWfTYM4C0NDi/29ixe6xDjEPRkXUqhyYmksNeofvJ+n1813DAucQRfjmeo5F
txgQXWjrZ6DAQ+7AHeatlSkmFPOYbBG/bjGVuSZmLW84RB6ucOEecZlQ4XA9L1d4yCTpjjO+CX29
mEm0wVe3NefR37JQ4i9DrWk50SRSZrw7N/ef/zDNjmbM/J0RWSjP8ZZ9tDfKI2K+g74ZXt2At4gp
b4bUc+0lj4w0BUw8Rf/BjqAG7TuJKgn5Dv30HIq3sCMUTyxtPouEG5iTaNdXhCB8nB0zNWHP4Fx7
ArXKphxhLZ+AJbbFHpeI8ABWSreLafBM45owMDkWS46WBhNatnFtg1RLkygP8kk9lVfUCyzmB6ws
lM0AiC80Id+UpAXtaTc87R4nyEC71At1wF+aArvIxk2675jv18+a2eJHCZmeWkdec8Lk4Vcr6QJ/
VaLophYe6glrRiYLgB1SVtetR8W6dwy7A9ygc1tDLxHJuHF75LACt2A4PWrbeHEuo/tzvMVIzXfZ
HDDirWQLNJDoYj8GL0QAKTdkwDq1dJw7E/PlVOR5ivch9pI5tnEaG1elVPQegZDrLjQztj3x9m3U
rRcyHEQq7H+O3MTgm160U8dCkBgWnV0Paj8/rY7i9CPYuatlBlEHjc+Yx0blWZEsuEbMYN2RDf/e
1jNsM/IeBN3RuIMkrZlxFkOvYqY4WhamDF3Zfu07l4szYKGbq9vRe+haejeQJJe6EJbpie5FEjfr
skVisZ9C0tDzca53VrfXRo4NyfyHFVWhAQJjJgaqkj7jEmsV/lH6izmFqWvTNRKQCD/397nwUimU
+uEouhXPZP08GnxCJvu3lmAJukdzTpWi/09rQ2Z+XXgZWtx2OSeylR26hFV1PyUqav8ZWCXJV1il
QdG2/97gmmE9Lt0BSrQRgOICFWCppf3BYC+8cCWq/U/lwfuT6I2IwHEr4oqfO8NG8FhBsQYapK1j
cccVIAfjNYjgAdEYpmt20ow62iV1Vi0FqNxSDw3/ttUuV56MoiBj4Xc6Mve92yJ5U2UAVFQPNt5W
MsHlfLTcwmvBdHh1JEUyOLir9BY9dRh+ZlM7L7u7dEBUMxs/zUsnYZdf/U95una6MhDnorsmV7V+
ANwbX7BgVaxEpvsF7w99usQY9+Vgxrk5rQ3ZXgBtt78u4rfTJVxHOFegNVrNenM/M/tCFArkpuwz
1hJEtCwICXpgIJEy1+jvsoNw3qE5L5KFkpcDWdWYZnMi+2X8azgbDR1g/3/ca21iW2JKfJWN2Nfg
07poAKOrMAGrubqSYYGApJb8uOimJdOLAijenjB/AgHhiPNWHdAu+l419Cg4eTBcTqdSEnZd209d
usD2h2vwxkmvYY7pPd+n4Mt9acULztUMHDhnYlnYBzDIc3e6DKejPi05duM2bksOXXPzU2sgE5BQ
pp0cqvIWD4Vce/pMbfTq+HOn6EniFbYi87q5/4ELnxFU79pU7EwfzvdLh5nlxS5Gcm/3ZvUCk7jL
IDGj6/5n9VJizQYL6PJNBzRJ7D/X7aLHGLzuYWsfGUY/PWiz99AuYwHpepCsaPtCSUW7Grt84Kul
VNFZXYEL5rIzPShPFLCsmPGWuNMaFUOAh5ZHwmAKiFWrd4VyUh9Nj5rpmYH2mjb7xGvtFTiOG1h5
Vgt9gEtmpEBPOdjikzmK1qqQ9tJxVMva/eQdaQR2+ptwfdivE6muxopqGtQGVYiLqojfdRFj5cYW
7+g8vf2k/BgnX8c90D60mVpHIURmYS5Mcsl15kUAIA5FBEs9xpRl451W7kaK3n+xp6TTr4O3mHtM
i01ewow5KUTBPVnsvr0joBxltqN79lDFf3TNLjGf97dpbEV4nTduQkQ43ubzMsUF9bXMeQt8JFOX
PKsQk2FQTBl2LaMorqEI+XS7Ii0+/LdDG8HcAHO2NzF+hWYRwMaqORYc17DSQy7O2pN0GyIvTr+1
0mRVvaQcWIFMel6ye1CQqXGrycInkz/K6sr/Fh3cxLuUtN5RYEnSSO9gQa7XNZs1oy3h9ALB9t3K
4OUQDMdVf28dQ92gFe+M80MgSssVyxCprXII6dwsqpXnSIG2uAMJPTO0WJgqcauLnY7LlQtxCx6E
69knHWB92b0Qvogqy7LP5V0NcTbFA8aZe4JNVXt9XiVxYDCkGhLCCojP9bx/9xgEciPEfrCYacrp
Grq0S6nKiATn4onQjjErOUpaBdVIKDQTR7ND36Hp/xsJ02e2k90yxzEXEVsyfycWlagWhNR4z66q
YWMnHRN9E1vfRp2HC9wKee/XInp/OHczlt6rn2Rrr5aLGKOdgSd3wFoH/+n2gtvoNExt/wxCN6o+
1WgcxzMCP+1FUKLECsKXcftjRds7W0doD/6U/2sVkTDQ6/Kp81RrIx9LFu1s/7xm0XsT33QPLXIt
DMwyQC3pKahfZoA3Pe9REYSpf4KdZaM7OziirAQuJvJO6Xx5IqGyf229H6EzglRqt7ltQGZLX0aI
9h4zDtg61I56zyYlo4CtxDoaycp0cxDwlglFhnxN89Dmv/1UzuX67UBfOQcLUCZXPy61P0sMEY05
wD2j2cA0XRsxjYBvveowNE1KBrtI+Lr9LnqQzFD15864uIUUEJOYfRhvIOOujlmHKsfbYjLi1iel
Uxv5c1RyqQasvB5hfbZRT+5Dcgws4JsrWho4WGHGjhKbXIwKh2tT8Lr6KF7V9qGw40ES1WyAakPh
C4myU9CcYO3s7E2B3gecZSsk/tnSbqaOqcEbgUfLVV+0ot3P6GePampj1bXnuizsnA09jCdnARsI
1fKk3NEnWqd41zM6naNvXzBrFBUiBKzz8BG4O6JC/bwehrhW/k6DVwQKxYKZmQzHLZsts+tE1vWw
aNXPvvRrVxTqWCe9Q8Oxnx06CKeQvXoL+XTIP7kmBA97L6vjvBVvp844uMmTuIrwnbro62mmnLvn
8rHdgAZB/bb0D9IRolDXT1K6YG/v3nbzC5VN1Xgmj0MVoruhWEcIyENsgTp19Q1ktfqZWOqS1hSi
yOsJaLocvFJ3AbseYuIQHcHvnT2M/T6FGpgr7UwNVbysbQ6BdEp2FSy3Ht/liIw1VkMNzQBhULgG
w5Y+HqLDE167SVHi+EhCZWJKRacL8A5aq/9lCJJjOJ58PcmVUcX5bMnjbgF5SR7OSkrTAy7sTH3z
jzS+6FOD1jnZ2lDI1vJk3jzULbPnmsvQ77JVYnDqcaK37BSQtkta0YEXryC6OF0K19vqan6VdMEO
d+7lgHQyZLa5C4z1dM7ByP8eclzc4tRPqY5uf65ZAe5qvB7XSmt1jNjSJkYEs3/fOvjraPzbmtJt
rkarJkGnhar6Kv7PwkDwVryF0UCBTd5W1Cs/CHtRfXmkHT7+4lzP6wb0RiZtvjv204fewCSnXqA2
vkqQiUOpO8HUUfTzum41yIb/ExV/97nMt/s6BOP4WdnSDXcfCBZUv8qzeASxEtVa5KkFUZMGGI+T
fo8gwWNHuwK0ospYClUqc9sejyWryP6cD8dTF+Fcb+VXBjGp0ov9DSzt1P5ix4QX+xSlZxLkl76v
6+ng6xo6CkpKGXmG1T5eu0nYIfrg2EzIytZP3C9v7DQ+zp6JjdRQ3fBk3QZdn6sCB0ohUL5JLZTL
OsrUsrZQhOHul1LUnjeLBJZUnjHkQ0cvraPwkgPt0vpInIuFKFvMCDRMq09Gt/C1rYKNydRtMF4M
Qj+9bxtt3VD/pva/NLiJc7k3DgMMEFZ6ZZJMXpd5KnuoX7ylMisys1qSMFqjG5KVQkrdLwvfp0Su
g6S9mVWGdNq3QCc2PZZ7a68JQJSxZlbcFi9jlGZdsZ5N9ELUJhqEbxwy+phHwVMN1BpLSQQoyWuT
81CAZ3470PH5GBHLzl/vQhZou2eftsyD8H3WQcAquK/4v7DGtzsz6iSsq9gCq4V111tjW5sVOuT8
D8WgRh/zXENsb22pQOqWHWGDkE/7cniTol3BXjMg1zQbbU7fZviB/K1aZm3UBTh3GirgD/M2a+ju
JqWi02YnIRhJbPGsLG0+WvXf125NvEtFd9DRe0S1yrc7KiOvifTd4z6+Gv8eOeg9DJ1T8sBRuZY8
3Aq0JoF2X4VwVAvB+3kz/3NLu8JYxQfjaV8iqShCzNJkU1jX2w5UDnhzsZ3pddahal3QZds2Scmw
d+GlRPUdVrAdpDwkVIHpI0510YMDu7yoSq98Rshkt4Yiqm+f+blUapz1P/Ui1jkInpKxOcBRJtUe
34Pl2xkqRGVJy9YAonkJ25IGLfyrRtcw7tTH5clBAVRiXR2KqRSIz9NLmuK72WW5tkEaqFYFBaAJ
UhpuUm4r6I1v/PojxhrkjSfwTPpZficLDpP6mvMNwV38+fTtC3TPNLNizxAC5aOKxKPje/4B5d/1
Pp2MDR3tjwIzTeTdSGptskVhHSvISPsN3XDNzWLVlzWpEntqxR4is1BYG9OmQhXSiEUIgcqX/MQj
JWJoO3GfxXhNZgdAnsMItw9h2zQWmv+ezwnLj4OvknxNvLil4NMIFTGTF0g16hSPl7AUFim3yIxp
0dY6tCUjHuryi6cmCPJ10aR2xc/y889Xe2kX1ZjARa9HbYN/cH8ZLAGkflzeonv8b6euCZqYNcWz
6NZVBWCJj1MM2cIZgd+AuKR/0Tgv1/+5ak6F51scXcVk+gwxkFuSptMHYAak65tGMsiYhaftLKkE
+FZLmM9dkPkyomd6GJh5jq3sTzkp64R1AxgWEJJd3zpwWo7JPj+klF6yQsCQJXhN0qiy7ndFfi0f
jrFRM93H2nQX0PztLYtuWpF+iiKrUmcBrlNpv3SjKtFnt1bVWrBoeGUloE8yVA10BI22dlf/3PfP
QRG0qSGgSbNX/+gd4y3bRMwqJjZTWFlZ72Qm4CxN7pqvelMzgyma2ZEhddg6SQE1PqTuZhTytJ09
qbLU9McnI/LrGi/wi11AnJjOte/yJn9Mwt1KESUdMoD6t+iVaBosxEZSgB2dLwAhAmCYf1V7Crpu
yperRRhdtc2E4WjE8SkZY9Mfh2dmZ3ePsAK+TBglrP4+sMBC+i73f0CWgvJllrrX3JzZ/WucfsJQ
6hVesSaakPirXMY8Hx6ceyQS1KWrtNAZpxgsjJ4BpFNqDRaKOqU5RzP9y73tiEuI4zuqDy8qDD4f
keMWei2DxjEmCxNfSYsY/RDAOPJmSRRThjCXdhsGp7vvfEP8Yn66UCmf94y2hlDlE7Ym/Rxhrco2
Fo5uC/yfmDkMeV+16pzPDuT9+vmdP2tBfWJoy289z+7ROHCd32NxN4K8tpBR+8U//wQfl4ZjDS0H
WQGnoy7CwgnvEVtZf+dL/2TOUfe5BcbbaXvXO4kUK5lpCr/CdMbed+/bxnDfPrKkb4VLg69XdY74
RGvpTu/zFddzV+FBdN93pQSCyfh7NDhhS2hlGOLZaZ93TbcnnoHR1J2PRzItu+MCvXKKEs4j1+bS
lVY01jqo1FHenjz9Yrl1Hsw4U/OGAw2l8QjjmBXPgeQq3vGNrrw/gRPnGtFEvWns2YHC8UU64h3l
UssOCPZ3LrYJwJknwKvFz/8UA20GTl+fw86MNC431H9N+pDbot29ZPLfR2uh0x+uNXJfQtuktCuM
yILp5kwmaWji5zQGa02X5PkMvcB9d8B7vEMYcs1c2RBAJRRBwyZFiJPmSIU0fNuOwTXWpJ0/LZqV
VC3H4kX1Vqsqe47i+WTt5bRL8lXB/Koe0HjvzpikRNJZtKHSYftVKzQV9lMP+xQoOcUw9wGyspoX
seg+T+DCo6cpQMqmy+nViK5s3qqVZpkXnYbSU1nZ5lj3kO8iZlGIXPTpKpPeub1NUBzXEPeGVqPQ
j8uksOMVP0smUHN1Fs4lwdh6/AD3tfPR4/e+Fr5CS+jHX1GlcrPN6UHYYut986CmYD+N0otBK2m2
jGmJ0ao2o2hikEKdz5BIcitLbb2Zl5g1dolNNSdWmGNj5fQwvSDNe+aX4Cjlw23OnA1jCtUXzzz/
Q6dsbUEJ/z4gw46+1FyjAaN531M+7uQXA3G/1kNlwj0SPzc+b6zmGR+wVCiS4KCeBsmnnojmEVYd
z1aeaPwRyzQz1HaS+YMrL3n9aJFq/2F9qynEd2QaatGL55m8v+1Czfd0pWHoMrbhIss2pULuP7j+
I8VhXJgyxnyLZZ851Bx5A3QMIKxN06egs/P6z2H3OSu1GqfLet3MNXqD44EgMhe2cttVywtmWNos
MNcMZeTj3h54bfPc8wMIZJNavUIy5CZb9I6Syeq1EuPfl+JZG2jCitgs5Sx1otz1IOglPV4kSyVw
0ddEsqX3oYI+yX9xWaNARnLJ/PoVwGrQ/mCWGC8KJOSfljN9ncTxNKlJ3RTgWfVpOjcY9BRlo9mQ
kI1g/i17HIPIseEW4nhBzLw1zdV2GcioHfIBwbUmQqn4tHbTPo3mE1nswcmkfLaeBV6PQLxnNxd8
joeA1r6sm5IV0czdIBUO2wt8RNQqN/94uFwLVEvq6fB6lq6RJPKpa/cRk2qpo8zC4UiLpcBO4RIe
GK2YRHvrcgCBZppjUBrlDVLt2yYPmDQMETNM+7Xd0YOYk3sRoAJOk12/N+3C7p0uMNcyvd3W4Z/N
5PiGbH7raiPyucnfrnSoUVFmwFeLnb3ecLxlg+Am9OvBw2cfBLb0WH74jxqsGCgOUKR7BKX8uhmf
IDFHJjgN2jhbHrfa4P1BrrH2CoWXI4VyFvxOYsT+QHsrU7DkyN/N3Vu6Vj6eNyZUgWSnOBOBjOlh
gwdvdlBEHevEjM2YlVJDBD8moa/QkkyDl1ROz9HKyZqdOWtmsk/6Ip2IyklZS322w7KJ97XQA12K
wNA77M4mY1Ne6qRkWaW0/fu7+jUmI20pFqNchf4KenYRgxvmDFQJPBorztG48EDFkb3qqqIh34WI
YRPrFAhj/GXgWjgie3Vn3OVze+R46Ra6A+aQBl4Sj6NF9YRR3iCzVDsZsV07AjLfHq3t5yDMGR6C
KPNWhNCPUOZW2x0FCbrxjymUSCFPKL0dAAM3/frbT3BfvLZLNMfd+FmiQ6FWLLiz/1FgXGQak+Zw
HHtapqYSPQYTx8JS/NBxXWFPRdlarzCtmXJtI42ovLA+EmhrdfNHvGBPvuHaDbj+TCDaPNQdRsvg
5bjIRyAAgANCklzmpOWHa4jI2CjeBu8TfqE1YP8FoLFLjW+DTPF2OUTWW6odnneBlE2ac0YvItN4
ZmgiuvdWBIka9VZdbAUHIUboVAQFsIxKu1GJar2SGdU2B4pR0KfapFjNMrdyk4hYuX0Bamxz3vNO
Q09DxidCuAyJu++fy2Bl0RZDj94KqX3trCW3SkoBJx91OwEtGiUX0mAwMAd4tMDz760po5XV0qMw
WJ7nkDRay/lA4KssBraWR0+2HDYP3s+E9nyzx6w0ZNZm77J0wOdO7AJOGEtpuwlT1+aaYbFc2ClJ
nb48cwGMWeZCAb0Xt++5JXyHK1z984jjh6d4uebrJgcvEc4yhpilxAvb40K4IzNHQPW05dLj6uyO
vxji5Umq9SYv4s0vjJEYKRkyu1HPWEH5rXKiAjXEgZKFZ5Hv+iChx8vjR+KFH9zyY1FLy7Srqd7s
cQ0FadM9Wdj3AEubAAT53gWb5LGXNoZlkVSzKq4XPX2mS8zaKM5VzYVxm5ugwxNtx6Gmlm5tsRgV
LsTQZwnJ3Lckn7CJLWrjk+KqX3+C6fKnibGuG5vP3vauZ7leopMFPxLwbXIsjp1C+nYH8Y1FMNHu
teOYszTPee60NhQDgsGi/ZghV8PWoO+OWWPtWg6hNUfsLPp14usGYCm8fJOtNzIjmVReRJ8rrNTW
yYcquVYJjST+Z4ZTnM/uy5hxQgjE0N8rflKTnp1Rz7y5q2YBkFInKl9yYSuQg+4gu/jUuskg/8eT
K7STHH/Ljlv42DkVoNbFZf1GowgbzbNCxlW35m3KG1H3Kky/RycMwjhGzKUWLMuCBMM1Zk6NAYBU
ybuwrdJP5L+ejWojdSpNi3ryRcIeY/U8XZwVNjo2mlop5mPUybBAuGUqsFQnNAIaODLTQ/gCEjP+
Tevx62St8v/8a/v6nqisNdFe1VGXzExpnOAowQllfwhNSMrEtwU/X6dAHCq1ALzVJ+q3NE/QMoCk
xcW5JDUfk/IVLOBCjlcolkCpaMNdFuW/3pEPdKjiEjM73IN/amqi+yQSUWwSuxe0EH52FRuk3tz6
31gak79jrIBwjyWQo9Ey9gOBOIxFLRjBuV9WKNySmhu6ARx2VUUo1QaVY+Gb8AWhE3C9OqunWUQW
JVNK8Cmh+XxD9u1vCoHwHdYyw2vjxfiGUaxpX6LWxO5Mwi4jaENUxwMqpaGkB5ArBpT3+EwM4qNo
gaISKcxnbVS4kUtz0g6YBJTW739BlkOxlfUN/pa/NOwCHTnbueGyaas+e/Lgo8CxXtsx2xg4vYH4
TtYO0hrbjfCg8pqMMaZOtHtl1a91yA27EtTehbETTEM3g+A3g204nN6+1lGJ8hZpWBnuoe5ZL57q
KkVnqNAAdmrYZ+xoPz3QBqlE+Z90Aphnxc/LYSRpjywoBpJQfLuM9arjmHdH+FWZmJy+SCNCU2U2
JC7rFlyNLViSqWcPoWNpURH51ifT6acmKW77Q0l6fsB7DMM3LLgvOVNT416zMWiCk1E3jyasi4jV
Di1OuAkkeHCvpOz7bttZMpXAFMzBWta+EwtXOzS2/HNxt8Rscwodne+Y/HuZkM+PfQe9EWMw7Lc8
TmACUteQwkTZdn3G0zkpDHLo2DTnhxyu9/ywKHCRuzZqSJgl24VwEEk2S7HtuPfjboVHWpeHDhpR
p5LAfaWuIEqlcGFK3gKqUrdZ6r72Ezt2Arzo+y7g6TP1dJIZ7K90Oy/8c+BL6PciXA2ArZMvBW0G
S74qcHLSgVg6BInV7nEUS4YOEzXdSmxCr0rEYRBv2VV8bz+u4sOQInMAAc+r4bMsKCay+5XGNwMT
wpMa8c/cxgKmaG5oY/mlZTQMMTn/XZjmVv9+784XSeFhJOFWpN5sqV+tnzlgGZM3gV8zkKpCIBpm
AtveKYXjvOH3NAQiyO8n3anUbxdfSLkIn+S9En2DSclEMqoPYl7hPW49XI8Z3EIbzpCGInrAVOge
H58aDq887sq4i8O1jaQ6WFLsNaAz5ksNrg2QKCVl5DNLhsVL8nHqCHbRQ3SeOQajm2CvEez0hHaT
6vntl3UdWHawvjklipGjYUyVPJ9Vqf5/UYvAVY85ByrctdeAXakMvFKZSalAwVD1ruYk8P/fv5KW
Hw79DX8KKHYmw+Au9FENytuYgBk8LTQNHYtewpdIKPczBbFkGkc8Ts0PTlvTJtP3f2GVkynf3RYN
f5jWoUN03sAeIzApm5KnS+drnHF6bj4JsfMqDxuobYm4haeaAV1LwPfrYitMVrUQjKeYUQLwkYUU
pjzyZQBWmImovEuhYzlBGF+sPxHXotaoWs8wZJjwhIoOkFKdp9vCDA+IZHspM/0y/kyQ5L5DrEzd
ARU8YHbPYXoDuOi1Z1Wa5bF5y+8J6Tiy7MgdbO08clJoyXrHmBg07UOUuw7OGSxEBzg2pzelu62u
lXJRMIObtCw8Ury8McOTU7KMvvZ6LZlkaA1FLigtayD2n4ppSlqZqGDPQC6H3JR9/mgwVQmZoYzT
Vo5bEwDW/ofpWb8zCXfBU4PXq3hT3MXiRJvprumCcqgyvA9E+7AUYI/hoQgM+xhpAonGYOfd18pI
npZJonoUgZ2n0l3I+60TnRZyoF7tvoTRStCpWbk98n5B8Pd4uMVE4DbLMhoKajYcJByTs6dTRBBB
rENnzmRknRF784ME8Ld2dA1cpWMLFadHHu1MhEm5tk+zzNSp5tPLsezgiUvxpGj4AfpMujkNgt3X
Z+6W0MfkqExL+KDolT7+47L0Ydjq2NIvR1gtyNbaA35ZAEyJy1on8miCkb7EsAFOcYDUA3EzsfmX
p+MF9plWnUXK9oMEXPQKo9nx9qA2i31LVF9+yHqRg+roJOf78OZmVEvfNtBb2ThrVFJsQQ6Ea6UX
zt67DY7HjsGzIK8hd2adNgxMDeV6Xoolxcah/W3AV+O6nHHYG0DP5v9eOhnhC+VplFc4NK+IiDO2
W51cBWlxhoz8Cl17ixRt58CSFbQcZaqt3ihLyBmrwXlidhpSO+O66fbOo8xjsLBmWgZWZaflFxXQ
Na6DaEz5F6h/XgLvoeB62Ws8TH8RrPEDiM2vXS1ZutfN0EjHZ+9cbscpfUSUqfZ9P8v3m4O0Hd5F
tyskePE8jMabTmwt3sOBoJPKb0aNglC7Bged1ZoRJRrPYtYwNCNRJPBd1IHX3kl3w0yLT1Q3OssJ
kMSq6xRKZs3GXeV86/LH20J36k8likypcEeYh2THE30d+pXW0J+CLWn+5ag/kYQRx6BXANP4YmmE
dGNQHIjGKpsV08arHaPSBaDrHTDMRo2Yq3H+oPcXnJ0PbqQgUeKFzOvp6rv2Hq8d1z9sIjkfgvhS
zWE25KRAO4wAizA8TSi/YZTl50e8e6GzsvEljX35SuR2SiBKdc4UNPluH9huKvc70YXzu0wiiWNd
Gj8NKYZ1clwQUiJyMgWIrG3OXosJaGJk3iSLdEzNVnMZ9R0+ovqTreTRrUamn0h/keei+5ae1x+R
RzQrLrIBBhrivBMWtToqqAyAcECt2yXqs2fZ2fL2VrtNcVBzqfuwiMDLTrVDelEEpmJ5SFmkliGK
aRHipCumOVm4K5tAPlYOuwcDdwrtfMzRMAgMxn8pQQSF18d2fddievCpTwG40NIo3WL25DnPaU+R
3KNpfXUUEbTcVzN/NqE6tJHSq/Gtyu7aNAZ/QIXfwIzLEguPpn4hVqFXF4gUfRJdoqj8If7Of+Ye
Yc8zIXBgM9iNe21297AyNTls0GDeXpKj4cYuRZDWbkvT19ZQ7huS/nP4RCGVT6ZzgwDP569DNGVW
p3eL1qjKyuryxiiDbKFtHPeQFbi2eKQMzVYma2fpdbkxXTKkCqreMDzekyU7Ad3vmy2F02o/tRmh
bkzhJ1wTUaoTJu1r0/5cdYOwWQfiAOJatjlVPiguHM3dh+GcSXbvKcXrYSfaqBVwWmr7EAxXyTUf
nw/Nx0tLomKlv9hqvtqI3Zzca1AygKu1WuRGm1Ya7f4AP/Cq62wrYydJBGaGuPcgFSZ5ubGnyO2k
wm1AeumTbb7IGn1aN8y3pTokrWMteSJd1/MbYk5R1BObV5pkded8D6cKKly9NnP7lYhshoGkuTjJ
NgLaIn5HhXXRhgSLF1hX5Z8pOfM9rQ2D6HXN0z+Dv8LewKuUGdnx7i4UJVPlgsDZifJkHY3TnInE
ED8vMEDRQ3q5ewmmQDLCQH1grzkv4Hu54u6hogoSkS8petFE26vFMIM6aJy+r34E2+ZqPZU1gloc
f27GB7lSWu2dZ5AHuR2vq3jYrg8oSuOQXO/kCJMJTYDeWdUZ4+c90VKjLbU2nnQNXe8iB+1YKYf7
Wx8qkOm1kXsY8AX8uKfmcweRNuBydExYb14ZJ9lSBTCAayojzy+BP3zNS67WPiXMn+vdnKnNBAEJ
Fx9PtL3p6VkQqPdD8dvpLXxmVEREAhAR/sFSnm6hOT4vysCrJzI6lA/uP50UANpNqBUZxNQ/WQjB
USUnjeXQwX+upJTEDMaAiVwwjWMWzkKh2pk50ULjpPo+imfVVeKB6dFH9mM4Li9+HfnfP5Ama2PC
n/2uZRWxMFQNm5BrTNn32TioRIiSFyIqyx2i0+r29FyE2B0YYWIcsKeqToSD9tPZiOA/w6EuJotY
A+fWnL0BWzrTKmR+Al7p3tmOe0DUiQiLzY/yAWcKiVhNtxy1Td4o2ugdjur+YjiP95T7dVkKejQJ
yi6Tdq9o5wNW1aMVd4W0A745fQYf3OkiEEWUdMuQCa7MgT5BV3Kx3XGMYQMvrjK4GgNj3u5sqRmN
Ft2cId9o09E5wNVEiW7VHRaZ8BdJY2mK4GE074JKhRFG3BOIrJ7zphikT10lpfDqrWZzGQB0cIWb
i6uCJVfmTJeP78lGFAOXG+dGBlcaCZ+pRi1pJ2yeO/B7qcb4syJY+KeCc0u2AANTDv49IyPGW5X/
3sr5jQ4CUyEnEpRVe5RRIrNWxAUo5RaRunhraYcsAC7UFInX7URCMKRW6nEEgaePiZrxj0+guyu3
pfTTSMZ8OzJebLC5CWb+Mxok0MFRN1HSE/mStojjJr7XsAETmjC39dFFPWwrvY25qtOv+82k0NjL
G5LxaSmX1WHdzypZ8k9DrAnTw7skkm5BbQWgtjt8lKtMawLVi4bJQGT1PBF3LpMmL/hcznP+zt9W
o5hcAvYYS3cn+EJl1ZFrHcm48EP/PvNvrn5jZYUQLNL2hlkm+kf9QBa8f1DFAhw8HHedGAE9fwaz
dU8yfK5CfgPzsJoR0xC7QHdofc8kxI019bf8EEa1D8l5EOPhor+agbU1adBBtudMV0KS1yxZ0T1E
DauE4BNzrusEd4/3c318XwYqXEwASJIYllFGM78lwSmvSdgvOE3cLX0xalaAm2Mvo2Av7oh6HjqC
Muu9fz11XT2hT/huyRY6DMO/rqV19sIubqhU6NZF5Roq7nef4R23HtJsF4maAzGEdhY9NscYan9M
l5Fr8TEZp8O5vHJyss2yUZOo/Sz184T+gvkBDtNNUR5Sw7oB1sKmXEgslKSkR2nmocrsNJivFMNl
uURa66fEJKZdufrCDGEUbqtjC/kDXFlrS1XyTS//UnfIBr3hlxvdXKF3LPUqqAClR9be0Z+FoJqr
GdxbfpiKsCBBdoBVkaY/nN/tva1QL0EeO/6BU/ijtNvKTkhhoe/yn4+hijRcY9n8b+BSeOnZ73Pf
b1xAfw5Fn6JD6JJrRjtbmMTBasVtyUn1sjcNa+U8OgBMS8AAJQxKJUqVDGrp1ItfKv1oOd3m0hhj
KC+TIi/WAp9rn30WsVIDasiN0j/hsePQE34kfMjfv9Kq53Xz67O9qsFd6oWXHAK40e//V3X9qD7B
ISDuJApiz85CsHlfN/XWSkc+qT/DC72lAawtKadcnlaBWQSlMq1OzLfdy7FpBkdpTY72XyrQPI/g
qOIampOwrL72vmN+pZIW84yLV3xwOTSTdccq2B6o8eR6BkgUhyJ2J+YmExkZTeIie7gLiUyjbYgE
jLqWAv89NJxk7t6I/CJhI5xAh82Z0W4o/X/yUOdcgIRKgmq8KDgnPft1PmKHd9+yoT/t11X8WKCz
qEa7Dcf/OkI2fqBu7Jj6rQD1ZcVqSTjYDUWHNdBJif67X2tuNLu40qyeR3qrODxkkMTSKlcZAVHe
dqiLn4al4QfGg56m/Oc+UNFE09ac1V0qJshYr9vh+ymlPYC+35Q+U7jkZ6jMQ9Il+8dL7BRjzP7G
bn6SQy8/cn3lczjsv877wH+wqiyHiOIsnVXQDpYaGk21nYp64o1+7xdIgqbZnZ5dWM8GQH4iGNx8
jHYmzRi3pONccRfQzAeQyvbnlQ7772TFfHQSQ8+XncU9FuRsLkr5SeME/eXG3qDZiTAYVERN1QuC
a1c3zGxeb8+5C0gLnUV6KhuBbT0Xyif2MQrZYqU3S5qd5mAxXuJQ4u7h6RCY6ugSGVAZk8qicX6k
Kl6Elnu2y9E404rgflCDvH/VjZUYUaeb4C+Pxf2sd8E0j1bXYB46+TYm1LDvxrc+c/kqLy7UjZX/
EuSQ4hKrCwHhj/1sn25+y8Sns8PEFVNhPMwPrgVaJl/oHmESc/JqZq9sx+9ovqnAsbe7oCFTD9kJ
JXGY9se9w6Zaaa5tBq5hv2KI+vpbTaCmH4pDOfHRaSUOWK2yXBE8c5aaW+kDRS49kKe8H4a5hNGE
CLddcPp2KXH4jLXvhH+o9dtqwJ+Eia6PGQzgUeeRPZu9qhfPxEPY4+LPszbAK3onC2/NZMisvXCS
V+N5j4GcYaVyVzoVL86FqZlMb49h0fl7Bzk9bG/EnkCf6uUXXZll+ZLIeYA/d8LET4IdlIaktRKk
3eHXiBV2E76HNJpF/E874okW0zxbe27iUNEJ8XjGqAgxnD8TF3F/QbOvoWmzO2Y2gTgWpZD2Dn6E
zc1Nq5Ce66U9yZgOY1HE8szh4Jr1XNOZJ72PrcDVUwo6OMfyaIlfeAIiam2mnlsLm8wf952c8Vh7
ZmvhXrGKatn0/UOG5zhfLq447Xwo/ayqzVltVU5Fa/52QTetJ5hS0bZwefppoSA2cu+kSW6WSjkL
JaDHVwsgaXYcH3i1hKqcD2xgCarY7gOdsuAvW/7uK7AeuBUYjT6L2CbgcVlzAbYbcoAMKSj8F096
pk9jJIlNV3q0tRGwbuxBxV56Ul8hX0QFo9I9Bd/TjeFwpo9ThzrJtnxJQVM7BQ9czLW/YM3IUahB
nlHUEiyT0m9X5NhYVojkxCD4nUOeRzjxGgLLxuT4xoumLuj6BkHEKk7/GCVFFQX3l/vNVyQwIcK0
1n/L2bksGfLVvzftufFn3FMjQ3q7fN4f2e1zhAv0q2MtVMQzf6wecSI0iFN36RHi6XhC6EfI55kQ
BBp6t0mYbTopUjT1OmBUU/i3QKQ6f7cF3YYQ9F4iB1tXBo14mvhvle0zMe2f7aM8OmCR3SCZ4V2X
8Ke8EUGQS+BG0tmsXxdTUep3w0K3aqJxNekakXT4MzfJomzEAKBKswq5CJWCpqSE21R1xgtymSuf
P7m4ysXF82JDBfdZkoavT8mOPa1NgeGfM1q9A8KUacM+4PIEmBsl+06osq8lBvYKoP+xb9X3XlJ5
fReOkQTmMwfLMXeZ65oF/P1A7ZwqHCAOf+Ms8OZ8J22Et5Dyd9svRaf+Q/Vd8xAPyYPMcc7+C41i
0C2e5/yOJmTyU2WBEBnI2WfXi6XU2Dg1SsHfcDSEepvkwIJEqmNnbe5ywMLA1HkstYqXBkQbsZ/c
dXqTb0H4rtHIBq2FCeGYUmtZ4IHN7VtW4UX9vUP+Yw8qSAaUHsc/kkIZPx8n2bo9MDE5NA/mqfcZ
maMOvneKPEi3MR/k0Xxi2SHDBAAp6CzsDad4OwbhJrTqmAvLDqNm4yEnSvP7fwcY5RJ4goEUV0W3
BpAKg2wGze/QKyI1cIMOPGwmjNvX3a59cPb4AaONSHM5yOnoe7wi7vShUNxn5s4TzIiMxnuYtPCu
IG9Ljc6hHhNaLtN0/aXtdKY3S5T1A2f3+N8jeU8BfLdMIG+b0hYNEHbWW2PsH6+vE5oAgz1+q0yE
mrirs9bm1pJdG6sw8hQfqZQnjp99LhVSUvjHlZMMrmVW7oqmPkcqjBbNeBS5fWAwgp3VdgwX2dht
rkXujreDXSoo/DwujwVYp1+j8U/9sewuxet1HnBMByo7kMKqt+fwxKMzYQg4Ts//bitM5eqKxB49
rkr1ZKu/6Z7njo2MS8p5XYydxB4PVrw06nwYqQ0Xw3ohuSklux46YPBhhJ85UB0dR4d3WejBdHBt
blC6Z4ayZx8EhUTBmP+ZKsqZnTJqn2+bbaFRAvnNr9YyQZkK6+K6EoweZPAHXfppCt/Ue7Q3razl
4c74Ub+yWf5NuyigzGl+on/qXNd2hx/okx55PpFiAiHLrsvFzUL4xqsyzADLMxYoGyZ4lPs5f6gK
9R7sXS3gNfzSuPYM4mEiAGsreU3uqKL4YZqtPBaSwF5QuesvgcS1wOf2z5lQhIdL8uwudF6PRLTv
KzzgowafUUVbdzw7wWsXAI9sijYVUGHWcPzX5NgLrXmXGP+hWmqYYQjPsZfTmDtnuoU6ozuvC6ms
t/xmZbgGEF1pxYE6ypldZFSxYCEiPEqbX/2i1q6ihlkw+hCdZllBCHKsBrKWFo87le8zZhPPqpvz
WXqcqOhMiXRJsiNt95AHzbkm3bECE81J5EkodOA3QymRDkwWH9OVXj/F+2nnZS4IW8egJlkH6Tyl
RYMyyCOzo7hDHbjTuW/P3OmuCvH5h+/qRHgnhatS/y7Fj3ofLwQy9tq89p7uzVJZguSxISqaiq7w
rahNZfGNRzmB+l0/gl+i1ih5ljyVT47xjzbOM7+E4CgcoBS8u5IPc6gkhKxVfxTARAwjG9KBTdvJ
BLCgxWmDtQRPYHp5oW6IsSDG7cQkylNIUliKYErOzcNyjSBHMvN6XLG86w9VEFnnq7uBTtehkBYe
u02vrQ1UgFsI/9lJlR8OUCs2gRFaMaCQg+ZY8G2W0mlrp3F7wYSTDD46Dpm5AXVmofeXLyB5+d6w
GsCbR27TMKV8+86AbmTVkjKBy2pyRtg9IaUyZlUUeBNUyFfj+Wy1DjX158zj/pQaI8lkmHDKiw8U
xZqDxk81c7RR/t+KRMTC0tvOUQF4tXMWC9PPXBO9HZoTdERo5lZkLbKR/IOfcWOE8taG4vYO9fvS
74/pulhI8/RSmJhq7/g5hm97/7ws8nrh9pNltj+oK32NnkQJmGKLA3/c37XYyjUYTDo4uKyY7dk4
J87tadAvKMgTXEADHJggclJcNzaV8myISsgCs04HrUlHkRmCDOyMoXPNW1OGcmMW+WEJiyciA/G8
TnaGgi2kg2A+C/bxVxi5Mlm0iPmrHOWH6R7IYbv/k6Zw7IE9VsMChF4RD6gS4lrmwDeKNWewxUNv
R6XmbstGxbi1UhCWyu26/aLgtsUtJj/XqVbQE0CTNihulN4n8AbkXpwgAFdb2WV5TCdAQSfL5jnb
jQJV+yxwmBV+bj4V1yOwJSoxv94zhnZ+yEpivPQvfSF94M6ozYe0bm69/zxo1x1hBsamaFfEkDZJ
giNq0khHgQhN74tf+Jhr8wWJqGTK1aMvdKXaGB8EGv074RixPQsrioriV9jIBp9sROReKDmijM1w
c7kwPxRe53l7/qnBfxuP+MVBtFxOJNFLhfRlRcEIGxrEG8300vUKITW8nNp8N5/v/X8HHa02/7Qt
j+PdwIb2Lw1S5lgOSYLJ/slMli/TnIHmaQleQPlpLixgQSYMUEN+KO+VDeUt5myohlaH6Y9cAnKS
WaXd/51g4Y5mVJavKammfSG5dGIwRvKbZ+xL8uI1a7As2H+DI9sJ4hRXJI7qtAqfBfa1FLTJHv79
b/Rftg9rs/7ZMF2lbTDnE9DCSEGlM6Lf0Hw/jgz7h4jhWI/6IKdrpUu5hXzQjASranwKVmrHDgll
jBDytNdvTZ2AXbxmOHMylaiPgSWOsRv8pfJgniGgKvXDN2/JJdGb7sfoBa2LGRdDOD/Fuj/a0iPU
OhthhlaHa02jPqZeAC5lbzznIDl2v9N/mdaV+BuChHb1CuWjvnd8n9b8CWZBnc+g9Zk7M7KrjIur
04iMJnZWACul1z1Stk1t1xyIXKSNhNP1ApymLX99VfJubdP3NCxZpbwpiTPL+x1PQ38dgW47zKib
dIFiP7JIEEtWLN8vGhmj6yFF6l7C+XqoHBfcPbXLiT6aNMR3UJCGSVqthMVr3LaYRc5+x1+tVpEp
LUxA/wsnFD3rvyDyMTSf7Tx140REAE/8o21EG5rjT5XD15iRuecjtv7j+4++GoJ1NeotnT+Q/UIa
UWDWY05gRGE4+coiD6PRU/RoEDd6qN+aunOd6G7cwjE0gME6WWN9LBozK7pPZB3pb7wzLRsBWv1u
ncu8m9NapR/A7wXVcjd7YO6H1LqAfDMqzRM9E6RWMSUKDHsTyvYoorp+YMOxO925OCSTF1TfB7v6
xb6G18TveDxV81BfbHQ3f3kCwWR3tuqGp0auUrFxMDKEdsVkw3bmK7HiegEMHkkJPOx8efZTAQrJ
etEKgtFgTcmvo8WDcen1b9w8ntsXQOEjsNmMEQSKoPnAQ3hR/UDm2YdUdjrxmzxMRwUJe5zstinP
uBSpEqhz1IJJ/bJ/Of1Qx0a19TbjCiX335+7kR2lfOZHU6ykEJ21v5iWjSuZkbDwFsCkgMIn1xm/
5OtsHIb0aLOffLfjb1XEQJAkpoxnPQULTNJAmd1sFAVUEiE/KNsqMtjJ9UJWO+KYcHSbHHDHxQgD
EoTB8+pHW+v3GWHe5+EvpHPqLACIW/2DrpUhQeeAGS9D+dhL9fNIU9BI6xxyNFmyqJW3shsSQlTV
WWypcmKrdPaOtKnTLu3b8FHRO8dAPlb6tAiTj4aKsiB5nQV6NFmEVPVc3H/UyTDTeFXy2PfCGuX/
zBLfZAuUTJ8o7rA/9obGDb06hHkVtqo4MMeyMCgULu8JQ9RDUaqDcJ5QA8RPXWYDQO7xNBqGiJCs
RKQ6aayW9GQymaBZwQ6rVygtl+8+wUapMbylVAZyPZMRxpH91qjiNNhYIcLTAKhzxXNYD19hXQGU
6v3/hHFAOfducUvfr7RHZ8CX5iJXUj5jEEsvHWb0Gtd1jlyvLT4gcyMGea7Ih9DAHlxcP3z87wiA
xE/SpaJKrMgFUSM2Dpg1tOAEKGrumvoZIOGBMJcyV0RosBHuS9/0jawJEODtyJ/asEFWqtPmS0Fl
oSv9nhX5ZplswwPhQp2bhQd9A9ngxVWkzflOvnIoRdOwjoITZVhFxquDWPuLU5zb1vap72C+nILL
zL2SDMKhkRvy4bipwF4zLfhOG3Q9ucGV06d7mfTIYejrb5Z0ksEMlGDF5vg3sdyNL7RWK4BGf+2O
SRiOXIsndOnJy8XlPZGZucZqX5rvdhyrZR49ucyriBrqamucmF/eJbEPekxUnUQFS2W8c/4EwYRt
xbpk5qrj+VPbTzIk1tkXNPvKCgQ4sOD8viZPtfI5ut0IvRW6koPDoyBY8J2cPy3XbTnv7WA8Uyun
O5SileulIUjQ9UBaZP5y5z0kXh1nasr35QAT1CwqU8vbVRztbbusLdpYdg+PTK3npoRh6MzbFKvb
WOwBKB38KQKEqclvl7aI3Su2rr1zVy7kuCE1xiM6ApFnaYnCMOhKy41nU5wJtqsbQnNkLEftKDST
lUZFBLoK/DeXY7zjrm7elx3gG00fgPBRynKJ/dzevILA5k8Nr0LC8TdarxJ8wa6b7LQlZEXO+vS+
Ve9AJflXqmPfQWEbPMWgslvsNxR9/a5i/fJdfNGdxO6P9Qoe78jNdeObzzfxQhGvZzetrxjiG/v9
jlFo+6CHE2EDOuUmc4djKGG3gRgQItMQhMCa/j4tBzeBUdEBCc9EHqbZYGgdWIRhPuCaGvf5sl/G
tV6S3to0IsVSZAdBK1QcAOJdzcEehFarClQa3+HhKoR/5B0tLg3TtCW3YN8608n4xws8vHOAv894
iLUvZIDMHRwnYY4WFGubS6NFg4W9yEXJbQ+0kP3ShnIB/2OLWIJt7Rryx7sG3C3PWYxl1V+r7fYq
NmOLwKQyrWD7Miji5nKQ5UXznikiK4K/6p8u2QigwLYTlLlY3CxHpXEUlOoSBuIUOIWQFBz3MTq1
ojtvEw7ycunmJfwbpsqlCRSZrzc5qiILZ/Glpp1xHaoJ5YwvBIRi+UPfbYCA65nlXmc3yHQflwBN
DX49IOLpLoJVuJB98tsIIH16FXKIdIeV+RT9vXQDaPkNnhFl4QtOPvc/JRenIdCuQMLfZGzVWNTx
IYTuQXwW8O6FozwrbaVjQdM3uV2itjgyhx+qylTOOpUiypZlkhK0evlUINaGqxP4xoKa9WWcMjWA
tq+W70rMgMwJ2vp+ijzWbdbflxDBEfxKSYK+jBIGxb70tCi80rkJXWDDiXZ4R62RCQ5xLzh4PTrD
W7eH4WP7+OQuGRfoy2Fw1LqA1wqcD/R9uMiVBK2BkyYfR4t2Z+iwregjDyLpeMdpSyn9s3KaTFYz
E3RQJJUYjjhH4MaIBkSgOt4vfhRCAdnhgQ70lnEAw4tsiwYj1QObM+yd16Zl9X+JxAV1Si6XofZe
BlTGd3i80Ja1zDyGTXmvWReUmw+aUv/b9T1WmT2taHUuRYcHyld10mmOrTHowKsKoLduBh4VGjPp
F0bBn1mcCbkP9AdpAP3/AAuNuTggX4cFde1Oh/L9IgeO7yTL+NpXbqwFQzH4PEirgPyJIGQwDkBm
yPFytbEmwHWszPEPCcTGBm/RnsFvK8HSM4njzC9pkUggGc065agCpbYoJEBGoeDlrNoc+kbrQXLB
yn3auQYUM/XeZvkLhZPAuegzaGCMzhKlH/TJzpDUb9v1zGvgMcSq0jgTY0kU0VMAyHiAYiTuN6HR
F0Py7o8TNDGa0LkgD7qKfRNzWZfwXWxdSpKFlZ5J/6uAMOhR64MSzRBTh1CQiyXw0vQs0kuuxe49
XNOc4Ulg9CGN5o3gl/7q6PYdoqSwp4+Qoif47Ka9QgDROdLYjswMuNTBfJcxcvbK12LckN6oKkTO
e5hwDulE6248iHRvY21YD+sT1+ywnr2GZxqFHAV10wOH4Zh7wAxdptUAjG8LKx785WLJu/ZruK0r
J76HPQZbObGRfIc7QuHT7+gQMTclkbo9rAb2vFoBGuzsymmZN9JYy/QwRXe9dPu3t5pdyMvoMOxi
s9a2VZ4BZ8Y2qkETZBfMiN3WuQep3r7bDHNzVWzELE9pKctKmw/EI5AfYQ5lgY3Q0oEcD/TVLGyP
Cb74+af/NH+ETgRZnyytx5BJTQ6+QJ6dYaqHdeLbKiIO7drkArkhVBt7lKcLwFGYullHPv21ZkBa
hJTdRK5yCM7z8yTUqUg6t0ICMxuSgFauwj38mmyvaK7Hf02LASTS2NTUzwMaTm5iTYQ4xE4CSoxU
1mj5HjHEI2QLXL8x4+4ErxvXydKMY2GmgyQKMIv5rxwUq1PLB5ZwoM8V49TJdp/NTt80PjIFB+Wu
+f9ouAUyU+YmD6LmyPUy1d+5t/D3gGDtYAXmyxO+AlhPHqBPQcoVn37NNsd4tAUn7r9lFMnVHtEg
Q3nnszC0w1HI7fPApRyXAesxi+OhNwidUKXQrB9by7ZYgEzq3AA4NSpLa01YywofmfYHuG/edgKB
Dwqgmp39Qj68d4CeL1X6VUn1yJ1FtNXYZtWWL6D19N7uB1d+1adtph+OXJiniak9qTXE3x9ktl93
nZHElKdsRVBTA5APHScPytqR4Ek8MWng6TZ2vLcRMwO/EVAcDLu/jMDUr+sVL9PdipOlWS6EuNJc
TY9FUMV7NjpqX7z6ZcGomJ0UMBVyhwzuT2vQNF6C0WQ0Sq+qQpYHVLBvN4w6iqh6Z0ccqHNDrHjw
dSOKL/vaFpBeqWz5YE2tJzagRpbULcTY6NzL8iZey+lmdFRwGXJIV2q//4IQDsxHrTJeAkgfbgMX
mTDR2pWrAaIPumVBqrTFgBuKlpsVZgiLIkA6FbRXeTcfoUi/dxZbuhwoOaPiVrz/508p+Ikhuuq1
IH8WWryw2voNDw+l7E3Bc21ucneWUDVcvcPslafbspQg4f8zXNjSH5BU7IjsjF2seYB0+CnhvAoW
1IM9ukipbvYiLuxXX8W9dTRjM9m8pQZwdlDLBhlEWKcTpZB3Trrwx9QXmV6L4iWhC9DdR2S+w4LJ
FYf5FIQ1TA4MQaU87zhOnlT6g/aro4a0BJqvDeLJUoGxuFMvcbavzvl4mw3el1Ea6E9HOjETsFCs
ZVVWWLmjcm3BkGmkP0KclzvgJ3zAvtggWPxyyDSmh7sVkXNwFcQjCXPj6WTYWAgW5howbuaiWgB/
zU7TrWXEb+LtjtRjpEL0078P7Hpv81ulUDXmA3BP6WlZb2Pp4RkH6Dzm83kEM/fKquGGRYFODCfo
d80DSoLsbbhIgon28ky5X9sscRvBcSI0wl5srrm1bmXvQ3OJLOJaCD2t2ibSe4zijM2888dnTdiV
n4tluuojZ9MJCU5B56kupLiZWNhS5d+96hS0MnkhPyq7JvU253WkLQq6OTVowHDjjTEqqjTOyQGt
A5AuUtvcQjiqdLfYHHZuKtnFV7MOnZCXcGew5mgn03OVv7P2sEhbryGZ2OhWrJ/evdPrM+GWZWN/
6nBRjM8iOeG1MskMvFQAlYvc2uEpHmrk6wmBPezVVZHsQvQc1Ve/ZK9sVN8jwGoEfINS1JkgjRik
COXYgrlIbKLmtiRehwo72RdYzaStZWHJjH2ul3XxtBK9vr/jCtaUZeKCAXaHzT08/xQWva6txXBt
aSxwC04sf1+4eHPK15BM04zgAlw1TXhYxZLoUBxQgUnFO1NUym/MTtOCgLonMB9dL3DSaoSr8d22
fsytSMPl9CbV0l3Fxtx+FmL4KtxmanEEMkr7ZnU+OOL3nfg3eNQg0DW1DGSTi7YER12OI6nL2dWg
IngKqUyx6necEKbPVAdk1gVQ0+AFc5RCF9XZGkFq5+koNev4Vwbxta9+CEy6xGEIY0ma7pnC7M9n
SB5+7+otKm9BBhiqzQJPJo9vxH5b8PPY8/td4EhctNPcvJqUODdd3iP1Argb2hS/cPkiS9exZppb
0/ZrAP75zQPwxNM5UtiW6EK93c7kcrfENjG2ywD/BwkKM79tabXiXSAcib/cSTlHNTeWtteNRimA
nOWQ5H7pcVRPPUT/WJ1rC/LE3tLqSfvsoRMZQEgvOs7Ugcrvkigg9Car2DgTc944P7HYAcftku7F
0fAB8X+VTeNsZnzN1wtayb2GFl4xcFxc4aBWeeOfhNq98x7K9Ixtg+1lvRCIN8xQj4cXJwhYSa77
zexLISyRFKS1Fz4JQ1w/0RH3ZRnSD44tCLnjFD1Z4OFdU649U/72FRUM8nDGQPktJW0l1SFSLYBC
lJ9KqKDbpgt+q/iuuMg5BXWxwKpbSNlSatzvAvDGJjZX3g23ikxN6ByoowGfoSa5RrIHhcxOCEp7
suuxJQOYzmlXuEgK/yt1Aaee6n8I1aejgcXzkICJX6dsBE9rtjUk766zEetfY8BuG72FP9l88E+h
+w+OmipBL2+JnqRCl7ff2YCqFbNSzpuRGm1wSQmZPJB0n9KIIXVeYYeHubuOmQdp6T6oqx/ttpzd
+X+6lINbEmY1tVKdb0BHgEjYkPOYAgUrGTozbs+6X0ng4Iw+Dz3Go4CpGGZR7m1h6+1S0TnipNDc
tDCemFVpt962r9wR4keYpjX9fITKQmpTh3S/Fy5bljjjbJKLCwKUo19ig1wxYQXMPwWnRN8Zj4+C
SLCkMdcMEZKkgTyy4/nCJp6vi8swtxaYSD7dvkx+8FAZUNsmO0WCzmRUdi1t8UUxdKLfT4PiJxqG
XyiYlf/YWSjA3pkrp4xX9ErRaGUNxfZnC9dUAe5wJSEW3wvSGivwmPsM6RGSWp8pY1vI4KAsniuB
jA+pkGsOTy+5+ztQEo8YdnP2pHNYLp/da4olLlnUx2cQGGtKc4gfRsMRIMXEeW+rAKIPT8g4Yi85
QWUwIFNNLDYAGjteycJu+f2HUk1JZuI/y75YMH1/neQKF+tSUYOYFXQ8OdoR/YITMangT+9AS86I
GhxsZOwsu9MoEsMz7HU3yYdP8WbURM3ir4lKRZowqvJktzlD4z0MceuMtlQ3L0sqIY5RL3vPJFUL
hMY1eI/N6AVuFsfVBPtdr5TQ1pUWv3SeelbDdki301IsjlW6rzRTdI3UodqZ+GJqC0+N7RK692h8
+VpcAJSYDtcRAhTjO7V22XKk77js9eNAo+JLhP7aNkQMVWafFGWZ0d5CO3XZTYX15PgqzYeWegMW
8QIcy5UIFgPLakyik5O7uX6VPvuQnWVsrWnf4diihgDVkQBrKcnTN9Fx/BNpaGn2Kzq5njMUZq3K
IRmBInYZ5auDjvOX8U7CuNhenQuKKQ9CzvUW4Cuv5jMtT+41//AHTqAXUakCSNxJoOhG9YbfSLx6
zqtsvjAPx3nTafH6n6f7uYtKatlZXdtzBEnwwRXUQhBFxa1h5prYKwHpQEfmguoRqtLZi4uDFrym
28A93clllrAVJngGs/GzXJ44n0Q0tzaRD5kweaddKyBvt+AkL5A+HY08agqMvdGWMp45qLejJG6j
Cm34a5ky6j83YbQwX1eQZjDaUCCiNAxkg09isT9D3iPtBII67yKzh22mTDxZDBfGycOzDASSLVBX
VBmiIWfNtsk4gba/BhIW0XBgXuQYddTqyrOddbHKcitVIueuz0h9DW++mAwtIfbfxZBtLYCwK1bL
G5O0G6ZBxwI9vPQJea2riRaD2EYAhGn7JICFmYSW6Jb3xhpiLaVNW2xQu8untgWVcRBDafAGS1cg
UrMJ7cunGYFH+fRXQJU4b3E6nqV16f2Y+3kU+5xiR2hA8gbGFAqFFMa7W6WaNOicig+4F2T6q0mT
RwVBuRZg0bQxfUakKtQkj7XHnc+AbXG8CzcDHGQDkZCnpcXKZao7iwlC11vSfBAeSxgoY2qMPwwk
FWCUp1YpvK8DNkMYRaK1wAEJOAh96tfAdlG9oXlTG9stlxH7ntrmWws6TBrGrRVsTcv8Ak+1O/3m
I17ytYaqvEnOQjQtX97qZQfKIdUf+67L+grJ+U3oOEdCUjW31Zp4vKhugpiEnN2Wdi69AoyGZY8n
un0KO3bi5uEgQ0KS9egzkgnNBT6cQULg0xwCJgyhzK8PlhLPuGebW1Sa4EchHo5r8rfQoE5RdnKF
G9agDd2+1Lfqh5ZL9Iag++CbSjPK3jK3bfo2s9As655VV4F2K20Rj1PtVcrheW+uH5ebopHYTqFo
Qi0MrmpXRzQQZx58pai6iZ8ImL4wBbIP2LqTZH8eCvpQM2oGurN4wpMDtPueGtgeRrDL0BKejfg6
F/oC1QZlnQMFxYl5b5GYpF+1Y9ZsiVg+iuz1iDkFcT5RsLte+zga3zIXz3EZV7zL59KSlYTvqhx0
oCvhStqn3rjjuIDgv4GVswTJ/9xjxV9SUHPO/AzkJWF5zzS9J+yKeFKKrbNYp0HpsgYFLm1T4AXj
3bO9TazGProVDYMhLEumqszwCedKcUlpLpDdSDnNUbup/f72qH6dLm6Wc04pUwieXakKOntUiq8Z
X7fnTy8FQS0CojQDfxurOk0WSIP3Y4phqUFUA/8HV/N9qKGKank9kWfpD7i/uYtiZwghqor1FWx4
FgGuMMzaCCSStkXNnZYV0zv8KHO8XYduv+0akaBHTH/ufjGCgdkb4FVeIoWCg92g2q2PzLFRVgOH
Bv9uIse/nphJnUmfxnZMAxt/7gt93t1ouHqe3FYJMoG1XlnThhLPhBZLMQ7sgn1vzTe8zuLNzANc
3iuApGG9frkKYKRcnMyhv+8qsZ/AhQHor8b55vlaaiUt85PT673CqDwjOHWJTw/fxvE06vKDIJjD
VfQmakQqHxY1T3SPxZXObM6gm7C82wxsJWeasEspMvczH2nQats/bFzvi2elwj/qMAlL6Fa8DkBU
euhEyjALMgnpIjNDgOqwS9Eys2Xl0IJh3sPgH++XHoq/gdAsNYPcnxsTg/FAyHg6mJKG4+ykapYn
GS46sbq/+GXVh/W0Gdtx8lRtDxd2R/TbZqhsOgGpWkS5suPPPQXY2Eqc8/afL4iwkAp6hQsMeCSI
f1G9pBJwDEDdFpJ/o84FKFQC4D3AM+x12gk13mSIiFaCq+0NM+uhknJWHCXwUYgJV2MOKJwVNWXT
614sJXJUV0gMBliCaY/CZGkfZf4AGPm1p114u7OyMKK0TTN+bhcRxBrVfq4X3rNBqzw9uZB0ROMA
DDOafRTiI6Ni8rrjqgrUxoX1fkgfEU1j4qn1oCDlZVDCExWswCuAPfaD2Az3jlmAV5F8ck2IC9Iu
rnWb8Byw6LZ0phzgPRP9opFPZWAPFrhoRvkAkDcdYfsDdnRWr3v70zEahwTIQnuh1zTOjW7QxpwW
OfyFQgT1WLx5+U3xeDpL9DSkO4RUExI48vpDYse5cW5m95kDPHyvf9bC2GakpMj+MrpsyaolZC+P
1lTLlfOCqv3EEWkwQgE5rHHCoO4JBNoNJ2nkaj9St9MJOBjOnKlt18TMTZzTPEu28bpsjkbJrlCD
Lt2Dn11n5E4Zp8CqSz7hlM4UxuPQtpk40qT1SmKE2TWXyA7fouXtvZLkYTlXvdQkLpLML+6U/Nd6
052kKJKPwK0dq2d/2dn6DAw8J8FRL2Deo0ZUCIsv43btwmeza+A5vuslKrhhhnPKEomcm+eFWt3n
IW8aSTBB3sapSzmbuegtPMtkeBLfyudmJXUxJeRkb+JMCf4sio6nCoQ9tx0GrBI2IFkBoaFc/cca
UBdMuPr36LszRP1L1575x3M5OO2armUoY6vVFbrYeCy1Ne0MNAaWcLv5IxTLjAC5sreXjuPTZFGd
n6ptOaK6m5BgdDH1b66V14k4Tfh2/2sWq8t056KhLEb+MyDJg/iSgxXc/LHIuQQy6L/yZprk+E+V
Vv9EVHfpg1koYbgmZ68sSmAlgsM29o7+3bfidYC5+/wud5zEy8ZSBRv/+Q5oGoJjVTd+H8uQsOj8
IMGC8S12f5tZIMqGWMgkigVbE+bc7YzVMiG2FrWNe23gFLqZOqegD3Jl7UMoMPyOvscF72o94dQw
slU5aaT1mxVJcVfThqag4df78AK0OFLFbHMZxo/yX01eoyT35cedhJ4lIo3VJf1uPSz6mA/efhJ1
8OcUkIbixLAVv47O6sLoDX81b3lf1I+eVTVOw2238+0pVjHCXBoSlpEvXouxRErBEpPZIUMFjtdC
iyUBmOqngw1EQton1oinnjffqo2SfOaio/D0yH0SuGsN7irqHvW+aTVdDE/1gnBqIGQrw5zcgH3o
Y8chNDxfnd2PuMB12yGfRipgFZ8cMs0bDzemZa+uRCXs6ADJyIaqgQVOBp9bw3CzukCC2sf1Gw99
9gJ1A7CHciivY/qCArLAVV77PINX0B0G2uvLthwRpET7ULemdJIybR7JUF3eHB2txOzKu/yQfy6D
PjZVmu+vguthWJvqsd19kwJjBCZj20ad6jVbq2WwnWwoiwuh/fh467v+b920YINEi8+Dey4ioMco
MhU6MZnQ5D3vBt0qvW0wOs8k7+Z8Pfg/s5IdZHAqiRZvn/KwX4BltgJ3vbdOjKEPzx55sb3qnpH2
YD+n7GGUsxPr3MT6rr2wki7IPnOc2xQS028R64Jyz/8n9/eqtBE6VjbMr7uoskIWuJMIkY/12vJZ
TgEJFCWAdNh0qX4Exawq0oIQ4FE4gSOOXqpKU1bF9SsaQhIdZQ2lz8pro0LGkTLGvnU2wkJWA+Fo
3bZbpI0ab6FL7LPKJwREJd3zKNScUkXoWCsucfyUt+96nkSge2pwOPOjSte/VSsNAPC0uhKgCWxi
slBDeQ8Td3od6JspkA9LEwMBJiJgaSrhKStDAoiseQus6lP5XnHapoI2egZwt0EnXPQYiGNqgYHb
dlDhmaZs1JUDw/wXfiNbn149YWydTkO275rsr/YLVilUZsdyf081+VvAhISjGMWmyd1ScFA2jCWG
4LNCj785gxNr0gB2ROEmkluUbnAYeeNgtdKI9kE81phDueKB7ggu4G+egb4xneyzmMz4VR/4mKu6
6Gq+fLKWzX3uHHIuaypOiSbPFpfeuBbpC4qyzVNEhhhs/70sxyadmHQLNJoci6OwdguBaFgTbfDL
I5ViqccOTiIOw9c0cZ4rbLDhki6Yt8ilzyuYkT20n68dta4C4A3VpaA2ikWNXuk93yZnOFpQ4dfE
hGIjTYyzDIDNMRanA6/6a2cqSN3M1QU1opk0WFaeCPZhMs9mqxSTEWsTESaPFcqbtvHYRyTzV/S3
Po+0uI9BQ00DpexpEgh16+Te5EjmJ28YBkulfnrFjbmUzmSviocFwEKfRnzczrAaNNa9XBCY8802
lH06DgznxP3qQ2Zkz7aCpqy//U1rkIk6ygcRhazNZUXKBxfIfBeqLpvi2GAh+Q1TwVzZ+VjipU/0
xuw9pATFMHvuS49ya10Q4S9lgP0zHmStHm/X3BjqFCO5A1gqO3PVJ+XCPTOriyTqSvck2d1+HPaD
rXTOcrpT0lP7A274qjDd3TbHokJFi64dibmdtgxKdaeZS2PxqO71rIKIIk9vilYnoSLkNXuzJ5Cs
Ts9tZzgnGQBIX5fRhImuPWumasxSHim6QvlJx7ctWG2tXXLScl1YKuEl8VoKP5uA8oSqtErbhV21
//ioBpxwIfbjEgXyyCr66TZOVjXwfgOadj1gRtMB7oFxjRTrVxrMS/Cilb2Kxngo50yvaQuypfOs
Fn1oOXBn+88VSZT2rOSJWBNwjjzulNrJQ2Ia3KZl5EJfD7CjpaZNHXMwtTn4zaJ46sOSuCqDqXcq
/lfKNANA8VoxERLuiyqEUmlEgHH7w9HRdiITuwixYkV6sV6NhxOz+qC8CLVTu99xSkidn3sOTNie
or4lYFncNv6JXGyJLbW/p2p5H/KOEJyxIwrkT53F0Ckh06BMA2YuJWCwm8ho0JBmVRRwzvJqaUKm
smtTqFDKtkjb5Z5OOY/4f2pY6AmL4fSDHgIDVNINtR8IdOzOxf3DeTr4YbjFgaC6Reclxx6dt9WV
Uly9VKnuz8V9MY5MEhrXRDhcZWYuIKkxmXsJJnqPe3fz6nQinWRbqhiSCS5NG3LkAnwM5QqZLppy
nBtwqVw5gjFzVfd0cF4s1igcrcGiKP9aVk3+NvND2e25H9aCJkh6aApZe5VCXDjf2PigqLAfPP2u
kaciqop0CIQUCQPA4Q2/CCTdO5kYb49hyLUvejzBs/NmhBlLDkhsWPXIoTdjXh/agEyGoNuvrMi9
VlGlLTQPskhWOuQOwNHT/udD/8rmetdHq9PfE0aFohY+RsvCJ4OXb3iM9PgNHekvUmVDZUz1YSKh
Wy+GOpV3mnRzMU/smeYYa0OM0xM3z/qMCJ4R4/1AipH1gG45nTFJl6bWWADGyycQvXGhPSs02bTe
MC6KWa6TYhrbPiH8Q9eA1sSNnjhH+eqo6fJBGjWlW+pcoSNH/CF1sk7RLxvY9uJOM27cLdKHJWUF
qkbxqkJ70t2/lQ9Ym7huA9maKjucGRC4aPWeqfz7C3oySv2ZDjlB0Z2gC3q5GMYs5O5nw72SpCvI
nT3aGnwxVPgeZ6tc8SVaVansLqtm53hJEdXc2qY/+YQUuOd1P11zh2fcr8x8nr5RPziC7AyKdoe4
Cw6raGIQ2IqRlbWbkjJgR1KucDe5FCAcquitWRybejlSa6QsId2owGRsVfy94SuIFQoXaV9ROpDD
y6HEzp2FPqUMLaZfzoivk5w2GvoZfehi+f/3I5wr1x3fBapTQ8dZgeUjowj0D8BsbexjcgW3qlIO
jFoamB+gIIVbYORxySZC0e/aC9VpNpC7q/4Lr++ulfEEVemBio29E4MglTAnSgbzWrkUJ9E2QeA7
PQ3EO7F5xpoMiMQ2+bmkd3UI5nxoZT26N5zqdiMk2njd1Vf3TL4KJJcPoAti/00AMaNuyxP6msxI
jizcwnjWPWXZas2/NRllN2213OPaY9Kj2HkJ+KyGMSYVT+YyuG+6j5XidAfStJvN7IfSEylJaJPn
KRY2Y853fbzdoN3Opmcz3bjTDF4P/Anzp6JBAfi+OKyG8jB0u07WznzPGV5aL7ExMn/ZsK31Vkvp
HXUURocVKDanbSDj8ZeYRFx2bowrDyEyRDGf7SJE5WUjTU3wnex+/UkZtTbiUABWwHEU/GS2SaTo
6y2ns9Jo7Nm/+PHvugNso+CPNqwxvx5shqYWLargyq6XD0pG2/3+NCPPGQz/r2iq7+/a38sSErgb
J0AbciIYg0EtS4lbiacEQ89QNB6VamVfr8vpI9AYbwliaB2F5a3Q69c7cmwgO+C0V8u0en8n+mBd
rnRkPnQBY8z2NyabSkjstC6T2Mz58KjOYhyhCgvuGX6xWYo4VUfVAniVL60t7t/D/NQYs00PgiGl
jCExdrn9WDlxWW51WMBq1gYY8RqIMdWf1ATMwGXNUDg5n6n4xeTmFuaFPmeKyc4Z2DRKJYWDCaR8
lAxYQoyJby7w4Alyafy2epmPTByeGw89Vtb0xgYJHad33JoLYYy2Ud7TMiaiAqN7iUJoUvNBZNiC
afr7vKON84OFqImrrR17qN2jU6lxVn5/1dAVdiu3RvvLhw+HWU5aOvYS1OWY7/U0GTXUgLWvCY/X
eJeP2F4MlGeuf00E5jhrxyIJbPFGkxKZSjbbK27oj+dw63FAt+POrxT2NFvfDG68/tlBkFH7YSSl
6ihRkSGJ1/R7DA3fURfv0jh/w0hMk6n9Wee+m4xLSK0g0sW4DsGNJ8SpVKk5ITLxgp/0dACbx1ai
IzbqPg1FbL0k7W2uqKIvJ4hS9fC+LMijo0EjoT08x7rcbp5GtQFfisUh9w26NpukhUqya/OAszWi
8pW95MXWYcPUjTMIVROfVvECXpuKNtX+2DANcZ+f+zSnRQqQ9xDBVas7psCAhZaj0Hrj5zCLrGjx
8keCZxw/c2J7+hmsb3DHE5YUAETGbrYab3SZIb8iP5IDQDSe+vSKzB1o/OQQrlTZeZ6VrZOjevey
Acg+tiwMcfk2hpBjXaHyO+s69K0Kq82oCvqkDzj9RvZ+cgGRTFplZj6ey1w5+D4Bu/vM8n86LoCN
9bfd6tsseTyTsBU2u0/KxIPZmL8CxzkgjakBLDPW6wWtxi92JoJNyV7ruE01A2p2PHMyPWYnc4zo
pP6aUBlYiS1kmt5jZXpYZseQbsL4kBkKI/Ss297CISbybTLvFwlPtniwar5vQ5Mg+0Uu5nh97eu2
cJqcLIXCTKzoMUiylmAkIr65xgMTc9bQLKvnt/F/LF5LAk/f10NyOlRVdTGqloBtfxMX+QVw4Wt1
TdnBc8rvqZhd3a3K0kf8Dq2n5ZJiQHbGigajReWvFhK0Qq1hP7/lu+1KoskcfVACSzxkkuBFuxi/
PQ74EKg7rK9+jqxOTM/hFtd1EYhMR+2KcOlGexKU+9/cPNof1SwXgBZvjTLYwWoyYqzk7LLphXd+
M17+2uh/qTfVLtTmfboo34lnIwpnJCr0o6Z0wx+l7agZIfCNU6oiYXFVpeJWi70J7zZvLWzcccx5
JleMqRwV7CY+bWtDagTzJppsZqmYy6qsh+Yox5ktvcorGt0MH3g8/TQQeo052QiJneUrOCgHfd/T
0ofGvFSOv2Xzix4UZ3HqMWf1Lu18b0TAkzgHMRlUnbyq5rQUOVoKoSaghkitSxoDshT6t/M/idMl
qTdpJ6OeSD2X3HA/i445PFz6kXKtSarExOFV1ZmRJG1SNJXAoP2W/R2oIaAfkWuLWCaqbwAIW0jr
oU5qfuHdCfpfsi0I2gC117TyA3o08b8YURncCqmXsVEYrhKuMRehoOkLcAVahVwgqL6YNCSZh/1K
InDoOxFhyunMwsmRQNRSh6+V7Bj8mCD10Psst8PlVyQBHJSby+GxFa4k0h9MES56L+NKcwXsI9FW
lh/PU2HYmvHVfsPY9URnsbQhSWoODj40fHAVSteL0OhQalmJDiTt/hI29EP9W4ENSan6WdsuFlGU
TYl/Qdf1B8fHFjS8i55g1b4xuYjbqwXguWnThQTzZ2ofTiYgPQLro6Wd7zmKa992po5OPVrcDuUx
noEKqwxiLlmS1t5xiql/zADQOdPTMecV3AM/CN4uetE/A/FVnmSIV/IuLYO7hXoqO2a0U/txRV7q
mat7uzPFxsCAaa1/R8A0+BPrU8BsxWClSGucX8+i3AlJ2F1NDPAVA5c/9+yXzQoqY8EiJxg3Ieqi
L9qsD59Z09siW0qtQtVIR9jtbL0buApMDXylaC6QVqAO/15xy6mN3GToWJ3sW2r4dAGrVfTpfSUv
jEk7d1W6Lvdh/XhxBBSah9PeYR1Nmkcbz447AxSPitTg0O2pUWuhxzqV1A7CjKZ2bRwRnJA/wZIz
WF5acAAQ/7htR2gX6fyiZNBA83WS3VD9r4AbGYHqvP9tUx1+e8+CLwhmPpM5Ab6Qld8t+7+JBRPr
qIGOXm61l1RYtcAFKVcxg8tkYXtquhnbtsi6zFfXFdw9nPNZvcKkwKTsOmR1SRJA2Xb+myNeeMDE
cg/cKb1lU554C/MO92eANX9gwEkCbYQSLwTWfCUVLyNmVRCEE6Oo+TjIyx0BCn9AZ4oPrWsm5mxr
O5AZlrnqtBFYSJuzI+E6NVnRojAtamAiJSgYxmIYn1y9lGDRv7m9E9ngSk0VUSf0W2vraS+vF1DM
B/yzTQjVDEBNMYAEMYtPkkZsKRzUG7hGNrXV8AxR0cV0nX9XrLlskfGq2JXTI+kWH3aMKeiIKVXW
I8QXBekkHvBmI2B4DVjubt4KIr1JqwfBkamugQcdC4kyqcUnzj/4TFuOXwclOCEhrnaQfVpnBh8p
NPvAMqTqQBo7vBDXqX6QEGzupfnLShMlFqccVUGDbyouOrik7qfulft7MQ1otF18JxHti+LcKrYp
vW1WkaB5knuf8bpA1kPp5LsDwNiZkFTGxwYzAp1PfyS3NStneiS3Y68nmmIo4ThTkoHMWRwLyYeI
k62+tpl3b6ZS1Z6Fx7DktVbm2bIfudsW2fcjXKXGo99lOs5LFA3WXVIvsquBmTiIZWCMBp8BZUpU
PopqTLIuEbInenkEqNEoeK9awcepvX6BKFLdcfLYtiSYRsd67oy6FIZ4xJtaPw7Gwkt3iyKuoR8y
sB4bpcm8ZXpLNJheEnqDgMBI6seFkfku31Q09moUoTPOEkWgip7YbeEVX7zM7LM28hxqqMmI7mPt
S5301+BWQY2jjcppVLB9iOJjQNDNf84lUvdqzxG1TGMY7Zj/dKAGSd99+YtkV5i2mVaE8fK7a1Jz
Ul1lh8s/ldfYyA6nJVE/+tZ8ibbQI76EPBqWnHojxlSYxqsUozCfHKp8yGXv4G0o5+/bYwmaBJ3I
fbntXX1G5JqPrq0z18qzopATT6ilqbtfHsQzvELCZz9Ks52vlMski1w1jaoEOBazFSRpeM5y3wIJ
RWFaK1eo3smJopVeKjnXJEJi+kOoMV92kvc2hcCusoWFzLE5FCXD5iRUFqNTRunYA/gaYcqnvjqv
1mbA84e5rhYZX5T6GYuC4gYIfVbS6LdcngSKyMw8UMYseTOldeTg0fsSejB8psaX+szv8TVLDsmt
15BRIwjKglTNyDOA2Ph3frJCseT5U7cuumuA35vK59wcloqGURgmN5Zez7uMgvbXnjZyxOjUvNXl
Kr3z0w48RYDGjk5Ke1br3dqzcbdLEFAsWnvq4wqScrE/euZr3u4u4OwYuSj1QEaRwmBQPRaArWwd
VRdKL2btU5jnGxLJS+tR++CihEQTrLQtbFxpl5l1bC7qr5XoQ9dMcoBFZyMm/x3Gkzsp7iQ2KtRw
7XCmnW2V5Zt6CoNp9Ac04PmHMMHsktIBI7yqf4eQIyx81xxYcHYpYmBnN7ttsXYKmbKahaoGxUVs
Ms4CGj8buP9KaLz6Q/EliYE4FZ3ZfZ0h0SmZK5yTTUHsqUdM7haFsY5BOUnc40+R2AUigNIbJNpj
uvoI20ZBeWZlVu75JhNDmDbNjzXKQu5MZxF7kCLddjvfapX5E/0wmTy/Fqc1/R7IniesFh/ntl84
gnwCqAXcVXuWV+efSDJQzRS7POeNebJQVo62XQkeqUrGhChVgT0ZWY8KR3cBJdou/S45i4qkC9Uf
zXFUzALEy4nMULxl/ojvcEGIfVpChIMlbqLVLHDcILoO4MgzFZvB7xIokGKcCqqAosr684rkwekZ
zibIlzXHPLmvuMyceNLQI1l1CgWQfHRhiWAbMCit3FVj3awdH3qWflpkI3Cu11tEyObIJ/ZGe9xn
Wp9jEV4hkmEA/LKVabny4jYTZt1yEkiSLgw6OtYesltO9uQ1wc7ueEuZSC3CWnXAN4hRB02UNmeE
hwY7TKuWMyrJPJlA3FkDhdw9GXiaqmCSd25clggNmP2wIQoo+9psFGEtHUAWbblBDnBQUaJm7xVL
K9CY3Tkkst2yF6sh6WoYIEw5fzeT1+f9kBhBnx2CKXtZiUi4zBMGaRPUXKkFRmzZ23z+WMyzbmG9
DQdA4NBYG+AyhLoAo4CtzJL2Klcz1lo1HEDg8bw47fqQYlAy6xhrYObGhVBDLMxwGtlYUF/DvF4D
XN340leP04YYeqIzNX8zme9/thU6l9+eN69iPO543vucPU1aWR1heBK5BTWUoTykeSVOEXksBP0r
ADOPYuYlYhdAeQnhiS7bJZaGxb9NzJh6ZWmuky1oRlTVJMdBa12x47bEmvdJAma97LJv1V4H3Ydt
Q4XzK/sLe84W2BAI5GDbZFXfV4MZEMhdfPVHypz6u3hW8NZQZX3oPH17DqJR5Xr2yAl1998sXqYu
OeSNsqQzBpMFCBEmQLZFr8EW+57Vliyc1/igeljZrm+4yZjEn167VMPMIsb/DdwfpxrmXAE40jk/
Fa/MBN+A0wo+g8yFYz5+P6s49Rmrc9De/cTVTeOh2VkoC9bmAeZndyy/xVIRsu5f0pfEUTW0yUnb
ISzhkC6SHE1HT7w2/EzQIRLs1TwDI7w0XBP7JzkU/sJqRESWZjFEHzB0GZRVBir0U2jWaf/PpMoA
YY3WoWj1u7HkALCou++4YP6hPq0y5yHW45/7uQbR70W8w1L/9kZXkmeGfDDQz9TI/5kpgcmGCC0F
IWwoa66xtY2GhIIaKPnM3ylOzWFF/qg+7iMc7cmvCzy5pAzOPN2UfB9iqoTij2WVyG64y9PjRh91
KJn42TPIPHJ68JeP9aTAGjeFSB8nYRV2IXovPqSDeWUgBH16+X+etW44CrMOhkYPkd/Uf6xN2aTZ
0kmhZimIOVGfpv8h+y0/9QLdgp2r6mKf1XpAhOQDw9N2e06McgHfFVtgJcVqgP0vhCBaVdTKT+gk
su4slbAvrOb++PX1SnVrsPGfU0MoobaAe4c6ZLT9OOvXIy72ORGLTfGipib1XXe4g9/3+gtXuih3
C93msixGOo0aiV+XJGa5NnNYr8BrNGlMydMacmUFKnPV8tKWloTf68g5l+9Q/NHC3MwcVY849T38
DMfkwZqqHyNFi7CCK9MYJ2GF/f+lFp002zTtTpgzBBtXNScUpbTj72Uy6zTrf6Aj2xSO3bGtt2R0
IyYSM4DjZrTsxBp035q9k0GakTc7C5pe1TzA8PMMHCVEzeRUmicszKssLm4Akbda4bmH+jYwf073
uydmzlKYmlNG0658n995BUZDx5zxduZ5IwdMAit7b/T8EHEB7oDTH/17HEANDc9RZwxlpvL3ZSqG
qaYAI63vyzftWBeegvq3Oz/OKZPBUmzNjrug//oaEChR6JSch4MB0HC61hlKuSH82KIvQ74fTroa
kL1CAdbVNKWi+BOh4DjVmQoGkTz2XvSt7QoQVXTxJd9AiMAZm0LOINs2a1Jj/LBFwg8YvCCkeSIm
lSm4xolA7n6643kCzBybDIAdrvaBOrtI3r9JO4oOmRBlXa+DCPSyIrbwsrcF+W7Zd4xZtGYidz+a
PqZqsw0F41adWBzgIq8mmrkmjm24gDkm0j1n7mh5s46XHNJYcEiC88SfRMbdPY44jclvBH7UU0cl
dtYYNUr8dqc+09kKFJ1jkQAqij6wSnqmD0Ol4Awu7fBtRXPTdFDvumOKB2RjfgYMvSsFC1OSuOM3
Ezpmny3aYRkmht0eG6ScAupZXcpyq6du9TNd2X5/V9yxGUJMuDOAh98noQLQPeXwP2G8oqkavZqI
9UBQ7kgDF3yyGRB78mmxHUFPPK3kfULyTXK+eVUp/nqOMCNriFksGpF4HqH8zP+tPgaegX9kxToS
ExnwrT7/AI0dfdYMRkB2bO6Js5nmWM0ttxCnqnLevLN6A4Immr9GKc59ERREZk7UdWNaz/2ub40O
XfAAu3foWhUBsgIPQY9MUTtbWqglyyEFE8hnPnmS8kz7c42au8dPMwtHgvaDxlNQPgCiXiGfcK6V
AMjD/vDQLjDgLc/kj1xD3TOmriHgFyl3DC1TwOQtz4KnCWD0Tke3ck91uE8IajT6+gSxJDDqr+Kt
/qDDr2GbbRS/OKcXOenr0JPo6C1IYIddKpbU+C1T1ccYxzw9Fom/SP5cHo66dQlpxWSyCGOnt6Cp
mCES63E1To7wCs0uKmJtp1FvjKTEILMICO+51W3DPFm/IGWz+qanT7JEWCh+dKxWRgxHti+aWvpd
6mqB8h5OZtHl1LpTMalV6hsD4S/f9f54UP6KLMR+9qttytxL1PxhmKMCA4zeGeQvkNe3KbNn3IXQ
R6EaRhDQJw4ozdtdKpzDhYndqgBergO2N6Xt/cqU7CQwlDP9gdvDTGKaC8eFP/FZsQ7BDXKGBqQh
NrwBH/txSzCKXgJ+EAL81hofakPBLBNCPV8WS+NquMQWnqGtu9ONhFbYj3b3aQiwlvDfNmKmMZ/Z
nJp/D5ms7F2OFF6uVgKRKy1H5C/u2vK9n2YOR0Tqydct4qgGxXbobsuEGMdWXgznyynPbHEoBJdR
qXTLlETJpgB6Droes4Gs5yFuqP2tHQbJWk2S3DUaC3OVxWv5uA7T2/FUtrTmHr3VX113H7+s4GTT
IEFpO7hxXkGLIii6moNvwZscXfSBM+BsZh4O25cU/FdzQ3l6+f5g0S+L2BKReN4S+azPMRf8MAV/
jywl9t/S6tKqwO3MCw8sp24r/T2NebIbxzu2ToEvOhxDyzhqXFtQD/RWl7Yu23lFAF0kVXVe9LuV
zpnRuT/v2ZTQhwhusaQuk/F/iOcgo20xW3VOfQujnYEqb6EW6VVF0Z9imD0n0VgE4B3JQ3q8NaAB
8qLLWV56WT/VIu9ZtJJMIu5H6wzb7dB0xoqjdNqvtCWybheepfXRG4hI65k9t2H2XHfgqy7KqHEM
/4jAffeBebEtmDH6eudYOAsBdsy133mqdBVjRIiU+bxb9scREmWGH8LUqbYtfM7YD2GjBMDxDGMB
zCsjjvjxR1h/C7FLMtSYfBi99OrhnPcUJ08YshAVq6tuqN2WMM9Qjm00G4Iu5LGJuStjpLWRoVVr
YmdWFqxf5QIMA01VOTSmdyUinFlGdUgS3fdchItleryrkc7/kWZlFDpATeVkVk6QuOvTz7uLO0H6
guODJTFYp9B3PqDfmECzCEAtklVE2q68IW8PeOs4c6S/RhG0RGp4xnMTbDboqoxDQD4A6cYxpq3w
P9pDK5AM2r5UJbZ0hN4I1ABvtiIlDxpG5kV/m07lfrmHxQ831wBItRKwK4FsKQpV4tlepP9/To3I
N2yaIOeyt41OLjkmhivQ7cmroAvCL2TURDXcnfc3j9sVGn64niBsHjwsZexpMvZbopIRz1Nd8o8h
pa0gBaAB9e3mQLm4EC1MyYBEakTpuE5BZ1P73o5GpDy5+g+lSOjKPaO2wE1vKVQgB5dvnHAT/RKI
J9kW38BdWb6cmTMHdGJ19d6McKVTQ9ZbH/scYOINILa9LcCLbmdkDFn4AsKrN+Hch0PuhirLN3Rv
UT/ifWDVBwUktLajSjOofji2VmT70h6YXfzwDjKml7/6grYcZyp0CVQylaFCkgtxFdblLn4oPiiS
yJhp47sm6WTKBXnbVzCkay3n9ouNGykkEXXOvGo2ERDg0r6qj0ZlSitP7Vaws3sJESqydT3ppkhp
f0fu4geU90W7OHYFDK/IXp49ngBn02vH20OFF+8nh8RTfZAZGIVntr3uGbCeYco5mEN35XzNfj0p
pt+FDFovWyWO7ZG/Dqx4LSysLWNkQZ/cNYBeojeFqMCGxpNE+Yc+M7OXOQI5jLIk+H3Vx46Uqee4
3NyfvvYBgOWfbL/Ir6JdRraBbcm4bCNtZXh6lnNNUPU1YNhk/VQ7G3o+rTXhF3xCn1P++H8bWcL5
JgGutn2lyn48+fDohiJipEaQFrOyquaTUZqWzRm5rgoApu799Vc2ltodcqns5szC4OuRuxF41g0Q
Eacw4SnVrlDAuWSgcjQnW/06WxCWCdgWEW95rixyGGaanGLcDjruq56ksFz2NIqC3ha6C0J+g2AF
r7GjQ47giYOa9fZGbKyey3qIImpGPV1U1gvaJJgPoREzebIxSr90ptb81KFNVPsP2bP8/YIDnQ7y
fpsZPcZp6t0w6rvEqJ9cW+5LLmg2jeo8XS4CdtRZHGPTPowcb+YfySa8yPEXTchO+FV8pemKhfSf
BK6MFOqlAR0zE435eVrqFmpEwadAnYGv/ZdXisUjmIplo3/sc+lrqiam3WGHV7gRfxLl+DiBFxKX
AYVe7gclxmwehW7CuyhFWEi4L2MqnEMSkEIP6H90My0G2IpKSQLWe5rBa3YZ0+p58Z65hEz0KBFL
GR6jibbEDEbwL5JEnfAfrN8igNYD+/U/snG6CcKHUJsWDpFKykPllx3Q8BGZb1vsaFx36vy8R688
h7D1p+NKldCqE3QR8kvO8FhqxXouU1f9EhYx+uR0DwZiM0K1pbKTphCr9FrI6tn4hE/I3x9FHpBs
nqCXiRNqAMS3ej1DmCFjDatsdfbc7rwYfe+1DlCh/qLiey2UXFDkTxsIULtVIOeFyRZ8Kwra6K5F
6C6fUP3cgnM792YfUck9Ly+7YBuGuCeEWCySxkT5DvNnQFiz0eXW3xAP1LgQZd4hEt/8JDLt8PEN
7LFgsWUjK5CJCMc856q/MLkXrrtugum1cyxFNTZ9Ch8/M3mXKzwcaOq5tLrI2YVKPK7p1nMRADUJ
9p37apv5wbcrM33lJWw8+SEricT3iOYiPIfvQJmfgCBsg38y+dT8+AcaG9yUIBhNxhpZ5Zztc4Sm
m5N98uuAU0dvlDPrWMmsHozq7+WR8tJsvKs2OTTIQ6rDsdHQB8wVaDT+kKapYtzLtkp2xU6eDOU0
MEf2alBp+vLizKNLqnxnOBNA59FLgPPDjr0WBs2zSQgckee9jrIAMpcjiEhRlKVy7ht4WkrvCv/I
rb5ZtwDdycJGCl9IYVmO9UtjD9/3EWhuWkPORffQerTzm64IFHmOEWYvGV9KTZoUmePJvUieFabx
P0BJgncIOmfJMvWRMMrhgOWw50XNI+H4bZHKOHZnCzjdXGhPFPfShtqPVAFDgtDjr36/Nt+Tpd3y
eh8si+v6sD9x2l555Ti4EsJRp6omqy5BrlNfJm/At1Uh/d/nmsfrA96bt8WorAfmUwj86kXrfs5i
aEPxFpmHXdCVP3wcC5vamJZt2V+2nUFLD/UhAVOuR3vuJZL/ZXrsW3ZGUk3HJy5byVlVWz254JPN
l+3MLi2WUlLl1+/jY8GcKiI1lXVgzbr5LWdoo4AfAmLaxl6spINOolgwILQtyWF1xCEjbzvccQ04
Nt08jpuwpS7OqX84yc5+ZqS+5TwBp8dgbXtMQHlzZ2Axc9Ii81qOlt5AXl8duv0qozVLdKqztHu4
3cgHQAlO7RdyDkCB4mQv2WaUN5EwlA96JrkSVPsljkDILG6mSb/0NZDrO2fGRC5iWiXObqpNjUyG
8rGutxx7CzgR4HmJmN+OYi77mG4kmPmDO4ab04Tn5Ma70SSQ4b0X5PvSCnX7d7QBM6RLjU1CkB74
HpXJ3GCaeAUrQym6i7BHZ+95/NxjtBYV+Uqf+N+QkDUdmUn6g6IaVrckUk8KSfbWEGVtZnL97Ds2
QqBbODLWh4+mhZ06LlGsKvjfR/0RIdWsEYe7wKIy1AhSiduRBOhSXWldhirBmjCCT6a29MeYUFKE
Dbtxqc9e5MW6MbTbRve0BMH5jrTjd3e44BxvoH8mtDEpCui0hQhLziqmor6PNLnBEGAt+cKzWDRj
ldwRELIhdJX76EMQDNBd3pUGyhqH/YA5dJ7TjdgX2sIpwyO8WU0SU6PuYgKVZVyr4FqIzmneTpKn
Tc52Enh22CAqB9TrIeJtPwX+pSYRx/hf9OA8iPh0RchAJUr66XbTiyu6N/kkteSfqNrTNP76V44P
BdE4vnW8FwBBhaaW3OEgV2jVgDCXbp1vNdj2+0veusxkDnjPFVYb+F943f6fqMdUY45ogLvU9pdj
NM7ETiDaWXMO8WVuX/QF66Vp2a2/9yoRjZhY5eywl5wMq48QVPH5PWsU6p3YGK8c2gAx7Nv0+k2l
nk4nkqzp08C9I8331Cc1Oqj/zzoAbDnaQTP9RAYCrViDgO3BQltqyILHCjrGl5Ji/yxW0x2ghLOG
Lp3vDukFzoEWQIQmW0RFcqN2bhY0nF5gOqzjSR8ZR10w/XlQljcYDnYruZeKTuJvLm6+GFIJW+CR
FgOqlJCHxGWVvS0TuZU0u1sKNF+T7H9MXyxpxDwLaXg3wPwazDfyzwpz0T9I9NvCPWZO2YHxUMux
Qm/P0XHrb5ekC6LiMKyWnTloEhqCiiXc3FDrT+05WvxOtz82nar24ff3gJNakmygOEDctLhuGxUg
7GEbycnV7Z6VbE3LaLgqYnhVnxIv7EIjubhl2KHLgeP9KDdtK0h5ZLzx5kkup6E7dGC/hZrXuW8I
omXbBpXd2oMAGDV8S17gRGeIk9CCw2xCE6x7vOrNv+XguIMBYCHkuYrV7xbGCOm4r5xrbtvaGgHv
1TYy8nOxPbH2+qKQUvaNrPFi3PU4ejgV6SuDvjuehXB4IeOR4y+NrELZ+z570zGDOqvliC+3Dura
TErJxqxY9xrwg5KXE8N4c0GLo4OKC5rMAIAONpQSySq63PQ25d3FBxYIDW+hdAQKbUzP7ojGQ6rO
GWevM6wrz6Op+Y4AFqTgI0shRv4+R79WV0jecu8RXckNPTcm9rKiK3IBfpw5UgRg+FSp90nB/wJg
7e1b333i9DwzKP4Bp+wdUoZI/Z8wcrftw2KAVxHvouZcKmgblN8q5j3P4+fj9sRWPICFAvFSdddL
FgjzSNvq6w8F/mO2Pq80jw74ZL/YQn8yQCSyOCLvVjziJgjuIa5psi9mork+c5fuTfLxPBPYT3R+
MyhAYLs88HTNHc1DUy7sJ/OFn6f4aGY5hcbFAAN0rKE00mFYb8KfC/RAsW9h06EGnZwZ7D0/mWS1
wa73N3rYPaY1+u1XjHeE6MSN0a2Y5UQTmrXwa3mdgLFw15St0PgacH4vMZG4qkSYLbFaLZlq5FJl
cz4JhE2StYaw4Gn8BBMFyp/Uurp40gbzADJkK1Z1SQWDP419Ul2AkUrb8TziFak6ZLVglL00Jkko
eIVCYS28P5e4qaXK9tnnkh6ldxdjaVoH3sycWL7Dg+9c4zF+m2wYca3vahi7z6BU3eWrqB9lV9LF
295KpfD/cl7rjbOA96IsFUgXSmYatDU+qLn+jQXbzZ3Tl0WVPDmwiE3PGWAGh0JHEap7E2YZNr2l
z/5umWJZqKn04morTe3P2gWBgMOlPCif6OfJLskj/FlARvcktsWEWnXCSzNgL+u9Re/9eKHm3VMh
ysTpBGXZ/M4CzAu6Q5D3m/CQBx4v7JNMFiHP9n7LkNnJNH+W+4UHKjcc6KIgthmhxk7HSuiQqtFC
SCuYzRCj0bL/dAcicSvSycYBhDZNb2zB0Ok2/8VRngMQlKmqcGeeTfP302aYtVIQq8Mijut4tUMq
BLUoj62Kl/2/E94uLgsxPcHp75lR7ifxQ0PzlBDwQGGKIqb5CAlmD3HL8JoAQwmx0HVBlpevBqUS
Vgctr8wiCf0Q0I6+SWgQ1EoshTH/PyqfeWe1h3sIkPoGu58E0NTPWriRnbT0O6LvGOr1dgn1GxEh
prkmkgz4p8XbLRR00/a9qoWJiKOucPadgoH1KUXW1umC0Z1gaXZCDnSnQbFV/GchadjROUmiAWrK
oI0XvAVA6626HaB69ecruwl01moRuYgAvk9menm5O/Gp/yo7tBrFOz0eqJ10tPiGUwXpp8Hzy/49
jkTJICKk7Nn/oEIb+XVV9FWwU6yVAd4rP2M2XIOxKRwYQSXQiY+4WhLfKhYH4ywlw+AdUijP4/Ck
Lf1aZzxYyeayeJyXZ7BrgIVOON5rmemfJBi8Nm7fJkTkYY4OSg2y+IAvc7mfDex58z8OzADqtObF
VEH7v3wKtj8r3IVMacYqEAXEiCSp9PMe7EcKJ5wdSsc4djCNy44V7LVKVR8+wVRM8YWXIE8PtyJR
cLikiSBc6PZp8q1rqXQZxiY1uDXjDQWFw1JNrkyDueQQdia9evtZfxikg1DPvrmdvX7A+zLMXlVz
fFMdx4udrzGQ6fVerZ/UVwqrOmJyYDZsJorHX77z4Lf1gDbfcJWBlovUr81tKey5Cfgztzd0kniY
qokzBi9az81sNYWuaW2XHI+vh3HhKzJq5KW0oKWe0GANkKxw0v0DKDHmAl1mx+ONHrXU4sJn5KVI
tPsMWVcv8KilWOfiay0RTdn9o1+mbQljg+fqX9iH498/FA1LMF5EtYv4avZ775j66wUhhr4V5fsT
DCtb2AvRtR7bjOdLwsu/xZieHqBx58gY8vu2X+6tFetzHVfWVXCmxwlJVjpjsyOsOg7TEa+Qtc9w
JOG3fA1vPTQYIGkjGtWxMtOG09s5tf7xmK0prQwgoR18ZoJEo91t1UNKkRL4ePcMPyt6kXTUbraH
TpZk58X/5gv+Z+BibIzDECS9pQxyTdcaXbFT9PY6G3fxOgMeEbJ27NnLW6HkZv2oCpSBOwpxm+1H
isVhpmjdb4WKqoQIFPoYBwUGG9HPdpqJVQPgl9oUjQ/VFrZhZL79qV29VgYQreVCe/bFsFYhthRw
Vqi53cROw7hcfkXdxfRj1wn0q7H5nsFxU6y+UO9hXbM5/TK9FsrHC3B7y+/Guw7ChMj0BQhYpJUB
dN/pLzopxchwdg4BMJ52VsRGNAX9hP8U7EzE/k5j8TQjL3EmjZyYsI+SfSpBFJITqNs2hEJmTf2E
60ik2ODjGkQ3LIgv1gGGs+NUmI6E6jTKyE5h7L9WhqOTG6R4IDjutNBMBg0TfsERTwX+LcXxKAJ6
OoMijmo9VxBYI6qM0AGUdqS23f4fNKJrP+d5Jd+DotWe6IR72G7VMvBR+tsDRDbT4mtLBxdy/U1H
mN3C0z3ySxUH8bd9JXGT2j9BCx+IQP36nujPX5LReRHYscqoO04SforALnbXF7h+K/D/yFQQV8x5
DVEaWnddHbRn5AWsSaOBwQ50kGVVjGxX/CIXB8YP0Osogq7Ey9nlwUJtc4rh5ulBVLSyrj/mcdmB
ZfFuwvYgMLbaJAyBgNoxKUASuw+4pjYp8ggyIdWawSvrAc4SDvmTk7YHn78t/XStZUPXIVqG4WdO
qVTIWVoUuPAAV/aNWT6WnXBReEChom4Nyuh5hPmvxShXq5wcyFhu94uD4D9Z2qcYFTLjXJGLF2JH
Wahi0ygFQ88JEiOK3CI/7MSAo+hivIHoQW8igipmNhHZ86y9Ec5MX4BJbEmiKhhijWhYSwbAKIm7
XQZ9q90iRF/3HT6gvpXo8uJe3n05mkTN60wmOg9Do5q/1oPNJMiUIENVtbKTQxgZsCE4gzEIyJSs
xJfHIjWqKuQT/POFp6N3cdWTAMIQn9ldLkgPm3/QQcSb1HdzFPCsfBudVCIMMKDVr6Ll8kzLq89d
Q6Cv1p4Pi0406ADDjnpQQ3c476sGYyKNgrfSEq74txRsQaBNHkzPvxrGzxGDLHyOxDCulke3+HkO
b792i6luSrA4MgKYkwKsW8m0z3hyNCUmm4RdSWu1qKRjO2zsarB2jczAkF9TcsbhySeUVm9mA/cq
FY//b9XLulvQiqmDhqK5SVajPnwzUcMtLri5IeWi7WZu/F4FZe81JcK8hWW0SwLVFUUNs10QwsTj
czbi466zvoUuHEiEyrSrfT8X7Juj4a9Ll20BuCgUDkOYrrBw/sTOsAvmyIBbUelxVV24kV+41qVK
SaxBLzQu6LUHxw6NyYawJFCLhdEpypqtFfwWZuPgeWK/mua2jdKBlJDKijBFcLjo4oGzWomcH17A
LDK4YtnhlLaZld+FzbR5LgTbwp7JkSyNDpOcdMOZrcS11hvT9I/D4Qw5jmJB6Pwp7enJqCHnrEsY
cZonMfYwkzqhheEzy+GdHQTdQ9x75xUSnV8uGu+874LzmroScd75GkrpisF3rPDur29bClebczvW
yeZcxyWmBeMcpDEuUjgI7kCLYBzmacq+qnHrpwPgxWNHlehHtGHQBozmYjRUYDbLO50AnRDZj6vm
Q/etdV0v5462Igypxm4kovR9ND/uUHFVG4UkeSHkQytzDJoiQThUdhhEBMyYHUCF06NHd2Bpp7kJ
3c+bdQL62ey0zaBP9qGgW9fMlkm44CScf4+EoJbcBj1HyaOO7I6cpARBHwQZVlK9u0nqb/6cXPEQ
9s3lSiFsM8CdO/CCq5t2h8rIryX9Kw31WhInBhDnjYMtIph4B0HwkPHf/WJAQ4rRNcB09aI0uYDd
l6Y5pPeSxzc4eXuBLt0hH96/IMS1eI9xotWpCbxnZxmtYm8qDKJ0GDYmD33qVdRuK1VERVQO/V2N
7hbSfELRrE70zVnbCLAZVjByNDi3E0qNw19IpsuRRNljb163a12tStz3Oz8K+qE6XdhesiOMgg+K
WVlqfXJpYrL2cm04GPgJ4Y9T93dcUgpJo3sczkWRM0h8BAVkT5unJHHg9NbYKU//sbmWtmZYouWq
99Rl13HLqSWbaosjgfCFg+xEvkgp+iUiIGtloY4HMim0AMG4ul8BDDWG2cdNHcqhqnvpU4XUpf6f
9aN4j7DK+6StRZrutQQYDpfnG/97dNIp/rzhUFGYDpCmC34ll+XShUjJaH88ZDIfoHVh9Zg7Xh0o
C0Pp+vC3ANQ+df0Z/XG8LwOVAuP/VWr0Yn+9hSokYFIYp41XjVd1BQCzlD+2SioYF4oW/+s9iOc/
p6yffUC/kFv9qXnX6FF5XE1V924HJTd74cmCzTXvHnHrPVZtkjyPknZvgpXqO2wcaJOWmiYNVbAN
pHAUvyRdn/lCY6FX+QPlq6NpAfRPDjOSK487GiZ5a5W2hOahYVDvqEJLxh/mXm1eRiqaep7ECDtE
AKNi/u7taGbR9MGV18lBcDWEbxJXzAJSqKVx/skSUw86B/owBitOzoIzn3briex8sXQ+t4pkKJQt
DZX6HUt38yQVySOgtFcEONLxSLXIsg8QprheSYqg9HuHjhzgJMaVs89M/A4Zl5IhNyrPHpsQOtiT
xCO5boKhkPCy/bAG3DUQ51jE8eCAQztRsRIH4QMDVefgmeoqz6lo/I3PQTrokaB7Zt0nQmG6SLCP
12N9wAJFCPwAiwJ+aV/3PpeeQOd91Zu/Vv4kt+dvoC2gxWqSkHPrLuHPni5Vr8j+F/Cq3io3x828
+sUKAPxO+wtpgfqUE+JBhZ1YBxmySGoBx20kllISsEZk6oIBv8A1oddx9faRfmSa1iCvcrjosEB8
ExQ3PMjKk5u05SmBMCS7ZEVSU9OVRsTLTdR840C4+CJ8V5fyENd7+KtXaIxn0WMR+g5bdsSmW+8X
nPnKTB332/jrGaCOr9Cve1FqFTYpeKg1d+AlzmY8cjTUTGbWzCRlxSNl4NpRY6NZMSa14pYQ/mFZ
3kCpSSvzi9CqDAGPZW8o2xHGE1G8pABikwty/JEMkVOYHTinC4YM1P7T50Vp8B7CYQMjBCixp5vT
8+zDI7LsRoz9BPbfbzvaHXAamvLF23DwAw9mijZYyyctS5UfxrF7q8luQvTZA4wdI4cSsIizau8F
E9z3qMjKPfRnTnMDTyTd+Y2DhZ/OtPZ1hgG7BvWSCstBLD/8LlDxZ8r4Gz2hDaV1UTwVpx8WbW2z
eOSBHeKNMXceWn0k0C6HPvH8n4Y/N1SchP3oV0rVd9GeWGjmW/7CP1qyzr37WlB+rMOs3J70wgEn
c8+AGNe9yH1KCTaRx3NAhioqvX6SPcYfvOy1fGoYAGm0vjnp3RjPLnTAzNloqPQUkind3biLh6lO
ugs+hB4x1F70hsK5DLdXjXFZOF2qiH+GGd6XwnRCguvfXlsoE8oc9Rmh46HHJ89hsBOgP6f2hRiN
NCrz5MvM2GW9fbmP9uRKmBAW0VzQqZ7DTcOeHbUO/eMB3hN12V3XO04OALqnkVa9pS0VpA4ZQcHy
HtWgAzoJUXdk5+NaSNU7BoGhxfJnOVBAbllup1f7+08UVQ7tyWmgQ7+1yZ0TCzB7QAFW269zGR5r
kQfMkExF3OYREU0m7DeU0y2t5NsZ0PIY8ZX4gvu4bq0/IU1BB3PygG0r2Rl5YOH3n2Gev+q90SdS
3ik24L46CmTfNyHD8w/O6odjYmEoRnUc1i8o+ELnAygy5RfnbJHvUZt/l0qNYgd9tih0klXsfPSo
WLoIFnzdEKfiAfpSnsLWWITHO/t29/nSrFlbnRJVUjLMx6Jy2dvxkJU/BSC+XPMmMYF3banWwNs6
UNK4Bdfrp9t8jCedyj6vtk7IuL2jcm/RTlsQb0ik7BNuAcj+i5Ua1+Z2Gbzlbl0diXyGbdPhouHT
Ae9IJMQu1jD94Ogq2thyYxrFTUulZUzUX60YR0+rYZOCvq+uJSwiN0X1nQHhi2sMe/5NzwTcbKfo
8WAqgL/Ep/cYmTGv2vVKaBM5KmsNOzQZN7PJxaJqFvTUGwC+w52JV6149CXekvRjoW1qav0DEsXK
apHR0VizWOXjhkGW/QeVMN2mZihMRC2NqxIrq9Mr+U7LS2rwxWq+rNj4YHJKRpll7iH2/XdWyW4+
WkmFTc0DeRSKqI68NIS2C6Q6XtlXzvDvkFTxfBTj+QxBPhpnK3bjA619So2EkV2Ow2on2wSHGgO/
g5q5OpnKw65uOzPSOEbA88UIhHmLXcNT7kHDEE8+vqmMKsvS8MPlvSJvImHeoU7asq0VR/kMOvXS
/ftXEUfSgIn6+9Frd+cu35hA5rbgk04AsR9+kPQI5TGvgVEZ8uumTHaeenDT8HnzpJXUtPfsD6Eh
WO35ZYRQovU1eaT4b4GzIqmfMJAESMu+JEQ/fxnf1LzZLAnN6YlmreqvUFiKBg6lwUziLaJNc9IE
pZrTOkwciL5qTbZjXnFu9fN5Sm1apNoWvF6tCCNFmUwx1zQ0IlAlYE7V7SJ98At67mtKQM9kP2Dm
8/0LG7XM7QIy4ffRIM+2EOtfwAUHdEBC4SkgiaJqM0XufXRgimJ7/0MBMVijy5caIGcH/fF+/IDW
mhe7wq5U5h3BFYho0mDojC5oKjrRGXw7g6iFyn5lVMXh0ujSUmApxGJ7XYUVpuc/W81HvihqiYx6
QVxLPCfvdGNxP6gGczXml7RJytR54ldx5pipRx1lS3q/fpD80mvfURE59zu4B3x8TK3xF4d70lLx
wRs+2BoW2hCq9xbwhXBqeIvwI3QWboy95s3n2L7unDRpSXEiTEJtGm9ZZBM1lgXIxxT6b6yXwbBb
JPGvLZbZbuPf/+Fut7PS35YSwM7yjUcbVau+CvhGsqdtAL8+3rL8E1TMeWdXQXwbWEcvFXRot5Iu
PkzTQ3lycMgdTv0Xx4LQlin3sEGYtR3AAwhTjaU4jFg4L7vTu/qzBLZ8Xr+mYSDi1hbMfufFdBC3
KfwRC/09EY0abLX5gW9t3675dYhv0lEC7hBrYfcxRo6dU5IngHWU3GQwf5i5QKMWeyUVfUuYDIaZ
Z+a7yXT8K3S4lUzMhbcGHaAoj9CI1LAIFMO9qFPEQ0Fa0/3cZ+/rFxQZ0QBNV9MsY7LkvqDD/Em/
JR4GzWEJt2NaGJ0gFAZGQwPzQLtFofiLbpZYd6SUclvsyhkefW346ZdVfeNISSKKW8XAj+87H/mm
v6TFQGpldGlLEVV1ZwlQBq2Jj1iD77T5Bcbeqxc+Jl9bCvbgVuPdinSutN2yHisIBci8CiB8LHvG
uvHeQnxdlC++pzKlyeUme8xdelGasPmDwjlT+Rpxany7aX5yQ0h7r3yldFhvOlxrl5LRyHezcVGv
ItPZVKMpGGmAAwgofpZNj0pfcM2Ux2rbseePIlJgGWjWMpjhdcjXfG+Smanq7U/NekQJGkVrRRbW
76TJ7WOD3flYM8kjrES606Esp19KKFnV3YShuxjq3/vTNd1kPyHpr1RxctVkmGyObMcRPRwF0YKE
PElamIrd5O1VvSDjunYpwsgBcxBu0BtIRklROHYKycTj00p/L+y/wYeP38WVqY1kE2NwvxyzGhp4
FuOpGKBiqiSqU+fJ49VYfyItJTldMRdkedLeIw7iZaZwV+zBwm0FaVMQnB2vX/FK0a6vA7l8WnCj
1vPah3MUV72qmKFKmhiD0FiuwesmJLjfppYWoOY6hQHkheMEoDKzmYF136HUvJ7FzXNqiJVD+oU3
Jg1GX3efgtCMHJZXgzD1YkayR3IoM/B6MO5AmbG9GXh1gD6+k+fv7tkrY7ucKT/7qPVb7q0eA4Sj
S1LvKQHUrwyPRRxn/pRdEZ/X999XJ4BbmtLBZtma4YwGiUUy8D96XT4YwED0Qg8mEnVyABcNt08M
ZPJm5rdbC9b5+JrMRStL5etG3YQlFaf+gR4Zddd0h4d8BDkFt6EcuN16P/0m9YZSqyUbXYX1X9bD
Qhr50r54UG9XCUlLQ87DEJoT/6/ul4/f2ZJHctYys2L/yAzTfPMuUVbO+XOmWld10hJbpoBgl+aE
Iwkzq2b8pvdSp/dgnfemd9cVQaxv6v8N0cAHi1+eybgaUbobfT1BSiSI1Ie3WcPZWsk+7YTZPvLJ
MK8XjXaI/rEkXKlJNy6WS394zgdrjl4QR3STpN62pC9hsqFXyN20LOI5ddrls5e6msPhH8+g6z+t
XPKZo0UirzGaI7TMVxmo37EBQ6mg29PAd9uONN+OLBvFBH26Hunw+QQzSRMY3RPdUYfYhwElnCSJ
DMS0mqbyLs1TeAv8FLFrKK9sAy7NCEJvdE+H14eDVWhA5d5PXvZ6nTISUmgmsbjbrYDI04sZZgx7
M3QF9sAOLOjJBhdLl5ugfWtzKKKYwzZUkEsSZA5SfcI4jMnNTo+lY65wN11M2FJJc7D1dxBm2b6L
tNS1bFR2j1kkw8gXxV2fN36BfIK4lEC7/szLvRnSn7SNgsfLpvsCSX2sYHiPsHk24pNJSbFJQB1e
tkz5MBgTT6HiZgB5H1bnM/A1veIkieBEbdAXoKpg+p76VwMZy9a7+V54fwyDA5oiWouowQ7SeXL0
yes7XP09B4PtmssK+nclaWSwv4raF3KGio5KMegF2XLjd48W+6+5dZSbVMIcRN8FE3AiK49LATpz
dVJ/gWJHToN+lI+ay39Z06Cw/DrcyTeS8/kTcfvoa5tU+HiX6YGmp6kngbHmwQq1oL0+CS/TjXfT
ZYTlk8jIEkUN9ctNh3iQWqniDgAabWhgAlTbnD5Qe3I8VAmytXOgI0Vz5V4Kc2SkNTALzl3v4cyv
GWt1Z19nN7PpsBqeCXx2y1e3m2Qs5GI6AHpVH6WQlSK7+jvD083LqVOQQsSTflHF3zfUAAYbwrv1
0PkTS8rglK7xPTy90BquXR18/q7OlEcFIsS1pff6bvoyIR7JKCl5OERTA7w1stJYUnXb79ZVa6Mk
jsB3ZpuWTj/LHkMMj11sPX8Qt2fhTG3fSqhb36qDhNw4M5IOMR9bo9ovSr6vNhyg0Q5bEeiI6IC6
f//ge0gRWNkl2EYwW1URXYPx0NMsSzqLlxCleXtWtpq5F8xz17NeuHGfIdbXMkCLCij9/Ji6nqpG
sfImGfX4lTgCW2BtpKvMzABGA6dkn87x5dOqFii8WukUh/YL+js16QCFrpcDKSVwMPWt76Rnz9iG
NiK+CozcosmgO7J/UdVHqrTp2wYlESdRq6qFZEFJPrpWwr2ccFCDlArQTZIEX7jxP8GmYaHlU5f7
/kol3LBe/U460EnXL8BF8cBhSE+pbk1FUTZsgT3gdmhKeVsw0wSjONSa1FDykXEUPCSuTyFFKF4b
0mvYaKD39h8p2Uk5j4y2JpexbMVTe54+RTaRuTgzA3l58JIYde4Wbcl26bmRSGiIlHyxhjsQSVPg
tT8pIOEgMwTgtYqcb0dB7a2AvfaLO2rOFcr3hadVQ4v4bCGOB2GhWwsGETrKHfNRy8OIjUyb/uUT
qaDkl0gY0tT3MG6cLC4zNabs7kTyWMXTQMjnExOHopcs4/EV1BxpiBGuELJpiJyFLfLtafJThsrO
MSQqgS7VOAHaWAxHYgdohhWh0PH3HsbF66WXlVv6VCDxhl88JZwkzGAnokJ1UfpEwaLF3venM+Co
WcRtfmR+i+p3ErJ9skrWULKsgwYf26Evj3JN3eJ1x5RyUwTXfrDBzNSuBgYCcxYDdT09RXdNqrlU
BFqi9K/0NuNJMy69WbOzd8CFWoyeFU7276N+UoM0KWbsbJrZLBOgeOGNCoW5yEuEIS7ftWyYo1H+
4/Own3rcWLgXVDIRmOUSxorIyRLIa5N13Q57Yo2cOLdC6l1xMmy1cUdCkXDX55fX7InlpTi0chgK
6pTSZ3H/lE442U5DqXsuMS+ENxQUcW4ZUoBJtEXon4l1A9s5168A/3122ucl4+hqFL5vWsoB1mYL
LbKN84HSau2yctdYqv2KQSp5NWE9VP8RaUhqd03rls5y+s8Z+IWnqp+35tAg80ctaXMAKMfrtsI0
us5TPcSG8oWPpaCRN+6kH+c1lx1NGSD8KdSbstn9HByH3JVvYESAd5916h8Zsm0c9t4qW6ohuReW
OCcbke4OuQ1AZiuc9vJTP/drI/8m9mpz2g3sYBSRK6LUIh3CGLDE/29JRppG0E4KHRCLvCYGdIfU
Zam+Y0A9HbQO9E6ihQXy1vrqnxBqOkpmC6qzbDJkMDlQh0cbZOb7S7Ls2nz2Z+zLuunI0v7gk7SC
gKgzLJ3Ipsx4e+3TtPibTnmN/lJ5KWyz3abHaJKwUU1ppx3NRoo7qdCRiMp2nO2K0Q8s95jvkvui
jxEpgnZVBlMroDn/cV7lsjSGNEhFixtnMma6847Y3foH9zbWNXcAS9ZBmaYXyeJr3uGpUyQZzhJN
euWkVyZ3zChtMX59iwEHLKD9Xc9Gyx4/+HMKBbjNB9z6/+eo1bxbWgisTvW0/C7gXhcWzSFvtKcg
vsBoLhkcW8ymPq6ccCvkS3NnoLSupRJMNMGq98B4tTSN5TzJHQRoHCT/p5/+jNpeu8eajKGsuu4U
mL+UhT4erADgy6rGpEGrjh/KNJxi1IUt4ti94W6uHG85SsTqHk+iwAhZEeLOIaj5ZlLB2tMuEjwX
0vaOXc52rMG8nSRG3Qqt5QUL9rEUShmwA+QlhLlb/AeyU+JMGpMnzJfWpdBwIAguu2RFIm/SsjPl
Nrg/DEpn1nLmGO8Es7vNPOMKChU26slVwIC7rHppG272RS1k78hFwvfBJ4b3zylJ/xzap/iMvUC9
IMrfwU/jLAi/NrC7QVuw5KEo9itIKltjBoINCxhGlMhWyPOapTqaWac0B/S9SavlDC9eq2FpjbqB
hQAPspleQtIc/UdkY166bT4Cdx4hKdg09UFP0vJEjpQKFvSZJFzPetyjCvjYXANUyaB9BblVAcDe
ykjzuFja38BDlFgIjcw8QI7+K7bNg5o4mpZZqOMSgie3TxLgvNoGLyo08fFD7QLMnDPk02rL6mMc
Et1p3MhzKq4BwdomVwk5D+9rvxGeVA42wp5M0F4Dtg88+XprqaZ8/45r+yWDEzo+tq8GpIuTu0jS
vK+gFM98VZ1xAEx3kk6N6LZBRtCOu2P6Bvw9btCm65QuTPHL3fLfqtIoxRQ29jAnhnFJsD/gxTPX
fg0JT3mkJtOnfONreV7yfvJiymJVipO1Y/pUlm1otx31l8MeVyp2+XKg1ZqrfLytuS/8rsN+XVn3
4SRPKj2KqnYCq7wVuhJd7BzxfUK/jQSOdlgYu6TLtvBZZ9fYneQLDicxINKT2cZdjKKGPsrApnIQ
SvCVQEF3splXXLWTJyr6IJnt3C8arIUAsWfxgy2NI0PNr/jECJM8IJbNM4a2EAuUSBIzxubKQYIc
bmJIzS8Rh0bmBPApBkxTNK82xoxiM/5Wpm210GR5AApvnJLLATaLn8DfoLvW8p4g5RNnU3dEs2QZ
WTwAHQfg7MSMlNJq2JILNZBp2dLtlRtApdp8o2UGXNhO1Zw0ImpOVYPG/wW66sNRwoUx7ku4LCtO
3F1HbUU3bNzO7Lx1EhaK5eFGMld5LoELPeNhYLP0NnYMUmyaOxajp2vqtfsO+gsjtc1dzsG5YvxX
eCWFV8IIqOZw1dt3SKzSRkWNdOS3LdTLMy8j0TBYnlsGeR6aywYDZkBAinc551Sy3WH+Lhwh37ju
GvUQObuY2eQFahXachrhh/yZlib1HHDGqIuDzmbIdHP6NDz0zb64UNrTUqW3Jsh0teLeICXCE7zu
KO5UcTpENavEiPH5uGmQt2hQjHTD5CQ7UoyLhjHqWT0TPgKEh/HnukBh2Nnkgg5o8va4sPe63le0
3S+vKg8buUlPdL/oqKGpXblwSm3M+nh8U12PKQfCmysAUcjsxwXy2ehDt4mUrK2bc4+q/KfSHvNP
hMWzmzGba6zVwprPGMYwy/E+5tcah+6DL0t7xl0UKmhBoipWROTgK0f2w4OoqRDnSejnRHfqXBkp
wv5eqHbfnYI7WSYH6vjYlLKTvhXhOskfqk5yNnTXdCmwGVuq7LDTdh867mz+IRzk/vqgjvl0mJuk
8u4GfrbhaszsZZ7RoXYl7wHu3iOiNMz/PdD4Rdro+Q4IQW4M7zbfzeWwjcXNuGjc2lUfi09Q2fPu
fAa2QVQuA7b3blf/eXGKi93p9VoQIZJOdRY8hPHquQd3Lpq8DYX4y2aIFwpBn34OJpHd6oEiMv6y
T3uIQD+mWQRi3jAQbmI91cSyLPuDqB7BctnKXAEVDguURudjcop2nqzjezMj4AVizGIPj2Sr7EFg
DDkoKuKkWBbtYzpId0SP//t3ym3K9TNK4Ak2tJ6FGM5W453mCCO6NvMcmYVO4LIdyxNLpMY/SPaP
oGDGJyx5D6umJhzbAO7f+Yj+0ePcD4P1qLjucC8Gv87S0w1AZ4MqKvIxjne612R2JAI3VYt3/DaA
hS6O6SYI/ye5ZUdHxzfiaJC4qXLiLX2QwCtg06BXCJRA6S/GULUFz8KUe6N33EES7zGDP76sVioo
8LRe6sTGX/vARwLzXTi7WCK9Nlm3NVThqETcwmcnSvYUHTIAetbTUAoBOzcCBFH0czDLY/Y8bfQ4
GnfCW7oUp9MON4DJgtcDGAL3tz86IOnHBf70pZ/WGIQg8uJIWlATJz7GTAgzarTU61HCk1l+d/DE
XOyzarDZfX2kw4Xm/6+Rctv5XHqlBVvAQkeG0AxEiOQJhXZAnbwusRWeKnxDU8LxZbr//+t6eFsh
FcoYu9XL7ekD7aYnSgIp8ZuuD6nL9xn1YG2epBeucM/GRnRtIodjxxlB1EbGBLp2c4hEUqqaA8zb
Bndr7o3H2uXRDM3mabHxZxMUK+KcOoAPYzrM3nKYYX/ELmryzWMGQb1qys2SOJ+bIQQTCDG5AIX1
xhLT7nFZpkJr2W4hiCEsfcwAnZnvGVdc4L55Y23dALtpv4mt2zMnMnVCW9aK0aKbIzqCcrv4A7Fh
90NfrsmVzIxIlq/OtylhUqU6ZCh1D7vaD1tF0LOS9PpbPBz/d0y+QbeQhAJF0/9eUA7qZEMjbSZC
uRf4w5vxNHreSwoQ2VMfBZpIVAj3ogpPJcmAUhnpmyDiD0qVkZyYRpaW1SbVUnhSS3BNWrFD7aul
vQ4HX3tEIkJ1SBy2jWaW372CkpuP4NFv7AbCDXca3FoI/y8gwRPVlf2vfvBJgerye464l+93sbDn
vcIg1OVPlF6eNdIym9TvaKHUPI2K9KAnCBNpQu2WhIZfdf5XJPp7NUDRmuW/w2oGEUknoryjSFOY
LWEm60O0GcsmjBCsUFSok6zAFe7j60ilZOrz+/joBxKLyT6SYEaFRg6l/oI1ImaZalY5Rcp0ax5g
DOTmTGsh14INItvSj9kh2BqRfzgAlKq9KKkl20277aP3jZVPuf5UUqFGc9Y5ZNU6R6NkfjgveUug
zEJ6v78qcdgDUZWa+JMzFaFfIpu79m70Spr7XAv7pM6VzSksHWAPabElkEf4tmuzKmlIrBnMxDuG
vhmjP4jTdJTMobKOl9FWfWvY6og1PZqLmbJMaxDjSbGHqVz3QfgOVLv8/PpZXCWaYZEP8ID3j3Gs
K8bqJLhx8vkPMHDsF5lqwspoL/OM3NEcfNthmWdA5z4xSBz9DeBQdlTVd9GVryckbexN8hNvf9Yg
6Lb5k6b+uDV/2QheJvZSJtJgIAZEhyPNavhV3CGTj97OdMg9xLzv0PB0CDV/P8HUiZ6TXBcfJICV
1mn1tBWDDf7qjv4N8t2dG/psZyf47i9C4UsEIutnusPaPcfq5IZFAl03tTPk0Mw3yChqGXsCXH0k
xyUCbBz8Z9mXpUO67nnP/7LJ9kYB26GtEIL/oYOkB4PeiU3fa6VewdV6SdWc+tzSndCVu5gftSvc
F16bSqoL6Me6qU7IxkqhXflDn1rBXj474Brvgbj8YVz5USjTFILpezi1+90R9Dj+hWKx4Cu3Mf5G
H+SRTGQThkmepgkActCFJc4BbrUdWleD3ILTV4e9I+doAkCrz7SKt36WA7nU0xkI8X9GR+YzCEnA
CvlUPx82Bdug/zui8I38+luV+8YR+xqzOj3nv14g1RHvTl2GfgJYVHbcyMlffPDTbFocjQni5QkJ
Tql5CcEU+sasuwqrm00pSofVBdSQXRffXSjmCEwX8g/NgK5AjkklcFeS/xSKBCJPqnsA9aWmBdev
x19GxYaZMSKEtSmlQ2hxF4+o8xcbdM/zj8o3gvGFp/stjtmFwlZPRfVPYXpLUoaKMrYGpk85A/Uy
8O90dtnGkA2DjrEwbZ0eQOZ00fzTRirAeMeFdDSM0LrZ6wD5chHTikxOpLNgZHonFZvNFmyZNUrh
OIxFjUQaPrUP7Vq2AVFo2jlfqikNVW+sWT/x3zwKV94mdJ3DokhhTBRZwZXVcdYzTfvJ75ntmf6z
qqNOJcXDQ9AWJuvqUbCvNCfxgypGxVKjxVqIWmFNI/4FtCUhA+ftvvP182R/1nm3lJMFndepGKJk
F29uIwl1fa68rXSKK+B8JSkPrH8KfYPV+Su41gT2sjNBg8fo6O9CxiF7oPPt6bEzqYPXwnJMIexh
AW31gQWmKUQbfX4WBJE2jG+qGPIIt3RR+H3KxTcdVKVWIUqbUPgOLFrU/V9bmtveXFnXi8gAAWKN
uq8RMb90uDOE2tAuyOfC6v8YBi0GLxcJljl9K7fc8WubRn9MadQWMF9Jrv26M1L5vGOHltje4HIU
MlhAtlh2t9U3OKhy1HkV562AGOV7nYt6V3fbZ/qBxeGgnDusIHcsN+xaqYMuYWccbO+bsVhx/61m
pCzgF8Cu9if67WUlhPMTtb5nwroCYe/j2ZrfvhhLv/yEoKJD20cYEMmDqX2v1oHWXrL/RX0pR0Ae
5ikOqk87FdMdfz7j8gRFcf7+LgEZLlebGAW6JgBhlzThqGUGJGhmscHnTHndaAuR0Zo6gJRqJATM
2Cx5IZAmjCWt2PXkbrbCJ2xSw9mT8azNnt7Q8Ht7G9pcND4YMjHzYCgxk4LGap8vvEg+i//Td0HR
jY9E/NKh38E9rNU0kwFdAVtgiVCKcHjHua7LIFpPCo2zlkreT5yKaK2wNJBc/sl3CRocB5UIapuz
iLczPaAugfqzLSN6+aGHPfDo60KELmNSuMv3RuHbtJDGUrdbKSMVOPX60eSw4+htwHq6NfudUUzJ
MJodGRFNGOxV/JdzuU0QBgg+FGi3Ue2zoqPl3SyGpojmb2P2O47nKC73eIAB2H2ZurJSgpGZx1jE
IozjnhJn9ColutX5le4HAEnD+u7i97xJkNJuUaabVObCBeFwl9rLiBLVJfXsP2whrhXJB4yPwIgg
cosT3ukehra/XTvPgvgC+StCda/YQbk2UCKD4//TbzzC20M6ssN1FkqnvlGFWCDvpYluXXe4yJnG
/efefqCGqPn9XmBJuwagLmpkgZNGTrUG1b0OYeFHkGHqbgqrCSuKCfMV2bEutbaCnogmE4ODSw4A
Dfbv8xApElFuDsGOZmEGdW0B1OEY1KKHdrIXubQ0gJ0+okzUqkzKhhDPfe2B862UgyS51p13ABTW
IkCkzDJy77i7HN6yetiWEJLVv8ys4BpJ3DXvMSYQPMfVLKWpmKI6YaSLZRmPmN5I5+gsw7RQGXP3
zt4ma0sNk/TMYXhHrpO5MuYwCg4W/RVZz+lBbmzuCMCTS6fT4gyh24bU1o0+c4noDNkcobj9NIqq
ikK1gLTHiYLDwV7os9ijCG1byqXVTs4k9hObVEECCHVD2Y1c+/3TQ1pHfM4yTUO0oG5MU6G5NaFF
prgqgelGDXYBKnw2cHxEh5IopJ9/mwrlWypOskVdjSi4xy85z81ihXOKWLnkPgdZLofJot2faZC5
tfCfFSxPxCxEyfvYjL6QkfHpTUtrkhL78M975uAeHvKpM/5Bg+m5u8npwbttPiEdxIAqOUR5MZXx
n41mnEw+Vt3rYb/ixfO4TtetYfU4LRgvcF3LiFzkRBXf+alFTmsd4ITR2+Vk9g1WDLbs2yH0jC+h
dSdtU4lkeHEdNIFI8cq44rOYDjuh4p5VMGW3rnc9xNRy4NzHIGIvJT71RV63pq5lD2jPKQScln8Q
U0xfBmr4LB4CsBdznbdOSF1jyDLgttAd+iFWchiycXtXqw3OH9fPrs8O5lJkU7gG7f385VhtUXjX
S0Tnp6Ek/t9N3y0Vdmso5BOSBJyAagpbXMnIExKtUsNWPo2OO9o8T1V7QjWoOKoCN4VXJ21Dq+jY
P89L3pFlw9WDFgtdfuFLs3GpOEJN9dahei0IHMS/DqgpicKLmiaJtRr9byvZgIt0qbXCHtC6NaUM
rIYEgYbl0B2lw8dS60BNuPlR3nic3HeagxQYTBEqJCrQP5Wq1+HyJ5e9Kp7phltOORWH8RYIv63m
rdCDMIgPHT5WA7xrGIf+o+sDN13GfS8M77kqRFmH0gruuIshdjXtUVbfaRdLKDPT8z9qMaudQIbB
7aP0lGM/DQN0Yp+GEKXFevzpXxQ/D8fcgXufRpJnnzsYLzNphnsyY/4LgsQ8GvI13tPWoxgnU/jD
4lvV7TKJzGESxlLlse8/s1VzPePTWMrWU374tgX9m1QqDkbwmQ5Fq3n+D0K1aH9sV+OXBeXxvRQs
GdLK4qIfu7+dzQuvh1wqRfc53mAwA5Ceuln7l9OI7i0v3O1QRLsBFupcK6U7zQUofFlE9HM/3piN
9Oi7NeBasaXOe45gIolaRCMAbKj2IDNugEOFbJnT6140Tgop+hdFmXmaJT0i2r41r0g9eWsaU7gd
y5MR/5383UIUHNc4aE+oN8CJBg9BQWQCKt38OVRE+OzKQL+hk8qADHh32ey+ST2qwyKPlEUefOY5
xKErtfsW+ieNLxMsFv+ggh8twdp6oO03WaboeI4AQNydAqwc3/GiTiKzVhqQUrxOEsVOD9Bzg2lY
Nsajznxt9FCKe0U2LXYHx4fQOh7KiZhX0/40YJ8Ons2IeOzGxp1w3WwfMT84dGLgZf0o28v8Lovn
k2fZKNyK3LxL9/RKWsX+17k4bOt4WJKuFqCAsDFGh1j6f5O5mOWWG9XU0eI+8r+JXl09FGGZIZB9
QYJdihCW83G+dEYGQ1aJlh5h8HRBp4qPBDIEtW9yMZjgx3l3e95+3C/bR/U4qGNerpKxK/rW+1rz
XmJDDbTcNNDFlTC0KNL/HsFu9TVgDn2xFDb/SIdkJLCSC2xTzvqMwtvbIoP4MPbip2Ekis48iEcD
mb+Fedi2Dshl/3bW6q/O+rLqET2SWaHnFjOip/gO5QajhZn4QOrXNhHWRfa7gCHB3AH3g2CMW89Z
DkmW9EMiOYfzvrgaEMWroKBEHO60arricI5SB/4GUy2RgU1iByud7ApsSkrnfD/HgkpPtZReCqdv
jbl+4OpgJ7Vsz9bxssxOu/mqb7L1xlvtSaZmrYwjcqsW0Lyt7gdJ7Qon9JddDFlguTWAN5zc8bLE
5La06kLVVcIX8fQS9uNA77GuIWrrMeXVstBQIDQirKWnog8gQBvKGwVjWHdPS6+kWPI6MQZy4zcs
5LN4uVf30lIAnlOA1+xr9vUKcdgGVErep/IuiAUCk7WFq09A6dGowbuyf0RfKvRCWdef0BM3+bYr
Gw82SQ3u6dfkdFkdHLAtMPZFFcoJBVyvKqHejFYpR67Qpr3cI4XpKxPle+Dn/TzXdSPTNETTm6Kk
LR+SfM0BkrP5KwRlxQQ1j5xXiZ3JrxgmFw0Lm8rEZQSRJfr2z761LRGupYXb/73j75tD/6IjNGw1
DaI97EqX58I+sCnSUtzFOk86quCygUH9NduH6EL27iWh+ObLHCQ2UHK+TFDO3/k1KKCVDrA0R2YV
UNjpHYrtMJymQCW8tqTjzz2jhot5iOdgPscP+rR7inN4/qRhsVkH5WLMOZDbC/h4KKaJhsWoYjLp
JAOTvJbto4zvNhw1j6y4YwYKKOhQk4xsVN+sH8iG4kK3O7CkLSzG3DZ4EaPFqbMLPAp842YKn7rC
/xEqsRUHfIUzqckCfh8T6aKqo3naWdSktdnTecOTnthXSFqR1tAS+7GVRiWZDeQ3k3ex73Ai5318
kMdPb7aRfQnA+gaNzNhaIUIVkVABB0fV9ulIeEpkwsqg4X2BymK/tF+RhvUmtR4tYbCJywLCvoAJ
er9CJHfpO6Z2zJJmDxOLMJEUfm2KsM6IHVfHejxJQDdJPBGcPZxxBTSJ6UouDDmKGU5n9K+mX4Ib
yCTcDUWdlTsUN4ShMAiXEjVJMHkaP5wF+6V7Znf7EWujIUXcWymVctGk/UTLKHHLdduoPIRxBH/9
3fuXNB1xto1YNqdjQJzRBaTu+HEF8V2Iq011C8ZOKxduYkYigk+k/RalmxG08F376btV9rH5OVX1
ns/81ua3nMxk1xxqjpKIWqOzNMxPTYgjX0xeuh71IXrllNy3j9TB8nGgakCgwmigSKoDg5yk3kdB
rG5RBYYDFxZAtCKxkdfQghLH18jxzEvukhWqkLsXwtTpAy490qMbIF7DADs2gDD285/wFRUq+R8n
orQoV8JkOSXgZTx6xbsPQEhVT/6uMW/jpk9NKQm2+ztvmzPg6ZXqPRfiB4WWDvTGFF8KRefma64e
XYXLg83pgZul0s67LJcPhgfWTtlbtZH8/DtTNGqP5cLOCxLhXkg8AtbsUAGY7lm3XQaIqGE60YKj
p3Clvtu1NTnAf4dtsKnlDtkTk9aCfzsLFz0csDpQk80jbCFbHCEcKlsi5d1tUNFKgPQzo+4r3pdu
zu0F5H4T7mlF6g9YK3He76cs/PLsMJko1LH4M2YpPjIVgfyc3vyfdJS7QRu22Nvt1kXpzxXe9Qav
huuAvRJkQvK5nKLrAlFQUM5MPkrC43h1w82xC8/GrA9Z9LZScczWDDOc8noJZswM22Y5ObscrpD+
DC7BoybTx/TnQT/WYP1Qg0I51kzJcGBN6rHkgEFQyFtVvIY918QVy3hEhm5HyXM2H4ZWCFvs2Xz8
0hPD04m/md1+LiVSkxHDL2JlV9hAXR7DXCFMXUTBypk50FqpItWavWfLYowjyM3klmGZ0RVnk+W/
KNlQ6jfp9hrDnQFY5D574dCfaBUEEkmicGmPxoWADkO9a2rQXYOwdcY9xMZTxi/HwHpEjRJie3uA
FLAFuncT8w2GBLtqYZoQINJR1EcNEuxLn1LkndRnOVKmI/pcq/bjCevWJGaBLBIyZG+zXVF/FU2P
SD6b24rv2UaGq5Cc+3qFUG3XI+hPw1+ptWVyEA8b4lu2TwZu15AWHnp9nmZqDGqXaQVmf46za+3I
MkFV4Lfk+TfHb5qW8y7RJO/5RFAS2QBtZzmxob2QqJHwCgXHTGnW8FBc3gGqqxj0yxYFX6WxIsfd
vTj4xCwz1nGlEgJDfo367hcf8A+AQKSTbxDBMPzhAFufJ+/dFinrajCPamGjT9B36aIkCqmmyHG/
gd14Wo3KM5gfCwIynS5/YSlJ2ORQ+nvRrzAaoBVAEGd+3A8Ecrf35Cyiic+U+uiVStx1QmIHvSbB
fzXWs2VmEfh2G55GTNUPXy/ec+oab6WS+N6DeyqiwVaYVSMDD9LLw03iQ8b1cNw8enag4j1Ya+z8
PrwNhu/sgtrdEH2y0JsD7tk116e+65MGwA59XmNqV1Kotknsm6766ujgAAUqH9aVW/Yck5ygM2Ex
4XMSJvQdI2EV8CEJD4v6Jh9LDDwKkI34TO/TpMO5McbJgJTMLNjkfP2ZW3no3WpS+6MPekMjBuc5
VzXqDxXK/nxkoG6hkAVqXRtOzuYsIxgLJ29lH0fBXOiH6VlA8q60OvjiyqiWnYZXaQxSGEl1ErcL
D5qkr9pZiPBgpPR9IwzyFBcbeWtRAPRf12zqCy5jY1pxnjl6x9XCrLbdrmUI3Vm4x+5tmB8LDRPH
BOcLj9w7ri+Mf2COjIh8J7BiMcykt3t0y9icdjJoSgELhjoTTyZiwl0GSDVogSpN4IzSi6vDAncw
OmnIcBXfaIk7xB9ZvnByLo2CVWK1ZPRudTq3VQTSG6nFiWjfDBnVrJhsT0VxAnfY/xc7aEkMEBlP
ql1Z2DtiHAtIqJ2Ticm6Ii/wDD+zDDUQcu0l3B4cV7rbP4n4/L1a5goaEUupY+HSu+eCBDnhB7FL
eyIk7hMOQ6VREFUE31ckO+m8uEyaFnNpatUiBHWXxqm+yrFwPlLB/hP6DXgMD/FvYeCn5jmQfhDN
4OnFPaS6BW1vwXoiD4+3S8e/fWkoM1lIMeYX2tEX1LcJiwilyT1bJ++lTEe5FEURRebM0FCoD4db
wWfmhFyIGSchuJ+PodKIzuI7/TdjB82isSOS00k4miIzYMb2Axc2TvvMCOj4L8ruzTXhUusIDGP/
PRWWcZhhScRu9WdttF5SqH5/9XLnYQBRFaAw2EyqPZJI9LxEMIn23I3zSVmnKHbOCf7GrT0V8Ofc
zYCxde5nqX+l6kZI/ZkVG6o7VzieCL2+Lh41AQkyAoRXVsud/at45kccQUu/gm58WiCoNnoiXZD4
M1gMn5SJnr3u2EhhNQWs+QKNxskKPo3mWEjbpdIacQpyOJYFmkqXBIgWjXiQMC4LzDI2sb4P9+l0
y4/qBb3fxL6onM3FE0SDIsOjWpbl7M/kdke2LJUSm7n7esaYCky2Cz4A5FqebtRsEEL4ycEbv/MV
8yfgr9WDK3Xm6IEtU3Mx0m7vP2nsUSPm/2sgrO1aP+VhWN/EtCbyOet8wREgddtU4NW/7FFaGeUU
F6VuPrsjNEJoN2wKraLE30xxt5LBPi8M/7oTTSHZHSEn3JmD1Wfwr2TS5Wc6wHtpfqNtaQwqAxdU
DgjoYWOH24ZCWKGfDHLRv+Vq3LSqFw0wb4oBwVHeMoNsG0WvUsVu9KS/KFJaeKnJQnBAiA1SI/w2
m3VF2k/CL8OTOvlPzbhNppNwEpvdFcDe3oj0NGcztQENJXHYWGIGKeNkZ47CmHy9+5I4XEUh3Uwh
XHYz5y+DxlziGXnvO2WimusEoUfoynHP/EqcQytyTT3L2b5LrufDT7Z8bg6eojjIHyqC6+LZn9Hw
rll4fhxZCvWVJrzdincJqnO1uASg7+9Ef6q1p9xcVodJzoWYsvN7Be/ippKC5HuMtosNhA2mO1OX
R7gvG3rokx+FeCwa8Q8y7CEYnwcZYmGGWHyP+XQh6Nq4VctT/ivdiHvS7VYhPUJ/HdCwamgCoYMN
dKp2zkDPx+tzk7xRKynwkGlXxEmeYYOpuWBtP3lD0+BhW0aUfTDKy3SwQ52HSid+FscMmkzcl8nm
OnzB7JmgqdgUCeGX4g/ILQM6LctGcN0yOEoxdDdpwkJ6IlLl+DvbhePIomWmrMf3CMd3MZPhMZmV
+zZII/TxhIkJIPEEEL/D48SA0uehaI8l1ElnC7Zcj8qujrJKBuFRDhEarWz/dILVjluqJEu2zIum
/RjYLbRht5Zc9rQHVF56InLfz2Ebdg2djv+BXgk+TuyQSLW9FNvj+KiPgUalo+kOx6qNRlntMy5E
s9TcH0ld073433roFcGNbrlxV0CevnMzvvBkJP0XKMqITqxHNsG4RfQXkKmIiUgOpNgHp4Wqm/Ys
0zQdJLAa0tD1UJnJ8/8+ee/FLWEbGZt96NZOZzpEEKislP9KTsUP7EdExqfwpYJArnZoAhmmZaAP
4A3vAQYfUu8uM9Y9/bx3JK+7Odgly5gzon7XmFc1UXvz0seNBxMM4z0QrNiKXV3DHzMdsIq4U0rl
lo9mrKSE2TFOS2QxxqhjyJwmZ45XulJVrKI52QjDQcDiIzAPZKwoQPD4KOXDl9w9Bm77KnliqL1k
G0fHgcR3w79+8u4V8Sp0mQgzQ/TRruENu0fAOx7my9qhzpNl19KB2RqCDapNGqWPryCOFYU7fjEK
zgAZ09lgMzBZsWvtGCK8KK/Knx1hMMiRDYb3Tf+eG9dnFLe69wELnEUKOgaFPOS3EXrvN8huSieu
6os31X9WVCzjlNVXfo5QVnnCTB2iPGDXfGpGUUpgYU4oSNiLpgj+4BN9god9cb+6xMFNErbPNziD
CkrmEn3p9vNApMuk/ak4PxtsLUJc0STcLzr7C5zM/W63I9Bbe4Hitwr+zUk5s7SYTcoXc4tMqyXx
GLtDZCqUNWHlP6/2CANB80gaZfa0V9UAqYn8YdjK4bW0i/3RSPE97bz0TA7qbhqq5++Hfs1hYxkI
uCcbWlR74dpgl+Q+62odzQfy3+rONH3UYstipeCr2O0JZ8lD8cSorjTTNdYoDlS51YWw3IQf5P78
yP2gS0q1DPB2qSxE9Pfrq3zVwQLTdqjsXqTo61dIORpO81D+43D1Ebu7nOW8OqJV1pZ+9yJd8gI2
asOJJ2svYjmpuTtPu54k6mevV/NWoAkXotrjZw7XRkzz/aG3zFBF09vSzisDt+HzhtWvQFuk9U5J
UOWE/vFCh9UHO6CuUAsY2WPJWSMo3XrkSstY5DE+wOPvXfVJ81/LtzRVwZv4U/P6ZOkXHvN7V7gd
/exEt1atQIEZhNK1teFeXM+rVIktj/Z2gxLRdi2ViSwAi6Y255yo41vznNGqqHwUIoI4ygVtqM4I
tcC/QbA7617B7i3KO1T2cjkme8dvooMFYLGvUAgfXv45O4nwg2qhfbggxWmV8puM866vF2yg8h/c
Nz0bGFkmuz1oABgCy7qzq2SQRgUrNd5b7homPTHvF8y/V91VgZZwm8t5bE6WoOk8eLQq8owK6i6A
Un37CjhQVQZpqrSgP/ZK4Xr4KOvI+SuW49tOzR93H3WNcMnPuWHO8REie/8h+Uj3RJSvF/IfOEWg
AooPVd0dBqTHGqg3Fm2U1wvEiZDFoh+nv7DAWnvm08n8oU7HFKCtPNvFwr5C219uRnpoSdqonCDh
2aVYFGt5QqDE4HDgNnrRrARddYAKNzWvI+hVZsooARXJMzvMmrq5vf6pfC85oMao5hvRUgzsULA3
/EZOGpp3aJpI1vsM8rgdjgKMevJMj58IGvwTKa2ZRTQJ0kuRtUeHwnWKgzHkasOKmvpEjc6uV2uH
BbYTh8LS+2lYKDsGy0qDFEYc68z4ElY/uwEFDWJHEkSP9LqYXRyYz5ps+8JxDlJ424U5aKz/mHRC
TR+m/93o3b1l3cydhayT9rJMvViOp/QppgLY52AeooPv8tlYXNxici6VKT+lXi6zfd/SmieRHxS0
3MzxQgrdhN0boe7bkz6U/vt7PKaD7CqDLknkkq6s5Vat66LNLldfVMCbB7dxLWgwvTw8XLACbVuV
4zTojkcP5+P/5szlbbV9FEh2JUwug/LsP+BK/2j+sJAWP2nNttZVhRcchpiQMaWOrHbn1yXp7qTn
10qHmOy5EXZapBsoy8LSSN5wGhkyI1fXqOHajZ+U58ru5f6htj/xdMfEu1kTHN89f78or7yWpsQ2
Um4s8GZ2Jnr4WQota5alx8u01gw5/iDsnv9YNIzBCcZKU+PcwZqJVCtzbdY/Y5kZYtc92FCGLrap
4Rz2F5sizn98eLdwoLDDKXDLrXtquBwa0Rkc/4cs5wj7e2e6qnGz6BhzHkJVmqssvROwlBT2wvtg
5muH7zkie4ZIS7cHeP14q9rRZntouR8NuoAuw+6m8He6daLMjlGY384AfkGXNR2L4bslCpgvdoKl
p/zcuga1UJGcofTy5zIKcMzJ6f0Nkpp0lv8+h7o45ZjsSxZAlrvjF/GTNpnptUKDTEkthbjJheJx
ZLQUhT6psCI4H8mZIodHvBFdSUhsNMe2RNlWLa6HRHW2NMKi7Oc+Li4ddTRAiG5jTtEljQnn8mm7
HmYBoAf802W5wczsH8RzKDeMPbWgiyCjP/EGBB4shrN2AYXiLNLjT1PesPBHDIPQEHG3CrFA+okw
UjSel8d9XTiGa3EtjNIO0esnZcEQmgYnAvo5ed67EunOqP7+F/eeCSryiz000zFtROrvEJPrj57i
B4Mnj8gvAAayfq169shFeEH2cYLonl0xueHxVtZ35wFMokW7QMqcMPGFHHtSvaTwvG4Y4vvvPlHm
ufeb5GkcSq73xUgW8h8J+DUOBhevXw2RIrmAbYx1yQHzsA0d2siltSjMtslM3X8AYZGRsflc9Jwa
a8UM4/lCa2/mEAlO4bykIMALCzETpewtB0LqfMwoclJjsFEKxTueEiKpFpmTo6D70Dgh46sHNEcI
ujg67JcLm+cinreOZGQ4muxdAB9GOdf2GxMk0hvDb0TcLEASQskiaHiijpa6PhvbNTSs4iTQZnkH
XDgJK+yI7Fy91XOxRCV7ByakAX84dKoWwCU6b+Dv+yZnsvRW2wtC9Vx0CaWyMkow/UIv9I7ueTQG
/QxaNkYc3GI6MDmPxIgn6x/NdHegYeFf/ObrWvnFlaRVO2tvXQaTT1F6Fa6Xu0B+oGVMweJNO0nf
n/pipDHHt3KtNO3/W6SYGND/QhTxLSXXHEVY0JXnBWUEdrk4z820MVe8RIjEPv9KEpiQmNymyde4
xq1iC2hFKrHQO9cR0YaHp62gdL416XCmLB+1DAmlMnx1ujM0zhcMU622MbG2+CgpVd0n7Pk3TXD6
e3v31z3EcFKKGK+zI2XS7ThszCfxL/MICDbFEohwwicmH31pTEHFeNEXDJO1Qr5fdoktC1+Ak+Ho
LAid0FxTRxbkwAObmrYtP4Al5lv4cPQMpGH/daD169KO/Bl12/mZO4jnqnb5CEPWCQuKeNrtIgkt
SsbINapO4wDIQCMZJl96yIiEKORxOlBfh/9BF1UrMUudjqc7yCQxQ/8tminfouc4JgTWZdCYXUXZ
3uBg51+RMKmTKfxTRhsFAntHUxmAcpfotez0uub5NxGRZRyv5ggASJKnQM9zJxlf8JBwWqUCAHhO
sfWnwGi1JGOjSOI3kZ+OPPe47rCsmvtE5pvAHg7EykDt17kQBWjIfHugn4aZq+vEVsC7SCNI4d74
ylAibcLrE4MNCzXNB3NG/OD5FKoCGj1uMIOLEXtvONPZafxMaXsCU52lpNL60ChlPVb+p3QI46l2
KT09/bbdOZ/UFDx3zYCqS99WK2niysOJp+YssC8ntNwpWLuM3GOpLRxADfwQdoRbfhozgLMvFA66
Ulfevy03TxnQnFRCxV7PxwSUKxBIFvdS0qovsSeqaQiGtBKE/7ptbJCNQ3iWwYjMak+T8NClkNzA
Z9FAlayZ0L7OZPVJRKGqVH8OAZ4kWhhp05NCyw0CHA78f+uzKGZGUFYgLJBCPWobXio9oi5+ARSn
XJZIkakH6HsH0zHBKCbVJ0V3FbMNrQJUU2ov0Hm2oKiIbx6Km1zRS3amAxtd22ZnqpOlpVC1iBbD
YaVghxxZM8xufh0mX192wY+YVaZOOyMqpBBeyxpr1+nwHlA4LoQRRjXtuXTMSyH+C5Qruo2PDpu9
uSeE2L6CMsAEOo3B3gmIfjMXt/SWtsbCgwo71JhWkjLPJ2idjI2AmiHNGmYxn4fV1ot3klwWJWH3
5zvZOi2ynzj+7IGj3Xi0hjGZyq8pO0FjC5SsRHmuYU+AAiMt5VPaICcWxqDPEavH/xEtJ06mVGlH
w+L9Wo70KzKrlCKfBRXwHBJhf2NFzWjLG0sWkFyDFmMeHkGJZTY6jsfyuR0oxBBkr4HpJypV5lrp
p521qPNWhnRTqpm2+G0sc6dTeThyWNwUIDSTy0Xq8YlReIiwPGwpuzY/y+noV4v8GdrB23z6SQLT
zBqh8nP9iO7nksU8gjZXWWzWPj3gzvpVcsiuiIJHrj7K+Jmpslrrf1N027mbQtQfbsIwh2Axjhkl
FNGwRLhScmyPwHheyJOukRHYxOcE3r11eb7elVrCxY3ldAcSXMjZg12MWVny8c0GtP7ptP172SLg
iKoVdtW0sWN3CoNwWJs3L+edun3WQpNfTmrPpbtyLBY7aAybbLNYMRZZ/r42OO02GlTXBMGP9yws
At43F5DqSqb3X7xlDX0HfBKGV+E4sAVj9KJ44c+niPZngMzf8aytD7W6/Q/eOjZVQZtekNRXIYAz
UTTWcfnD2YjV1VnkgIMlEAPdOyiKeFejd3m8grx6WAGuMwNsTCqHgZxftbbDecGxHQNLFjiEe5Ur
yl71j1DImO841t7NQShZ4XJnqTEpJ4YL1f6EEjr0a10fXHiXNYwdcsJ7pNaPCNCoeVYEAHk22uky
/Sy4aDTUSun57f77d/Jcw/4xL/0tsMxhVG9hO4aGhQRtN4LqUkFG3zEDuKKgGY8JZu+Yb/+1klI4
ueW/bC2JnNCEgrvT/PRDr5UEqsh0MaKAJCMVBgRAcn77XDKvwtFRtqoyw2jvJ0+8Tc1KWRlhbrzS
8CDCbCG0ieX7IhNmU5I9HQJQDJr9ju5glbiBkNcM9p+TpNvtaUT0xaSWMSBdyMdXz0O2eXyQgXPi
4owStw2gzXHO0xURiGX2H75r3xq9yNr4wP1a33DSjF9Jjvqvlz5EqUnK0T7zGAelfXYDF6nXkUUz
yxU5KLqZWcCXS2g12CFymFjZY2Krb3zO7dV1ZQsQ5vJXs6yf76ivNbGEMP6xYi5egkU6Qzasb8Dk
2CynoyOURxiBKJC3uCkpNvMUhwd61j7yepgSSE2csbfYtH5HDzUs7kwSJvqgePpCALVwvG2qt1BR
abCPPUNjhKOaX+cpCUCfavIxyoeDg/pLgrRw33hs8pr8KjZmEkPVJgbdpj1u1Yq9Vu2Q5NJDiQE4
K2eyh1Is+VVDMgL9/q1PVAsc3VpT4EFcZm8Q6xQyreDND9vi+rWdT6aukeg4TWaFEvzlPNOX75qg
hxn1Di+VS+UfHhAxdWS0Ld5q+gjQMZuYr/fPVKpIQutStQp/XFq4XxLfKwSg1ZV8VALwFar0Xaf9
2EuUUNeNaZL9heK8p2mRqIiaE1aCcxt4ylw5veYSYeQcTSBm6cjFxCKYf2xC5enbQTsAmFgiLH8G
ZgZVovhc4AzZ0Hx9raYRg+WjMZiHu+RQ1mqz5G3yZsDqX3a1UmO/WO9WVJzyZWG0JHksG89V4QCE
RzYz7hyL2UOP0nnlDmfqeZx8VKcfacfi0elMSu/17HbBcZPfgauTML+kfpRwykA+FFU/9OMtARaG
FeTAXzGFbbmJ8DoixNlrbNEgQRxj07uCGoNv/ZwrwZoRhBN9xinNXVBMk4MnnPNT1SImt63wnHJ8
E1UMIDxuATVVF7h3Z/fqxAGxWjt8OadHeT6AOr/K9guNXEgUbeRfBuDB1Fs0pcmtEujWXEmAZInv
F8KRrQM5/zOGRLQZaBhP0EoCk3WfQrfT2IBDw4dC7WFAxpssXa/0IBYsAgOI8lzlXch6BcqILrWb
H0+sZ5DOI/Kc1HKNQvTAmcKXetjL9ywv66/k+prU/zTHy+V3XoJfQ/ADeTNF7qt98ORwl9vswc0G
1TxAdQAdgIhSz65CYFHmvVitCZa/p62vlDCc1dcKZV6LMiZDz0D7I8FJ3Z00EGF/oznPDBYSLFh0
7GPR+wJZvKoD4+QZzSZhOz8SA9Mu9jqqYAfcnciWtotRudU0p//QqyomYr9iglzQi7ySOUsIbcdz
TTUKx82B2AAY6M/X6W9wgWa7Ny/YlT3UzVUbAkz/jsDaBE3fKX3ERuGi+msIe7egtpLKJi9FCh4d
2+1xSxp4+pQueOnFo81ioLe1DHec65Aoor25VUQIs2Ah7B4lhuT2mN04wO+W2gT4y4LOApWkv6tq
2E5dqTgqrWkIizd70Yvwh7riFc6qbRFneJ2gFB00nsu++W1RK3AxCAULsM9Fbm4X1LqwRN5aO+6K
aBEoj8lPizP+fvy1LkzncM9OtOftxSrf/cI4/QAk6W2H0G0NjH22J+GsDd2HJd0s99Sx0X4Hp7F3
JxxOKw+/zsO3VIThSL7+Yj+eLkoFS9E5sJvlREIINPI/UaZMaMxEk/OOXPEcdAYfCgq4pzrQq0dE
u7iXV8+s9r0+MmmqrxHmOVwEjH9g9xr/9Rh6vmju23uKCxyDguRz3jpQywZXAU64q8AVoo+jMD14
dLRk1+S6em+aSfFpez43/yagUtzwPdgZBe7dTz+H4GbVD8vq6cQ//+n4DmNQzIURmAlGXnqv8IRE
T9Repiocma02/P3UecYDYoBJ5tgb/hM0g82//wfYGVTW3C/dCAL6rr+z2LnBYUpt6EZ8x5LnB4K3
+O8QbRbf1Ak3chWbDgY+X/Y/cI0gD9otxGbFewyyDtGt2xEQWsssJm3mwx1rNAGJRV9On2aWjqFM
Damf1h0cH79rW77xhqffwiduGucEZSZRbbv6i/uHGbtQuTb56yEKnWQNcM4+v2DtCzTptR/8RLVD
nHnzgEf/+Gt10ENEyhcJjoSfqDeeW62BI0vRBUWuKlRXOPxKrqz7Fx0mdzwt7mCwkIW91aKW4Lu3
drHXBwNSatApoViLGIuiujBH134TD8MyExMhTPbDYECm8qu1PF1smufiFpmhEsw0fS1bd9NLzVyO
4XpUbihIYZhjYm2HJ4/GnCchcd5x01DUDEjP+G2MK2lcyM+cz4QCm4QI2T9fyVteg9hl7ZeLjl27
ngxG0Jw+bHOaES8KROThSUWSZw53cgZ/93aO8+b0SoK5xZpxZnQWsYC8BgUYfvKOUktGBrLBF32U
vw/jumURHVpWOAC1GLkQuwSrktwhwY1ncdtaaeTWW6paMyUZZtqmBBhUhgZS7rfiL1ljs9jsQYSO
o/p0+/GjksjcGSSTlaE2DUNoiFWgdQOonhzcouJYNWQetIxX5WUHtkRuXYwzl/8hWt9eZh92qfG6
3IywkggygkSUagMzHR1pj4KMywb9vqFc9mOGAaSdILFVDTA6XLovHX0ERFgu4NUiRxGVD33eVSP+
+oqgURv+j13pOW0cGx+zZ3YcQkvihsaUSd/Z6zq2DfZ2bFoyiY2TDS18waRXppuGi8wUYjSgbBXk
eGVjayN+sdpNK3eN0ipdb+vpebs0E8+fGq5iyzaEPnv/K8XgNOf/HeVzq6MEi68kENNe1Tcr0nkx
fnElRi6Zm0F9Sa58AoOXFG4qXL2H/BWTq7jCsYEeQ3XE2RysqPNpLZX1H4K+EJa/QDpqqmp110qH
HvHFg+/JzuuXD6v0OB+aL3ENEsUAUa8TT27zYE1eHoU41moJwVOsMj1z1PWoo4ePWKu473SDYClm
gEAWy7nMy+CeseaJJwHmI17GcRzrpdllM1wPb8nOEk+d/YXIn+xxC6Qln683Blk0sTc3QHcvSNya
Q+O1P5lM1WvWN3Y9f5A1c9knW39B+HT/aJlBHtjktbDDCD+rJRh93V2fG/fhMMqutYfv82hm7b5j
/kift5K192AfPbBjHjehFbud4wybfiN2gdoDjwmqTEH0Fj0dGhdaHsZj6OEsAfodf7EU3gqObU4P
1r0bLkpkOC8CtVarwjx/1TJ/mAyZJKJhaelJE8HWMXEpeTvowL8cBa/bl747hBIFHaFcUJGd039h
h19+I24u1Xfjeuvwwt3yWJrLQ3fe8LBoPVTw3dA0JKP7PEU2JiI+wPlzY7mSulGh5+hzNKaleqFo
yoMNAP9amqntebo/t1/WgpCAQs5GfKyawM/zBaAQzGz4hwjC1xfO+exo9KIbVd4nOsq7JYGkAbWT
FpG1FlsKH7VTGkBttjFGqNjdFVR4gWVH4mCLU6WJTkBsc4yF0gamN7O4IoTQqRwe1a0xf5kg7ICB
Mkd1oF2tckdRIyF6Vk6ZPAHHiL8OazWH55z/BQ6fsnQqpV5pn2ld2zrZ+p6Ykj+FO94V1GySlXrp
OQl60G7BI/ln7nTjxkpj83B0y27U+cqlSG8obKjc7UfpOdc8r2GAJXVewKOedkPuXnnNxuUrx75L
P/PYEscfO9qkWKnnEgD2c+9SXD4Id93VgQpYN+ctypSfVtNROiBL31+0gWzV6lBGpA1uPR96UeaX
rTfnPcxQ9kMWzibaCx6BZVuTfwkTMzTTW7mMSKymXuAo/DmJZXDCV0/N3JvGlUj3jmCehN4wsoau
cl9d5dwEd/UHSj/KTJcrNHMDJYrEDHQQVdH8xoNbM2yXCXeMQBxo6T9xb5cAR+CxQpmRhOoPxXPK
h2ltchIuPmCFjvgV55MZiKm5YL6nGJyc0GmBViErtNRXIDtjxBfB3Squ5ZikwIFllLj7qvVbcb0k
P63HBEO2RYMifGmCiFjk+XsSZLTSS6U2Ez7KcBhnzZUyT0YuRqHDbPa3Enu9M3H5WxMArESGK6nP
NInosGBVQAEc0UIyFDEscBYENmczJGsKnNWxrULjddAl21UYG5pitEHJWmkcBaH986vXLheMyrD5
rgvmrOnnnOklfRJmjjbQu0ffG0Oa3gIiAaFlttbGYUbJE5tUxXJY6MwMYhbclEDrKDlBbIaJpypf
Et5z0WndumPK+pr2rDU9O1gQVq9W8fMMNE9iYyUyfA74MZE83lI2al0TBZlQfdD/PpQhb6iOscpn
uXm04V5RcV6LbhDPsi6Rk6gD6g7x3QnxCXBLzDlF07m3WGmRyuXPd5aVuYtk163qkJpclfpZKG2g
krAM17/rGEzgfjOAa565UjqjnuL2s2nNJR2ZXeMQj1KN3ZpQZR7KkALRj9Xl84DONvEBkY+XI2zW
JPLxbyNYoD+OQRK4wAeWd2dDIWJq3Owsh1oUVQ3iJtHmVMnEbvp2+ZOWsMl5FzQiDdEtJ+UTJO07
ow4zSYxr5OHB2WVhgBDHXVX6MR/1Jtbt/mFKIYnDwwHjdqqEyUMxwW/1qimtqhgfevQpSR9zPbC5
q6+FiZkHgvh05hImht8OdAoqH91gJ1XCSch6GrZUC/Wkkl/Sc9p/fs+6VaSuDWWG0cTmgyMl7qHW
e+c6xHLFIYk1/bNaJ7z8+yXmw3At3WAccgNJuOVI+Toa8/cWqQzP4QtLoVrcaj62fMCwIfZwBhLs
bIHoAQMGY4GX1pUeTmSEjeBuzR3b/p7zJXGABiIRdn7EaRUGgoRupP7mWHfkuNjP0OKFXDQtGb6+
PurPMCeKAmzPSGeHSO+FZiDxkbxv26pgZ1/tvmdLbyFbxtldoMJUp94q5q+MDTdEB98MMCSswdqS
kcHQaKUiWLCnpJGEPBPhhYoLfbMG4/dN5OX2qSqn/NiuFJGGqCUHb7hOclfBqVzVR5ec1vSHxWHd
wv/PwIcbFD58pf7KUJDfMYACwav0S3vxgnaQJMfkD2fZFpWAKO8U2GjKbRI9j85HrIJxnK+XSMhj
tOX5nAxkm1d+Cy/o0AiotXa3PEsE9qqRP5gxXh/UElKr/pHE0lmHf0QjiEC/Mu3nL+Zt+csGtnJS
e4RJzDFtHwL6k7Qx9t8HlEPJX9eS9q9xie76DqrU/kXDN4ukjX1GzL5CqF4r1O+Au2dZKkrPKACm
/FM08tOPQcIq+K6PF5pwv1ngN4xg+jJCLa9Wm5vwXh9kTXQ9BTrgbCynOhtjMvc3mlx8bHX2BbUM
vaMhjCbDlhERvqLWNjryr7C+/ZB7tJ6+b2hf5cOdrpAvFf8Q1q+V3Dp0YnCnq+NVUyhMGR/1o7Hg
bpP+NYiTXMKzOfZB6MijW1fhTziXk7AB2Uk0BdppryWL2BdSWgkEGha0gnaLzMVxqPzPNTE3UAEl
krpwIs1CdOea493EH0llIILB8NWYdZaf3hr7n5sTECLVdwn2IAdhcnL00nSZ/5YNI46yAsUxv3bK
BVkmkr63xa5R9jHX+S/ZlkPy/Nf7LL4yLKryVjRDcnx+xRpKgqjsIP00hV6Zrv4Jv/wrtAtCTEYt
uYPsGfupvxW+UG4jQFpXha6tazrakBBEXsp1y5AGUQ9VrP+Z7ZMscauCFBka/V5V8gmYdS1UF3AE
RYxVsz0Uktdk9dV8e64+Y5uwuoYTEpZf+53qjz0ma95589yc5Z4v1PIP0IadcswaUsJB4ZftBoj1
Nb/s1g7g8fMfh1p10DxdKzwM5oZZK6DyHVp5TN/qHCOMemtKSGQWW8K8KnFH5cjPNtfj6gbV/zFv
Q5U6GcYvLQnUFJHdROEdzDVIiMD+k65SYxzJImGBSK8e1j47Fb+/zRqyWjjR8zmOar08Bohfnccl
iYWuBOPe4SYbLtcUTq8FU6KG+ubrBfdg42tjDA7CkNmD1QbQyeMAIQC3mi8GLKjkqyQut+qDYkDR
irj3WRPJuqoyM0PKbtImeg+Hx0t8R8nDMz9xjK/StwiMn078Zl953uEgmyRGgt0svf0CWcgq23bf
ggk0qwwto33H6NmVGQ/GVHD9D3hY5PjxKp/CGrlfeb/EL85CdYJWclhaHdoyHESl1kr3IxLvfzc6
IJ78hC6i/ScAvGwPMbjQlavRyL0LeEBRA4JmEgkK8nyAsoac+KWwT6MTnaBF5QatFyniWcqfcEkF
65Oknl5lwjvHUM/BJI/J5CkD4CztH99jlUAeuyeEtGqS1MFFTCB38oEeb8Fz50noR29p/dAnjPXI
v0I6aQRSQbpIOGUjekU351FdQEDoqU8pQ00FJgWeYstadhi4sXKlvhvagS5HBD1jtiSmP7zEo8xC
OBAnfcDM/Dg1JsmytVEL6K5JVv42RyeeuonIShaMBXJaCAHFU7vx/30jeyhbPvgIBqpiCeDzWRBl
2VYN4wJ9NurwSCmBbBm5Ek5/kNhKsoh+mjPg2EIJBU4CjFt+kPYOZ5HhYP10L98EGBiBk7eETvPl
9TvwNy+e0THY+HUbq6z6hOlKheK7veGDi3kKLZv1KhZ8X0ypfZzebNR9AqMKZS0lUGYKfoukXm2k
4n8sGcdorpLAewt0jI8f2zY+CGnQuWrseJUCLyfSsEjLqOReN2bLo/3+EOEJQ2nZlCGjkhap2GCS
tqpLoAK6G4jd+WjiUdOfF0JyPBcoikI6ceNtNZiXxToUvZHhDc3OPSgl2a2eTDQa8HpCB+9XKhp3
4hiKN1fLK+NoH6KFHuQmaC9r6La3/zupfD/91kY83OST4d1LJJsAopea/BV0DgOGi3AawkedVBz7
rCxb8gxzRs8FRngXoE3Xz/FbZQ5q6RslOH8oB3Cz19a+rNtDIHszvGxCxOjOzoHb3T/YjL65tE01
joHZNsa7Fw1DPqbOWsKJTXpIMe/zHQvNbOoRFPBeMDsMa64nj2ciun+KRR0+8XRdP4roZcTlXPiW
SlTu0YKfw6YS/zk8Kmv6yacFJGnnlCeKDzcubJx0CgKXnr1YVrIWmbXaIBGxgo9J6Fv0GX1jDGch
mXvZPUMw/b4zzUsEJSwcuEHJF0cCRJWyc47UcVACu8EyCSnX+dbsGw5jsFp5QArnHKztr5viuIdT
30feOT0CdArTPcxx3oVSMQBla8FQ/d+gU9ESLZB1jyREY3XNtZocvmO0k5DUgprlWwO+Qy/Yk76p
kNxftNbE3LWbh7+8RV2y4vxAGOb7xkxZ1TXoPCM6pHcoWnWzb8q49spOekk3sGu2teB43gqr4K2E
GVU0fRakpF32NaQeyFOQR/wRRltikXmORBF8oDE34fGE/fidt80ToxGRli4tAE16yP8UgUsTUBJC
z6AP8cJUbmeLMwQI9+q/NosLfKTyXOKXiEdvud+qboqFROW8oOt8DP2VwqpPQx5qktDEaZHslTY9
ZBO/LfWGd8dpHe9hFH6stX4eiH+XUYGGsJ5s1fxFf7rxXFTWumPKU3FgMyU4xN5OZe/kEHIv0WLz
NnxsqWQM7pNsjcsm5MmQq1iO6p//41NfZcddhDomufU68zWJhMbwkYT7elkP/1ta8HVDyu9+Ml0W
G9bADt9xGenLWiy9AAEZSiK40TdIh5Q9fRo+Tzzbuq4ho3ocDmwd4ZVB/22FstJiWaDJiTZl0P3G
d4bnZSwS4hgvAA75MSwfqUM1XAwCFm9SepyIhAX74RnAu8mWjrQacSMNhcjKjy4VO3Qe/ReLwyBy
/cG+8Y9yxI3CUPYoBn39B0E1c+8vDQfn/4Wdxg6FKcJJy3V4r4PSPBg3RqF+F/IPMaK9tXCWcLWM
Pcxaw98BIHb8r5dDcRv76Ow9Z+LzphnWm9mkOUpwzvF7xGqOSbYlbTGsAxBmHNtYfnyXr3pqvqg5
9Rd5Go9zJqJPrrl5Zx1xqei+Igc6j1YrGrvxmPNBpBXdEpFIQRHSqvxZTFgfc/beV3lRww+FV+zJ
W9RqHQnVlzVQQanCjqjU+0JxdCpOFJpRcUAA6OeDOetjiesgfL+xh1blj5b8VRy93J2kBdq425M2
covRABkOiGYFDm57h7gCuajRfBA20/vohDkqumpCYT/5O+fYLXPFk+oz7pEc0mQ2zZJWB0z3SnQT
PQTNt7th8mTxnc7C/ZOR7Gse3YlWRsU/Ozr4PBNf1Zb3kZWwln8umBJtH8Vp5b5jOFH6FeKAP+ww
Id0TRx9ps5dd7BJqEJJ/gVOiqR6jCFXwWF6g0I/404SF9qWgvi1o3NPNWdlmoBthTa7j0T+Cp32e
zMIPpM3zu5bRGliC1UfOhEtEg3BendOoIDi7pV4x5BQy2rUq1oDPDcUgb77MGFjEr85HPOlRsabL
OXGAaxMkSgMPKjHYbVqo6zOwF6OD7am+BSjxFNE4LZIvvGi9lqhFi5JG4qOwb1RKVu26BUU1wBAF
JvU2y+8lYchsZErjYxLg85qjf+Wba36FpHCDJpE0UxuKh610ekyZmLgXQuL8F1jZ/qz4qB4qpBvc
qSIF+Kw9y11vvqY2cdsR4MB5vtukbpGmhj8nfuxjNFK6SbFsM2nRGXwv43ZscfcTp0+E7tf+NJcS
UjlMH+l72yOucBIV3Dt3JzMe0SyE8zV2vjqi2dDD031pcXUiGewwbKtxoG1X9DOG820wgN02Uj5Y
9/rnhglXkRdPBk48C0NJuYiaJrkyJgpYjO2+xALg1yfc9xdXojLNVcS00cgti19KcUeMMlMy9jF7
dqs8L75IjmecfLp/MxNCVImGrG6wR8KmAvB8EBluGgifkDBKqKQTpnkuXn5cXWuaQuWV8JCsLqGO
PGI1wgRBySmrZ+FBuwiWNmmW0pVau8RuKcPIGt5Vmd70mAYlPZQ59Zcvs+wXbTi0NkaaicJ7hDhy
2q+2gZNpxSWufhjLITFHWS+zmJqDuU+F0zISi1lKC29Jb4cKAfisQSG6X/9Q2XMfxz+LgP3YA6vs
+Xb4oteMMhkLboue6uaC4fT883zE+f/xGv/XYM6t8MzUx8msdT3bXPmSCM9+wIiLdBBhVvaejmjR
rq+3fyJ3TM1kOH3j7qoVzhbLLQQ9a2ZIbcCwa+vYYgKHBVqizNrphnIzQR00pSE0YCTQQiPFIxCm
r1AcC1NPp5h5iJ3lvOYwvjbv1vhNTF0682hFrEbeiirWHzHLgB8Vidjcjpn4a5bc2eCf2hqxLXQm
ZNDYGDp8bzfOTgADcrvudVG5FfYmYfV9sjusO2Cz9NS4AhIkyhWpAJuYh6zY5PfMOmQ1UeMflKgM
8ABHNmOEKU2mIldbzbLTuAGRlXM9/z8wbeBRHJxnOEW3qAJ9O66sRbG+CFvHvoJ6GvImluztzJPg
doKI2FZ1X9kC3HRIdFkGtbGdqe035FbThdKInz5ZqJjFHool687uVsL/d8rJk2SlxqsbR/5aH9kD
iUKsM8xoaFx8pwLGUD3t4SB8k3jg+J37S7jZKaaWhHAE0aGykDT7XgVaFtt4xb9i7625M0DKE/8g
qowG1v3pBa3hGB4wYMr2Bf7QB2oaxjTadWrc90+jfE0zRYaEh5Of3ZILF3Cy/lqcUi14pUPIgqUk
qfIwr6m2FlrOdJmvn5OFuLjzBp2bfBYBwajpRvlK/0En4U1S+/crbZPhP4zA06+nJqw+cct4DqJ9
LEDYkWcS8XixGSo6SkP/VzUBh0kEAwUxfoa8+BvbeP8ZADKJ0owk5AT9QSCvzyvoQeKZarvFkekc
Ih2545Gd9qLl+FLzl0WK1LViGpSh0IyeStdC4Fal6eVUEZBvz/Luo+H0GeryslyFrNFyHLXscPpG
W22ZSkzFtOtiitpgje3dJuwBGykvpj1T1hYN/IfTm5UPW47KvQNmUeNmZstZoaoaihaueyTIEqMC
laLhYeUbhBXBWwoKXMT8kBiulApwIRLFuNQb2huDkSSK7aQ+Uq+1LGmLivTB+vDFQWo2YPj2WrLd
kW2bL6/yr8+eweg+XfnQK/UT40h8KOf7FvQIMZOWMaa1jyXg7t5zkHGpaFnHk9+4RWin8bOT9Yo5
0zmJGYeivq2sdOJ9McQhszG3bUdvSb7V+w9ztRLoFbn6RlhXAg19m1oMasD2W7hcyp+7oLYlL13i
+nd1rjxvvhEiOoTlnh+dZ0czupUtrixPxNz4dilRVjgGJESY+jU6h4z03hMT2Nz2G0Fy9UwcZ3ZO
xcVVAfa5NrEfRuNvlQcvdb8mgi8EB9jvpla3MZrb7kQ4kYArTWWFU+Y/WkddmCG5BT/ARTqD6pAa
WYxohNlrJBBH5p/9CMxYV3F0KuzNfNPvsK7SljbLxGGZf+CV/XwDqSWXPqJcIh5HxdQxJ/Q7NHfZ
tFlCXMbLQ1PIEzJ80WZa99Ax8dLBCtpS8M7DFs3nLpCoeNWLVLWxqHLF7dGs9fXhf8CwGNxzfK55
PXzuL2A7DcpsKvgoR1vGyokecVrQqvMUNTpyE+6H4erf5TTCNjip/U1Zl3Q+4vcdP5NaR4cZQk0J
P44E5gwqHnq/MP6mcGOlvtj+1D8Q8oF16AHfM0ObWGi8W7VEGCwC5DHbNt4HHm4N/8vN9YdPrPYF
N2zA6ajOWn11PwIxo1lzxh7iWI+cYPWYRzTIbKb/w6AzCWIZ+C0Dh6gGhxGf8D9ngqXKA0m17kBg
k7ZcHjjTEmnNfRqLe2J1uSin46scMTUiOxi5y+vzP62/J9PZV0jehOc3nO6KbTH795NeocFmnD7c
UAfoy8xEWbMjUpdvr/imMojQz9yU1rY0n4MK3qgS0kFYGiYaE5uL/oddYS06X8v0useIPvM/4NQA
zDEgqfypf2s4l+pvvTTJAw8KmjoFxXijnXFahRnefNdW7yqShAXhOhpkP0yknCJNvcQXxp+Ztfvr
2GEePNzTcuohQK2+In6+/YQK5TVh2OQrrd5SeeKkD9mjb7dHq1OkJODS9ltu5yNf5FgCbyZb/cNy
JuKPNi049eUSU4B8kF27ptWEbGG9z7zzG/0yE0SUBLUSChldtZDG5h0zHSTfI6m0uD+xxdWKv8wj
f8lZ1cxNDs+n0aMKX5l8etItiwBcM6ovZcsPMeFGphLr6WNRW55cRnuxReuYc+ThZ0FKm9IBddFE
FZDorYcEB1wxiCgr6eu3CorvisVRwKVisetML4fH3xDaHFty3p8Hgudrr3+hOapH1Z3gIQ/AGJLt
mI+zPuE0+8s8dAYI/lHuzWFPlajW93xU7Rdh9TEMBeQP0E/MVWUMsaijo29L/BX0GqiDshN3qJD4
mZd1oKoqTVm5FXVPeGsNVLqt4LUqYSUnWwTAMcDJoQG82rYDryy+M4FXL6EMeeXXVAMR2lwnYnuA
Yof0C+bmlmJIUN1TM62xh71lxpozOAJvA+7BJvqELPtkDfT8D9Ej1K1lulMb/QuTy3qgHJsfv7E3
OVr/AbD9smKvZ3CL7TuSygZlVyMy0uKOVN8zV14I4NIsHeCcntJLd8SgQbreXe5sXd42mvzUW1GM
B23vD66HcjvhN047D5W0gQHIXllSKfpWqv/4aJBfVwEX0mzU/VQ5XiTr2dlZOdjw4vwW3nc1JUUu
3SAYwYOkEVfglLy0dsCzEVXH33VCDjPTHytqdBdd3J3EP+PvpDj6pmHx4hndlKzMXsX7lrKBEIU2
2lqYIlB/7aTmaMcivf1HPjLPaqn7iuooVFogw+0J7R6yF3sxFKUtSwL9gM9DeJ/XD4tsaRS0c5PJ
ybc6a6thubZXGlrgFmXk0fIavndEZRdTOojcJPqex8b+gYSNzSCuyhHylwG3ClKIsQps36PEuqQ3
T518/EDT+0UsmD7jsV02aMZfJKKsGe82+4oYFVJO16v01I/KCX5xD+Wry5B74ucqs8MTs1H3nZNn
zExvlnSaFJLs9MUE8Ey6qmw+bzNdejzC5qLyricbChcz3hclA6goHI2jP4QpcA6JiAExqNi5uP8C
cnBITKVC/TlBCV/lPOArS33+ShRBIfJ4OfWhy/MujhRpZ7dr+Y+WsLmEF3rqaL97LQCB0fR0wE8y
rUxgxWBisgEnFok/AoLygZ3oRPBsB3R4F9dMWaisQAPAOOIbBiZe3AzSsO50irbvVKYUe/VIANm5
lJBq/k58IyU57YrkHA3NIBgd413+cwez9U4F/NeduwNOENw8q2hQKcNKSKU7UFh/9mFCa/zCAUEm
ZIim7ESEhgRlynhVeRP+7oifoc5JkHXkzMb6iphU8DHEclXVQR0nIT4mFy+DIKYu4YcPpKkB5+Gp
0/rYmrH2+xQS5unxNmfH3gdkojr2DwiZQL2y8AAGZCvFrDuBZr8LeGjEW/B3HtD7YToJ8gZ8E/qI
3cq0BNtSo/izVmgoQE+L6LjxJ8Vg5vR7poBGjd/6YaVwgsaIIXFwqgfGrvCFBm6SAboY6ByBu622
LwIyiCX3JJK1WrpXe6n0rn9kH7i8VsmeYrBQT/K1QrUXGcdtZJEP7wURzXPCRIxaKf9btrIZVpXl
OU5/wF8DtkvPqLEG67RGrGxO+vwcygjkvA8UpnvjanQGcOP8B2cgLJx3YZgsAxFO7C+SjAKTcPRy
fd0aRjWaOg5PS15hL/6iVhCeMlcbunhsj8qtkb5LxrYy4xjAS0HNKUy//stc2UGBj83bvYodH1sm
jw7NaagkaOJgNpqGcI35h6rRcIee+pDPOGHyHVHfSxP//WHcMM4Nx0J2mjUgFQCkzYAKf3sNlKHk
98J6ytYZda/wMifd3zfjQ7ZRONC8N4jCkY3RRV1JLPrMdbRqAqr86sT+ZppKICQBoZ1cA2sWfSEQ
+t+zSfZJqscqDYyV3deFFHyHcYvXnk4P0ME+7LtTgX1lAHEIo4H2uZCCi/P0SGQsKa2bYMw+6oy2
ie6RgbNljUUaa5z71SGuSvjhrMQiFTWJcvNLDaCw4HhX7IXQislKaOVSS8a4liFhe//D1rSJ37DK
ZP4RYNgfTFVldyeTGJZp4RH06IlBiinCfN4StNH2kBaOWIsgHt353Io2go8nUj7xLzIRo/7qtuCl
aa0NcgG6+ebhZgqS0DtWKIqFHo5pe0k5uzNo6BrQz1FFICoYCnAY2TybOvTXlVRWySRTUGJ5l2dD
gpi2hkIgK79VxN0T4hzsWgCjJe9vfWN/My3oNJluIPfB7TQzN5BFpLU7rIAbfqBRyN3ugGiE1vo7
2lBWVIEUm6NNwWiWtJUPfH7xGonT8vCu29fsW7Ry1hnEPhXUnfX8P69L98UTau9jsmKp6Wd0q0su
Qu2qkozURZS5K9KSqvNdK2ZO2ffOJYIkjDXita6SGQBWtihPYQBqIRviOvb9dnGrydBIzop5S2Fb
qNOi7aRciofH6SnEueu7p/qltCQqFx6CVdaVMBpqIsZFrfIm45Yh7fbuund+u5ED6a5HrNhAyvFw
kXnVO1N2fbTFTb/tHZG3rKsjInwtN2UTuVdzhyjUN/wMvYafvu4+7X5n2dUrvz10yfzEUzS4XgwB
HZsUSqFn7T/0aObTYvqd1krvH4hU9yy1HXHSbSmdNAuijx+68LSXRgGkUU0jcNE2yWKSFQAGTe+2
MUfW6n4Cp7mFi8XMFwjKrb/oZkqvY+SUZ/cPWb1CUMmJZdhDt4aBteXt6ZKEWalfHsvZUaFHFuCj
9Eqx6WkkKpx6Seibn70VUfw6jYjRf/1invoJE7+H4w+b6pt4pt3vdnmRRmGay72NLiXWDE/W1aPL
HiVo3mF09LMkwui51PWedpsVnowgaL+8sq0NC5GDfbba3rFDtxuwwY4vyTdihXcfzd7v+1Re6kx4
2llJkOqk3EXlizbtaqIiRWB+wyBVolIkUzW7sfRjGCQ+hl7bTv33nECOAbxjgRY69Dz/4LXeGeJ0
F2PUgQ+0Y6JWpsUf1Avn0LiQy+muvGYm4aiGcTRm1mRX3qTfhs0Q3Aq6XHwwH4EtFb3eNplnMYSe
7Ee9E5QZeLBK9eXMspVdvXz4G0Bjnoso7LUwHSgIr6+vgWLFnGy7S42Di36Lw49A3LNvJDwe7CuP
nlywKmvHyGrYw7hNWBLxQIoWuH1DT9R4anCQPWfMLSuGHI9OxfwOXx6hg1hfWOPhFPK2FipIfRfC
OrUYPyd91aiHF17jeX+vmCvBR/5COXwclPpAHyEIclDuoBxAuR8JeLDC9+vRxyFPfD9Eq+5dGH7w
TMPDvFH5HtEm+3fnP7dF1MTaAn1Oo2+ylTJ+Up1Y9yfOnnlScnKvkHfHKqNMZxJhWF4DOGUk5SM6
PWxfXkwm5tjvkwUEdMR4pX+RNo4zQHAXKpYvRDrm3fJEINfGOxUwzdqSBklHqO21YNnskJgE5e5v
Pnq45Tf2eePAXj4oaJT0c12B3iTgxXVPvkYLBhwVNV2VqEJueLhizxhX/v1asHZBCNykL7aReYKi
yc2d6uefFiNcDBpk1NeiqEjrilnQL2X/eXqSLc0MQIOkW5AFxXo9AYvQUM1fTo6qqfgrabeX/4no
5TCSQIGbJu68i5T/d53IQmtmP64vf859iKZQT9iryCTu1axM1Ca4jXfVKxVQqLnUd3SRMKlTCTWO
hwgZonbW5mIpyKIndFY/Q0/7K6LMCLu0EyDteo4SCVpdqRrkjMn0HcK481ZL1m8aIsyXlHMeJ/9k
7o6JKnZxYSYCogbkGVdgKETupqFIRRdf/S6vt6vG/6do6GNHCf9F3YzdcnVKpy7TWmoherCD2oph
+kdpcjSQ37bBlYCKeF6tz1GxY0EQOchW9sqznIAYyKftg3+MJLJvOFnnfT2z10gMmC3aujecPi2N
3oNnE7tD4Vpm2GltWuklNZ3jFsmPZ0ME5ZRLQsLBeZxcPBe0nTIqcCHqSNWOFP9FxJZqGUGImMBt
5EGM1lVe51TlQetUE8juHC07nCBXay80PaARbnZn0KZRiDUfC8bmECpe8mDLhmTIFbxZ0ZULGlpn
404yb+HHp2xTu3haddqwhwaRchMPqhPzYKPHd+JS1HWLimq1PP32cVK926T/HhJB1BeGd73RTobC
Xsa37t6tW5Pzx0/kpb6fUTUPT0Hi3AwlbZw/1D1pg1bmzneJ6SKQomcKcuRFRklavkLd6Guhs0be
h9lpVmh5o8e9xvTk65EHIAhbrK7O8s47znrdzvwNGT6eBK6fpulFenr7m/GUgT77gzuqXYcPF67I
OkyiUIoxFA76kenKfG8XFsJNmmUwqLTq/t7FRPlrXgxmomiH4p5gIRZLfizSb5+oxpsQanZjXaVb
SzfPqtg3oiXP8iQMEG1PPGOlfED0lbtKvHaapfIAUjzCGXjkBJkWLLBpMHSdAc/m+LUD6V1IBz1Z
sVouw3UbkRqRaPRrSHZotRlLZjYg0/xbPYKDBCOzM2mGSJW1uHIq+iBg9izkIj3VFhrD7z7xgC9P
UF9I/50uL/627l0QJd4GoC5Snu8BuvmxfCETlaSWX4kaU55RFR5G5T6Rm4dgB97I4r2sc7gCIAFV
2jbQkDPrgojz1S+3/Qj/dWBPi5sSENuZhHbbdMNoHjyFzunvTPw5/6qxXq+mjhgN3//T3X9lSqxQ
6fLVirZaqFxVSCCgShonBZfFmRw5lIoz6MujKOHlJx2YgwdFD8mJicpjBQKKwHa/UZ+H3bGjE+NR
yYGg3k+bYZZDnxl1nkPzQg1+iajwfpiHPFCx7T9H8sM+oxK/aX1dCMNLVXtafawamQlKxqf+h0AD
IJniRWu4s9xX5cCv3ARQ1j1/VDwjRQ5TjVuZ1ujQAIs8t/zMIQfrL9Cqsrq3Trn5zfPEOQYoaH2k
2FEd9vdXhrQj78L7PmoXAzL/Q0ngOBbJM4TRw38YxY4YhaPpgLtne5NaWIzBcIepsSaM2SIlpHSp
z05CUrjGOAlbP6iPmFzmGK4nuxJpjZA61UrMkj2LGgsAAKFP2v1DuYQ4wMKyNt4WwMQCI2A44THD
0Y/aPiX6aqI2jN2oLfkQrAnuFOMs0LFQNE8eWBoyIblzQy0eOnrlQTzsRzNXQlNVqNyJfRaUXA9F
4mzs4BPEvg0kDtxOA89EixLDrObDhplNz0Trjd75hbS87WvxIJlhYU6zhJomC7gqXXLXbpWi1DQ8
E+QYMbuvR+rllPzIVrE3CgnpzDyPHwBoXjXzYtH0c7yriG8PayOayFA5Qx++3fag9L2/ElinzK6I
0dxwOXCrn75/2MjXis0zRg62ig9ioNiBcX0HlBbwzUXHfobGHXB/iQPgQ2GAoIj1+Q86HJEdbeTC
Qv8FYheLbiD7D9Amqwa3fRcPwfAMbkwEPcwCePz5/tPedo6t1kUiO2LmXoM9AJ19RtlaTxeEPkVv
tH9n2rvATtS6KybEn81itnPMOOi3qSEHTr6yBFIerkfLDxGxT+DsdUNsVzIYXNbe+Bkeoh+MFEku
LiI4WfX8Nlp8I6BP0au61RmP0rS9OvjkDIewdtu+WMN/H90ME+8bAjSxNRP5InnGPZ27pos3hIh7
Hn6MPo02dihL7uT5D2ebxqgYKtZmC+yzDd8HTzFEphcmQVamTh1bvrZEjDJbtbNggWyCvkgUes0u
6SY0BkSnfsSzY4lAT1DfjMxLSB8OjgmVG6zNbNM1PYso3BXrsgb3Pk4RDHg1V2Fcd7a0MrILLQfI
W41rE69sVN7TbUmQR4LDkuGqDbGUttIv2+yN3DrSXO+SbTlCfKgGCjPg0bD+vRWspPH5JJmbZ4mW
H1auppxO9SJxQJs6nZTkoYqbdgZLhNUrIooG6EcoYINv7KIlod5BEZAaIewXBQnMAXz8UY4IrGTr
8/kaFZWUhSmdsE72Le57WRtXSYc1/XMjNU4Wq/yMeBU9qMaHqacblEq18zp+qBIUJh+Iqdvhx+Sa
RWCxrVAozxfyLm+tYGA9Itiv3BbYyYSXE5RL7JG2h7jxd9doqZoITGMmLkcVPOWlcsjpWrzJ67fo
ihgLiB2iK3s+PP6aaiu5dKmB4xXrlNeNZ09ZDxlDhabnd3Ldvai872K878QM8gRnsY2OBeZ1Qmb7
vl5jD8qnvjgiTdRu6pflDz7/MREgHv8yPlkrbW6qdvY1IV0SDWy+cGViPrY2936NGMMbRwmZHl9m
xvAu7LJIipa8ESdH2VAdj6TeLl/4W/evEwyFQDkppEm5ERIRQVcuD5m/hUymH58VeafKx0L+0cVf
tMLiTvzpHbiAiqUEJkHZKTJ3vfMqmisLYfOK2BHbbFsGhi8iOn2dKVYUniEHkr+HoDISPLq8V2nT
jEExsO//C7+T2XZH9o6c0V4pwmoEwooLbNiQUh9MG5wkVXYYq/iPC9xQz4FNsL1mnYr59XB8f5nm
SN6eu2LvpAEl653AAjGVVP0fmdKM3/T49NrogFIcm+lLdbT7BBLuw8/WvgLKn9WOSQLZMd2Kz/yl
vHrfSEMn5uSCiOctBOSzgjVWjBUOMZfLzhYRwhFxRFE3sM5RTgoahejJQeTf7OvJygxmMHr106dc
9uCC0JrnBqWSkq5j8eW2u73v2ealpZqMW6KRXDCfSw6JZpDp24op7DJrz3nxI6XcQHDpkBKEXSjz
Wf5BPtUYxGRrvuQi64J2sNY0SNneKC+m84QAbXFnYkSK9jpjZNS6K1vVeTLazecmx3rMM6Ijhitr
AO/xdCktCcxd50pK6KwKOpXESnBSY4E0Ro5n5FS1CDxSnbM5K5pavFCWxaJSS3JOKsaOtCSWO6pO
RdmG0bUUNglHrKCfPveUgEbex8pVNGL7UaSw4LrHGLg4GcFlnd7C+m7DdS6s1T6iMuRFtOVPTbEz
lKwJhSNev8L6n01hUwuyl3dVRPLTiAPy6hupOOe9ZGPREt2IV1YwfD+7WN9KLF7KpyG2MfMcDp8G
A4qxZ/eVMZCLBYoRXqxaXnNZiPWaEOAGhDh7bQKZMSEiOXjM0F/rXQYfJL3SlgYVKa9pvGbGIhPn
tIHFbnA6UDBGNawlhzudrTiUoSsrF6KA/ZuTF39jBf6HuSOsJKGsnbFS40P0GwS/PAL6bp/DccAP
xB4MRmsCOeTKcS/eoaVavR5yaTKDL168uD4rW0tbUgQkDFBu/ibo4XpQHbqaN6+nozeDEOrq+pH+
wNkyknzljXxHqoWXNT805W+QTTnQSjsHPrI0fjYcADOG1JGMxBGAh9p391i1BrV5uoIEvVWp8mWD
mjxlmuRD13uZzTl7AQwVRx3jqpLFWrilOVpaQyzxPApjVjf9dcaFxoqcuj64/dGS80IfQ9P8mLrE
A3tocWHXiZhhEv/4Dcdb6eWBCyNCtq3RUhzizqw/ZjJoJiHrsCWxUd5rBH/km9gQkp7gDv/1KbhN
2YAqAngcQLCB5AT9YaTbTB6WlsRh4Yg8rVR4rbPf7owX+eo+N9BHJepvg2ickXlioGNtLuOfSvKh
8oFuNz5B8Xpd/9HAMc8XK3cZYhzfEgGz+5sN62z5tGMIb6kOSRLI3KV++CnQGNRQDFC78gol36YE
2iQDM4GhFTRnPcg06QOR26Cp75acfC03WZ6+kkjC/8ZalLv98hIveJN1FEbTRlWnMnhJqF4SdkXH
dz7kEa7H4Xa83AdL2Vr6Qtwyr7GDXrWTvu1yNHKfYF5yIWejYYrCJZhvI4UGBLuMUkU8EA1ONFOf
/tzqOVQBT4+Vk4zHfp9zT0fs0HEe/29bhv69BwXtAYVtoNWhPbhYfOvk1uAm3uTyJPP1NonzLw7U
2W+ZUTLZyDSivORm/y2JEvGeVUtW9zi3bxYpdYN+qmMbHwLqWisTGJ9f+3Rypwv81kRXVj82ca6Z
8TZneVMKkIGYGuVSB/NzmWpqFUGYPJCDFotTKxfp3uyo7reGXbmLMmkUfQkHPbj4+JltLm2ISBn8
5WKvApVmvLGpPfNDOk6ARvJ2AcQgGu5csEWlRV81tTQ+MtQsZbJLOB2YLQYwcybDjQtu4A+JhEHo
o7D2mUbFMqCUrihJ0KCGNGIg2uPvGq1i94W0vsOm2R+Nw7aSlBDRh+7zpfhao7eaqa6UYPTy7qbr
5gsVCOrD6f0ZLEZKr2VuObr8xbOf+jv8CzfxZUffg1AMJ5UEQsM3cDKAWsQB4nA40A5N0YfulBuV
fSie6VDRLK1+VwnB5c5WNKYWIZjgg/dKp4Pg5QDzEqHU8WYHm9v5k8i3BjzGTRDFEryFA5yAhVCs
YVqzS4StyqiQAysJ2Q8DATGkHmTTXJmSZRYh4PnCWqB3iSb3oxluCg6ReJRpg272JeAY1AO1KYA+
H/j6V9q+13HVXXcgnQAX2gRQjha73M/kLbmFsHZkLgPv5X20JB9P4bvpC2jViZLzHy610JPdo33K
RC9xU3QLEFl4MebJmtOtYLopEKZI1UDAviVIdJOgUspM09C2Qo6hjwKDfq26MrznMTdDSUr2xxDH
59oj7rYDSxTHvcsGVfpGLrwrmUiEYSDdXTe7g/ZfGV6vTOKpmCU8ECEo9jPQKMVeUi+43zrx+CpX
It0jjugoIRt9GqlKJb8YDKOlqQp+BP01JR3k3sJLRLc/7zNmpVDQZP9RzlkJv/sDpzktvsJOuKVx
3hOYJYOknH9d3/Xd6rk3hWRGhidSCVo5sfM4iZV9TOpmyQUfleeIncG5AjG0mUR13VXYqIXH+jl7
N9w/nqt+MY8j+Jirg/gPHmGZyAhkFuBq8v1SplUVI2woDEigDfmvS439aL7r3fp5ZjObAPo4aIpR
ptvoaQsFmB2Q8Xy9/Oy7kiNN/lCRbIHV9eQwXd3Ekz5ujHXI4L2hA4psuMs9M24tP2xolXyhf7sa
XM/DjetmrAXwmeblz7EIAPvoNchg/69fCixQZY5XJSnIrkqr2wotMyowJplu4F3xZw7GTdiluQUU
487K3iKW2mffNGdR8j6ijkJrTOYRdLX/Y6YOtYZg7GZ550IKUOlpR+kUvwWxxtOxyrkSyQ6X0BQf
ZdOwWpK9TbG/wRFvj0n+6+PoruDaLSx6dYAmQa9gj3yR2CCkL2QjGExsoCDQ7Lu7eLmv6n1a09Ch
CbhmfIu8HUNW0tHrTlpjxd124PQFkHolxQs9I0g1+oV1jPl4gj+OZUOUM6vBueSOfKzFGSt3RFM8
VPVjiaID0pLEHtPW80vGn2QpzTOT+jisVGnWudpqPThSUvWNVE+tyzApZ8jHecPLRu8EXRUPcCAQ
uimRnRIiB7kV+de4RQAKdf2tjipNDGa1bvzwFR9onzO60fXIJt/j8TymC3dep96VWUFgoQUMM1hZ
r0KVhrlS6r6ydoV4C5giwQ3Ow5qk6nBaiY3cgPJRqD4+vuMp7ez7dFYSsaglo/Uhdq2SY78vv87n
Bf+D61bynGCiOCsXF6fvrhQZ7aIQTPpbNbA7Umn/wQ7yIGZnNfeaei29uFizbYZb07tmY7g4zq6x
KnT29sbkxbu4wFh/t7lsWaZNaBmRWj+FNGeCpTMBr+F8nDpbSl7uL0x8tYAZUKeSQ2LoprspGZC2
ZvddPIm+cv7IIKzE3i5NpgJePxb1XqO2K9DEpLYj3aRfsIhkW4Dn+D/WyTfmuPvabtSieciTH/B6
h3tO+csjZrJ/00RDG5vbrIeyESdSHyO8LLFdkNcgYZZ/GdnJfokPj8vbtTUNVP6j8EkuALIhDmwT
3mYj0gxSS2Q+xuAMmnOOEpVFu/yS2ZLSz0t7uQeSEcfLbGxVsTbeDB/1k200JlprWBeU4ibF6vex
tETjuAqhT1pNqheckqbKk9ObyY6C9r0w/7rHcxe/g3/E8qaRW173cVQAFD5YqWbuRn+HsPLsihRC
dS4nhzRYQQhHRySj62iUxslrR2PpdHSFTvu0d0CHmTk7EkPQFQbBBWkP6Z0BUrjRZAcEJnDHrxdi
kpUGM//aca6vlLUXQw0l0S5xsTBApjDnehCPUZxctWCQ/aRC0qlBWd4wUYK0O3YXAFmU2I+Hn9Z0
+iJZGWNgrxRST9UYLs67+hyOv+eLOsTZjXTq3/II3uTT6yDyiRX/rcOUBDOl1J4tcglZ3k52VVgl
G2iBPCb+wWap/r2Ce/EIZSHx9stIMgc3u/hHnCNdkuEyuid1cRDVzo8gB2NME1hjphcwY+nUM7vR
m5amhd+26iuXxu7+t+hB//I/n6fiuUz6VoVPN6yHOCYtT5U20M3gTNxH0GwwH8nCHKwyp1uhOPYw
KjksFQS6XLM3kkoyA9YZdMviUTlqqnfi5Iyn1EJ1SvhmIS/HtzTur+38+KLLkaDgrXCds0B3DexU
dJwXla0fTBK1GJXwP8nhu9cdlzuKj7w/26jlqecdFQ/GFKQTI4qBkNjZBIkJqaHDGe/oTDo/fqM9
QiD96YuHjDFGIgk2XkdpoEJvJ7jlRWObq679nl0qzjx1/vk8taxMM7mfnZ/d1YjRYOeYdCyaF9x8
bILC/E76Wu70qW5LMvAGzljuGqLaPCgYeUsdUfAqOJ8mRqO4eP5rGA3ymbCsvaX4mORHHVOaVowg
h7aTpMw5aGDMRoXHT5G9c/kwH+JpJJonKkILiX4bIZkakE8JimyjSOc+eMQwo44k4cYEgYABh+9P
Jng20dd/cP8p+SyQ3zkScYqcnFa86OanxZiLjbczXJo6pOePueU4CGf3kj6kTMiPH44/XAUCq5H5
rbIWhI5g/oJO3cjcL4YdGOKsyskrnf27+RtPqA4JyrtrXmZj/skPd2kB36dUrdTe5qYMPnxnhOX2
2fOC3IoaDPj26g0UNuNpVwaOnuXBTdOMiTdikgzLZl0rKaMlVTwazuXgq8obSV1z99yu2nIArktd
CnGBiRD7q23nWSuH39BG6BEg9jJKVkpb/3LvcZaWkZE7vB5kas9oBdr2Ma7kQEzqcx34aY1fDY6l
fX9h9IQFZvWS+IOjBTQp2HqAiwXNDcBjpwbJf19rxP/VMF8mhR3eV46m2ybBnjtKOOCb6l1z3odh
4GM84/6ma/sHIF0bKEVliB9s13hrKtblAox0o1/ALhCpwEgF7p7k6DX2nHE3g/HrH7sHm/+tdtbt
oPihoos6rsAB6xwqFk0EO5uimCDObyYGSE+06gsrwlPu/NHWyk9xpdJMnT6bXWYKGJHyWZMUrIEk
xNyRFpLlTPbb/uD3BN50TGDyOHmZ/eIwUj85nxvj6uCZQHZDDEkwqsZdp9JDQ4HGScVHldJK5oBH
7PRbZEeiPuZaX+I3RzqAzKO3+xYIgH/q20vsDZUxvDoUXmKPbWbRrVTszdG6jrGF330sGOosn0pL
eNEfC8Hy20nbsTk7r9rsEiysfeFsGKm68RjLg/8bIYAlEtc8guDq13HLNiySQiE8sn5SIujn/TsR
IIOTlRB1NmISDhQkWQjRyLsCwQQsDziieqdCji+Ed1nTDou8et7S4Z1nUw8TvUQ4ggM3TLrI7ZpY
zBmwbjTCVzc8tk9OpzZKH4ggFtyGU7UO5mvtqOGr6QauisyO7ej+8OVd/+4zPqTH0RiDFy3ZF5mD
x7NKh1nGhzqs9eeY/OD/SO1E+wvCTSdZHM5BU7XIafEx/hZRUY5GMDyEQTHKUthunr2jb0n+rFTW
jkqwDFjQ+yTKe9hKPliuBHXzQR/q3Yx5u5YTGheFqCuywntkdqtmF04GREJ33jOaWkpFjTRrnyS/
KcONBr+TrIXQhC6W2GefHTPNqPfqKt+k7vIHRA8/bMTfhdAFiHd1VvHdUwLBHoo/owOFq6sRExZj
+Enjvy8kTowsSHbgbGuzUuFpy0Iotz5aUGP5H/6UPtui1Zkyi2QddnfQ4MwNiCqOf4lGwx1hB7Kp
sv60GbQtljOMUtwsN+tEF76Sg4SMP6JGUf1/DvUJ8M+RUsN1fn7ekIgO83EsUrz+6eR/Hw6Pz5qk
WxRc+izV9iokCq1UIM812LMYb6WIfAzl4y59QWzpazi9kCPTS4UPuI/4/qsxEg4WNSonYGC1UClN
XVJO8ibhxpMSchQ0trEWjFCNeOxrXUCL3L2egoGhYrBE2NmNbsB2LSDAqE/WMNzbmdPEI1jEmxe0
iFIKEVoEGdQkQ4+ny9HJOP5XAHvjZSYvTEzPpli6uVPx24NNWu0gOETar9FKzkSWOnTTsmbU1Xgi
80NK13DSuFeyF25NHRroUXyOW8fJ+ooCmirfpff5VN/BpV0wugiOu1DB14/y7v5jxO/6w+SLhrLP
Ij5Rz70DmlheNiR02hhxJ70i+N3sc9C2VJEHa1Wv/BhJ1JnErW+hac9PgVOpldVeySJ0OPexY4E7
GSImB+ZHnpld8KfUAG/A+D079ak+Wyzn9EXHBp6YQ9n1bESBmIOJS7YUNKQfCHNiLATUQWSadSEQ
GkTiPw9rxbgYXUnmfg0cKeJR55NsIeBHINFrd1Celfny8JYsD8P30lWGck+hkB4GTXaiPsab7uX8
HZasMlvJA/oXOOiZWl/KdHQ7mGiiBAF2QyBHzinyxP0Mx+p4UoHNd5jEBCYG5BybmhGi7s3jfKtk
t8uBoDMAA2kiVByVeBAAQe9E1cUX/o/UmjdUIkOkXzdCM1UwqeNe8phgthsvIZ8hY0DkGqnSJlkC
FdloXBrZeB13GLyjNFE6sk25WFAYubc2vuyNsYf37D96/nttXjS0JMF0g0a/rByVlNbkEq4n17q+
9goQQU3r9+QCWtzN/GwiVZ6sE5yy1RtEMuPPaB0TDK8xOtl9yEx7puGhxUf0yD8z9BElY+F48KQP
OeJIByzz8ACLuDZWn9NJuP64Dp/vp8YNeCmkEeFjVe7IxoZqM/tIaqNxAi+bI1V5Fm6NN0uuUWRc
e/TYNkl8rUEWp7/OtH3VpYAjXfXggTAv/I74veqylsn8iVSS5j5FTIi6bgPKOfjeqczJ1IEns7Wt
Z9I/35Q/uGbnCtiOk7uNNVw1eM70ldFWMJ5JhH30ZshWUD2mTRRxzuSTaalD8AF0EaULegP8BkTi
iBBIfF8wQqdx5ST/G46Cy+WsTrrSLJWjfB+fvK7aLokTNagFCvYM3pCRkJF/4QpPdIkEdscBASnG
E4VqMenIPaSOlz1pj/5lNCaas+hq7GF5K85VNqKvvIquY3OLW16oyuc6nlsu01vb4geYB/IoFx6G
M4IvtbVb+F19vlGgZIFX+fs3XSBlLXn99iMEw8IUu1ZcSBm+UNzAkFrLkfXxxafcjEwpxsMg8BVX
coA6kSJYEIKSXHOiUP9z5Ud6k4LDlnKFon3mKThUDQUFvQ3HEChKG1/umMED69tzd41Qn1nuoP40
zhNbV6X/5PWglmaDEfSDwc6Fj5H31nSAK0iyw561uAPazVEAsCGfqOinsqY8OQ8Ij8OeiAyY7rZJ
emwf9MBR3hTtRSmPApCknZSBF1iltfGPo0gycqvVcejybmKSM5otnArT3UoyaP7FuTWRRJi092s8
kBlMqmutJBj9pH2VwT/LCULbmHnocVrZCbmFRb6uDPZLUnf2rSul9F0oy1PzoQ7k2QJ4Hm8Ns/X8
aqEzO/UfsGnAVcrvjnoSwRcqCKK/S05tpOtWqlwxujIxYlXb0oLBJm+BRbpHNb1Ulz8pOXWeogeq
rjz6beqOLk5vw+jBFYYrRr4R0mKGxpK4fRucC5/s3kaMd2DML3Llb6W6riZFy3t17HboiqFjORXm
HYt/fc/OYw+4FaYSEVtQRsNRbUZa/h4jSHFSVU2Notl5G/sbNV9wG1jzw6loM89xYRxlgJhFWmbl
Wjcog0mxuh7P7JGtXY21gqfp19vweY80na1x3FOA8EN6wka9P/Uq8NlUXU9Jm+9hZaiO0wHi+UR5
Or4Gwjn2svd4KKl495E+1VuDlFujTiHAaZDAvoCQ17en3fOzd5PVzhS8L/BDgN5d6KHTAV/ItCVF
eB91seVSrl1KjjzLDAB9DNxuzfNZVtLLX4/oqcWyREWHQ+N8ZtAlwM3f7B5lWSh+ttKrOTM1EFSu
WvL/yN6ip1qNKsgJ85Y+P1pP/M2SZtMMPTOC3AbKkhERB772ZDg4rl7qz1BB639LgiXukdupJUBr
0i0BgCMBCB9F7D4056p4YJx3PXLFFqlYbaoGWBJoBIfsVhjohDMniCoFM4FkV2fP0jP+5+pxNr7L
Li6aioyLDjWtVS2bXyC+zJWFXB1t0AKvxeMrqmzRAjFhWoCm0ZVboKduiBufLq+YwfOel4QAM+UE
7C6QtUST8LivM4N3WV9G8A1NlUKtilmNbwosIQb9ft2K8S6gm4zs/Do0x1hb4ZFSC3z7cMY0MwfN
RUCyAzoJ6tAVSd69q2StZWTiy4oR7uAReRYCyuTjwELBO4dBpeh3Uii20fR2XyOcOyixZ+bEdhJs
ur5V/fHZUqpfl+WN2gxxEfBB9Ux6KRklTQ0JCnwYCpsfYWrRaZeAzUUDLR8zkZPqwy+xLBN1xhYB
ncX/IR4NItHVYA68tydGzML3TqvHEggv/vTE2DaX0LME9t56Z79UxcJiV2UkXyd4YvDdrDzvsH3i
VmSC7x2qq0R1TSss1gBWEZESPAzivAjZS+DTmtU7lNRZ2IL+KB/DYPp6sX4OIr2XHPQM2kUfEqoZ
7scnrdCZW8WEnprO/p4ANxhU0EiewWg5pkpzVRP6kh2cQ+vBZcUpp34Vmngkc67E+daTaq4A7vID
49omTohbqNEY/HSPrJSVHqDkwVojG4NL8jcxJC3FWPJEZ2ScbnCyP9h3big2mMGGU1pXeHGxhYts
MEh5vY+ZsL41PDZyq1BD6wCrJ4c2y96M9P/nf/XwRl6oTZ1qMt1pzyf1gb01DGMiWjQseiswN/Rr
rn9aOuiqQh+3dIMVSLHA0hQMlJPDK6ZAKmEoXlVA5C5Q//IjYXog/ZFtouOP7KxRdM94C5hR8b65
kdrwPssnRGf4kMloFaJqs5Oh9jOZBGk3bPclkRN0hxb1booo0YY5jGqFkNm4U3J2vRHY6PIJEfw7
Jemu+L8xFh7YVaTMK2GZoTR5h6oAC7H2AOQ7DIQjN2O1AwTt8Sz7CWFGuIELl1q+ed/XpVcFtJ5J
x1rWYHXmGHeOtJmCgVHU58DCHIO4RZThSq/zHQWO7WoxZH4cnZGVmt0hIalDHa5yd0BL8H0Ap64H
NMzzNOyAkyDIZMXigPJG0RduS3HKhR5JXGHuzPiExX65Ui5wieXgwW1Ju8lKSBaBG7AquhN9fBOx
J5q6AEhqzHUDUyWI/vO0PE1oSZCdpuC/eWmga5jtOy0JMjnQc/6aWXdlG6XYxBW1ie+nnKR6e7Ue
6okgOiYnP4qYjpoN3E8BEzvl3xctC+xHLxPTGIaAh0E3+6bHb4DJ0eWWeloDC0oVLEIJ+hyN4vQp
lzqlo5TaYCqlsAwWo2pXO9FdfoY7TKqjQji0RNkps2vSygsJ8aUG5lL+++/4/8wzEB7a7IAt58+H
7SLc12XEV0zf/jtTndmG+HO7cGIsuzsYXQNP2rm2Gxut4DSsg3ZkwSThWDjzHqhP7pPY6mEvB6e3
Vk63VBz8dFluqNRZYozEm0+qnylVcxmGUOOnZHlOLG3EqA/792/7OvnYuqlw+3BrNXQyLEWJ0+lG
O6i4dObEUCzbnAG9cSNoFRWU57ARf0fh/pLxCbt1JHYbhVft2BPnnKbw5qqEaTEjywObdOv9ybE+
56UrKmcHIcs0zQkHYCxALalws/4Huf2GNQlJ08NSK9WqhLXtoEfsA+ZLRit5aKHqzAMDel7qrsoI
ZTWMjLiyj3fo8s0bBNR8XqgeySyzFQPA93vZai43UFb3aXVyoAVPsR3eGblRv/vEGM4jOXQ8g85q
3YIK6auuBNF2EY6yWsdNJhQiCIjifFw6Re5761OfA9ZAmITlouEt+t81yZ0yZFJdBsRpjE4cpP3V
PDaZoUYcGhR4y9LjAqKqr0rOTL9SOZP64Wegte6F3w774MmlCZ9DHFfhRl0iaz+cCQ208Lw03R60
vB5Q1G4t69/O+2bERuDVg5enI0WwSIJsWz7plRN7gxuil8OyIeEN4tJ62bRJDBbk9TW7WaV+xNHN
W+Pk7xhNOOuRJHguRNQnEjS5MlxcosVSsz2fL0nzvJWo0SnOKm6kFK//TrH3duMYDZN7yrLNOLmK
ZmKIddpqj1mkLhB5YTelP6Y06YBrQ2yJIGZmvoDa+NhTkXJaPvRSL+TOqTE3YWgXT2328GdVclJN
+bA9mLlPLv6mh2HitpEvsAW056IUrFXLKN4lUtTU6pwHiO5o7VOp6ZN+1Uq7TBeDSRKTO1swEUdB
JQJA5lti2jPW8VfYwZFv/k0wUEx0qZrZ1aDakr0AvpAYG7GsFFKmYgZrWjVyzPipuIp2Q150/NhD
sieIjG5gb43qyMArbD00IyS6LojAN+jYb1nfaQ3OApFWLTGtOFxkxnGxQHG9XHT0w1iUp27XDAUq
lXyH/1Z0GAXsXpsf1mBM28zSJfw6Cqvmu8lmlQY5M9iy3z2rBxXpSSULNVVo02dS8AUrRtbgJx2B
K1+RRR/cEZBUgBlkTLJr3E5qeTq2kB20gjfFRb+ChidsV5tzeE+e8dwADKUdqNyilqgZjp2PFnno
IROXJ2J3Y7xtrFlPI07e5oKvI5u2ElWEfR/6VKoDKpSitUxW7YTqBJOInA6lxQEiQABSbmv1FfKA
4i4gDYbPAg9tOFCd6iQi2hv0BLf7Lb46Lh4Es/j14OB1qLoLMru9qVnQwEAu4MRf8or/WZHZoT9l
vydvl7e01wBsKYhyCE8W+UtSg3kGRq1rBvwU/DOqpYjVtZcn6SbxY/veHQgLohvjj7gs3yajWJPs
0T3iYITdpHYLIMt+pMXE/AmCG4YeoFkyI5X7gXWJPfVoHmKj7uYGt34luE8wLXzxt+xfU/A+8YbW
un8I5ESdbAsh3LqgY7qJ99aem6w/uxrKsa+I+8X4NqjLt5MBEN770i+PUVgl3AG3EMoLCUJLKZTm
6vOitxJPowvEMhinUa2auouaiYulAV9ErWpek3B57zWaCwkbjPCdku1iw671xKSOfpm0hyVs1lZc
o4ZztjWG/2LfvQkivC4tFney7/NXSU5BEkWU2JsnAf3CrgMLJrNvLIgKtBWf8JS9lPnLIXgrUZF7
xc+M1r3mszJhw14lqygBuMHbM2QMUIeDblwqIaMGSQgEK8qgseir2DPISNPNv8UgYv/TgI43zCgG
ENCdwSK+97J8MHPfx8JUELvDg9y4jG9KG/n6HPYYxyDNaXKmD5LplMJW+dgkTnbRhmVDVhGFMQ6W
FVnj3W2SHSVr1c5xRp0Q8VqbsHL9tqx9KeexZZuhnymfi5zdj9d8NL6ITnhihh9yiL+ziWKc7p/X
va8wA44LYZOX/12FQto7LCcnz6uHndn+I00cO7tC+w1b48shvtyDI7REk+x7EodAbYGiVf2tAyY3
na76530tXuH1BY2R7rDKIFfhiAiu5jTQwBwbclaVaANvfFBbm79ZW+eyTTCMwF91slujIk90r2p0
y5F9BZMvybOEJIi6AW7ws06Mwf/ImqU1cKtxaNSGeCdrfAiMx9E1NKNH2kGQjRHotKDTO3IbfSUP
/EMMEU0kelosYhOkS/DVfr2aw3ipzrDckUj/V1n9zx9+cO+4HqVMXJ5Qwq/t2J2yIrWy/FlNK4tB
y70bqBRivYP9RrW/UtaUaDIUm2AVs4gsRGVpFf4Bo6QHSGmdoQQnv7p0iaTCkTkH5ut64jPsrIKo
9SdstcSQn9K66GW8uoYVlJWFR2GO3Cf0K7uU6ImjiK7+U1O2rnkqCIG1yUP+xhb1CLwLo+Wx3h7p
3Xd32T7V6xW8OpzkqP6Pj/poATy66Qe+gNztby7uBpDMpZkyyrRBT6B3JyJrYKc8RfU4IN51EDhg
r04NyWpN6j3GLwOVbA/4JEvQ9ItEq6NfcBP8I9xqbimV9/623ESP48G+TR7C3yNwaVVaxSue4p32
K+tAnvxg33dalfshJ/W6u5V6x/YqSLExZ+1Ep/n/z+WWL8gXFhCoJAdLgDX2eyJmEmMGlkVXXapS
4BeiRd09d8ca8KzuGK5m4HnvA+DiBSS1Jau/MfRyjMLqJFFmuJcuJGe2hkv6EDLvkcna34U9mpOF
HMlnCWLTuwWZM8qCCKJ/YGpiUGC1rhT8qDm6rHCDOkhDUHh6JtknlAl0FqA+VGc85LPEDYb1adan
tGCUlNeNeWQBvg71BWTtfMA43vsCeCeP8It1bX0twx3K3Vvm1tbH3rq0aFZuFwXQ8+r+QCFwJPkn
dCaShViZYrLGbyRT2v1L181e9WmJF68YRO8rcu+l1YLCK3MVvsKmkDzBS2QnH0c6XJ+yZCKfjA5z
avuz7UXEutwXS42m9ktbPa/FadYwCnMrH/qXR7+5HNlbrEduS0pBB4kM7FUGTFpxgnIxIFakutPf
NfvKM9cSToNEfsReqIMC9pjEgQT03/hjilcNgdfrNKIhh0Pfj4ft+w9AORAgDpdTLr1RfzykvgHM
mXXkL/rArPdangOr4W0TsnEHv3cp4SBuV0LdtxkWaoaRJrW+cDJGo6t2+wTTd5hKxc8neccvu4Ct
ONd92f0nIs1TfS4YKc8HnhK9bbdc094nD6LgRsgiO2WC9I8fSz+3rYKRYCPKe5lN4v4Pc0BmQadx
/qIY+09bimEW3Fqo6bMhx0o+n8xN5inv59WUCziahy0+JoKTructRjTKdqWfZwlvf0KspunbMyFv
F5FGeZpULQr3FKMsfBJFZIaabX2FGuBTMVWYphvfNc4ZqyWqXfW17tevSUhnIOnk46Am0AkaE9B+
JMSAnn+8sBnbPf16MTqwL3JwyDuFW4Drh4iVOqqntqblvHt5D8lemFJbitmU4xt/oDpzowJYHgek
l1VWvM0sJH1PYsJ7DnRMAxsPrJETr03I62Jxax6PnsOkHBLpgHok0I9njFsr1SKFdOAU4iIXJboS
apuSGaAqkDfn2SPqm4mQ83kS60/v52Ns5IfTSgLLSWwJ+NC85piXyYBIh1rp12j+xFPM4VdfurTR
m0Wte1hWp+aa+9lz9ZlIcpQHT6Yc6p8WyxeQO0edcA9Rd6g6FNvyMZjk9U8RLF4hbMo0R+cUFB0Z
ZtofqK4LgpbYH2fOtnMOgNix4DwhZfjQ5bbnrN/N5qto5PZIb5EvJglOUfGeMXBVZ5hloZAajdNz
/Qxg4bEtx1QA/ST5FI6BKUaNAJYj4tnDBbP8lZUxDMXZkXQ+v2tZY/OS4bOiLOlORiOcPxpi3Rth
wI4j8wH0toudsMrFoN6nkbCQbBBqEeK3F68B3sDZ58I79l1CyvBhTKnnKdfm9QswQ6OgMyHIrJDn
7IP+iH9iuw891JMk5I4vsS5h7iI/zy+txS1B2yG+YuBcviex/NIqbpft1XusQTH8ZAC6KFGEG6AF
94ym0Ypz1Pdbs1HE/TxDJQSUM/E2g8lBJEF8a5vAgNziq7BNxn6OgkRePfvXlKrwb1vuyQHKV92Y
3c/aCvhT4TbsbuM4/RWMWTR4rPSQcS/aoBFj3+njwkngYfob+UtJ7WUaGPajXpXHfXMd0+1/0mQF
TyiWTXuVHZwLMZ4QIbsd3lWpP7jj9TWuI1tAGdPqojANf2UvV5zB+M8xnQv7Imfrax+aZNaynlgP
Q1iNc5FL9cgNlaaMn7a3WO+c47f2yyZiOAoItyKyOf079LbVyyym/xWGqlZAsCDBmn1duTchZTv3
Vt98LFyrBsvmqnT7s36gn1eiwl54HsQsTIBbK492oFBDsixYh+VThbrd4FpVUhltSRO7VaaArWi/
T8QigA2/P6jzV4AWB+l/TbBxE/dZhsBYdiurnjuK96pTSWAKrwo24nEcqq5lrLSH7aKH7TsIdC0Z
9eigOP1OypI0zJEleKss1d4HtAciV6U8WrTZw2aZJlxXr2iGmbzDnlagM/jUCq1yphdbGUq1YYfT
aKgt4xgvr7q+3PSqwqxlgn+v+q8L1WYSDDykqDOUpmIJWMLwQHgo2jnlvM9CrLcrgvkz0DyJmly8
XlC8j24V0cqMJtAsVugd9nI5T8OvgC/w1qYNBYe001MAHsQYUqMUv+/FAoPFq+6e2yCMj4D/Fsvh
AN4UNy1wY3oUL1KcoX0zz1ti/K9KFz/r66VGmqFy9otgJaa0Vymzf+XksmtjE3c5itg1w0m918n6
DVx/HfcDaXppKZ2X+z6mWdwgWqg5BBj1CO3EW3b9vVNqFHWXPZt1RtWWDalvr65iAdz0+gx2OfvB
mXD3jzTiV184L5aa33BoCbTrfLz7sGV2gts0P3aaHHCrohSGIrVZCkCvUZAzLvK1nH+zNOd9JKuc
+SUiNes1M04QZk6J78u97c7v7YJ+XIBxOt+bdGvnXAx2+B6H3nqnsdliaVeJOVJFm4ff0dc05UKY
2/Ju0ZCuaqs76oIDEdhCQHV5xOr3xHG5E9vObSBS/rr67ZgxcOZXBMQ0eNrcNOTkicJc2d5SUH/X
CAAMPyq//QTSmifygWMkiWUnwE/OwON5CeKH/Qw57MxlntzB9LSsKnPbXXiLY63t3GgSO0keSaxa
fouH/NE31ji6a/uI9TE/Jy3uE9/OcUZ/DE5jk+bHdQ1zb+WYK235qSN5Ug0oWhnDNlKb8TFnk/fM
EK2FtmeF5zJcsimnPR1pgUYqLO20wWZM7HWw8idODWbESDW4f6SywnyMUbQu2zN2jJjt2gv02Pfz
JxzOPrvCBnwChSIt5gZ7s9Y9cI5S1RIzkIibh2Koc5/diVcfBjWAnKTV4fdU7csC634/NDEV/w5s
JM1s27f1Qp5JeC0mLb6d/8YloJhm9SSwtYANMiEgtfO3WFzHMSBm1kHj4j7frKII9J7qYDooIEWw
JuYCHHluvooBpX3QS+nStMRMvLZs0qOHniJWLH9c0iaY7TSEwaOIt/frQQxhoP5R0UhFeUw/E8SA
yEVhp83CdZDcsbIS2uiCktTD4W279vPqok97RyCqMmyDHX75t1u9aspIoo6kdEsrkklyT7dgr08F
UXZw0J/MOF2j62oGkN3uUSpmpi+y4C87iZlv+GnpgIUj4SguvHV/AD7LTHSbFhACsAz0MXgxCbqO
M5QN4que/xJsdotW7K9ejtD/K7HernKlLa8ojVWXivEJqdL0R8z7eEbtuIkYJKXQYKA6S4qPt0oa
LHHuvlqPe9MiEl87JT2McesBM/EZqSgCveXxQhxCdYSCkwcmCnHoq8VL+wJKmCNjG75v41CL1Smd
UHSxUVm+C3+3F6Ut9YO7WDFHj/5efwaIbgBwdPy+7NKgEUQDEb6djoqa+fVVIcWkBZh6m7ii8Ch6
kE5fd8Cot5f9DGnI0UUm5J0eM6wXMzpnXaSnhEbfEcpkPg1EW0Wngd0m/OIAkaatssILcLCNsop5
/FhIZOVf0Bo1B6lzm5cwqvCfnOqr0hbEj2DE0v3G85RysHwr0BDMzAPjEZ0VFHxbpjcBVCGL7Thy
WGxPGXTY/nrFkjCF0oCOkOFIKHymJLCwvO4jZXeZkiMyoDuDiwiiqzSiidluw4NSOsZG58Azsj5w
HCeWIqsEVU5SNCx9h2vdAe8f/WB8RD7C1P2fVaUxGu6Xk5kBXuCQM2QDvCM8R/mXMaa0JQ73ebWu
qODaZjL0Wo/WyKUsDHqSn4+ehhM99oQkvejJQrEaTriZDnVyte99G8gVf1L+HaCaLwrSXZj9DGv2
1gDKIYyJkZ/uexCeVxBSLivzHtAVjUUvbiW5n39HFgQYLP8i87K3gt3phFdVOkclvF/aNX7PplyX
GGZfbzY2ZOTjF68r7yZHFJa3Br5z/Y77HQgPhz+8lFhSzG2fbH0BUH+JRbs+1yC1EPwmIb2RA9gE
ucnBA20bciKjoSdfZbZt90UMviLpPlWhMSjgjVXI7OYnZCyhxww3/CczvCHy/5j+HQpf/SAdOYhL
XAdrYR/Ivr/DwtFh7CVnizZ5niBay/Xj3ZmaWtvFBdDYpCZi3WZ4CBxq0Cl780rEt/QkW0XnZuLz
/pSVT/whLBgSEpc3V7cS06ijVG70SAD99clRiNj9A8yEh6pF+WcDf+MQ48QIbRBDEMVeKO/VmwM/
Uw8B1imPz8fwWulpSiMEdQaSKsrmeWoNAzyXFXjsALM8+Z8wtavvU02faYSJsHiguPFtCH8DU7aI
1bOZk6ZPkm2LKV6svvh6dxsA65AzwIQAniqLb2b1TzGslYg3yfEORZxICOXZQazw+xNghi1q822b
N+xqxzGnzjfAzuvC4UMXVZdPbg+6/hjCQIF5AaadawCm+gAvk6/Trhu+A5IQ/2ssh/0EQ2sXY20K
WfU/NaDdRhqN+xGAKNHZFWhKWTSshpvRj6J8uy2GLOXmKtKQ3WU+7iY3SeGmtzW4E35snXsm7vat
P4S6bYs+xUqsJViDLxa2PyhCUNn3WhkUFAbPR5OPBlUGm8Nt4QVTYlbp+oJc+ZtrAqrnxRFe3Giw
I3p4TbQdB7gN8mrB+kF6o/uZ58Du3j6MBz1aqwdBI8dSMGEwhtSZhzfDN2qptu/ryb14WrF92l/Q
jURZD1s5QK0pJs8Fx03NfNM3dglyUxBbZsMNv8X8gVqqojs+W3lYQC2GK98kWCLYZlX2cxH1Hwjs
4yjFgtrgyj65toQCYXUaC7dwM9+m07kqfSsU0UIezmvP/ZUX1Jl6lMM5Ia5vTXr4GKhfbh3xyrAl
s462Wu8y7N3JCjauTGZOuWuFSwMlHLtAGg0Cxj/ngGGcXiFZfKWTAlvQSaA8cB4cj+pJ8Kid0SY/
SzXN9fBZkJTjsXKn4+tovBrOpv4QD1rTjZ6bKBNRd3GpsIt+1cGHaaCx07+454fnouWncqgnM9YK
fJzI3M/I6mn5MiLxSIsiJF5lwzFber7u431skU149RBdAwB4vE4KNpPs63wETMzflGocGVVmsBIg
aDlC6ocO2HOAd2ktVRfAMtuNbSEkYZKzOKxZe/GCDCVLOEaKI120caK9wv24sXTAufxPrIhPqFPB
rZKKrb4MDD2ac4ephdI5jptnQcIhfr+3fuXhV5RXSTRsxvD+oL9+vtXa+ZvlqSP5HowjDKH3glMa
mEmNd6bq8eieZDh6pzRKGpL5ry4w33EDO/asA8g7Jflqlu9tf357b2H6y4yWLCQBpuBU633AuKhX
SD0Jheov6k3uzd8yp5T/cTZNXzwS8qbl1ptWKdU01FtP4B2F8qXOXhHhJ7V5cxR3Nf49ZI6MNEPU
fYXIGB6ZSrB9FnVWNzOs7e2fM4P6sCWZesnFY+9yDsiZLcdGPbNZa9gkZwd/lrdhoWwsR4j4Dg6u
ihADR7sCesIIzUz/5hOQXWfaJMfBlHBJuD9yhn0DrgHLzena75r5LLYeZvySRAold2cUFwZTEGHQ
kRW9cB92NwDIY3yLnZNjWqT+GnFuwefjS1wrmxxqrXCA7qyL3bcQPO+XlSiMCIMWA/TEmCzHrBxP
120UeVy+wAt+5hASlHhtjLouhSSy8hqN0kOhDKvMwUZC5k1ncwVJOpHKQA7LHmA8OAmGZkxctPWR
4aCX0uvUvX7RfZekbj43YdYTPNWdnoV9F1HKDUg5Nf4pPpA/Ox06fhj6zWc4zmAYNo0CpvYV45+W
YW9zi/5FNyRWN1+ePlFV5qgpSJWTvW8GDn9lIrmB/sXVRIvXtlMb3Liva3NsU/akekIZZYoIF8BI
pRe1LqeDgPOPw5g1jrY92L9ekhnfplzpX5zBzLj+7Ly7rrevVHwT6bXlnYK4KrRRQghjK/QJDyQK
9st1kASHEXXmWx8nF8rhug/TwvB2Nf+LGZdxAlmQKrtJ32ayzFS2HoOcpSomvukm9pygLNuYrR6E
ir6Jd4Bf0gbkO6Tda7V/k7UmdOVVKtMNB8dGCO6Hx8rHw6nJUFa6LEGuKv8ndPauTpIqWhAPRQAZ
HU1gX5dXINDUdUw/6afb67tGCzH5va8wnSrVGhp+LSh/WjEuB8upAW94sUGhAgfPeCWl8v1SecBy
3yTW+KwbnbewQmVDExsGp2SgQLY6nKmNQcXStVmhTo0osSM1GfUgEBEsnJZo8RCxh+VzJU/ADsDy
EMCsOI+/13Iscr5F8V6EhrpAOeQ7pV32x7gxsZ4xW+z+AF0uiAIA3kYzOmXzR775NcvIpV3xK0ab
EbG9Gcj7zjwNuiHrqp9W9nLjzR6xlQADGEw0gxHFrWysUCTNC8CwErKUdaNiBR/pRDzwKtSjyV8l
dGRsDaSxCHtuQRgGLGDNTMGdkU1JpH0dyItPdrLzfd1+y2VjBm0omZxp1Xjz1NwlOIOrkb0JGmTb
0EoOuYpBcZJUkkjMs2NaHd48Apvq23x8msL8jhriq4A+kBPVRJijtz6qJvZbOPq0Kffhs7NaBpDw
MEJggiys2CG5+h1i1dOiJF5vlGp3xlHPRZYc6tgbWr4Mmqk+2vUJr3ra92XtZLT0P4yy0IcrK04D
q5zLDv6PiF+NXS6EOhEvP5SPG/O7pgSle4cOfCNti8F6Qcsi0MaVsnIh3TInKOE6LUq8EhyrDiXN
ZB3edbo4WOMOjNA8sB3+36MEJseGdt4gBFKXm2oXra7cR2yHcgVJNnv7JaJBlrs8NBsoLk2gnKzg
YG4ZRVJQw1dCyetNNnXgqDEXvDv8oJajYPQ855Wm7FPygq0uBxpsNRSYqPHJulWjyavR5oIpRPBc
Y4Ra6SaCFR0VBgGh5UE4FcQJLeRXu43LQWvZOGuAFSS0GiR203/kRkXz05o/U8BNzmQrqICpaykO
jn/ODe67ehQdaafxTJdv2QjICAixXjQOTYJVL+peIh702weLH7dYvVzef8Td345+C+9fgC1xgJ1h
sHNG8sxH4HbatqXnLPDyAB3RnjF9KK2QZLPXILKPg3vO349O3FRfyrFwgCO2nKm46e+DmRAbOcwh
nqFEnQZZvw7Wddpsg7DmvURvZFJM0j48AOer4TstpCnUq2VT+XG9nAhI1FK8RMtAoHdLFUI8C5Nz
zW8HDK+tg5j2EsXn+nWLoyGU++yjG28ZznZ8KHF4kq8waCh6qAWfqBytnwRUlboEY/QYUlZr/rMV
VP6gTiuHIfcpvGiwSqhe7St/2sj3zSiPCHuAFqGC5/PmwiX09sH5VWUxjTi0o3qtB41WV+MTFB4/
t8POENI5F5v6Mbr76pERjmdAnmFPim37PSSvxeMumQuct/+Toeu79g0JXpNZ2Cj0Y0S5l8vQ7gV8
1lG3WRu/QSmY+Voh0LEr+qVe7xqD0DvTKQS9Kqm7dspbVty81Hkhj9phptSZLmBlR9Dd5ilJPgIL
VyJYGWnFkYiIbdqB1nDRnGXUgkemPFTx7buC+qWIaWZsP45b2TwAXKW8vV7WMGhXkYz9bW/9RYSw
Z1GC9ig7MT9Md8N0AEt0YXflrT9xtuVhn8+APrti4sbZIGulv4LoE18mxUdvLz0EPVZOl4xWq+ps
aM1s4cUZgsop4mtMn35Lm+5NOmxLU4AJZ7GYOe3T1Gor+uM6ew2cmLztZr7RxHGSx/s4erwouEHN
5vcEnwoe2AOkmwIaIbvtubBF/rwH2yzHhzlWuaJB5q299pvZgjUvlLZ99TqE6Tk8Oc9PVk1w5lLM
ucu7ktoEDX5/MTNF6clNsrmGqdB66tq9d2ac0AqY14gOV4K6plbvnjPrBQXiFQiBBN0gamnygGPs
iZ54nsRisMR2xUT2Ghc97MM1z4vpQLsisaFhQuxzrmPi8kWqeyaM3tWTVjEnEDNnWpPHw/nYJbh2
9R7e/42W5pmUvpk77XG+NBZzv4nzOxaMDSygh59IjqLZT2Kek/oS8WXDPQdgOZpDG9Kup6ybj/Sq
/i+Q5XEWs9HS4YstvqDI+OhAQGaLODWSVurfRm5TImvyMU5mQLuOz/xXXB6lQg0AFapltOAieIFa
miTO7KQJmHiTFlJL/OY2LErSOAF8CObKey3C1buBs5DNzYvGDA1IlpPA0CJcU8SMzUm3p+WwqEG4
WWtbHqLGiP95fhj2Gj1s+KkVTgFX096AOiBC4GuLv2i9c5GSlx6OHGePm1Y++0nvKYV+B1fym2NW
Yft9hys53tv7uoCuUNipc5hVGbKh47ilK8OJCBQKI+VDGyMNnWAH22sQisgl65q48vb1PWpgIMxW
9bZVHmJx2KzJSQEWrolScIskDSOSJ6w5fjGzwxrCLUC9YTV7AIfKHdiYDdBQAlmFXHEjZEhXM/BL
qdSytFL6VexscK6a7DUsEhBgj9uiFbCEfK6/hBNmRwvAcJqlULgIze4JUyZbFHwLBLAiN/l2l1ox
atz76kihuYx8nw3DK/f7lFaDmb3TgEtBIwWAhUszvM6VDHxLrIbxVCWqzBYUkVCRoHK5wySY4TUb
d9G0UC/mPSB8h6Pf1/bjX7IKRCHp/jPQWYkDzPp9Iam85/WahtdFkPu4Wv0Y3jm04tbXWQtDM6ED
Mt+Ntis0bSx1dUnxzrnBrjaxCzn6NyZ7i3/rPvZ1TtLWsZGH0pVHPNhmqg1BlkvQ8w/jwnohNr1Q
ZZa4mJphEwosWXCfu0sS7UYLMJCNQXumD3DKi5kQRuofCZCqt0XnFhQpRQ2c/oFjr2hL37W4qjE0
ZlGzDfdBGAbptERh+wrZ5/+7+mXpp7nces9ZF5feI/mI9E1FZr71osCaSwmcwpQfYgTrXOxkmkUO
66aqZNgot+65gRMHzZMTGAwEYtxMh012JrqOm+3IlhqUhD0QaHI1YAdDvrVyz30+JcrOqYIcFLeB
FgS1EY7huRIXsiJhgLQ5/rxnqsNiuC0/2bCGJjuDKOkz2m6SSFuGndQHlrUWRCAybzhKN3uQbzUw
1q0qZSxOcH3RkZv4TnZo3CZ4aOQTifssrws5a2jZyjxh8E3qE3s1hRfPXOaJ8QjpZdNFwtH0KG4A
ZNctrRrVZNQXoc7AnDrW94X0iun3NgQAmCJnpaCaHHmcnAiZ2mtuZdhPd4TkZeJixkf6qH0tn36A
ZHzMmXHf69ih1mM3Wd+wI+ovY9Q+j9mjceWgSexVTGnX0dk1mjqbp+MeJM0tljZEuvfB33OJoTgr
13PxjZdISs2lud8L7L8+9A3JKkQW3c8dHrmQurj/5ccYwsulKoUT8I9ICqzgohetV7vz/5QQ5A0n
yyd4t0gjSvqIteVHGQXO4P98NAAdT6lFiYszs9z6iJG2pFW78ZRIGMfm2sueu6V/S8vgeQ/RX8AP
cTz4bwLVyqQ42f4ckHoxMBAmOPi9ouY4IVocblVEDtsLc4x9efL2Bb2M6YyZqZ6GsG2s1FynQsFQ
+dBnWTAoUw7/3+uwMmKWfRZOLUoD/kq+eHp0Gx44nKQ/HgrxlCeuncZEKYMI9pw+N4G1ueLcYeHu
sdyboei70SOAE7pm22WsK75CTc7+aO0tMJgqlDyC3mByZ0/uZgCZZ6PKYb9FnKCeHulmuGx81i2y
r4a/PSkNv3m4+jFy1N3Ktj/v1EJlkP+JAsAwL/e0Sj/j1twmDugSTBfPAC9WK5jVrmhRboQbzdTv
hld4GYdqKDYpo7vLQwJQwq+Ry9BlQT0oiG/EP0UefXx/0z9OiS/8mbKAoWfwGLbJFnFXehQY7NW/
xV6VADEAHicwmO0qYT9HrMDVfBqes2IbA+SGokJIASWUQPUKp7MBFKAJB6At5sJwAjWDpnF8aYqp
HkFtwh9UEK9JQHZzaE21FyscufieCN3MnQY4Su/6uBHCQvDIXUgaPSCC2Z6avMZBfudkadIw0khj
oA1ItY7+3bNRfDaAmjnEh4Xx3o872auv0/+UicaNkHEQRHDL3bhJmS94D+EK1ac4wm99xveK9ewx
ISXBRndJq0bUjIbW/qzVhzG04toWpOy1F0gHoo9fEzEynD12QJjbnbPtnloCVejXOCdsDOBddWfJ
yL0dq4est5Lgqu49AYeZ5THE+cTmYVkqnIYJjEigg3yUOMq23EEAyES/+fMRX8t+xT6vw8BNbkt6
2nzsGaUS37gdUyjFhlDGLBS9rxnAAv20rmlH7j+Zlamp/D9ndI4+WxbpOsWw8Li48ya3PEtfXbqe
7PkgDi9I9Uk9qeYWZlH7bsLBKSyFxPj5+JMZd8wYGMMBMWUTmmLqRdFQUPa/1iw9MSm66r2HhfyL
MdT8fs6TU2NGpFG15Dar0zN91aN3/kqYurhF4PePbIel8joAssL7AE4Xh+U3FqpQ4KTGntavaI5b
UTwgmPMFn25hhzkuDed5uT2IDRJ4HWaRqrB7HHUWviAcWqBcoEw5KJjwG8nlRgmJ+BAkSuOTZg19
6L5NYi2MFiHo9WZDqwxHsP/O5ZQ7WmhAdbc9AcDEXB9APjgDvRHmNqAzKoD1ujHYDxB4jmivQYwf
I25dA/LfxxjU4iaqJ8ISbJynn3iGkAC6JvuSKxBjHzyga+uQ9TMPX6oKMwUoXFzP7Up+ieLJt0uT
39nVVXeiF0KMU4m+N15R7m+Q+qMBvPGD7c1FYAqoLYUbVho4ZdHclaqeUAfZuBeNpN3XjdgW08Mm
FvLvd+5sjCcebl1g03xAVw6c/HRtuXjkj65yejdRqQzv5BDorhGusfyXJr0YT+JPWLvYB3xW+n21
3wrY8rsC1+3O2ZKwGb8viItiTY+ltj2mdSoYBq9LEgMTNY47onRn2xNqy4f+3sXp5lJXxJRP+qKj
9IDFhu/wgaAyoB1cJXPCF7Q7owJU2NZFatYpVDUsvMWDVKPAw+IlI9zMh+T2mrQ/O3l9TAhEIiTS
ppPBoow1jB2Xmq9sTsYTr+H2jDiO6pfT7TotrXtc1FB9EyxawUhR6x2ZxP9mbta5aJ5MzNwFzJcU
h03i2AWqA6v5vx/XWj4bvNuj0wdKSa5n746tMofPHeTcRkCkt08mBoIFlffy2nvP5mE6qACzhrlo
iFYN2sXQACLOLOSxbNQlY16Elquk+EnBBM8MWIt5O2ot484rTaOoqe9n090sLrip8W2JdRC9dBgM
ggyfj/Z9W/7IgOccAt/KjlNC0hA7XdRindql1TytwtJQUDsGD2QpMDCx8G+RLOq9MhKLzXz6Uw9T
g/tJ7u0PKwxAJDrBwHCSGCiY4v30SbPItUq/OlZYR/OIKgEILgDepSFCpyebf3X3NHxq2cYLO2Wk
hYNVlXPyu0SJgTwsDjIeunGdHyEFNCk2REMwbCpLgio0jlNcGX4f4lsllBq9nriL+76+kUfJxB7g
Xl2ndOxX1BDj+JgHwsibW11woNDdYefuagixpx9mlUZ+xVKeQSRHSUCvPwHT5gGjsWkF+nLX5qjn
7THbw/Wl0GoOMgEtiBvT5wxO64ghtdjAsTbVGnfp0Cx8rKn/kIfutiCTPa9D4uMe6TalPudRO/mG
w/e/UyiJw/Lfzpu65CUUJd7ia8jRvIgWiPX5heKEuVh+bdJ3i0ZeRHd9YcEeB554aDhpKGRtkqKV
8/vqxU70MeOAqci65q71ity84jvVVSk8i0qUNLLXhQJYpI1FXHYvD6MN4xplKMvGAu0J12K396s0
vUGa+tXJIVV2Rm1X6YDPwicmhqHeoTYstaY9byoajcUHhcOxgjr3NMLph/g8Z8N7te3AUBWz18b9
2JqvX+SG8xOt5IQFWT4P6nGUyg4qEZKWl1jKZbjuD6p4b7F2+jZzfFsyt7yCWU6wI1anExUwic6l
9E5OvXVFLV/MsqRdyGxH3QUUKqlNehOBZoNdHM0v/Twpto1P517qIz4ANCfM9SYLKLajwJVPa/U3
l6tha7ohmNoi3y5DAxtH6A5wFLomAkfRt5lvLkYhHfa4f1sR+Wyuk+RBhUuxSBCHjrVWf6rtqj7P
nlwyZaXRaVOIhThJb+IwgcXMRpQqJsJCTC8Flm2QEhIJ++H/vCzgYk6obwmg7PQ+Kl+0pMjLZT+V
4yt09dFIaNL6HHx091gi95rErtPiKnoL24dZ7iCU0s1VrOY/ui3U+8XYR5KwPaFa8q5OO4QAOR0g
UJUJz5Uq//5Nyhk3CqZdq5SN6vZm04s5JtWxrkn/mXGn/duvhZLU5aRrygXQSJG8RxIAlZlDn7ik
JITFEZ7ASTO6Xs7tzwTmkED2MYxiKuyLrzvOBLHom24l90yT08l/iamnPGBPRAsXcWt3xZS2HAG9
kM3u25w9JzO+lRxOxHJGIOv42pjHiXVG83BXnge4WAn0leSOfNF5K8yJfDfQYVnLXCZss7eA5pmr
KSuXuJ99sWLm6EwtwBsoaVYDbLfogyqAsatt8LuurLx4CXtercitmpvJMxBCnIMWgK6BiA/KqMkf
fI/S6jZD4LiS25Z0mCfTrD1Fz+fR6px6JKdOkDjG84+UVJ5wqbVeaAOaxVHHnVxYO0cKE4U2d9e4
i/HW2zzkZdllEb8wLFdZYy4q6ZSuwWJgkzwBuMKyK4y9eyyEiWKgDSENXwjPWCGa2g7v1wdDhS2f
VUDf9wxvkgH0DXyEY0+cV6Ly6Fpk3tEWDmTQWfGCchkQaXUv2NpxmYjNYwZ35dLPSpIVWpVUC238
fx2LA5MZ6ITF+b+QqJv2SfGw4MdYrtJCJ7MoohNDifFScREd7BkGswI3pQF1SgH7Rp1NyeqeHeth
s1i9c28poJOYy758J6WVgIFAb9kzN0cRhAFXYSjhFthUFfpZ1eSRNoZ1GskrzYjsqTTB1ZRhrLmv
xRn8FHAyHNpHRk44pl/mlUFKNHAAAikMJUUQ/OGStMsQlegjICo+l1NJ6DbAR/OKAifYEb6neRdB
oPUdxWIF5r6EeNxZhN05bcmk4+vQz8ztsBsLwxKfWuQhukGGEFeaeOhCyMGBqtMsjK814PM5Cj31
fbf6/jS5LN6Q56gEulgb7f1rljlJeqPdMBOIxZ/L4X28Y8RA5e1vu+gAPAHNqjny1ytaHJExMXx+
pEahqSAnjm5LxXaMcngey0K8bDZQFGuDL9FLz8pNQEItoPKzhVGCS5XqFU6U6JrT4ixe7PbHvl3b
JeUIAKHIEk66YifNTRRQalesXkYa91lFp9AaHr9a1eexEVoTP2CORQ6+xe0FI4CpCwETj0Lkmr68
MfteGj4/mGGPa8wJkOrzpt0kbXLUfLFtHeHkeXfVceU2oMFXLB09eR8QUDEYi2cuWP9vqrlrGV78
9Jegfo7rHTimQsUciU3+71GWFlvDlZcLK2T3YtjzQx7r4PLcAhIA9Jvp9QGGxVEY9ZtCjFrKW3ov
+U5Wqnge4zvhywttCGZi5y6jIGpqtc3Gn+Y9EPIeqv/6MCm5iIvSQCyn0PtdjMXOnlLJRXerKDUu
3rn0UgzGT/JL5Ri/IZpIhwa2mQrsPcfbH0ACOTazQpaP2zWN09n+uGFn6h6cIFFah5R4kBxOStXi
svPqmdTsBii4FFTg1llVeeoioZgoRwJXGa2IdxbnZf7cqulb0X0A7vwjIQcTwSvmNgR8hBUfQEJY
oGlJ2LfjFtbpQFNepQWY1iJyKweoXBCB9dRLprG47DLIqQxVonJ4/pWaeVeSRuRMZKXN020ubD3w
KRkXBk/pQS+FdbPBoR4vi8M04I2UqnUvefRxzPctENsi9Zzk3NbKpkQuxgbRcC4CFfatUt8zo3Kw
M8QQnPPH3og6vJGJ3UBwNUFJ5m60+sZGhMCsaL7w/IFy8x2ut+LpAwhKcFRjUWRNR3x5hmSp82UK
TUC5YJaKjvrIA0Mkoe9a/XLSTI6CZoces9s1xqkyMX8vi82XUUGyM366WM5GSvyKAF+Z3jXEiJ7M
MVkqoroI6r2N9FRyU38sduIAAez6lh7wiEyeybFVhIZTdIzm8E+VpNtfrQp4wNF8PAUNQQytslqF
e3Yyu+RtiAmRSkU99sIdMMSX1ncTlsGdeY+npSo7hMxQNsufXukngHTqeuQs1EPtmyPBAJqTB7Zy
5V0PcdcSB4kPZS5SFQ8W+KSvqoyqZPfxSnk/1pwhv5UWBqSbzTD1vfkYbfbL8ryTS87DkFK2ypJO
iy7Cx7w5hmYM18syug3hL0uNzNOp0XPDA/ZzUoWAdcA1/qD21RPNWExpMC2Ijj4siPBXU0thrh4M
1TeCUvt2wwahxvZS2WVy9oflk64uOxRcWvFuDmoLhLgbMCUsLGcKPczK7pG6UbIkOb9bvgfK7ra3
3grc4ec6QcZ8vO0OU6R1MEStfBDzQ8U1TJ8zlNCTe+9W5ifIC+kkPXgAv657GcRMYODGL2j2PEBW
I1eql2G/fJnQURbvjx9sZAHZ+isxDBFFuciMoGO6qIo+TuL67R5HTyAuxo2jHYa0Eh6aPLmCldUs
c+DttHmdjZX6RZ9jkcUGjzAqY8DNaV2on+QCYJTVRocktw+uVUZPX5E6IUrkufaAd0JDQqnF10gk
fu/PgWYlJ3ClkyEoQ2ahUhC6M/DTe9jQpsy6s0A/E0+NUUr/E73Wfrq6hboS5FF5nq5GVxr+oG16
DQsF9nCY2gvd0Zz1O+pxvK0jyDPVWRIs9IwSnj9dewB0BxfXuN3+kYQqg3oNOQgs+2XEFyiLSH50
zY4kbwrYA0EliNuko2yB+Fv+0T/81Vk1fZ2UYm/zyojTJ3P34hmyAHFYEoSxO7sSIN+LKj0HQ6AG
Q3ZXxdVPWapfxWD4fIzOWH028PmR+jGZDOrt5aYdZ2NzaO0FoJo14dA7CC/H8/a9UDds/VeHgj8v
0mrDSUm0W4DfwJwvfaMrK8LNiXmNepN0flaq9TArV8GgxhMTAIrp48XzxMA1MxgrsXVI4eGSQdQO
DIpajc0nG57mEYShqo3/U3ip68ZtVS2pB1ANM0wfnjmb538K7L0Lceu/Ta+beWTxxDIHX5yyH3RS
rSO2+xOn8WVyt8J4TBcAlxF4U1pN2/aEbIdloUamax2ssGTfJIXocFJwd4cTmhy3rSPMCDk71sMg
NqOtqo2YKd9qeYc1VUgqYDDy+fW+Iuo+ZWtRcijqujUzlAxeFAG9ak6RuWp8n4N1T0ioxuSxYVZS
3Udhuiu1uL5CC5rHsqlT0V37lYF5JTRS8gpCx6KSiTqY8q4xWuchFLCyuJTSvq6NYne78fU3viUN
Q64yzOZDsJNUPWSTJFVCb+gUEKB+Is0sOUYAC7VUP5wYYoa9ZK6vPpt7iLVi9oh85KddXnsGHghQ
xl7c38/h7GJluamgY77gGZeDvIg5Nj6us/pLZEEMfldzHogT9ksPXqaFfHbgxhkI87MUZ61Wz6UG
EUnOnF3yikugtMZNmc8TmbTq20lFkK19NE3QqmgFubIgmGRNVfSBhL5CZbae6fbUl33aaME3xgAQ
FvHlTtlvAa8yhcMJ3I0G7vHC1yfNVOXtmHhQ4UGpagz+1LCMoN86JJb9I5r2Snu1FrI86A4t9BcE
4eGr7oirnPvUpJyMCBvVhAC6d0+o99cbMHNtfvat6WKYyhFYML0I2uubDyJfQdq2GmsWxEfxzbdL
59gPMm8QNVfdKQvg/BdtAP5mBaDMecc9i1y70jc2CGJN8NqjUiJvuK8aJRfGQsi5tuk6sKeSsqnT
YdCrCUWdw2PqOsLUiCBJion2xkD4VM4aJF6y4/b7iCGmCAvs4wCvn2AwdDOXW+HUDQWT6ZJI/jXl
7TtKzzT0onsPRDUfR7PFdYHc2IDot/5KWJyO3jHrlejZllXZanyYP9ey+VWR66y5eplV7r+HbEjR
cQntd1u/h2PI13xghsxV1jsn4RO0eXJGQvk4acbw8c/+4fZM8Jb+rcnI5jnJAfPg6GHK64FeS4ZP
i1tygY4vajupRFpGq5yP0A34ipXb09PVD78ZdEBdlxnkqa5h5yrbZ7aDTqXjOyVL2mnzbagzuPXg
/MoewmpmpdpCSxyXkM6s4+ua8D/F2B+TPqkjFynV7uOWZ4jxOIrWaHfN0FiAZkVHHadjfeDKd533
25kyrvuje4BKi/8FQNjlDwho4S316w5fxxYtr3XzhKRipkjKRgPb0/gjSIbtMg8QK7gorsYmdGjf
YKT39Ny7rjy92qGh22jjblVLC37Cpd8MDE7YWlDUtlj0qL6xZng2FS3VI0wJ+1sdnoPdlvjqoWAd
E8L6MD5+Sm0O+2IJwXojg1Wg3kvAhZB1qGltvrtvXrueeV/yNIrajjQjz8UnHu4SohXYGSnwHTbS
8AY/J7wY8PWW3za5+ePQHD2fojyL8/0+WQjgbftndAofdzXEbvJ0wX7mJy8+2/sQgZvGeMZYOJhJ
ZummSyNZ8AQAe4ebN8O+dgWV49SBCYSuLbjIWtZ4CiKXlJ2WvMnSwDKM+5TUMJcN2AJrUt59T+pP
Zi960dL6lZ0D1kqU2TjAlSvbVT/A4oc0Dc8C3zJB6fKo8k4sVomC9T4SlcPRpmBIrUiufEXSwlPG
Q8+W8AKJbuQrnAuHt2gazGBhmwQp273Hjia7TPC4SXXafVKZxfCBkwLThimv5VJJ8npsombs2gbn
iapLnD9dMRyUeEEV/PKiwGD2DdDdLb/7rd3iPPDsr/+2mFfzgHjf7tAWjDNtFfSZQqVE+jPKObyf
UGoY83Lwr8LKHkkofcVzzTjGH7sOjOJ5qUzHbYABgUP2XtYVHFNtoFTqOREmGLMgDPuPUGNYlELi
jJKP3yK7B71fSxKzvzSpiM61p8DJ9j7uvVdjecAkkb0+BcdR5YPzlW3huNZdjIi84k+zPKFCGORD
2tx0kkM+MuBUQHEw72fnStEIeK+zTpX63+5mG592C0cScS4BZTwyODIMktmUKm8HCeUljPXPkJ3M
E7mBmzrxVTu/FbgP6xHdNbH9/5QcKOIfj4CVOiaD2J4YFmzNzLUmpfxHLBDLiFsWOaymzkayEOAa
6MKj32c6pm76CG5YvpwIbnq+ut1HLKkHGsE5BG2uhUHV+VQWzaY7U8rHgUbmYpw+PpwNTODORcKQ
ySQ37oBRVwoMK29x4b57bhsvrOokqf3mr7RCQm0zbFdcUuEKvJX8uZv97Zkcw2PkWz9N35xWtn7O
n8tocTq06LoMy7gLNG0PsrP4wvD1Mp8XcBW/al3nzNvb+82DhO8xeyCTTuShE74M6vzGGqKW23Xy
FTjloKT10lJGvm83SwXyq6kPA5akmk/RdigG8CH+pnROlMm34Z5ZsyzIFLav7LuZ5zOeDNKC+pDb
lwGIjIC+nxksOF1AmC/DZXsGIeG5oPLJsoEgSx0Ewd+R6chmEUMqyueJQiZLYesqMqN13IgUGG5r
Adp30xAAzc8TZ4L3kAuzEOoSNza1kCM3L5GsuCsUvgOAezlBJMpxPRi8K43JexZjtC68NmvKQXlf
s1+yJjy/kMDbERjTjACF/0uiD0T/gmPJntCW5UjOEo1/boMpsQVm8qofQRFF0PLZoCeAMG+IDKGw
jwKPUJ8EEmEdhF3XI3+knwT/eV1cQvdvoX2fRyfwKGl2T6GPyOg7dfR0imh8Jz34EepoF+RbrBEx
Mm8pOJQzHvWKhfi7Vegx7pljneaKtbI04bBJXI3RUnb0hQTvjopRXND3lbABU9acg1mkmewyImVQ
KgZlZBgw4Z/qVOrHHxS+wIWQ204mysexcmnHcylG/mpXgpMi/f1HMc+xRMcqAEXNAOW5kwbBEFW/
35hiiet+kTtEYEc68+yN3hoIXr2tRqrEowMuP1MttqKtdYmfummZ9wi96iwLdtClpJOxowkXjRa0
KeMB9Vvt//aKjkhfs1LFayWS5eDqtuFmtfF56bgAeA3H5EZyOtyhfy7LwPXzpUlJEWzpuEONdFa6
7xL2bB1i9JA/IJw08c8nLo0A5QjXX72ndaKNsU089YzHPiVt6jUzMYVWiLjRy5mV5PW5B2cnLK4g
liqZ7yfT44k0B/Ms2ruD9D4JP3s7ZfKp6sPekVRK5pxjbz2FgyvujRbXmkKdRUFNEHHcculZizLJ
xZNhBmGM/RTzV0ELhDWAWElKFWM3P6cVvPcJMy574ygdlDd4V2HYePh6QQHVkMspfoLJGxlo2aOl
GlB8cvX0aBpsqqOlNuWs27lRUpoaj9hGu6OxcQti5y03sBfYTXtArTM+7JJlVRdgfUuUIulb3LPr
jQiU3P1Ubg05SQ5kKSze8Xj+FbSiTJHnDvcicODTjmLu5KkYPye/qYlAMOcCdZoBrDGScIuBMMjb
F3hEbSQqz0EO2sjyIDvv3MCH1u75L1uUI/r6/g8oUep2V0DmZ2tGhxTylYNBVgRJF20+DBLK8yvI
yB4ZwZH6AXzmRGzkWS/PA7JWrU4ZnIs7dHxxRDeWx3sClPoiMoJYQwfKZ6dQQDWjj1q2E6CG8ztj
YRzQBURv9bK6eeHQbNK/wc7bBTK36pMV7CJFZyh7EL3pcBLL7mEg6cPrqk6duUoxZ4WwnJQDcrEN
kB4NKHYrXuIRkszxknkeSK9mvRIG8dTcOyuSP3C7qH2YKiWVaVNV4itUPQ/whOtgTeho2blkncPy
oqaIMtlHYxSGLwiOGPiGu4Zmpw8N85ooYSN7wwdRDzNnzykKo6ZJEQXpi7mmpdNMD8E7NDl3UlBp
o/7suirWhyjUxrJZjnRuiUqY7x8K08fOCoQhWiUa1CEuaZOrtSY9HlH8cBtguevZLGkriSyGFOrj
Y9ux0vu3w/4vhk8KX7yCwbY1h/3GQCxoY8I9Xezqq03CPzKXcsoPqKNnR96EpJV6YFCru3pcUhnL
E4VcHDn1HjV28FAw5lDC6dkQabL0xGsNp9EE2LWLJHFL6s9bjQkZOK41YP0v+43/M3jNO7ePYjPD
77s/Tjql5jJOvqGq+Z9xfA3HDawgbFXZYAaFXl3vsLAZXBI0Dxa+6Gr85nVUZHpy+R+xOVTyXTMP
Ibsb+HuUhH0XkLoXvfUzyo5pPfHTyACcSpbs911RCJe+nKnYBAQ8hptN2O6sr1g2xwL3ytt0U2Ms
Vcc504zn4VnF32qGDEnV1sBPWCMpAiltHOUPSlOe51XoxvDNKBKzXodS80V0uVYXlDbp7ARVSv4x
fzkA8xPyZnlHc2SvTKpcwEEHr3MewzMIdDDymFqMcGoe3/Acvgc5F5T5l74WUHxrQD11Hc+Hlcqt
wRc60MFCn784kSCb6/HIdUBVp7bHl5HWr7JrkfRtnfKmU7zcIB6J5ONh9uRaZI80UAZJwDFE/KlE
alUeBN/4+Ijt9m4qQZ2eVeXQ08sOWh8ImNMUsn0L4q0LDWdokVeUQH/e2f2Zo1WaK7qOfExjmGKB
8zpx8Ojc/BJ+1Bjab6nqYqe89qJe4R2TRn0XiBa2SPkwjT+ILS0a/jwuerIuk16+XRE5sU9ckKsk
ADv/ZO5G0D9L3iYcyDI6ya2rYAtTky8bc4I7ucD+jF+HyB7cLXDVRtztXuubMSdCWwcdcEaNVtp3
F20xFr6dznWxwHCrE/wPRjHV/OhwgrT/oLp5bAafzz8ewnV3V8ebLDE1hXCP/JD6toFZmzIxGXT4
33seIt7DXWvMoaelWOZFaO+fysziwWe1yWuBXylmLCLVrfHXQEV1bko9jxUlyBSQg7P8kYe+TmGv
9AosZA3hVNoYBHt9Tr+7X+kpW1yCDW4IzwDB84QDYmOZWGO8NrxFPUXK7mxq/1F88TbZ+3j3kgSI
PVcgaQX79i82C1DoJWAfNIAJE4mqR3lYn90ErK332J4stqRLgztXQWEqXa9vYuX/S0RCtFSIDVw0
l8m86GS+0/UirvoOi9q4xhP+uvG6ahCDDb0aqwz2oJ7spwLGHzYyzgJAtDTQZR7OytxMql24NY3m
fKkDG876AO5KoJJdwAPLv/kiRq9KzK7xVqQcqUEbf7s3ArXt47PxgEbzAzMP0xaNzc28BSK4O6ID
hjSQhbfi/5p6brJgDNhHfivpnwvkWxZZuA5C9+jtMX60GKRO3w/uNgUWjj4FEl2EbJSZoDpB4pOS
quFd+wt+WIyNFphEY7V0Yp+wbXo5qKXdgrJytYkMCXC0yeyXDPAIlmRBnCiZ3iO8k8ZZFbH7jnju
01fgBpxOcqu0gNkf2XnX5D741WR3q4cDhrC2WTg5SBIfU7iJ+4gwcJQVuqIm0Nrd38X2JZF1wD7b
yRtSc/uLDwTZRUIvOzQYLOZDs8AjBlIj1L51jN20BUmPBokHuPeUiIOXlZMwVp99YTV1e1bbBhbl
sdo7mMbavdAQc8EVlPeBqYKg7xsZs2l2HuX4gNltWPGQvK+ngSarVK42oX15Z6hFs5w1YaB+Xa+M
XeS4PvenbRShVvOPvIcg7XYzjfHvruO5yjZvpeQ2s7FPME7vumeBzcGTUoF1C3H7ri4Eysti2Qv6
Psv4g+KPZ+a92lKUke8NFjuvRL77GnIeQHRujebOgtpuSqdOdh+viBSVkkD/UicD9C2Cy9Mc3uD/
He4eAZiJfUcE8+v7VK/vmSBV2K9VXxMfdBNAyhvc+J2Vk5cFeVTFKY1W5Xhv3YSynV+NkXmCah9T
SqVzgF1tSyacOThff6wA8A8Cj7ifNAp3J7YhYJtTDvQwS8smpewQn0vBr52fS6wEdrI2Xf1BsvE2
qU0c3vVGTOuPK7V1gd973F75f7I6hzKllhfACjc2stsjOY9WPQ6B3URj0INUyGwOHwwhyieci8XI
Y2IDj44fUqBVrLPKdww/coI3EkIOR5hymLUwOzZ/zjBqPVuxo7hLEerbj808qeQrbBLuRuLQvGA3
ObeSkBD4jTjutB8MpxCIBCwNYsHZeaqXX1gyfz3KlFWWGrMjR9Qzm3UdGdEnj6JNxSgUm/A/R8HQ
+Ay5G3hatI5sJJLVnYJEr2WxvpZDtY7naV2t4wZYZGnxLtDN9IVKqqT8j0bzv0AxtMMEu0aBad+x
ROb3CKFYKizoIm5NeTD7bvHJgpspIQiLrAueysyNkgc/b4i6/TLGR0m7sLa21NL11WLlJvT7FJE7
TsRA1qBQHWnrtlTFSb0bn+2GSob03FPzztI6tMZBhFNReDa8h1lraab0T6JmhZpTm/upUWQgRor7
B/mWktIvhhX99A1oOcAgWHcV51hx5W1p8dd3wY0DoyYpHiMNLhwYb9fk1GlXKPQGrCK53/AV1BOu
n9H/Pz1ExFLPvct9CdcPj6fvMgJRYz+cZ7PuWTcpwNmLZsQb1vGEe3F0NjCT8GzODXJDjbWrSpVX
HqmDWWwXk5GLRlfPvk6WFeXILOmxsXoXttXvpU8XE0XrpusH3SmtW+N3/xJAM1WKY9XFX3ZIpZM6
PJfOP4lj738wHFQXA66KlHhcMQtVw2KjT9n9Yj7cvmxwN3MeZOlk1rL8p+1qQhKF8FLIYGgmJDT6
MxRE0c8aaaf553A9BPF2XCBShsTMgakV2UjxZuA10La7b/j15HxZTNQtObUX023jFua7wM1NJY4Q
lBUt0zXbGPiRbt5J4gthuRIAIqE5bpgu//jXSnfpOVsH/m+AfkeiSPmrrpUcaqOuzkrGXKvpU1Cc
B+prT9h+MtuoBh22OyzmcEF8y+NR6q2gKg1M/zhxE3hx7KSwuAbzX0zZkVrvWmkefEsbZtKIePQ8
NmlsSxIewAtl8+YhqPyFJUrJJSimDe3XbVR1mDhdr5ZwzhVb4P9CCdulS/Fjdlef9+j8gqaeoc6b
nnVk3Hku3KMu9L1/Yv/poHaFQrLqMm+9m99RB/JUxjvawnOGypZIEp0esTLySF0Qj1F4HROw/umj
348NxV7Alml0eZE0v7BQ48hQe0TluAGAa+gQAer/bCO8ooJzLqFrzXkzLosNg7Byl4cYxhLGo9kB
jfARI+j6KoEi8CVxc+iFASwjcyn5b94Hrb5XOM+nJ6ZaIjr/DNJg4N67vhxi9Lu67ajxVEfPNq6e
zX1oBSvTpxmR5Nsd61y+VBGfQRCyrJ1vh5+UEfbwvPDlKLOJjgW2Xb3161nFTVVIExxmu19b4xON
9/7VQ1pXlTKnrkZU3d0BLrowZfMZYVZXoe/I3mSkMuqkMUW2BvgkE0yOKmjE5/Od7nDf+JX43DJm
09JP2K/OAlaYvnB9rPp4DrhQMg2f8T/VUZvAQlZy6pgNZA8l+pPFi5F2uCQ8etnm/wR2sstx2dWO
ha8MQr07ujgL0BG+Mv+ydL5/WSemhuAmtgKZFr1JQDg4EaeN8+8kOfojaBzfWrOCyCa9HBGsIVE4
BntKRtl1L+QU0zoBWnfCOorxjEAZF4Rx94AhMoG3hO/ScCWDmT7vmR0ZERqMgByxNwPpVgIqAlwB
UqbQH/lRz7nOpeYN9TvuzcE+Rt6ogZ5VNlAbB/1wGwlA/6XQ9S0oYtpv1UUbYN4TPyxC5nKQ6rwc
g9f/fCUHc2EyDt2GFlKDVwvjocsPn8PWL3vImfGZaV2BYp+RCg5h7tmTl+d0Ro0YMbniSQoj44eu
oRySG/PrZqIuM33jCQ+6xuBvk/Ohr+85eQvMV8gqUjn36mKyjlKYvU+g4CBKfUrJ6qDwr4qhHOKx
0S/ykYv4SxV1Q/+Pjzs9vgZra4Pu/JXZNUoT/s7+SwROVfaC3qjUKR1uRitMpwLTZUZ0iyZXoNWk
NEgSnO9NItER3C0dC0CPDVFj4jXjl0KOQ5AnOSnrJBb0jYx3iaHgeuvNZqXEdqGatF7UYnM5Cnmg
xs/s2v1B1tGLZofA2HHl6cVFrO9tKUk7A9N/Md/pDavhhwcVTpRzBtMU8OL7p2ls+nLNKbtUtLxG
k8pSZltFgKEdmToy5Py4/i3XJNakGCFGJZ61qqQGbRKCtsFvy0SdVnJfgbCpmF8tIo4Z5WadaGX4
j6xZ6VhOsPPcSyzgs5RudGUYIzKAJe9+55EkI4uElpQ5VLl81ynd8SgX4YSSCFwHTfF2hLifH9gR
TGYtzCy0J5DxrlBALvjy8kXu6xNVUljoLntNpwirqRAC8bF1ZlBzeDzooDEkBMgqB3HSM3MlOHOh
WeF1r4gY/7XGvHTHVEX55dKArseFJhz2KNSbdWpuTp00Em8Uqrbp1sHk9BBzyniZMkBZaVfmFzGG
mWS6Ms6IlC28UmLDBu06jrUwXc1y80thPAqy4L2ha22RQUOjOBiIBWJyvftQBjk3NisvfvfVHtUX
1TOqsf8zcwAjSfz/si/ShsaucsiZ1Er6T0kNKT5B+8SJnUgRrvXXJj4lHikY2ANYrnNz8K6gicO9
HmZI/2ldK7ptipiH9/rDs9p3aKQQ8BXs2TgPcucbzl2J0yvBsXyLVGrEZYGbXsOg4etqnhFyKVTX
TozeDfzlWGHsmWpuB2K6WAYFAC6tJ04w6jNUqDWibcdDRQOUhCbxBh3BEwD4XVqA4hMiFYJ0x1GP
9xeICL2be+/U9JRlTTlCHWbjNIimKumyLOqrCOn8mjaexC1yh3M4auKQn3E//MZJTDN2+HiPw/IP
41I32ZErciuVCOaTBexN6kLBp2dB20ItDgACAuzluh9XsBW7fyaJuOtM8mBvyF1p7JPMlFEYXu/j
17wI+5Gk1SWtgNcLiMn4MRfpgTH9CvTD4W8G1YWwfcfhgIXffMSQI1NPB5PCyYQY3M/2avH4ZpKa
HYvPSOCD9A7yj5bfzZip55EyR8U+92quv+XUMIVKx41ynX2BgjAPgcEFZhiAUUH7PF8mNyGvnjEN
mYWsEA8SzH+uXf/zZCyz1/ygxbjFXUfvshSFi+zRzOR2iGD8HzdWUlQEhITQIzMddTEz6rX9pS9Y
ovz+H31t11Bo9IBkX0nOhAjNPJXUrmktlEW33JDcplSU2DpTYaVGO/Z4Nd36hbTE/UJGWde5X103
NnyOKPzDPclt4JyaZl1s/sDDH2vYA8r/rO/U9sdZaGhSoG0Y3fj33hWlF8PW4X5yg0+09D9iGKFD
SIvxT4Ms66BGSveYoBxdpqhylTIoq4iTtd5nAChUlXS+SrudxWa7KiWkqDhPlWwSX96+yLo71F6L
k328EFsZPtI6izF0H1w4R9hsO6y02p26Sq/OhML7pua/UDfkI3yZNFwU1pyK6ItljncFHGRJKCoP
VfveSe8lLEMz2w/DM2OlThyowRB7nAW5lcKq8L+LS6PgIMFlbI/Qcbg1z4maOgQbKiI30NPgDWNZ
CmdMqH3MOxz7p+vUYnLftrbTEdp4pdC+CUel0ikeJjK80jO2cYhQIq1YYfmDcrEe4+sqTCZYh1x8
ipioNHhs7nzy7HCMXzyf9fCX1cBmFWn6FBWMvj2R9OZWXndTSHe8jzZOd+/GL8bIsvcS6ZKGpQDO
eaRcAAherHcL3QZpU6xDNsHjigewR2WK5gPZ6KxwA9TW/KLhAJbUVFcIztb4Xxg9LUeu2/3VKOHJ
gvrFRBoWuZ4VeGyjE1974AUXedhTemG8m/JHW61yd/jm3RRbL7taOKZWRpppeawMPUVGEOZTL5r2
xGEQYwzWS74XUsyyb5azZyRwmpmGOSs+uO/Qfd6yxLzgLX4lA+vlnGXOyFofknzhGByoD34M1pgx
uNhgaOOUPM0rEkO8M+QKMUmxHCdzTrho37a54w2oBI8Yz+BBf1v77Fs68+R2GwooJzdMtXILS645
3TlKIDnCGYKRHbT74Gws//aNMIuHQjN1vt8bM5MiK4e9SxL5YIr9VJt8AXqfkfOfQZbzZx7c6S65
SbbFKR9UKZov+eCWg77TAiHcImgjOrcQ3GaD4yJlUzUyXxxQLgCGoDvVF86tWUwUW1qInoVLz8pL
t4CxpNvphWIGvC+o3juMmBIiZdCwfPSm5Tp6GQuvOBNX6h958R3nXCsa+vKGS8zVSZEnFevFS8EF
fCzXsxG6FKw464sFXifaCSjM22Tz1lAqp6N6VPlmiFEe9Zv0hdzOm5kxToXwcoaAvCmSISo6CxMQ
uJwjpglCSXu4+L65X7NNiKxWvD2K9LVD4vee6mfO/VSDCenluUQpX5oMB9HctINkJPBoyWU9XY+X
KpL2hHnBCYn5wCUxtcsyHI1QFABZ0OqVZSrnvKp4EVhbRvLgagKqfPo1LqzjLMxvuD++cBbAR2OJ
1VkFUMcPHqd4QhF8SCIngfy4tYwq2LUFuZng99QbyWm9PUGoZTIAdeDJraedLZBpIK3eIXjUEgLI
9e2RoLZlLeqsE0E7ZkUk8IM1rtIzqEUhFycK7ZngAOHK4YdMSxRbSVL7RGJ4/f79cIjLdq8YkJhS
xSN6fQeVY4hYiGy4wENN0zWKgfYH8SLthLeknzBcsuPqQYIpRRJTTzaDDLFmwfkJa9zVYpZLbUDB
0N9NScdabtsizexpvq0GLbEZWiWZAf+9O3VFx+gsDdMcGy8qjcMKYkgDetUHEBwI5QqXVT8OZf69
KyE5/ow8BTiAu1419YIJSU9fkUdDJ3WZg8nT3h5xD0ISzj8mQpq+HAQoQdPOAX2N48VDkvDgXNgK
Ul08fKIso7MtaoH70e9kKacp439GFRIPqwVJVmbO9OXRmdbPpTEEE+mDvUg2kjMjQF1ZAwtEVstM
1aT/N3FXTYUd71YDYDG4yf1kbF8m9Ta40nb6jlc15z0Tzufu3+8cBQwTnnRXgJQrT0PLZ6fMs254
Z9o1XF/hhxyNpZwtk8Z1s02UyTGIOG6LGjYvTWClGOR6UCdfwJ3UtnNbRfzREywUvU46fODOsYMO
0N2dotkIm4huZ+xpSFkCjs9iKWL7v2xhSfmzc06w8+QiOaf2ydsG0u/3vLoWtnCs5M6Zwv+zMsst
b6sdhNDuKL5gsVKCLwbsi5jWXHtIas2s+nqLFD14Pk5qUPQJFxcwyWvYp7VLu91qaC57kf3+YY55
Jw5Z8oQI5UBhbNKxvFLitZ3qIdSNH4zJxsW7r7GBl5OVYYE2PFl6lAe502rmCwPxVyXRZRsrcpsC
Pdl65FElddRyIjGS7OlGB9u+/o7EsiZbo6LQfb0rqFvaU94gsnsLNs1N4ryNWgFLbvRzLpsRl/sg
3PLhfCSDLkattlzFqXBgCZJWrStDoI6W+RnNCDRVvx0WjjrQEbc0WbGwtLb+9oJ5Bx1PrPTZX+TG
thc43rs6yS5H9HffULJc5l9ZVG76K4kVpYEReD3GqVW0835qHwy9pyXItQdy0rNTzWaiwtGO66oS
BCEIgZeNoyoTj+3NPuZYpjUAZl9W7x96nVaucEc4GEBX9krU+bM5q6NPl1DeGYmkWsBUViZ6Dtaw
eEePR9t1zIIs7/+YZgpQQmtVJMgJVrAfHHuxRjYw/c9weBxl/X1RJ9i29OSHsrAaJJlkZdixynYf
pj/O/G+hyLk/PfD5UULGsezmMPILRfPjtuCxdXd3mWpqu+6ui3KtY9O3bLu5WAEwNAAv+5OAl6Rv
3oKbyV1MSsIBtp7uHbW3Ry2c4iyO8sCnyAs6NwxtBHzTr4E9v3Y27R+YopFUhER13ysgm/PRK1XD
VBouljq1tkIX8NydPnHXYQh+ugCBbQnmYT0+Ppn1eS7XtkvAN3GTZi3pisqvh67MTnbRzSUcbpUK
HEIn2XbbFKf/ZzYMeuvqJznqHMEzz4jeUGwM+yQ2A7Bth8KgQ1Jvn+0I8L1gME/R9ZhRklf0U1gs
XTyfWVM5b7b/fFuxccblrkWCeI+lKFfIN9rH6DAyfvAaXhYO8RnhpOjcg5MsHI/0ugoH15y91RW7
6Z5Q49UY6BYQ8G3k4OkRayL2Ss+ENQS8l1NDCdu+ynw8nnOf/q5//MaKUWyYHeBloZt3mO4QOVd7
w1phSMfZqPq5yI72dtme+Mc5w0mzXO77AoQqG6fjrJWnc+mFOQ00JiU0YgTHzsDvBNHcyr2i+LIX
fboOA/giMz2J10Arauluccj+qYnbBCXd5P9dpuT7El0WbgYZLrraPHis8dA+yoYd+wH7yPMjP0rx
qFNe5BOZBFmv/cIE6DQZhQrJ6v4bGdFO3MvrPJFb997eykWVMgg8EquySkcMyklAOzh/dqFsRSAp
FYLOg5Bu3PsCaGv0PGRdrUqVYLqdJ+ucr5ZCc4hTqZMykFFm2wMVXjYX3AYv4wtkjpEDM4umPJfX
USLivlOGcJUBiOC61EBcCRiAMNZaA7vTWa0/wsN6sO13/DIdDnOQax+IP6Dl/opTWxAJ7vcy9uKr
y1zAc+4dXNzqEeNeSfp9eciS4vWXr3D3x6DzH2AXMjGjBPryl++U9yBRls/kEVoK4abguv9NeJgD
+q1/bmSkc5lSuv2VXZvfDmoVSN8DmjT+4nm0MMM7hj8YQaPOqlozV+fcBDKHJdaXoU6HhJ1hml8y
YQ4vHK5yJ19IiXHTigughYHI3tzwXd7j8usMB2+mHUReBjI1rLUCzwgQDsf4q3HyPFaGRhdDcQlr
QZ31IyB2bwPzodDir5EodJDJsf2s3Gy+xHMKxphyjpNcLf3JE0424yYV0Ko5pDFjNZqQ73tlvrwR
sm/1ziXRfALxcskbECBfC7eOxamKVfea+GvaxdE2thBBRxr+jv1bd7UJzxAN2KBiCeX1BSGfi3T2
P8jrXAF2+wHYlqNTRZJEs5MKXPRVe0AL+A9dwIVT9gGVbPDB+CQLUdC+Y3eN4nsyHEAp5TJ2iVrA
zmX1i+ZH4xpwEFYvDpG8AOLpH6d/D3lJ0Z80V6VAoUtB99bCuE49YIMWot3fWoW+LcSsF5XjWkvM
Ifg8vx7crJXy0FrSS6grd4XfKqQbUWzH2znrxWsvnawpcXdaWz1W6TXbmVNoA2q+NpVisgMOPPJq
Csr2gZpFfSRoE4CtreV2QQeFf3FCjca3DHDFfr6zMCeYnjdRDYuyJhZq/BCVglOkNfWnvpSYydPc
I/bkgch9AlWganDj236El/fEiaLX/vuMtiDIcEhpnvtrOrXRHtQ/VmFt2FlMOGun7+X6IUPmCizP
9s+JSoPxg6zJjq+zWblShM9BfYGJ9wyaC1RidMcuIvCbawdYs74ykuaGgSF7N80WnAcd7Q5Gid9L
LXl4k83iesW7JQkGUE68MIDgcEkmMvXKdOW9lXrg5FckmulRciFDZk7s2vRjEwsCKn7Db5ILKxMB
J8NUGd7fBDlRTTKWraPxSfnIhWNxsgXi8h0zEDWSWKMkkbkixoAFkNGAcWb7yNwaxu8ETDsnBcht
Wf+SfpsD8wXoF6LZza1P5dwj4z3AOYPzBtL2BK0KrTXBW5HLp01SJuG/NVeBwrdaK/aC+D0bywf5
u//hIvri+6hIgqTqHRyZXj7nKl738piUeenadUyN1VgBpjRZrhu0ADTbPFMOuuCwotsBciLreVMa
UvnRtVoutK9ii4AQrNWORZVh/mmRChqbBJKxMv5674xHLF+MCPFQQIizwK+RmwN7tsc5UijiojSy
NnwOiSzhTYTkVfa5n13nchRzpRlt9y9MwI2h4ZkHq32uxvH9zDO9BMTfNeY8GScRYsODVKp4zno6
ip9u/qOlrgVKRXG9qkiTVdw1wktV0BG7oMKLQcr58nXrylYhn3Sjfh9J//jm3MLEPvpOFB17YnI0
Ds5qP0RxHInwKh6fPlvq/lNTLoO2lcMrs7NKL1xdf/Ebe20XG5WgK5lzsjrRWdOFIYp247cakypU
uhV/PhWXpmTZekq0CmKBdGULF2OgIAsNreUQqzcxq+n1FUT9bjDFyEzEvenWxSatyAG221ME+Kii
qkIkgWbaQDfgpnwfQvMpZ5toRCoL7shoMJ2pv9TOPBvcJjDDZwP/jFfjZ+sBRBJ3fR/Ge8Rt5jbZ
1Jhh41v7/STPbNV9sfLpOftcbjy23Ed2IWhrC7ooz88syzsICODtot+I+6wMtEQYMQLlFHZIuvE3
hNKWQCQ5A2CNkrCxMBycwcIKoSS0GtUqmu1j3DaV8ks/syhwg8mX3kNcNQLSj+Z3lUDgBpTPS/1s
/0Fh+9GlYxdhBZRkpM8/qUsivH12Jf1CAZAOAGrkqAtc4CnBb4xRktmo/mI9IdpudT8U/CqjLZwS
LBPDgHXMj+6zl7w1qeo7OIeJTpbEZXCu7rSUHxa6zsnaqJQ/Dv8iRs2XeQwCY6c3HTpAQgJxCucj
P/Eb9x9CfSY8dc+qC3yRlqRoAQaK2bVUY0slZt/SE/36lOGr2tB+BF97yPuErKgztiHW/Bex/U+9
J/QXC7jwgTq2idKNTDOQey1tVR7Ji0nJugkKNEktc6w3H6M4VyIUZvS6Eitjxrnd7nnOEFO/ZafN
A6jcxkeOjJvAKqHtludqaFLrOXi8qbs1ZnvlMN4vTZbQp1UzYNX1BpHnb56brVXbOwfCgAjik0xn
YGEp3LP6T3LQGu5ExTNFpZ4LVzdH6jb0KAutcTUEaExW7K429wDMzwNGikFMxbn4EsfgFzerUq4u
pxh2bXNNNNsdxJ1r2NNqHX9ehntcaM14G+ovOgpSe+2YeL+9O8qdINouPFzaiMJSkDd7KbYC/spg
M0K4n97gFAYYrnJcNkOzKQeorgrlHRxoFY60Ll9xKlIFHNVNlhbrLwDllANJf5WZ0pKh+IkMFQMN
dKwpXiz6CEqoCdVkPQ4aiAnT5F/JRc12G8VdlASxLnGTqPZ0Ex8wbUhNO46141uGQ18THa+v1fLk
6vyX+3yBmXIIkKX58ux6UNDs8toxKdnZDLse//sf5kFumQgVqfdwHQ92ajy5AHx+CQdZB5G0neUc
ELMo3DEmoQ/3yPbqvqMOePkAl17b28eOOhRtT15xzjsr+5tVQlUhRB4kXXbpX3P9FLet3IS2Q3x/
lxryEoKkPDFA4cNiYQ7w5g+kg7XuUyy8I3hvlNd/T3i4WOO//0kdTJdFiLP5sI3JjPZXi7sQYiky
9JcK9RbYU3+PdvnWzV0bVn3B2iAjhhE1VpP/hr/28a6iv+qbrW6wcghtz7h49G6rtBw6eQgvCQv0
j6ks9cCdRa/B4bOnGcUa1qsMGDxy5r+FHaZY5zk8Zzr+cHjGo8bUEqv5FUIXvBsq9CURxMLoO2r6
SOy7wnq/AANdutLRSiTa6hhwoucOaKuA5UFOGjUldyWrAnOo8c9GQBjrMMoCHIg+fNHJN77eMSd+
7HtT51h5Qr1yB+qJSHr4IxjVBpQtX1Ryd949AQhEKJgl1RLyX2o+dk0gg+Fvo7RF0XkzKVmiQAJQ
0YTeotsGMRhEok9OSyfze6abTjops/n3vMKdbEoUzIs6ilXbMLyeZdld0z/8ptbkgHRCD42uaUpk
pVCnyWakwAkIjzXRGPR8k7EgBxj3G/oOzAWDZXTNdM2v4S04WXQ3Zy6XVFnN127xsrrkZ2Uz/LSO
bemYvIgfSYXn0Ai06n1tF3OGnI5A+Wzju3iWWtdiAhxhxmnA+7usDv3D+E+RQ9d2fymPUkgPHBfo
8qKMYIrwFKi5/cQ6/P/74xcxK7sP98+CuvHCXzCpjIlewIcAUXq2FkLOE/tmzb789xld29TCtiXJ
pejd9X3iWEGBjjj3yUt/0w0NfuovbFg1k7W3MXdhu/PPPT3OjsMD8gQje7qalnpEgoMkno/W2oZu
GyHFkdny8tCT8c+HN5+XvUybwb1tkxLVMu/n2rEUOy3sU+rVnKpTZnKi+r7J+NSb7/SEAg90xnVH
UdscT6jjbtpmOmGIJKIwcnnoH8skosbUTTOc5gbRpdkIZtEspr7++dLLqVVRVpv5mZvGXcDKTli4
6Rv+yH8fDDD5jv/lGJJiEMdJ6os7w8k0LD7BFzbVSe7EIO4KvW8dyjZBdwW0QCoYSBmdQi0XWuA7
YwM3Nc+TkOU50WtKbXQxHy/Rp4xI0bBF2TfIeBFojZdulM8v+Bx8NaNYVntItlG6NESWDTyLLpd9
RSY61Op4usGhxbAAMOLdSwSYXZi4cTetdkTADIusflOUGuFD0d1FAZCaptn5fXpKply1aSz9zH04
AbInOQMnY+cXZB2c2McSH3G/w6Z8YIcf8fn7YweZYY6rSzw9l2eaxuZIX84c6gk0cZMY4L5g2nqg
6aI9kiXrXkQP3J5/5bjdN3WogsC7YSlynuF9LkslBOI5hHJ4ncyrF+rhdXZsBpNpe8prvc8P5rRL
RJDIthzJvgjReNSLMesH0sDLyNzvBfEqoXOs3udKWPYlQg1j5ZiPTyZnAw9XO0VcJZQuAZIUbB2P
hEoiaxQesfTRDlHSbvvcjNjUOVcXf8ToUMFZzHihSU/JT762aqKjPXxTwBb4VyC9Mz9IGDNf5+eo
aU+3N3oFUSbXDKixykVClDTHWlHTVWCFwFPDOSBnaMpSbB4kGgXykbuxCFOQP9B9fbRe46dNkbtz
u38GOa/Ny8bn6xgTm/RGoOvB58jf3fUWucl4iMKNHV+RMqEDYn/jov5nwzfLBbQqGG/ptt8b6598
pAcSdO2fGxv7Plpt2+r8740Vk9Dn+HHFc+PxI6TeTfRIJ+jssHxD4H5ww9XQuBDNijzcfQTt2Gsh
R95oNvMQTUCIS5CFiYZRdM1c19X8F65CrQ132ls21D1azrKLTB77kdZ/UkxysTZirYNni9ficDLB
tjmyjf6jwC24v+wPPQdHD7tvq5vUMnXbfFRGd+G4d4Jo+M504bTKj0hDE6SYlwCuchxftJNhiDto
+kdF8rWVaTgvALPGs8xbBPAd6z/FxHxnsvRwR8WDoRs5Wvj3woBb7i5Rk2Tp5bFUvGa9gpF3V4yD
QkhMXnCnz0LQlFlOwoFdNEZYS27Rx4Xaw4cuihdqx74+MrdXbBmfFnc+a2Y77gdpx6dzOWEpwuDs
KlcDCgKGbDlyrg900fp9uV58t3LLL+ZNwlTs2bG3WflPwa68Q0dueEQn4Uk8Rko/01l81bi2aiy2
ZUDZQS7YV8urN1161EChjLVAPqqMDAnsnx2zEj8atBu0lCFZWGJVjC65/HeqPN8Rbms0n3ignp51
LhhOVpvYm1NxpRCxix3yxMHP8brEOed+52tXUo5wikiQValAIytwGOLd1z6SxUeBYSbukcjJ05IF
3h9+S4a7hQBLwVTGvCwzZoNFn3g1TZEXmmdVa3TjCS1eEI0GR7X2xajsII5RWWtpvMf499LeGiPd
yhTjyaymvJSTNSoORgIWKmf17kwmPKE9FpCY8mfvGldQv0P74PurqfGnrKkwPGdUa3MrSTUrdw1L
6yI1rDIg1q0eESN9fZ957DUaR2exhNotQZHmlLGvgMb4p/Emw5+lioqS7l1bedJyT9C+ApkeHHZ9
y63oad2VboOvdDZ9/+rV8fuxSGNN4UIEmh2/42XdWurXGmAW6lq7DGoQCSjM7V4OBdSv9CpBVPhr
cyVEYD9JlkIUIWt27aNR8Ken9aiHVQxxKzUWl2J7JeTafUhHNF/9QjFPdjN1n/r9J06dDTLQuM+q
zWfPwxl+3AxztfWGLmV3VZd1iLLvORUiJ4UHejTrW57d9oldx2JVS6/WL8vhfiMGo1tg2b3sd0G4
3rVnvsb6bCBZGaUiaHqopeziJ82WeNeiDw57Ue0AdiBhxH2zFMrl7Gd1z1txPkJ9kEpC62AMDXWy
FxX4OUCJWIQfxvT3nfGeHcwLC0YO9Jv6dfHdB0S3D0BHbfRJ7kRIJTr2UxxUM+AKymYNwwsd7eCn
L9qDDdfbWFYi+bcY5GdkOu2x8/axiH190c/a5N9JkmqlBVEoD2laiyA4gegSTbYZHZoZVFUQbfyO
7pOpZI5brzW2zYdjn6QaqOd6kkNTvAUpItOsrQ1cjeCva0wmZnQjzzBUBadUwn7wbKmLX/x2ZCaB
9oHu12U5xrKIYI8hN4F83MSADdQcZhe/4ioZ+D68/s9/Z7os+eNrq2gsbbeeljfJmIL5YYT7Niiw
0jplU22YImIeRsSm3CmvtZ2pORqLLJfvGgzGUwSjwljInhYE3XTH38asZckcdTqcMSIiRp90klxY
J/qZ2YRppncZSy8UMNWoFKTcA4d7T5+EvKr0T2uIX4EMpS8HW0GcqG79HJsjgGfR9Nzgr6HlCiSx
tD5pW0lNjE7jyoXLYScR+S4cwGVyXojt3GmWsVPGixzumLmGhly43aV/UdGNMn0Nid43AcXZV0zA
sVB/emaKOvGY1nmFrZzWAOi1QcxOKZkQf2nVAqs+/hRK4uYozC+XugeTYNU4LYR4lZ/mlDOsNQH/
4J2+x6XZeaFeMH6B0M8GXhN1MKI/JdPV6UM7ljDU98vMw5ihHvYPyX1TmSJscD3O9+2aygfy98l9
ZDit61IVz2Bd/ZrNpcXfYk0V0gcz76kCjpyFRNlCzDRJjOiJ8Ury0gePD1x/PyayOF+qIFhgD9sU
K+Ks+rfIUwdV67PpTPYPzBYGKWsZ3j322ffBY9uS7De/AJ+S6+qvJl/uv07kZaIcNFjpgPMWJk6S
3cig7UBec+tOk1FHbYyegVNnvwh0Ku0/kxKdQsb5H9tozDh/LLB0slLi72ZPTenYkR4ZMcFHyDyF
GdTZQhYv3njjNUcrMsL/3YG+AhUoNXZUBodfVS6dzT6iuQETrcKblLNyoUdQVo3yeqeSukEDqx0k
fqH4WvpFREbu+h8KwXmoumDiavMfHjVnhnaVesdGZrT2ZRRK2/YkwvWiNDaVhmbHtG8+A7BxLoEp
CXycj9W5QxYGhk2/PKT+aFeRGuqzHxDpaVwx9+jdfR6JPicGV0m1cLMZtQp2iQFln9zWBJAjhDji
ooChc0UDrCSdB0OVhXowO1XHpFTLXWQVfIK/PwH14m5U5SvYoUYmTNsj4HV8jK1IYqZcyD1hPYn0
sp/JW//thsFZkYgXZcOINSBmMJLOpVCGjcrLtCYkCLDUdb7OqpSJ6DmT951qgKkf932XcB9l7wnT
BPRjgjRM9AYayDjzMEGRSVJ6Jf/7FbKc4YLtAvpFujE6zFIEfkkV9i8ZrLZZkrpaQesv2uvIelUD
NN0Z01nvzxGRU6DoRgdzlN6DnaBpPfSfRvqximu0ooWtNPS8Bkl5ZbvlP2av1MweKf+AY6WSLfHx
4xqimXqvmYcg/wvd9Ozbt//BootsKYeCgZPCb2V7KA0NOcEBiYynLjujhTPlEbKlUT0pUePvEG74
EqbPL/Xeq0A2F8znl/oNjAMdn9JlN5OkMnhsziigSxSfYLYeswMTOiM6EfQMtyz4E+8YzyOcK7du
sZaYZ/viH9DUqJowPDiq1cpUqgap7QCTPI9AtbmX51TOCEUz/EVFE7sPQq3l+SZ+1fNU7QfqqdPB
U1J/6o/ccMQmr/InalmLkkYrOTa8N5GCF7fEve2xQfEq+Zep/Gb56hCaOSaMyuK1MHKlFg61r+1o
gRO7pK9GOHDzIqJ1ccvbiH8fUBM0CtWARG7jJb5ti6bkAGiKhHO/iiygzwtebe8hIu99M8FITGpP
Jb9+sarEcNS+eqUqFQCSYzqFsTg1FUlAl1XS1IoSrCDnqiLcIzV3YcYanSbA0TG3bG6uosiUCk3h
+exsIm+5ZEx+oE+kNBqkqaABe5Itllur+p2QgyK5VV8K+6oRb3oHspcm2mVAi8zTcaiMT8UriG6C
oRgRwmAiH+vv34v6A7V5f9v/YWOxiPC0+DNQd6wa54wG90VA1wxQLNtcNI5zOGLaTMNDyOZe7Gvh
w8BsaIxNPK0fX7AbD+eDm8INyFukOZgap3XSyrIDS6lr5IdDng+fllGCQok4QSv+5NOOhYCTbDsm
6grpByy7GO+4bIh/a4/JPQ4onGBFg4z9vqqSie/nv72WAkKqr9NuKLgMq6xAu/oqWOhwv0wcEwZP
R+1I74OFtiprDU3hlhrIO9ySv5BzPVZ3Lz+z6B0t2W+yvwgqKguXFlJGgODFRCR6CmYh5wxhXZ6h
05InbujboA2+o2tGitQ7nxky2Mn8blcZKeW+0YX6Z4byQzf6jElAwxAS2Njy7bMEFWoAw8LjtrXA
zyJHov4DuQ2QHwjIpHWaBe23e+aKo0WNKqlYM4gK9agY/tK8nmyJlxqGlH7Ls5AfFFp7BeyYmvDR
44z04+KiOWbzQVhIaZAq5X5S6zVaP1h/i0u2gJmZSaZ7udNSt8y+h+obl1qQLsQr7HXQcS4gkA+4
peuYChHuwGAYk9C8+r/XHqro+MjLtccXR3vwGVsyVQ0j8Uh6Kp/IL8QEpBxQoRxGSC3B8mrdNP6/
mRk5ZVuAAS/mJSA33syR2MZijqWc5CPxiPUuK+as23Zj3cPvn+kBrxVjRjsqpj8aVrEeI3MZMEl5
/WcbPAJXkOzu09h5bUwmDyhYC8w8EszX/P5pJWtD/zQl7sHthBZxYpue7gxnLyRxzFzfcdZXyYZ3
hN0VUSmtBRITkpIDnN8gXgLKO43oqetZV/HSG+ulCZgGO/ZIngC+/2wALcc0qd0Z1h0f4+XOKD92
WCYmLAq8fNuF1ZJC8qkN6kr9M9UP1bP7SLCeivQLxZ2yAxEjF8WiAWiIoovtHVg0CQRjGso3UE1n
Rc7I07y1TUK3T4Zd4anH1/D2jmNTGvWsGLVVmyzmtXwarumrmNIAiZHlGLVcWoYsHLXli6QD7CvP
2R8wB5C/OLYetAFD1Ca48PSXqXpNDSCwoP8hZDyuolB/U5Vmmt2pyAX1Q1rOaE+znvcq/1uJbSe5
8pHbWVKy4wrer6zp9nCl3CmLiX/FZURaWlhGEIJLjHfShFQhZexux8Dq/Qqg4CEKudDzhR2IuzKr
LNPbkxaWZ821NmXniFlmoQLjMnLY62aPFt+S9ACNMoAq8NkFXOzeWGNyxNwno5Og+sUZ5Gc2fw0e
lQbm53ib0CHbhJT4qnrKZ1nQLn8IFtJcWEIMgNtZDTyVfimx8TtQRT0YOwQXx0PuOwdXPCMXmyWS
nqQi55/00R0eMFRfoTxcuFtqLGl7baxGTx1mMU4rkbRtQF5YHq4e786vMicGK1grZq96VVZSptk9
MV8cJRaDK78XlMmERlDAp5iZSyaWHGnO+4297iPG5R5W6VadhdQyl01EeePWRQeZObS+KPE5vQPQ
yArdWBvlkhP0Zs+wuogPtD1zwjH8D9JQb9AEXU/lR+hG/oM1e7P0ifk0yJNoYZZjK9f/FMPr9YYb
r1sV+sV/CBwbHgZouj3AZ+t4GvsvwUoECqDunM1bjTSQeXUjLBJofXIoefMAFt1kc7sAw+mYltDf
oVMl9PhlDI5+WEhaug/d1FbTaOfd9NyH8G+aWeroHDSUOJtRsK6YZKGP2+GE/7facw+IG13F5RXR
SW3oUO+7xq95iBYWVqf/ZqwhueJYygCj+wpPFPhCxaZrXSX/1EGQbp4o+haum7pseeSD0/d8ulYi
jO2iU9fgDQWoyc2VIqYTZCPsKLmhsIuibxaF/GkF3pX3rTzWKUvsucRh7lYhC49/ni4cddkiKrEg
niBoo7QBxF9aUAbXW+sgeC86zETVPzCQB7pv29+dljkpUHQWPtyId7pav+jvmRtM9v11gBkTikSG
errFxVA7rt2j8p687p2cOD0qqgH3hfegC9we5TEzi4uxj3BIB6Lg3s96JNI57boZOSYCtLSsBD3Q
mujl1xXJ1yl5QimPuKRN6QGSiFlvBuDynu7FZDUrKQYD6kCIKMk0YliCOMVMFu5dGsdllGtCMih3
cxJdxdqcTexaIvgCGN0U6vlJGyxAlShzfeB1mo9T2Hn2d6TPJ4m1TMtBgx67wkMFy3Se3ZrsIHmn
atEQJ3OV3lZwBkWR4nQztSYZcx0ivMDgx7ok9rnyBHEG8H15RzuruQhP+TxwF4XpRuKBM+h4bj4i
sgyB/zEiH9Etjmq7s4x+/7DRozgnQQRMOI+hIbmxiwomLUeFtEBMH56wlpt9+8h5nz92ge5SxDmt
uJ2i1uSjoHjTfb08TVc5v2SvU91sEIP8Q/4HxLe35knEg+EqLbvvfNwucG0VMq9kPowyZyr7RYgq
tO9b+tYEPg/6dAkP1kGiWEwyD8k0Qw/qz3KyPcuUWkM8P0HEQx2MT7qCnryJS6QUpwC077SbVrQu
lGPtJ2kKPH01rc7sGWmWmawHYShmNmYYG6RO1KbQhliz8a4lMbkTpRF5AztESLaAmFL6g8Cy72iG
oYdbGU1RtokhGIB1P2q3YrH9fxqM3R6v0An+MjRWPYg8qWvBjrb7gM3NHgraTSVUa2wajV9fcY6P
druXNeAUTmzbsdAQf4FGgKtzjY5yGKcs2PcbjiM1NLgnDnaKB2QVoCF5qV4fM125xD/qs7/wZ3vw
Tnz4P2xMJFcDWRTAJ9o67tQQitXmP5ph+RoTBdMhxKlg+7hDGr+AQ4WkJPVBTgWe/WBXtBJkMWsr
4F+SPgSg7cs1DixiAeONsUmRf2id2OaRdUKNe8jIEwEVhmnjLWuoj1fPxzcTOWIFn7KN3IPxylsf
pnAtRlae6j/PLWyyq/5T9UxpfYEDplfIRxGPm1eF6n1ap0Uv6C+3SWzvwEKdKB2CwuaXX5IHFyUQ
bOXnkd7TnQrFdQ9rvzVkKk7KZ7a2KdV0BS3f6zyjDavMCEYuY5JVs6O2Uhj+/pmoalXAzHGsyTc3
b5TRdyGFwWeMYnFdGQZ2VixWCB8vJr0DEdSa27FAhTQG8SBdOvgVVZw97dySjYvx5ErMkXb9hNi3
VNQldyGJ4Dq689o00d7Asf0vg8iaUrPKM+Xs8acJ2wXuTl1uviTSsPJb0N4u+j30iGTnKLGBPZqD
gfqxjiISCA4TPHHTr4DEWhWO/fyLiB4fy+rd8tWmEjz9uu6csfl+gfVKXeb02/QaMD2gtbwJ1IcH
PvlqQl6y21Tf6Z4Q6f5dANYHBsgFLwfjoQolnNML6TizXS/VQhnzYjb8gMv3AQI3ygNVaCN8mV8d
bCyc1lFKJ9QNYJgG3oh8M0mshl94/e6saq6c5NxhQ7DNhNuEXBYKnurz1GxNp7n5bsHGL409q44W
8Mfl6d8MS9BiYQturiG8bUTqiP/DxFuq+DwuSjkX6472OZTymnMGz+AS2VjvVJV6wuSpuwi8YcMs
L/fYEc709UTaStJJAsqRw5j/qgKOzxM9vNDvOvl641FsQkynUKjOus76Q2wXF0mWpQS2v/7trUjl
bGNCRUgBRT5Go+qKJFBwkHakUO9iXvfNSD38f0WmRQ6MEWTuevZij46xqQt4iteQeWBClzZhcbe7
BPNl4f7S5zVjSsNY1v0uxoic21uOxm6mrk0JsnxhqsGRTx254vITBSqx3zZw0jPXNn8Auvg/dLr2
5r2IOQMZDN68dqr0CINzI9EaOk/HHADfi19j7PnMNvexahklFbS5Up0AOZSv9B9n1xOxHJKiuvdO
zFAriUtS1KwgjPv3Z6tbxhgGybT0rj20pgeVixo4sWuIbolgcBMnKViBxuhVRD+NP1BDa5WVeGrQ
lDJXjfW5A9odYnRCiVJXu72GuWrE9W+Qx7eiSwqfqyu3sv3i4zaw0jlykJ/EzMhAoDXOLRIzVnwI
GG9QznhZsRNdowv6KBHVPkke9yfW0N4Zxgk24OFWl/2OBmC+azpxcaysHD63iH4BX6b/uM/bVDJj
X4t8sNLNc6iNYeXYtCbGLbjHt25/3IL3oPq+a5HWQmy61PhbihIkjI5wE16R5r618QU4LFtn8uLF
3Ugzu/94zvMzrhT9QxyuN+DpBUQDYm1VV6r0vFYEBaBbp3q26tJybP56cZ7mPOz8gKUs+282Ya42
0CNYlXmiEmbnImoWk24nSpGu30YSUXUeBkBmoxjoCEaib4cX15OKKdQKrfdHIUJ2t+mJeWfSYdVg
cSiIHnQThqETqNZccGJUGrMiDJwiKPjIa8XAl8pcQiIXxYZF1MVg+SxnPnqu17J7zeloUQgm2y10
ewIsOYiB2zM43vGGgPyGOLC3P90f+hDZ052dBneHs4mPcPEJBIemo7nopeSM7XGZ4PTPQ6lNJ5oA
27+rY8/MFxqX1DCYOTOYMjclEnVnFevd/dRFKSflPNXyNPI170Nqq6679sk/szEGlLNZAN3rP/4x
fecKA27gzJGWV40Zh2tU4M+IXGY9r/OFuP8QkhjDFnYCAenAyfbw+SERtnxdHzNcqkbreDIfGLaA
VTZp1yhj1B8d31Iqm7oW9YEa0ougrh8hXlr9CYRkyygTuRMhbJEJmt1fzOh1lb73sW+SM7XClsfT
iVf3Dc8Kz1eQaUySXo8WE1/nyjXzbDGPv8qXoYhUaSFhAUk+4uLP4wY1W9OtHsipl1sETkKxkGsJ
LgdBs+YZ8ux6dEHWaBtLJ7xc6HZh+Q+fl23XdfezWgCTe5zvvumMaEoAYS5wxU0FGRqnxUyqPioE
ZklPldMMhakKrUCr+out/4s6Viw8D3thZBE+J8/YWga0uDXJVkH58BpT8MwovBTYohvMo3i9eDDr
bhLBkFavJIr3i7rL3oqQf55KGF566LI0qHBGc0ixdOYu28ZTY45L6UiNEL+axGAmHhoSIwvsietO
+Y+YN719/qtf7xfm1Lu26aIFXp5bEmxHVu7aFU00VKKFpb3H2xeCRu16TG0lyXJ0wwJWrBubOX2M
gZGL+Gzg43EBi0bUHztyfWkY2Z9mlStvr48zZtwCsbrK2An0+6qQEhT0RbsvBvwVkGINIDCnyMQL
tMUHzIdwgm+Va+3YARXLtUhWj+MySDy0wSNxZe8hx0YacCEuDWYAAzVRVfOz/r1hwJHVXJTcDKqg
u4IyIIRqxuPmQaRqQGqYaVbCYL3DN4D5UAJpWCgPpTYya99jpM69JkLJKoaJkLgO04EizzEhwRhp
YaGfm5yDOePA1sSofHcNqziJ+HgNfVeXLz7o1faAvbvrpx4QMCQQ3Uc2wAGzp7YH+IuAfuC4BefD
0hF3oaD1WsbruveyeC1AncV3qu6O2PeMfnTlKJd9/PRLS9PCrPcD/8bWTJ7zmqNc5o3Nvhy/t+5s
lzGHIG/F4BH+YaRaKpA2thNzA5l4qICAPSqDSmw2kv2D6+x+I/WDkVK+6N8wBVQcHJLUwz7mX9bm
T8WVEyjzrQq80qCQmHG2yQ8gv/jcvPYgD4/HMQQANSHyxMLP6UtX8Bo1T75GtbtymulJ6MPK1KZj
teOAE9AN3p6DtF7WBOlM80EV9lLJfKVnbtg4U1PeOXVi9nQHOcgUHje7bmFr67j1aC69KUdlKt/H
0CdiK92duQiN4QGNuQhM3r0Vh4jcWxMcwbAT7nkwc5O1j5TmUzoQ/bECZ9SXtz9sPLnYoe8SPR8j
LxTb68W6NRJ1GEqptlC4CUeLWUJf0EL+lCqzTkIKGTSE4Fcgvl4BhR6ZyTOpD2/BgH/I0SP3BO2b
KqBEDRw0i8jcxkXwt6ucAFMcnSTA9BN/TUcJddWrFfRtuCH4919OHKKbrCjlRw2BqCuM2Za50xWg
ItP3Sx+4lMyO4YNh7zux/oaiGIIFkVzcsTBbK2hYGtVcmm+KeuN9IIyFvUahbpKk3BSc0EOioUCz
x+ljZLCUzkXCH4VW97OVUSEQyVurOdqs4dH1yhDrrYlxOo1/Ic6OYAHIH1SCPZZb4U5e1famC99v
0t1+wne9A+ylMoK5tIjW3WIwQTWOfvfXAl/l+VfbGRC4OXo7Yxiy9lXTbKSpncAgfbNgK8va4kzd
hoBBvn+r+QQx/b+5N15nKmkXrmzMGpmSrVLj239WyT4FVXXNOo9V5lOERUv9yA8JHFzGBufIVHPu
6b2GfJysi6kUmJ0y8oiiNIC1nIPswiKxd3f5wniTHP4mH52WVMz7x9ZwRtFpBJ1/xJu8f1QCoVzD
5Vr7j0t7OTdV4+sRgOVucV03AR0Lf77B7eASmt8E9zrnfCtp/0xwC2XbqGGNr9gArzv1z5Lhk8CQ
zTwigAL/7mHhFcJwT43XSkDC/CkBpCCNpFxtm/6Ak3c12I44ck3YF12ValikPXDHgfnjVFve7Q/N
ps8IvuwwCeqd2kskSrynJrjSmJiaLjl0MrOApDyzXK7OcaE/ywxncOJb0n/6dXSTsrxAyim0yyua
wiT2h6qjzP8NILbCV2JRhLb7vX6jhH1BcsqRP4fzdaGY1pc3W9xSVJ9RafVEJJ44+RboxKxwyHUh
e+fFQEX5uV9jmgYLVMbTxx8yNugIJ4nfmApF1nODLqrHNw88J/kU2QasNiyHLlbKf5frusI8VliL
nOVvYBaccSswITYVZ/LEuIoHg5XwREhWPsfHU0hR1S0iF+pOHeUXyVmc233FuZFv2y5hduLBZh/7
y+AQi5imhnZXbNH5jMDUS9nQmDS3BVjD/ziWznFUJj7w8v5Fq/kLltQ3oN3LDwE+/J221/TSYLmP
8pvo5BoHsSFz118C/m739hkprCtLDPPPo7U57s8UmGcYllxvvRnmD+ObarVZwuI4/JQQvqcPZaKf
b+WfA6hZLhoE9dv1EYAYhr8UiCsgHBj/ccHxVbMIAEFDXmuynCeDbkrewRcxsXMq8MJhxM9KDyIr
TPZ+m6Y3otnYP50kysKFRz1SEdk/1UBMeEez0I2r02pL3QT3jho+0JpnhumG55qoTaVeynFCfMVT
Y2xT/jvWlyGgqGBUytN3xgNFEpaxuLxbEfFwvv7D2lI0UuDPvwB7kC0wpdxpZLkTy7nxX/ynT2Ot
MjcyRQL+sS6lc911iPsY67DjIzQmv6J6uwuIQFE9XRt8V7H8hZNz8HjnCYeFO0NT/IJCGLYq7LCN
uTgSNep/+zQlroqLWyEyKilX9dR2zlgN6ygVZxiQJA+iO3L/AgLtg2dVbYS6dWqpAONA3DJ9guLC
XzuMEOd1d9ZFQL5OYjkI9T2g+UF/ivxO7VI/6Upqazw6gpWSdQsHU/ZUfIgOwaCYSHPASfNebRj0
sEYUTVSPsHQeclR0NDyWqgo3RexUu5heJnncQSvVwCdd4JRDbWo8XpE19qQXi4TWETKhcxQMcc5R
YgkZ0WS6rBgCCU60dh4b2CWQav/+I7lKTO//85MxFkk65dMM6yl5YSqSiqeQXS0uexNefbzf4gyM
8rRpf2t1KoYHbs017ZYX6xQzi7ThAs+Nwu7n02UvHaVqqJ+MNGrE4iMx3SZ8w3ifrT9a3novxzE0
pU24N7ROFGRw8LGaR61y2CorC1eUn3t/ct92XWLHHLzBPL7BJPHXiJ0uljrQG0gQEGze74Mc+Z6M
QAxpZibL+CNsWDdyAxeeWCA6AXT1O4dvpTxXRPJMCmW+Fc4JgJFpQ/idyvlHKJTo/cxZfm27Knk3
+0FfqRnOEyeoxhlR8HjZhsRd4SEuQojkNYO2AC0ycpV+RJAqDl/o+rwXqCK0SR86E//d30nsQzSG
6UPFR9lI+1zQgCF3MuWm20sitz+nTvn3tVTY7trfQmdimWnwD5+x4hlkbgIRm9qrjkyFqDIZR0kk
foWpYpsOir/ZmXcK0HN6h756uLEBWEZs9+iralAl98iJm97hjwQpkYHzUW/bftjhAjy2Jo2UCuab
jzYRSMpq8SD/phe1mV54FPTBkLLQd3+kMzkgRjCFexWdyN1XS5Q6IKXBr1GOiIuCEyqDotNUfjuJ
Vu4BAvHs+83kziB7kIEORJJw8uJSZ4krKDIr3owhnzKggQsJQ4W5yLaeUIcTvCemthIESuv7hUyh
nsAsClxHDH78bsdoi6l/iP4zUIsWDZnRW7DEEaF8F/wprefsu0X6FgyYtjJiVRgEI+F/u6HV1nwR
z/X3jJPPOActItSAYZdiCHOBOGfNzEnaEP26xV1OuFSWRXTaaNLVp8MsRVbFlEmGWL2HlJto6SgB
5UU9ckFXeKTbcgfV9xm5/p0qjW7u+glrO+z95aMH42yCdlEO2sS9mGvZNItLyfDL8FxTHRf1klyf
tCk9KnJ99CJC+wIsVL6fNNoXNZ7ob6BF11xu7osFKqzgWj/VTFgS4XIa1hRfy2R8tKD364kU7rmk
0WFpd/NkOflhl7n1kNvtB1isZ2XD/85OnJo2UditcJSbD4M9MnYYejUoJgu90E2+n6bZyHR4LpH5
TsiWjgJluDopmDnmN7rTEQVgCe18PceGJDzftw06Sjqe6Cl+YTzaE+/4dniZrngHPkpNN78rEu6f
IxmLodII7x5X+PNVnuxYXI774Gcp54ly6bBtZYX7yar9rz6i0JUWDzjomLeLAZfR80IPlMYCSVfN
aW6d+60pUM7qyzdSXeljGawrqPxGcOzw4/aAR3RYskI9IspXc86J+82/N1LuyeFqfiMKnrLEDP5i
yHiSTjvJ+txN5IUKwSKBnQD+lMmihJWqW9sEU0UtJUFgGBXlPJ1vo0gE4c6zuMzzDZAC/gbZLpwZ
2kEMvlnNiwhBwWlNbBIU6Ppmbun/B1TTT7q5Cg49hav6cEJGbxm/2Tc/hwhyYkKDOLtn/SPyMzUE
w6XAUlHD56lue8DpRoGCAKRLdss9p9K1nPcg7PUMUut1EK1EuUxakXwm3LVftZ/NVV8CaLJeACS0
gaZWn3KWZahLITStZ7XSyuyBPiSQ7lS0ClE9c0CaOmYukfzYpCNErfbGFvd88GlUJEPGJGM8jju6
nJep7l4vPP8KczD0VfJLEvf6HyaYzaW9rmNzu2n3EyclaaJ4QpITtt0HjHOKFngsTvozX6Na4HsY
xwZbOIFp5HJ+a6529loQafJIMXhXAky+8xNKhdgC40NcLoerqTOH/c4rHKkMyL3TsppxPGj//vJe
9Hoo0XpSqTzwQ4bVZwVrlqJLPxnsPjURS15aYAch4SgJCRFvGcF0PgEjofzoV/duuDzasxDmBExu
43xdDuXF3pPntE2hGXW04NJywBPl4IT5XrDrzR8ObM+w6R7g3tdTzxtZKX84oG62El5ikMji9BiK
aBEZNmjTS/R5kjKGkMCR61IkDCqYKOzzykIGQQB4wRTd7fCzcO2Nj5NCLUD2XrohuUaQUZ6MGzII
bIIUE6kx/eApyhHnUka7NUwZQSUyrXjKD9jtsrcNPvfMdKBQ/3jUWsR1sbPqNx31/2etofqOSneV
MyakgmNKaJ8YcLisgZQhZNr16SfopBtH5vSUWa0ufP/3WLJUqBA/VlvKw1uH3i2Od4G1OvuJzk9R
yN6cMpGHyZbRzKof79QuAK/W9WMkr7QMgaEG8p++cTKb9cjRtuwiB7f8HpiLqfQEuZHFksK01xJN
VBTj7gvPj4Bloz/90o+ZrpN9EnCCMiFiJk/Eo26QQXXrfeu8xE7gJrXQtUbVUreEAvXfIDsxWzad
X3RM1fi4OHjvNSJ5AcdNMCow4em5jgwf41wSYzRT+4gnTtx5KJgSK98vGmcHoLJllaPPPtwSfsNp
cuLFVj9tS2lo/iaOILPvfLrUtbDSnrVHi+a2aM7uaVkDoP5aynmMEK3m7CM5FtK3plpIIyWZh4JV
4sguGbmVySp5KHd/XF2l3TDVoAeYB4UPM3ZX/fj9BZrWM84Q/6Eu6mSB355+4z9PU1VX9HZhE3k2
DJSJO/yD/MjPfy4PtEaj8UdeBkfsXGlobye3ge+x65z9488OOvpHLCVPdYIZtielB0JXEZx2Jj8a
yzXJbeLDu/KbpLgzK94unXtXZSoyh+xFdQPlxQfkxBMWOMXziXp7uI6avaG25keSy/eQGtqjUsEO
UfwAbwMqbO16Ds93a1A07xZSLNPLSXNdo3BgPcpWjLT06t63Kzmd6O/QCoT/Rp12HwEgPACctC4O
FzHres7LYzkkJKvCqhun98lceC29v1QSO5pC+dU3La62OPPbnnUWPMDUcosSZ5LbL4Ku9Lv8YNXT
1Np5ddRjNqYkNqpMc4bPH+R8F5iPm1RqXdV+araB4pqw313FczE9sCihIcEsgnwMfdrvetrv614M
aAzq0YWQbYdG0F+QCkJxrJH6AbSKYvDKqgVv13MUtnZ1EsBpDTNyHbKFSG320nL3c59icL2psc6a
F01k6ZKypeS4kSXUjecRQN1JbOgRm5ReBnIBGRnV+ShcCtBG21h833ehkBK/WO/1BwRwrZTgwkON
02Le/Eg68do7Q+Zbd7ACt7+XdHkaIU/wjH27t143erOQl1aau1c5W2YMkofBQuUhEjlapEhvtFjy
K6LeGCoS6p48xVnDkSZJdoIVtLp+tF7p6QHP1rxxY1CH9Gog5qG82d5gjDoC1K8eqb3VVmKAXL4r
AOMr33IP9CGAXvXhuPhogtyYo/q3E3nEmXQi2WsXy3uwMOrxzekKan8HDounxMo02MaKN+R9WQVx
cBwjAANd15jF+7AhWUk/5wrSonpFgTVBp29Zq5dUlfcP4ye7+vdj5BKw/8m3NOqRY+V784+u6yGI
PYH9usXMeYezq/HdjZpCXL8ZI2GvwAy8jpW/h30JaVZhOJta84ELm6x3h77N1ISrwv10sjs8fo9a
aRggLRMN7I0CnshLhvRVDjUUZjc4z82AqmLat0ANkrUA0xqpctZlk1pHJYxIfe6EDdfMswG42iVH
SjkoQD8xdzIziW/Gai99Fykc7fXzmVM0E6VayS3DwaHV8mBOcWshORjeqzsuw0FHUOWsx1/wyDKP
eC7T3oyMjHCP9CUhTVH3XopsX1ITxHEnbl8/up+LxMjE5oEycPMysipgie++qarFu32+j0fNl8Mj
OzO0MbXwQvyLsCg6ZkllLKC9hmMrx0pHL4WEGjbhcUyFysWyzROXl2/AT4/YzISuH2e7bSGUkCZF
/nru6TqqaoA6a4W1Hlz5nI1VDQWmrIvRm7ed/pqj9fTGuIr/1dsiK5+H29f8dBdQQJ28p+SiDYL+
p94PbZ43iHuaDt45e/QSx2VPWP+N4Ou14n62YxzpC4dZgiex6btm6zYadUyEPCb3DGdtPxZr9K2w
2Q40XzmdQvTScFbSc/Vef5jdOAVFAzTAcwGGFTCH7RG835bVCMO+mDmCLWM0GS6CE1YeA4KUhs/Z
uuE8ChYYgJEMwvYaqofctvSiEfBQ5E8sja/INAtAy4XxOtoQwq8fuXjoEnImwJfBbnsBgbPcX3Vz
04gcCEpVutAvfUjhbvgmd+ci7j8uUud/arlAa2lvsBtYSu60JUWqwGkN9tCDBTXgar+IrOydFkg/
h1XHE8oFO1P3UKCGLxn+Mic6vOY5S3OFwUwUcWjY2ydCbxi89FnIBCUwQlbk7vfj68yoaDwMNRbu
CF0GumKnVnM/zMnt/4OKjZynEfjxItA+NDvUTX5no0tdgXID2XT1HtGxLEE1M7J0EPS0r+/Uf0Rr
otbImFrbV+1uLEz/p+wee5v0duZkhI6v4R7kkUB1YwhJ9wFSlCC3xaAUKGGMWeVYfLknnnpUvzBy
ou3UINo3LZATQlq0Ewh3NV0l3VJSdDyyVRuKJaPpop/zB5rf/twfQvViK6bFi3dmRxrfhnFvYBRw
zwXssI8pyoHhXNSs9I8NK/Jy86pLrU6PPMcR4XCP6wUdhAMOOKsocC7zsX0JlJq7ueFH9DseFtVq
5y2E7z/feTG3chZgKOGS9YRvNBGirWCi+U7x2pAWOBtnrd6SPR9IeMV5nsBNuF16CXVNhgAAP+JA
EY0K9OsbafcB9SusSBx1AFhCZGUf9yXSnieY8lAO1zbSUZWfMcn2Z3DOAQwpFeBOABnkCXB4NKFx
C3mJRFBLBLMg6yAs8HuxKq6ipo+xj/8OS+7G2hy0gjuhr0QcQttThNA1BDMmYhkPoNMYT9cp/sof
S9WrHKVtBkF5iB6kBmanWmgQCVSvHr4VkxQRmTDIpLlJj4QwGpDwb+Ypz5iQTiITMxUUmJzwjY93
3DDTyia9Tg172Lemhzc3gXX0UqaxXLJAazOqfoEJ4TurI3WYRLBJVPprB/YtOCzYls8fFSVP7QLy
cZVxJ/IfpBd36HcP4vdl5QU0OytjbQW8Ss3H/jQDHpE78W/8pKkr8n6Xhr81DdOSp0+c8SkS6DiD
0/wGvVeXrISfg6SfMJncQxoo/lLQlIa5O/8MW3NAMHGoWkkUArazDUkm20rrwfVLPDsAGa/8eagO
B2JVSkRTFav9ZhdvfGPjTCTF1qrw0CzFGl5uoZLuoZJusJjo+VA8XVc9K3YWvo94vQ7P/P8MAMwX
zLTvYHfJr8e+Wu9/vq4nshXqKaJVO3lMYy7G/TG3yfuO4itIOC+QWvDQimhg8CVwGGfO/uHTEjUW
s6sbHfUaZ3U2wgafJRVvZDgS0+2wCY5yskpEtBOs5XPoWG9SW6g6jzy1EkO3BqqIE6b3qHmKfq4D
0EmQYwDdsssiQKUdzC+f8eNyBIW7U1JXc5y/44DDXMVNX4L+s4XqmMIqA6yx+tikD63c8bz3G7ZV
yNOUxz6qkg16XDyTYdjOqSqOXKfFKjmGPtLqtd7HMM3czwIAexGWXA+7YWw/pWnAeQL1LubC62AK
906hRfR+/edz203mXg54ao+xOaCPxCXEAW6QIKeEFE8a1d9sbdR2M0Xc5seRtEVR/UbXRyxO3kSD
BE4F2ortGusl4n8LxlxlnTU+NCELBdj6e5rbS7e6WR2PN1fWOGjeUCxli7d9R5kKwTMcHfOFs4D3
CLcxw4y9TgyGNJriq2PlnIovh/ZKhUzsInaWP8IL+hH30inEVccumBrCjbOh+bIOYjqVMcyT0UcI
DZ7pIxZOyPKSAVVSiDRcqRViTTAvLVadTbY+XYbb7fateBVHaZWbnZpjSilqigbavULQ/1P8LDWg
gZAEShmlhaoY5czNyw6Nawrck65FAG4/NUpRR+tyIlk3ytFrKJVW+axYcVXKrd56eR9OO/LV4Qno
MVyE8rhxnObmOT40IzkIYSVmqts/orVZQLpsZttMKdGgTH+FVxkencEXUnt3Rie63Ami0wz0betx
rmJSDsw7IDw7jzvhTgFrIp9scAW9crEPy5gWVEImTWQ9RJp4pskWKYnr4BoZfb6ca6hs4JY5fzdJ
3fyjlcJYNtXBbksFnR164a1AUp37A9cssuzP4kfXj4B0Y1HlEeWWOW2dtMDbt2Fymhyf0jVLdO0A
i2IAO0YMRnKBk1V5Lob1aMow14PcFFY7KGJk1Wh/m5mIgKLtWjrFaasHkEzgNXH0pzdiHwtb2QZe
KJOJ5+fWO/OkgCq1JH+ilkzwwgoyrafrwiBv4UE7oHbspPsTGWOVcee9z9SbDD8jEz5Yehz/Nnd2
B783y6uKBYGibsnSGUqsj44fad3XGYmg9/SbUl+EFEdolMNfV06RHGFaB4dJ208kE1EUvc9xR/bH
9Q+2f12jLds2+GwsHDcaEVzdxtF3I6YGkw0H+W3AJtBBN1J9QhU5n8GhsezX10SFyuby//0p8akN
YlJOL0U5m0J/viqslTZ32/Z8yRUqoQudzhLPFgrBPqplPPUxVpykwjTQrhC0PeaSqX1xoGiMT2GT
JKYZQg0wqXwEaJATY+mhFOBt8YUM+GUaxjh4L7mgVJQmaLNFWluhzhdRlJtTCoBsQBOK70WiQuOf
/UAtLBM83b00uvYHuOEFf0RXex0AbnFfTH+ZOsBjiVnWFYAlhywHVA1BSxPI2ZGHzsTxSslTgl5+
jWC1ZDF2RLQ8za8OtXE8EiJhzIq68wzeo93teRIzUJkPThDwpGewpABQ3wlUhG6HUawvn+gBPHKq
Ua5/YrvAW59wQAUL9fZemioD3dKJ5oknlOvPA9YqmNq0uwayFLBuAA/fuepoU/ODEeRC66EZmUVE
Yd1s9wcrQoy6gcR0GGvRRlQ0fCrnN3nN5O2sT5hGuyV22Ksxbv6oWoYfHC7ed2/yBumKezniL9Cm
fKGgZcQjulnmP4slLSN1fqY5fet+JlHW+mUyr6bGfA0FxbOERLmqNMGZyLysU1Mx8nOXS8ETJ1mQ
LNJw5cRpS8pCyDH+FWVUfytRb/inBxrsaqfTNX6v+parrgKeUPm9TfLXWFCA37o9dDtelMF0c4YC
gre66s9lJGv6ZBlWViCL7vDWs3nqvHV7ONNph1mOsk5+zWlOITD4/YEOVkxZgDmy5LdSdOoB8NDr
ewvgpkZeAFzenEyS/XiRrs/f8fDnTf/qdjuobfDt57ZXXZY/zJ8cze2U1LjK6zx2V9/UKVoANDZ9
jUb9MGVT8Y6HJlsQeAUB5RgKtkIRL7poXHVKOeN/06i6MKwLTaZmgvlszFBMZYxvxxvdpiz5Zzk9
1v7mck7wEN8f8MgSIne9Z10SCbeZZL/6Vzd12Z2SSldwbDP36n+7rUkmfugTaI2JPJ30h2X24YiV
db8zjjnvtWhr+GQA0AhPnJBB3xDN5vyjdwSPUuf8Vtdcul63W9NxedEMH4+rMAfZrFvH0l1ZwB1M
pVOamLDOpe1e3RKQmc8vma3wqyGfHBEY9Wyi/E6x77mfOXlPfW8Y1Qhn9y0FJTHZ9OGz3P5oTdYd
oITzoBR8NI4H3BzB4indrUfi7aTBHo0r3rcqoW4WB6plP4bHfnAXNL4E6nYBbVb5g/oJvR1uuz7l
giTmhcGPQiu5cP0TArs9gQmODZ9O++XofU29LuBrQLuBRqP0xou4bYSvmu2IBr/HRLiDBK/yPwca
2Y0Gt7sUs9o7Kr+vwt7xYui7eNd3vZxL20ujefAGTOzcbG0kLTWUrxGMwLP1EjnSGL2WVyevLEFa
9388ZcEfEwo5s9WqbDPCkcEwCLlM81XxJWyHm1ihzWxYlIXQTZ2adDABA56g60EET3qh4LOqvyJ7
gjw/vd6jNey9OcbI6OQgdlMCz/BFk6rpExjMAuIotX7+4SBtqgx7LKum2/wynho7ObT2sST02Lqi
Ia9gv4GnKapTp5ZQW6reEhlrLkWAPQ4TofZmbc4ZwfY2LZFYigkv1n7vpqjOQeHaqyZlOPF5niBm
m0oLm4+rTK9eZXmgLavVbSb1XkHPPhEPHebZLmpiLxNycqDlx0OlGI2SjCtgMtsMtZhehm6BhAeK
0HBXzAc6Zsgt3LAYZ+xqtjbN3Jm+JjYc6ny5M100la4Sm/0IiEr6sOAoozjJEVsgPrA8hLIlDctl
RszwuJLjtz6uuMBOBJOqLb4Uy2BokkEH7xZV5o3GuabavCSkotpM2Z7dGLeUcAepuWncRPUJt4hg
ORNdamTPZIwbyUWq8jaYW6WsG1Jk+88jtvmHLrS+jJy2r7Q0JJe/iLboHVr0dMvvKFkYMyVOVJ2/
4YjbkYlDMGAFL6zPo+RyhS/iZW/w91dnL/yRREHpbzO2JSddTQC31lyMDFL6PQcLk0tNjo7W6v5l
izRXmWptP++PU5ACdfQUXbcXh3CHOKRlIowqRxUvLxQhPnMhx2Mn/IQlo+XMbZRW8XRviMLOgeCw
k4BncBL8FL+u9YCCDvjm7M6LBgHJgXyXkuD6/FsgvC+FSQnEjSbIdkdbaKW/y3dDvxgNpfiLQ1Qj
1ZmhiFY3AcCNoXvQIAajiqJDnx0GEfnWHha4LjXFRaCxTQ4kauib3+uyeH9cjqCgVwKuz/m2ANDw
Iz5jyMTK4c6N6oWRzzcW0mRDp8s7TCDRlQNZa9KSlwlL0EAMfgWDV02g2xKXOweK5VbG1iqimCii
71PiUpf5Qn3/ICbGCydTLzH9ucniUfIkwU84DKw+T+pu88vu//qoLK2fXsW0kW4vbVePJls8KNLy
EX7fmTPd9X7PCKrztKH+Jh5rqmAVBFfZIcFmlfhev7olsBV3j6zRj9w2VLCuNNYQLqSglaId5JhP
h8N13uqO+zKtOeyyW53QfvoDbXnGyiHLGqHYwMEwXd+NGNojbTiBIuk1tdzihUTa93wM6Pbj9Pl7
WeS4PkiLY/TstbzWQqVFyMv6KJ32aJhSZdYzxQWVi1P37eNKbAvTxAfLSeCGLl78To0RKe1YYM4w
85d59aPgrL4kzdH8DTeoHKgY8FZsoeSWqnmwRa3asX0/t15DQEiUN1jzctEdAwtvE5GyxZp/iuWT
rTkZ/5H/klSg0DBi2NyPRAkSPQnTPMqLmDSPnbXmRkgCKw0UpT1yamjClHxZTm7Y/Q0hWON6kw19
aVzEB+D4J5C8zW9Iy2njUbcL6Dgknl0sFFBdzOyBKGsGU5SI3+JTTd70T+HgX6or7PVhixmUCFOW
B0c8ZTLmC+F2E5TCkg2CiBI/j1zqKl7wWlvkS33kyYU3XhFMzsAA4T6W/9HZSjZNCNbpQ5lFiJd+
X0PuJHRLk0AExbjArFr6RXW6bUQGU0bdRLzex1D6GEDSj1ZG+nRsfpsjTPcgnUPl/sgVU+K99snq
y8sESMICvVcXlPL0W7qZXPPM6OKhvT0jdxjF6kqdmwacdqtZhoZ4VU/m4J9lHah+JPCOMar959FW
mVfkdN9mJ68lsri4xDypAY/mlHXo9iCPPk0wraI8B2TqiZ2D0cLpcN0C6EyF1i7eO+s6OvLw0cBQ
H8lXUEtu+GFbwXXSO794Mt/37MtiFc7Cb7TIewsYNu9Owf/tD5H0mmL+eEQLRDTRJ1mGxIukelv1
AqaEA7tsn7Sv7Mveh8nEPjPDkCnG5z4RN42CcbhGs1Ryl2veC7vAwXMRmAyPRFhKWFK+OzkWbxId
F+nrBgU6BpaRbb6l/S6gp1NTsNJGdy9B5eDd/4nv1HoktAcnAA700t3shepdYhHZV6VMgpoiyAYS
seqVheYl7UBeLn2fpjbU6R43Am0X2jUBycLw9PQhBBUSIJuaIybw/BAVeII3EGzs0zYxqtwm/BTM
dw4OswZuy5OlMFcWiDxCXfuKadEz/bzP3xEbNUcPiOtWwKvtq2y1t3NrirI9IJO/tQSJJrmmu+9S
OHSS/NpW5Ei+TDaqyJanOmyZyp6vtrLZU9IJFe1RU+i8U1ozZFBygKxI00Ml1DcROnY0iVyF571F
6IuX3bjSNom+fPXgM0lmWTy6WuLtw5znhXX4AYJKFHANmRXLycabx3ESqylA4/PnNSA8/Q/AXD3e
OLuDWrl6OWLhK70lKW+6MGXm9cchxvJnVX0CSod2bBlLb/Oh7H6GUOlfbNFQyA8kQCKbL+C94u/G
C6T+E4el2tT9x+sDd7GczlSO9w31N03mS8d34aeLcwuGOkF6OMoCXjZxIDet1oH/wN3VzJ1n9iFI
OTumeFEenlnE4uenxjlpYo4Kq6c5bzthtlxAGTw2IjqeV8cl6QahoGon8rlFWJzZmZzImj9Tz+wn
Mt1wWZ8tvMgqkJty1rrcmAuqfmPfKwRPNun/ktlaPsTtADKa5DB0O5Mm/dUfj5ZosjUC/gQxDMTT
OycctGcO6xt8EzJTPQWxZG1/ouHCfor216ZTD3YQ2yZeduSf7BFNydEGbH8AGyy1lufjG6wiho3o
ETiOhUh/xvd5fwkMugb6G64juKECB2Bu7PB4UVQ7V9W5S7C4T1clV+ZTLrM+YhYC2kytmOhp+vC4
93ebARvxzar0byX9DKm+BjJz5Ysb53F0tRSm3ORtqj9lrtC6+vgJwWeHeXtG4qrRRo7eWNbHfIcT
TCZJfm790L2pIn5dveiP+/TeEWlDpi6+N0sEcgu10kgjm3ttPd8sU8KzZGgsvvtcaIrMn9scy1yi
+rNETzLvuRbmD5qSZoOrm5f/xqPKzw0phw40ww5I4qVdTUhpCiGT8WlLZ+jcL4J/D48woRxuekxi
oNf1gXp0Dt1h2QQDLhqmxDjAsA5bYYZvhkhZ+mG4MMR5pbmpczmxZF796f3p2Z6+eWr6VB0f5fLz
AmmBHLaTh3JBDnuFVRMw4lbNKqSJ3H4T90TMH1jxAH3NDEZpfNtirYG0x9ck8xyMw4fTUZgaPMG6
pv10jwWjN9b1E4x+TQlgfVZldESVWaRD7sAXP4SfI9bXQhdNC6Darzp0H8f3jplnWoWBUnpSfj25
E11bSOAaV43N2SQDfYWwAEAYyyvRIlI+aEm9HVCsMtEzwOFAcs2GJ0WPzEd9WP01qHbS8nADe+Lr
zqRHsENn5X/DoOKwKb16lLk6KROPollHmOGQB0lbpiYtp2EkKE8o+Ni+q6O3XvPgKGdL/VLSJPHf
VruC0qhSBeUh4kgEqIXi9tVvXbKUnFsYzjwSoNl0jtSV9IM3UOj4XCIpvzixX5wAbMuCyNf6aCa9
H/ghKCPOK7Cpo9KzL8z6NmAHQw3nmcjlYB/sOM0vbFqdqZmAnObYeU7+HFvV7EeUVBXdqeMI/sHb
/mrTfrSitg9J3WSUSO+Dlkg7QsrT5gv839oAEVIgYbdrGQOeMrhYr4cR+9lsQ50aW+QyZ/MCUOCE
9ZNEg9IzcoKOzPcnIOEKkaTYOE1lyUS0TZzE8eJ7P9KJowIC5Ai9YWLIPxH2DouY2kYsPYuQUI2C
/lTNE4JR4JB0HHJaAJklw+PasYDdPNBZtogaC2PMXp8reSkPndTnDjpy0MBMNgdHgdqylOZ+JORH
b7lMNy11ijPe1sVbg+7VilG/Zfo8JLVY/lUaxdZ9GvCHLXBSGDrnAQZzHCTcRW5EJYBiQ7m2ZrAO
a5QtxpUnP0VTkJCD+cPpDEDk1lOrwUe5CYJv0jvHwUmxR1Glf+df5xLmeYnnRXzUwAmhy5wjH6d/
UM9zCRw8LDDuM+ts+mFRsHNM9G89odXcVz2iB8xV8jtb3bjbMesOL8wuCG98HGxQwRhev40viDKS
Pne/HfOxfd3y7G2AXcNN1HsfzLa2DQMynls4An0DfD9hOUqK3p8a+kH7UN+KTa/JB3qE0BsyVnjo
Uv5mAaPL5pZUwYYZ8vf3FPsPCmUQTZtQFc7RI/+jNWeuSCUfzyLpDnOgibUmpKECGNtaIg6NTRQX
/4AjVmo3LT2uClLx5w7jZZiJjo8h07LGsW7HrzADv23pfb2kw0DfDFnSl8zR5hnZA2AhLvVkXgOo
GFaHl4Dvl1hEhJAxybSNUwXYWpZ2Xs+B1mhLBArBSeRPcShNtLcLFuEVEW4yL5sXxGfb04ev3iNc
S+uGrRzBovG2bW/1GFplMM2v3hxOOiqeNy1uix2kQ3ieCBdKO1U90o802eTKjZXjAieJPAMvIVVW
Hg7WIzWS8zuyjEzB4b+rN17q8q1/eJclJsVGpx3tNQMYqUgrelA+YIXWvYeiFJi3Fkz3OS8Sq4/7
98TEEWONTEcppzJ5wztkqvI+OwcvA8FEEhKJIwUA6XfLMnvyki68bSI5SI5almEP1SclXGT/f1hD
HFw+Ufvsv7V4PaK/LQjutwxGI8cX2+O9MzEcOymI/3FtJwWUTz/0RjGojfbJY3RrZhrBAUvhGMLN
clATZiLk1tYcyyBeMW2oZmL0H8p+0NZ5itnrDqHB87NNwwWRLhfrXTOr04QniBnEeUSvoklGDwTl
kOAgRv2aCYcQns+sQz6LR5zNbGTXCHSUO6gTOPqHsEw+kHIqTspjclfQWC/GBctCsgIC1/W4NdgH
pM25YlBegp74S16At9xzn8TtAWR8hux+zbhcXFTD/zJlLTlBA4rgb+O2IAlycVyjgXppvgRDF20J
JqPZ4j2keNKPzFBhukoVKk4KW3eN9wD8xaOeGnOU6qCus33xJ1aCtXplt6FseRyRzZ19usecAr5U
j70pVNFZMyg4vSVCHIXQaAWZPrB2IAtHRq0Libify6Oe2onfqPzv4AU74nW68dP4h4Fh/+SpypSY
3qESBqNYf4CTWeWyTbOZaFC8pyLwaTz0mR+4rYWvTt3Cu3yDqtozxdv4cbfngEn3KDdtYLCXdK0U
19vrLCXGoWW/Ixc1xO3R0n18QxpKfvX4LqMSHT/2BHTyAWVKsKT1iSADBZWGLVFo+nHvbZjqCpdv
jizNcNmkJywry1ugs9oUQLgspxGxK796x7f5QbzwUGcDzt6Q2Hfj5eHxDayqPJtTBZ+axY9LC7f8
0lgdidANYWHk1Emwo3OtBmASYeD72DPOwnjLJqK0OE488zfdTAf9hSZ7C8325SbbKKRdVqyD5won
biQ+gyn2oQS281jJjGKMJjqfJEX7xPsK/tqOUzJVZVEadZZXt41PiCIpEdoBQghOimI6NUfH8XI5
jxpEJ/ejCZAn4cTA7BmcfPco1y53WSDJ4hnxcX9a/BzpJsw2vwkFhkNASBAow46lyMH0IV+sSfun
wbg7i547eWIgeFcTLFVdSYNMzTPuH6KZHPPoWr9R7doxRvZUbRuwp4mQaW75Q+DDhM18FmyJwVZS
v/nVtSUtwxGHs350AF0oe/madOmZZHfgHA3Z/y28k1urnjhgEigTShJnSYvqCwfpAbWUUZS80+xl
nVKp/MB92YS6qARxeR1GBGQL7bSijeluR8cVVglcGQ4fU73e1sfMbJccKMOiW4AN0yWzNi5Ou19F
YESDzA2NkTJPRBDHjdZyN3t+kiof/h+DrkjyUXE4DN5xJrycYrq8Gyrb7MhmVcYlWoQ+FtLQ/W0d
iDS1oyfUvm9JMhgNf1ZBtQlnA54REfpKV4ShvfKE5vhQaoRpyadvpE3r3gvUBWr5RWe7Lv0pJd4m
WGRs3A2xV/+ZDAfm3IDYgHS3YnSzxFCNmg30e6D9OUCMzK/EQMmbZ5onP6q42epIv7B0LTWjFs7n
18jgoGpUsuvBKKvm/jwXWtAdOmglTnk7lODFzFVFRCvIehp5azZ7jEGkZQpGmqxLmQPaVFT/3vCc
tSbFmam2XdrRckzquSbOtOagq6tYzJDHeISahzoA0h9i03/txndoZHeh59s+PTvMkTpVknoAYVOn
+d17M6K18g8LQCCfamw60mwyeuSGQxLIWQkxP0t3lm6mpEL7BEnfRtPMwzQKETI06gbDDdySJsBA
84EgVGI5S022fKsLddJQwulp30NLM/T/7zJT7SqVeV/16FyY9e2gTQh5kisy4rPDBPsK9AQybKGY
V4Hf8xhEP8niHIhOBATNSlZUA4mSXT9/oABCdrON8RTX2ES4Vj2LB4ASgbUdYcuXCTTPHqcvnG6O
vr6/G0YB4WCRj5q9rJcjgb8m0m/sV8kIwndYQ91rDXQHx5KLLLt+r9b/TpalHE+Sh3dXic5zyni6
Tc/o5HgoW14zntEA1xjhHCR+vnUPpJ0qZbdvo1m/M9AWV2Edj2l1jFkgk/rFQAsKF7CotSISw5mB
w0/JAv9U8O6QS6XJ+mR36ALnyKtvzSKNQOsNcgiiE1yIVL2RY9slJamu1lPhCHocUB9BkfwkE5bH
i8ghXBKm4hFIx8RkwUUSoc+HvOFd/m+EautPjCj1d2HrFLZaP3BzSVBWzLdAfP18/WxnVm27L5k1
3WUunYJLCOY1Y3FdNf2r9EJlF4IOBuss7EDTyWvGpAgfGn+PZxIAZnxdg4d2vkjoMZXB2NFOigGU
5SDcpzX/wXB7THWittDDgePL/XFR0poBgjSbABNA/DZCZa9qAvwQSy6wXryqYVLWvGZr8QiBt43a
0F+s1U3yR8RwYg11vbHFbA/kClYqOHANJUspGjZTAChXrch8Z01FuVRFbRreDmriptvonLX/6Peh
7sOphpaIjUYd2E5EfA9CrsVGlvQ8PKyz2yWuejVIJaSHv20fcJwiPY0nPo7jJcjUjLFw25JH2QED
r2bM3SN84lOIIECJbdr4qu0tjBGbv/Mmo8NAiU3LGqSmU8sQrfXpZHSeQHOIvbIZ5XkYfghOhtNz
soal3YGLIagDrE8J41WZaFaLdx810c3wBFR8jhnkLrr/ZCvtQazc9Ny83z8gzLlO4X6pUOsi5NlE
eydy55SVJ0uRi0Rr8B2N7hD85pq4oDRR/GCdE6iH7D9huF/0zG8bcU3V2k5V/7AC+JKkT77QwPRS
gHSrNI/BUvHDITbjl/BGoN1Y+0VBiglTSFmXodYk6/GOVu0sN8SaAaSIrWuQWE3AHtQFYpIDh25T
aGRiqOxk5K5fh8XPIvZ6NWT29j1kGboNI0dRcQh0QYhA9t8XAyopSC5QOtWMx1pH5nPc0dhlXYY6
GO4i7e86wmIzF1mUVFOQVzwYCTZESOtV32wncC1cHYgtiIRAUABfEtJyC+EI32QmssLR2FsX1AQQ
WfY/nzr9CAVuZhKwOPsUd4Tn1s2Y+3LOt/h1IyzsS/2KlLrCVFX52/slk4rKJPEMSxsQrVI97+zP
P3iQjZfjf2iVSwLxhvMqowm0M1qmuAyuxqOUAvzsvqzjTYa/9vArb+cVbXV8JNi0I5pRb17TK1mQ
MgdW8xO7D1cj3MuBt9a/1dP0hMwZsPZPySJBaI07VzlmS4DFbtyZQcysJLXyM6v/stwzr73ubdd0
WNZg0rUWRYX+9Oze/xeogtvuCAlv3efdXOlaRKFDAzxsVpsdq3LutwO0qTRyvmKEFf4wJZfRuRle
PrmfLU5uOox8YDwKgqgju8kCZ8xTra1k3X0JDfGpbKilfHQWwEdPy0AJ/ehDxXy2GN6CuhLI1qO/
8ty1pfSEKFxkPwmQebgGI2iHdMWkBQFHfxATGKdEC3n+sFU6PT/Xqy6Y22R1mh/siXZFfT4R06XI
Y3kpL856CKlZ3+uh3aY4WsdlnpCki5ALOCvG78FVFtyitW4RgK8zlaV0OdF8uxqif3ojZggFTHqv
P44eIrfYFa6MsEnqse5ZfH+umZYw9NEBzlNmXh5Xlj1Di13F1v//9/mdbCik1MHnWQZ7Q04Hzzld
LOtYg6iGoqsVPzHBHTKUg0s0M05sBQkaixm2H+XB0hAjAgZ/tX+oQyOCeRi4HVBDTFJx6/CocI7J
Rx/xx/bL0SXi0z+L9vZ3YsBWtowlu5tCnAREC+kp3JEYynPHIhSdkwprmj4D8YI+pBn2oEvWfUaa
+b1Us5RsHLcLW8UvK5oa42T+voWl6Px2C212n79aqRZnu1dOLBj8PFbrkDseX59APnYpZ28Y+nAq
Igob9u+0HhAFJ1Og6Pmj+Q/O8Hg4spTS/nkQLN8Ei+2J0gDCpFLLKLGkP+ItGv4Jiuj9n+5S6O+B
cj92BLc/vyD/GJJz5SCJmYBwgt3vpP8GjDmPKVOBZ/wuad0zPs+J/Nu61ORw0sn2kFeEhxxIZDqd
Y2GIIYO5klt16UosFfNbOrOHm7e98TNGsjcG9zALIcTt4HpZaa/XkSsuK+jGGvEi8KPwPGq3wxeh
IIQIBE29c5Sp2vNQIG5st8+DIDvWg23wm43j7v785F37KVU92NWHvr4MWq9ZvcO9KWdzQ8CELiVm
0Nsb8NH28N7XCYhiOsfB289E0h/aaUO1JcMfkyiz12hCvaaKVBS1PBOSiGSdV3j+1zXEP2fc6INL
e0ar4Tm70ubO+h/5DLGtR7SwyaBQhsIZ9vMrKSSlCf+rzqGgDeDpTrpUJW4Fh86Iwc+Qo4jp9ln/
dNgJUcxUlEZguYu3XwVKn2KeAbE1E+1Z5yTX9oAuvLak+fd0/NReUu7Ja7yEFP+3SBUUBFe8ojNK
R5RbDGZuBVxQsOyJu5hkdGNeAvFg6AnXnxV3CxZeo3NVp1l0ZDm7bNGvCOYwk8dPRv+xCNYyPGP9
FaiIXadQl5Vf1L1Ve0QbMrw8fHuRfzhogoZr6S8FvkhiNsPT7h4OFWnhqGS12wVTXP6T0WCRp+4J
shQX+KmLtJD619wbQmDZaFTd7FRDH5Xt81rHaAM28fBtX3l6X6xd8ZL1Y9/hGb0FMgjpXST9sOrW
3h189ij4bXHpWP1GEqKNFITfQbU5ryFTUrJjBUkCW2qY21azXJqLXqV2daZSNb6Bj+zNSFLlNinz
JBQzyUTVZvfng6I+KCy1qAqZB5tXCglvT6FC1aOr+7fkUi3SNm/0PJhRvnJySOFE7j4Jy7Lg6jxF
Xhs6PBmbcW63nwFRf9j8PhW4b0oSVfiyEaCgBtyoKKA8KigSWyP09hbnYuzKYrIig5LPGgg2zaJw
ezfd53qw/RKJUP76Jma211eAeBU/qRNTaaYWwECgkFkEM5j/5LRKUELYbJuMIzM9qJFEqFocd3ja
LyyPdlAciCtfeOGApjRPYn/qdhhbnyaHpDh/wzyu9O45+GjCyPw1mqNHpCKN/FYYLFlWQJYU1+0m
aG17OBHuzPSYe4xAZHL59hqV4qury0QNXfSn15MyCn85jQvJv8cTNZI85SymvbKNhotNMQOXEP9Z
ga2ZfmaXG59BLpeiFbafwvI4QSof1ERFqNHQVfOQ7DAa3MYaXn2e8ybqgwhSJQspblaCeA1TxrqP
2oL/1nSHXSDGVkDjN9XLjojlWBpHIeXdKFGIYk1vRD0Ap6y44wnS+vTdXDt5Y/FxLW8QEsyxtoQB
MeN0Ix7xD+Kfz69KfS+/W5S8XYZRSdrttq/zfwmb13Yid1gvgbGtRjoZFel5sgP6vYodT1XB1UBm
7YZaSGjYIa3ioiGgU3kvCbI1zQMd8AaY0/oSeHtBqQFJw2tPgcBXHx4YIogyZfnTc4flSl3TIQ90
NfjfFLv33NlGn0Xk/qZ6HjyVQ645/ZklH/CsJvbiYI5CnZeSr4ofEu2aDtQzrlbQR9Ho9t39bkeq
YbOuXQSVjt5B/teMoIfVIaeXtvaAujbrGwJm+McuFHtG+nIKe0x0Tny8Vj2MUHgwrONuOhiO63ae
jqO40Sui+QBweUovKDNwR76hVcE0Y1ofkO7UtohiaCud5MFI+BMnbp7v8EC4qk7kmXZVNfRzT7a+
A8MnheX2k/ySGVJzIk8qp+Ih13tO0ObI1lO/YYQ8r+LyKzlvN0BbqPo0ljzo5yyGE/wvO1HRll6b
8gy5VnxkQhSA2CesmSPPe4B7w9TNdcp4qOf62rMCc2hkYWHuI3Z4UfKtXBzL4pkiKbd6HvvWcOLq
/owD0zfHI9nfhW0ZywVKYLUxa0bln4dPhD0e7ZPqOot039ylDwHEws2k/tm9eZM8UHillhBoo+kW
PI+inVSssvofjO4xlVrb7O5c+87a3PxhyVT5OA3Xt0VhqtBwiJc/I80S/bjXhozeDyK6a498ZiYC
tvIduBXn8lS7/twt+gni+V0SXQ4DZYwIEAIzK1wsshEhNfucfZ4SCjgbCmG+8qOsLxAhPopttoxD
KdJxh/JBDfQbq+afSRQFTmMNDeSdWwJSQtRzOjFrN14zliHW44ygBTFO7E0p5J7xcedHJ7Jc685x
WmBxQQb+MInpw/mY/6eGZvpz6e+ZiwBmFdF3rK46hpj54zQK74brf6YdqvssJ19Y9lbSFdAtYhSG
ek58EnYAXQTkiO95OK/htCGm4nGXmvPhfAdKRaWzKRNy0oQq0X3K8efg9H+5Z0DUoxxGnTDM+xkC
67MFWbxn7ImrjBzvBX9r6WG/C13G2hec6iqey8fXhDh7sGTBi2EJS2i+psspDbDqtLeciK0GCVtB
9a7rMCASJmWNPZZmW0erkUqPTbqfF/AH5L4R6RX/hO33tY1/DoF5sW/apu6nguR7aX4fQcXaEDly
J1a3EeK1GmOLU8zETzFjbGseIwM1MuA1BPJW+fovpLTRoucf7LjERs7q1Ctxlk72jKwt0+Mjzbkw
AuDebenF0bmVXI5XPJ65pDHPg6NOHLsSK1RtGuMVeiOOqCmAcqvfUFWZ4Qn7TMCuJaVV4jDhckeu
RMGtAYLvnjfS/FgTFep0J0i3kUhxI6gvuSfDGdIAkCL1UeEOQ9PUD7rtCx4PGbTs+5eIBjiuPpQF
drn0zapMpmtAj0bSDX20cuIcQVEq7hoMm3Tl2AMTP0V3IuzlrVyyTHV7/xYeeRhQfKMZAdDXeAdN
6NHk+fMPqEYSm/KUmFj4YX4QQYQP2oYgkx7W1TXA0+IjxWNaUd4vw6NAllGbmEqy64RhCMT8xQaB
3R1KCGaKn9L7jFaCakSbVp4DbEMLg9FFRUrtJ0o+7MqpIw3kNIW7RVujYz75n2YwnRQ5MAOwPXFk
WWh38j8d804uHgUJqwWZbWsNOROlGhQSZgNjdQIsgUONkBaLrXLtVKVCwURBVzcO7wcD+QV5MORv
naIWG0mAE47xqqFAFXur+3RcILUDedZfU3vhyqTwm8XGJK0hPE7Mg8BZ7KC2cgHUCyreFCirSXUY
8m9gv9Mi11RhH+eeQ2O07VZlMiZ6z9jib/5LW6+6zl4TF6lxHOP2Z67ncwl3Hix6WL08iO/3snLb
02BM4dgpT3GK0uKrsK5Of/lC5mMs/B6sL/SvoUPVyF2cexjZCAqQK+fV+yoDPdTkY3igmB8Yskwh
1ASvHJA4ehVRyWYyHiCnQ8kzcJLQyraWnmhQXeUo5fBWr2Yh7EpifuR1G6JbYbRCVMPwCUHCvJNe
bEeL5sbiFViHev1aAnz1qjpexxGG0YZKzcjY8bdwM9GD83BQKk5Wv8SX1IajVF9hibUic7uXVcfu
zbUnOH2c0PTFs7W/KyFHM/Dblm9O84HS2ykIm8pKERyWaQtal/YBFCuN4Ym4FCcEkN7eXYdtTVGD
ZZvTaxgm0BBGnL8qNoQsf0rRjNCHZyr96VQzpDNGJXpbUMqf8zewxcfvq0gHvQ2xNDw1BJGjNaPP
s8t/50sDcbyy6bwz3yulJnjMAvHSJ5ZKMBPe3hbOsrBr+ex6Z9/bS5aAK9OTDpfACjohhuNOhHkn
3IYShK0fDqPgz4xdT8Rrh0UKON7ydp8UoynaIqqGRCjYchIXmNIF2OEg2I2ZesuII4pp40O6lgCP
5azC7UYBkKQXjYBg8azKouW7Q0cGxMXzaqgQheKnFmStGQ+62WIBW7IpS7oLwwFKjTZMLFqwfZIH
xI4rQMbHMwaghZs5fakCvtB0ItorePPPrhCtQhNccrEzdHVer6yR7gqlvC4rOTdDi2BlCR4w5WIt
nRYGcdkXANlnat8iu0CZZ74+JKr40H+6nXq2H0viRVhUtL1zJiIxsrA2lrvCAG7aP6HGvoCwsJhS
RW0O19I789SqZhPSIpg8cCxcGTr2qf3UaEgNEfxEwLWvD8Q3voRKkVBoVoz9Qg+5d+aiGlU/qaUr
ifTyjt0y5wWkdiunhngH2Y8ohSXWfQI4lbYg3QCiqo5JAvmW5ZztfyWHDTo8+erwZ4WslnvWd9oD
cAIVuRZD4qJ1T5XQdOnqDiXR+KvtUCyDcMGRC2TUuk34rVFbOk/LxXzSqpCqw8K7qxq+5TH3TCNb
LU2mzFsMkMY0BHue9+USBEciB7l33+1SlH0+uMxu7e41dQhlow2ieR8bXGco/oJXlq9R5d+SAzbw
2Qki9rJNQsB7M3O8qPMCNQ88wwtvu6DMuYDi0VlOo9ZRwlGG9mTwP5yzzxJPA8ouJ1kpydFyXXpx
ZR7Rdl1GfbEdysop9Tc07j+umnozdAYq736HHvQ7/1HRBGDvHz9NjFcDR9VyQ1R7VubaQPc13RiO
+17OIpRxLOdrHLTFvYpZ/0Of6rTXl0XBdUlF4WJT1rWqUALTUHKWVz3LnIDL+m91mz9RxRu3QhoZ
4FaXXFUW9zZ9WnoZfGnt/S7PymyaI6KOQIlheLdmt6gZrlmlfDa+O2KK09+lHHKJrA4L2wXBxlsG
bY1h85Ohbu6LThCbNEV9SGk2+bybNu0dLLKdxRjfJEyIwUcKg/ijlPPDbjrotHiAUzJMsJsfABTj
s/Lx9LPPd+giFq+GQIaB52o96hLM58QgZIN325P6D3oVV6t23lMhGFg3bViBBumPG2mXdGaPs3s1
XNe5frgcqGlCp1S0yLDlD6qGvpVIZ4ahCqw/dJTDarUn1G+kkAQex2PNIy9rlLGlJWETjZ4LGB8R
11CcsVO0Q5oC6OyS22zcQ9ZTIAK6t+lHxdo1f4iIWfhj6dO6QUq2mrZnGc5RvsSnux1dqA132LMR
1QFhpTIWEUSJqYsOvk8tCDVfqOsf3lCfJRT/A21T56ClbbgxlYGtLpIoYx89GWdhKV0y2bWTst+G
/oh+X7T83PeZB98NF4HCn67rB9EmVlg4lZAqylSz9Rd2owFuCEw0wHed2YiUZZCkkwXXab9s8f3r
QIJCozQouYCy3ihiVoiz+1f6+DK0VNrC01J9cvM0geFQSgq/20hETeiEwuYxM30S5KIz+7tBuwCR
bosM9aB/rMr0XiHkG93Se/lxmBrv9SsQ27z8NvnXtHAXpKAdeSKdhb72OUgkcLw+TYcExaZJregY
i3LXR2Ka3NYAox5798X3wX8aRxnW2LzaQMczfayWTzHObfFw21xMuxgd3sHJS1rTntYFjnemrv2e
5JWB/whr6dfEcNuywzMZEH8E66p0xP05XrnabD43T2Pyly2bjdbdIs+s68v8aEyOac5hE6pebjJ/
sZbcrNrCvDKDlii9GG45cIOM1AMq7mwF2EJ4QzefPnhhAJHI5r4vHBgCM2E7PEK8rAsXkmS423S1
be1MvwA9as5Vs+yV/AkxCBxBgNYkOqjVHbCr0V/zEG08wS5kJ4JxsnzzEtihPkKEtByTn8gDoQyx
VwYI2qtGO3LZJfxBP47+Bui2Q86s0lWxdVR60n86+QGnEKDpeBhNiT4mEsRk8USwyr8jX/f9uuF7
2NxpqtVG9zqVTfQXd8msM5KVfRZsGSv6RKynECQgH+txGkaBjeMYi0vu4/khAGgpD5/y3im1Ad1r
xKWR59L4N2OAlVQzS7U8YPGYVhug1rPKcHvrIfG7isme+f8+xM82/VQDsr8V8A5CIwz/NGOQMx51
bIoOErNlHHJE4OveN8uhqNKfv/U9SNI2UKVYnmJWiX8tamL0YNb0hJzb2oygA4luyT2cDL7JiaYH
oKubeXUtpjKT0ZgGz+NKUgAVvP9JY3+zqtdFOja0e94vYtviW7kg6niLzCYQG9GRoDTdWwezoPUS
XHygZfRNLXw1zcNCBLgqu5yvPLCmsZTN2kEGti74qOb5Bh7ZnWHIECHFDlyvEZ04+X7ut0oTLpS8
l4D8cKciokHU4QXNtM5KYR3rTwCAl9QE3eJd3t6i+TACmnzNt/uOAotehhBh8owShNo+zHGlMSIu
lWoikiE4sKIGOHsnufT6IDd8ZCS0vedZ4tHNOP8TvRp37jETcQZ0ZalIML2sG3imJnGdKafT3hDr
MjT9r82zztMiICj7nvaVgTyyMF/+rOIFECWp9sxCxjf3PonTMFTudUwfzQlk2eH2LFw4tw0mtAsm
ZP9usisltGU9LoUquDIAXmwv/C3rCD3F4IbULZZqfJZApyAv6qACiEc8UbqZEWbnw2fGBAidHY1l
UxhE55NwHUaVgNgaaPvILwvD04Bl7yFp4oE8OVcElRXV4rrwwB6f/AzgN7bIr9Vrt5lUEa0+llab
mwqAnHN6TuIVH0PFSwtWPPwxoUoTVFOMdfXCTmpLI8LKSilEJVArV7GuUgPcL896FhzYROirzOcx
4rrb0pcEQinjx8P68Qwkrgp3Qv3xGJB6+ajaCkoIH0g8ezRZD35MRmCbM3Zi6F2tFVty8cg5My8D
p8gKNwtEjF3gjnpFLf6cbhGaR7IdHB2udpF8Nl4YnuZoruYyIpPyHXEAyzVFvQCNkF0Lx3A8QgiH
+k2dv1U/fLoUj1WU83XGcwrecOz9MlIP5P0vPVtAa0R6q9JE28HmzbtdGO1fvty69vD64yHR7qIS
goQVHapFh1fz1sPyqbCvT8uABzerwLPgpRSJqxlz9AHDWznMdHBMsAwOQ5+VzzUTkrqFz0SfLjWB
ZiWnbawwLSR55fUwrBQY+TKvQPEuKaj6oVLnW6obJCNKErPa6NstjLkmQHeihyFHKp/Y7Pf6qKCh
+LoTb1ziqn5VL5QQeY6UtEqKm62WRy1suL5aE/d3jp04UkZs+jDRMHMnPajUzqDIznysuNtNKIBQ
S1xSm2baUMXZxU1iRuKjfLfr4Y549NgkZYgqTrTiXe+6Y5mUIIc9aRFM8511MlCl3tR+wSIKXvHp
5S3ZoOlMh/9hVHXH+SSqplNJq4woQhhuEe+4MTyGYOxNlMyjdtALfoL/NUiXazrftstnpVA4U+YV
bASv88PAsnHFV9Dl0YmqG9r7YSqxQT5aT7N/TvUIB8H9RYWJMXxDzD/+iKTF6uiBASnLEzvnAOiv
BTv8tKWpq4ck1kQqNFWx5GQL1P/NSy8bNIDLsem1N9658MB4NeAfaL+4mPE6usLLTtmkgAMYqZZU
Zv/kni3sSYp1GjluPlaQP/yJmNSDuzev0b/1CAnC7fOMSnSl338kaOxl5PgKeYw+FB0q5Q8KsdIi
HQ693j9Nf4UMxC1ncZN2gTdWzZICfLrthJDGu/uP7t/hX/ncr5+cVBsSX3Xtwvxey854XqdEhREW
8ETPrakP7y4HFrUdd3u/CX0NzqVP3DrTRu9QOxC5d810VjUDnQJM2G3I5Hee2hlU1gJzTRtrrSTE
QTWgzZ/A+Nk28isH414VmWnKBvIum1/IVcfcY25iYJnVkKQLHxT7TKcjNW7BQE/mOj/gjgR+NpFz
htqblahzfiGD7ZdlHR8ApTkjguDf2sT73xtrajQMjo9BgJTATSBGREkNkgy2N1zklfYheqpQAJjc
aGffcJbiYLE7SWq7BWTa5AhXUVh7p3qvpAGb1ie7sIK3IygHuq5dmIg1Uw1pXTeJyQgWS1LnkEb+
+czVCcyfleCgvUAL4SPmzXk3CdmU/bjCf/VzJngTfhlBocvgyjNk7SyUngsqXr6S+q//V9qYRGKx
fSkK8gmWnAXdsv7BoO0ZldYDdFu6FZEKnjMdCci/prPd/xsPCGWUjSUAiCKUNgKUJ+ditVT6I+NC
38qcSopbp+sviV/qp6nMaKBhrUAU6r3Px+YU4NG4FwMnA68mL9ZngRRqseLpcDyHpY1qWfH+IbTM
qgCIDwMdn59ZN+7gAGo17x0B//8y2E/kPiHuUkRxG7ZyO2gHwboZRapgmLYLIHr5W0FWXBfZOau0
tNELMiz/13mp1XcN7d4ILGzR5nceN8/RnhJMkEFen88ZzqmYn54lAPb79Lv34CebjuiObj7Hs0Jr
U0XZRKV8XRnEh2evKWqzzVsVv815zFaAQl/Ib35iLA8NfK+bEOVyclsebEJxF//3Cl5nH6VCyNzQ
VQ3naHc5ekowBOsJUdvbuoZgSVf8mV8aalW9jr7cz0IoB24qqkDya7CE+Kof7/NHd0Yq95BMFUHa
5ptIX6IIaT6lGkgA4wZx9UYycOHJDhVZZow0tTHxQZKAXh/rqrrNlx4c1bS5DLK60THcSG5g5qWk
/B7ScR3COkLpFM3BJDTuw9h3SzIx4K5fWH7ABfkj/TJfQl0WAHjkDwQyMdTh/dX6LkqBVwmFWyQI
+urYhU9n8eSK4zSAVV3eN353N58hW4Ep8H1KmDQgHmwEMjhpEGFsgwz+Fl+DSSNHqak2lynOnlmg
px/dusYux8pOlTFx6eksCG4LiyPYd31KG7YbL8daBySH/oJlRUwFkMhVvSql+qQDSHl+UXIHncsF
n1uIWyvezdnOP6W4kUPdt49SZfiI6M6kGsQMEACZKmzMm81yg8E72NFG4dovugeKndkVjpD1ZtsU
6voI7vhojaCnjexKpmmdb2PMbIZxXGK2Ce9XlqplshZwXeO+3IkOE59uNa7/juX7vA9tPO5kIxJJ
NuYPT2fqxB09qbRbEjjPLwtw8qtqNOBNrn7RMVqZ+oieLMnPnA/LrD2IyRR2v7i4DFiXsrVkPKKz
CfIa9m0VzVzNEiTs8/6GwGUogEUUleE4FAw9sjLM7/6QrGaqfYK19j5+BVxgkCpnIFcDK2DLPHjl
cqLvxy/Fyj++unBfSWSDyRp5lHRT0uA0XRc3FOEi+0NGshadlBxglqA+DODlIsWTu063G/3K7oww
giswPayCqAC7QoUS7nI7ZJthtIUccNEv4qrsuVnXfCLVIvtdI7b3+5EFnJfUvTDYfvUntuznhPPf
0y4aM9QuRNJWDCVceYxJh6p2mEOsztGBqDyxTfQBj2458R4Pf5qLecY6bcACncgRerxPrwy8YRm+
vEVBfLtnJVlAKcTOYt19Ut2/lvGB2LrBDKU482YVFSpd8ZYumxQ2Zt29vnGASm1xcCBlTonCNn/v
OIcgjl6y4xy0S7XNzFGkD0R9AU3zQF/iPzZLAm7iXWqg+cBrEyMw9Aqj9WrIicJ83j25so/YVS2Z
NTggLAAFiE29RBpnQGI6CnWNpWpy5vVnf4sZrQIe1pUiBK1YRC8WvPXGTb33NJgz9t6Y4ugBI6ca
cBTtqZVn1VEZ//ymPEhDK0z9vLPp1Qb5/zYQKOfdsTwjAo9Fe4AxqvhJaZ2/3QRjnZlpnKb4BdXu
ctOa0eUD9eSyz4H2RqBhlGmYIJsf3pUsGjUz2XJg0kmcxP1UH9Xm7mrQU0T0BumgxYyXgllsdb66
DinApp2lsh2SMQx/ZzZ0BbNYEKxzjSdLLGkEoQ+YXN8OQ+J2m6+Xv3KdHArVC1aTkeQhtyyTV8LD
GSbEQH2SEKNXb/choXGo4L2si8AMgAu+Krb50WkMjGqgP/WIfHW3U/J5z3BsBlfbIaIPMdzvcPXn
5Iylr4qov3gJy4lrHadNX3ExW8khbSgtJ0QOceSYlsumDXT0Ulxqrkt6M8W7lmt6k+a075/eqb3/
ED0sM69pPfErCAfEHBgThb+JaCTRYzJv5VFRDalGQYn8GVNdP6+ByuPidMumd6QxAKdWfiJ+bCet
35iWLoyWef10x7ozMlXYw2he+R3oQtBzfzObmGbLZ7Tj7LLR2TQyAQZh6u7UP/2tU/ATR2NL/YBU
J6+dCtXFNoeDDrSKc7cTTI9b7PJguru39nqk9udgzXKm2Vf7beG6JGD3ddadFnvTGQmg9XRGfBlf
H53j/YRHWlMoV0DX3bYVrFCULBI3WVwfS6w09K42x3TjB8T0GgZ9gNIHtvB3Ys4Xk6u5Q3bN93nb
8Ww9kJWSWyxor5yqt8vs+vFeya6Oq6U7BKIOO6FTLuIGW36tZ0PQ0Or2uK4QZZ+EDtt/A5uQhDvp
cma7PfyLbxkP8L4HxYroRLggz1bh350nFovwunTCvJNBnhjnsa6UO4tBw+Q3jZIVYJcLCJFrweJy
VyNdclzu/hQWmPqLjoCjY/cWkbL99CcQxdiO212xdC8lj0gn7gY5fk7dCjtxeNjGHyijhHrY/raJ
3bEkcg0dRnuxNFYxEHOUi91QNAiFCZMLaxYdo2dbH8MC6T9AfK849HWwbtUi0nSMiE+ozkk6tLzO
NQvifqvo2ja9OjgQvlCOUHmprPECo3LjvoOY7Z5VRZmP1KI49S7mGxx6e00WVc5Ny2U8YJ7BHVHY
96aa9ouPZDswxWjXQTKExD3PKdMlmiag1E6pWFCwlARro76UZPv/3QrRCz8qcBeW+/v3CSMWbqWX
LNURvmVBwgF2A99+RCzJ7rFw1uXEeJm8aI1Kft7DDG0Uam5cktwRM8Q3Y74OLR36c6fsnD6OpCcE
3og+TVGvHEfKVKCbn3kMhDNBj/S+agY8iE1r+NoZNoD+Uf5aaWraPWGZrzJPvMdvNer3XyZiX194
M0io761+ME3dmFZh/yAresb7uJcNXRxUFhBhUM41v/StiWUBX9w1no4Td7OwR6C5CynCgKRjzu9c
kPakyreW67dgEpjcZoLGJ4qHTsbkeT6m8tjKRwIlf6CZBASjHYtHjn8qn4sGgp8Zsfen7tKhwPwL
Mx2lFak7HcknHirnFWLzuEQgEw45XQt7tXbJM3gcek67qOdcJzCUOntBcAQZ0uDOCielOj8V3gp2
NkWd7rw6DqeA9b80Rwjrt3Zj6rg0PfiDmiMce7xt/oOGgBN3l/gDuGuHiWerbCmK5kk9IqebSgzJ
jJDdLKRCjfCliJxJW+PrLEWlGmm88pHrJjyEd0Vi3F6uofiutE8sdKUnGIkQqEeiCqPqiEqUqAxG
U9o7L49RMPr777RT1+iiVjuRmdMsrm3wiKumx3XQJlShOzLzK1ii+R6XTgBlkIEz3niFrRoteRYm
QOXKXEzbEaNAfVRedW20X1kcv7LNp0C8ZFiz8/Bx/sSmaFOLLPXlgGErzCkP7KNQsxJwIIyA3T10
Y2ZuHXe0X78HhkhwDZhbKIiNYw1vTP0PtIi8mCzAxJ8+rNhFV02q1zSyDzuTNoUG5OIlJMeKVevR
FMv5ZbWxUetyyPKBm1bZ1YmFY06Iv2dGSrkX/wElWXUElRmXtEAxaBIHyPf7I5V/a132OjXlAu95
XrYpECextW4f2Yp2Q5yKgNZP9hPzxt8/jB+Em6gieEGpEDKJoe9zrqo3SUJnnYQyO6k1ByngRFNN
palrbTAyAKDrCr4hL3In+aWaES088JPlsCQ7ZzJrlptCJrtgKDeINo9Optx8YdcIKYlTG3ULOPqY
i4ypCSfZq/upBs16pI5HxFIuuRBmUhzMaU0pYJCyp4IHMpZ+s5dSfXTIwyhyFa9ApkdaSVrm15Cy
lYdluxT6zP/sTGp1TorrKJyAFRlfDF8H89R/7Gga5bD18h74LkVNB0ArMLesd/UtJPWpNupdkQTj
iuXSPj+E6VxkcXiw1aAFujYNH8JiWCGvyC6ozMAHCiuYfz8CY1RcUgiO7RKUJGdhMxkVTQoPM1gl
YOBY1r/89P41ZsVsAeN5NPl8StHMtLUjXVow/G0buaE8t9uO1iBsIzvRTqy0SxDvdhy2v7sdIY2L
9/IE1PWZmMlVmubkcmxTlipky/ww+hFQG5+eggvvsIAS7pf3+2RSXhDClO4x50NDf2kViadSDJt8
GIATDBmMIvKgJW2ZAjNkYKFzTcakkil36UTimo5umna3l3HqAvbAZGkokY+yBJMersgSANhGA2m0
MJZSVMr/JNIxgEaKSfvlmYPWOJqA7qzoFtSg9issCJHwve00cBKkB0Oi4eWt8z/4f9naYKWJim0c
638XIsONYwPVQr8Xd8TMF2VfrCqe+/ml9fBKus2qYVVKc2KGXPjOb+bu+CecTXbIgH0D0K0klBIg
c7WRrF+y9Br+2lBDaGxt929m7xnVZK7/nb63au3NuuO3wQnvjig25ewpH8T8LodbVqkZNP127soC
yCb70TTizp+SeL7BCALtuKBFzyVDFZ+U/4i3iF7e+qsYO+K2JuvjGco8cpEUOQQqNGqJHv9q7N1G
mVOHMT0iiUPPa61AVWB3V+Gy9o7V8A+dJJkVFEwFKC9++5rpK1IRl1Vb6kC3y1fQfaoGI2/AKHLW
gFA9hJQbbYfJNt2G3zywhI/0JUKq76S1E5JjbKaoypFgchv+4+8zlNsGFJFaix0VQpUf1RQSmgdg
azccGjMTaMlStB5pJrZEWcUg3jkQcKQo8XgcIe3gYseav+Jl2FnEvjQ3fRrn9BcgGJjkAwZfzemn
3fYEqdFwJ01pbv4+aZfPMPQ4Npqif+QMkfIDJ/ETXrE+OA5ESCwD+bVkISV1zlOGeLFWqqk9QXVD
wWG5/dGoCtRsUaNhg2v4YIgpmQ10P8CVAEecrtxntvTfgB+E2GiytBW8giWHn6ZwIxkKJqCCwNJt
5WTXZlZ62e3iEf7gmzEY4WKrTqO3IsZZfK3OqhPs0KnGaYQmo4Atu+J2+DLY667mWpbYrzO5ZOlj
m70AaDyIvW0LUIQxeZXKO7uZUjv+gJ+hvQ5vQNDLAXBAlra0WfjKHa+6/MUavqlof8s7IauQkuMF
5rgspUTjYvOdh4aG6pN8dKV5NWNzUg8RNfRiIcLEn5ImpI7f7mEaRjteESNtjphv3jJ8op70QLUd
qz33Rp8R0pPzsMCeLww6Lq4qba47oQDSBU+9j75cdG0n1PUICuM4sHn7rPUKoNCYZJwKKIf88zuc
Ta9OuIB4yz2mm8KfU4ZKpEIcXJyIRUBL5dyTt1VX7pjlJ1vgxcusaJocX7SVoBqQOtpsuIunOLpA
bn+QnPGwD9oQGciDFR5Wtw4aLgTEPT4LLKBAxOwANSu6bd2OQgCoq59vysjnydOAV/cl9pXk5use
NurbBejgnLFS0i9eRX+7CEERdpA0luNSCpa4CgJl14/JHY/EDcxHUzWDxLk/y1uVUMSga+gXRka0
VzEo0UDnhM/yFK3CQTzXLCwVOJKI6+AfUQ96ZY2WiwA4Z2SVN5hHZX7LPu15JQJBcBxaNkwprUNh
a/n5fqUtqYS6wWuTC4VDcciJ2l50tjQhMmfEm0B3gTriT9SbZkzzgkPztodLpXyeL3og3lk6/PN1
43/EUHyMQ0gEVfReRKahvg64uMuDn3mmrSTwKd1zzgkh3eGoLGjQpJLdm+SBhWxxNchskW9V+nql
RNAhTyBSkoq4XUnn9FN2Z8H6/jyRzyJbxmYxi4UW52Nmjppxn6dUUiFLMyXyPfWTY5oquH7iPKni
a6Db/1P4zPxTNrY2LqsJDcjrjDPeBekdqj9BKDVKqQN5KN4U+YJFZNaSqq3Cs2GVMJmavd52k1f/
4GxYnqw5M8ePKc3u9mjYOpCbBEU2WoYCf2aw8u5Ez2J7A9haXkat8Dn1lQtefesu7Qq0tuQC6r4R
0ZE5DYY+ZCXuORrTrPon0EPfW74ZHoS43UW0rjcX0c6WcWLKyj1b3Yg0NZMex+SIlRF7DRkDJ90O
8icoqw28nmDeCDU1K+eTzJFkojSXH9H8yotBTymatPjXiFlYixsiUzBgFkKTd3Pr/Zyv2/HboL8D
BsDzQy+JAIx2ZCnjiwYyFwZ8mjRkFZLfHJb7G+QDY5BTxeRqD+iXGssiJCcg8Dq1Zmd7E+pDcsUx
BwRmnUFH7+5I2pGuLyZgImRa+DEGRduwCrny3pnyX2KCQhKXk4o2tac5zAlyOI5ChZAlYJOJ7iB8
ULDfT8qY7rcglUgAmMfv1+N3U+NczGIyeYkYtlNTR1oFf//pq/03znSHYwBSxnray8e5WrllHtPR
r7df5oQJlFBnSWxgzkxK3m4TCx/FgNm1TfZrmJmYIp6CzkMkTRgA0/914ep3vkb8512sOfbtCE4T
pvI41kow7fr/LcD/2Eo3a8DtQXcdQHbG8dZOQTQLY+JqqdMv8nn+LcRXpMfe/V3QQ9uYKooj18r6
8jT1+DMQi4StdryJ5qlilRX4Y7U0PpGlgJAKEdGTwwA1+sXewlTx9ICaYHc0Ds82T8yPin0wOKDD
50QtwQOHNi+7j+dXzjaQCB7DzQnvNXK80siVI1JVT3enhJfqMGtQ4g7ihIQ4UtENTp80ogsnQVu+
HsLb7/O86zYe0BPQH1m5Uw0ZwgzdvzDxBo6zu8VLBSQA92isMUTtBomwucsDoncsfrJYnYGaFYm7
7a+MbeCZ2e3jpaoeIMXhpb24OVURgPJO2IXICthgIdWMD0GAr1RUNucQxgTWoX6s2yddzMnudFo0
vLO4R4uuvtZNtaGBu+/93PwEPybchSXnilUF4IQwTVQv4pzXvKpyq2uEcFNUOLeu15229PQ71s5J
yo1VVoDpl0ECiP/sMduuqG98cWVIoMxqJg6ZKy4+ELZnA3lZo48UUUxE88Gfy7CY6488EgvuBrba
upKueN3riInvySkh8Ae1/nyDxx0YAvuHuqZkp0oXbU4jf83w9LIxLYmaBfkk5yEfRDjZ4o1W/JSp
MyS2zdFPd39CKjwwaSMSXAZGgVzKKpStqR2hCHof95AHE7MEYtj1RS+Apeb2GfmhxVooZzVxd70C
FgcMzLBFKA84sDUsN4oynDslouf/INs/wzeFJC8BlyJGfsSmOKHWOtTQGlh43CNA322KENK1hStx
iGbUiFNkiE3MiJdOT/e9SgMijJrvI+lpWFHCKcU+QhrOJcUHZvdomjlbyHsNe6pkUOFnCrrxjzgJ
naMC6Hv0vNDXfDS7ji3m0GoZGbFpJDlO/YUcOhfwxmAvxlaaTCKoRghPPB3RR8sG8VNdwvGpdtrA
UytFz5UVMBID3Lj2Q+CQgR23WMN5GV6x0jrPvyDQ0e+HOZDnnPHG+VGVDEvzkYx2aC6rmbZzWBSw
iq+he8dtlWI9zmmfA94GzB20FdEAQqpD5p994WrlzB4dBkZ/Izyjugtb3x2JdqAq5tRXe3iP2qdX
8h9t6sL2nadrZa0aYDBsWjAbqSDSAvPfVfYyfHwj70Gd+qxCOx0JOiip3tCfMKS7zVHT4Av9CSei
EsvkluuXA/e4H5I3sFBsRNokwbDouCvHKRv0pgcg40eGp5KJCTZGyofuqPdgVJJu8ObtYVgGdrkX
as5QW/VuV/HHrk37OC4RaDnGQkz0EcK+T6G+xiUDxFE/deX3Ge5Nnac+b/9pSjWEUU0GCHQS5Wnn
/ZKCLPJoDKP3wu+ZXqKEssQLgNypN95R9EaDojd+wLNfiSUyyTiBCwLgIAzAM2BamTUNM3ZZbQmR
kJLt49Srb17M2WR77NO9No7eoOJWs6bErt67TF7iiIWDwL/FwafJEHzZtfXwcf9DbsfQ7BeRDD//
gO4cEtph8PZO9ggheJhZUV3+E8yA4oN08ABnC0r80f2K1V6ca8qlsR8qyOMAi7ONezMT6B4QdhT3
UtitggK9TqwtHBCiv+s7X6J8t9iXV58+kj0JhTJFqFl1S/9l1joo0+Rl3zuC7DBnr7X6e70UONaf
KtAEthFsoo6aIDLhZHc5+CT3/RlutBz77TGbzjuoS7GFYQkKWkadvPK+YgPvfgn4kUS0/D2ut03S
/UeSeXYA7hbG6HiGhTRQPBlpY1wPpBG4qFzgk7z1Vic6JxiZwljSyN43YPMdpWIJrmcY7/3sTcRj
wmp3lPtBXMYhOXM/f8aRa6e2W7rpZSCZVoYIHnuDi/NAsbbOoJYsbOUSszTagSzCoA9ySAIPQ3SX
DVajES/6i9CpoTJ+7ldfvKIzDWn4NpFTKITgcIWoE1s2DHmUVnTS9IyNpqiZCAYksmdDCJwZU86n
K+lseKb/ULzw/FHt01ymvvvzV43e6GbQbsCi+6ZEJ4jEHP35jOzy5UIf2P3Rm1tQqmrbhiJjVqYC
oJ/mYlliRW9hQjfvYyVteQNqQUlu46RZBmO5EAhMNmVmDaUTL2Hys0wzlgaPvd3IJAqJgeiS2xfh
piMxBalKFrthXkrCTOOoOCsRsjPfMCBjTFu+1aWNhXfzpE1fz/RlcgR+gNGfkR6mC56v1FVnb7Yt
Lwh/V/AT1ISuRP0Fgxv2p6oTwOyIsBtmppTt5PbyRzDSetA0ZJVPWF1PUVgYZez3H9bTgNZK+9DZ
aXZtBlbpW5kLf5cpEoUYsMzewqp1h7aTHINkZMU6s0SayFcbw2g6V1GSwDOrZNzoZi4yhzo6jMCD
3HXpeZgyxBlj9ccEVJYU/aNFVZfMoXV/wiU5L/U4fG3Js4WT/yvqzSaJVsIipZ6MQ01Vq5ZFQFrO
SkW0m6OmZkpyqSE7SixOL0nTGSNMOshF5bDwoz8dLsJZeqtbGrHIJ3Dx9vA18h1GueKHEejbARUc
veAXCY3/IHGC09Y5ioMZjWdoaaKJ8mKIkfBpyTyT1lRMB2X2CPyDwZUcJEtlkw/kX5Y+ujTQeIIS
TUnHUHkkfT+zk3pJ5Qh/0asLFd9CqoXgdvYkxcH35hdHCxinknRikO0DSeXeyOszyiku7APN6wSy
q8OlgD7yue0gBPIxTEa0Wn+3Vc/4O+8/K9aQiG+CZTUEZOV7+6Eduw1zkvVxb6SJbj8kh8yTag7z
w1usUfgdEBTcW+0IxAVQsD75szFf+iC6y2GSMX1rZ5KsWt85KNBnHkHT6JcnJvxc9cw9rLR17nSH
1AYL2moWKFQ4oRdxXqKHxuZ0znSYeNCXyATV1FcMQpjq84XTokNoaooxqEk+LVgHz9gqtwHIRbXE
0w6iWKMz1nTYw4qUsoOLXQZtp17G0wWpWQdh6HgJvHzsSuZXOX4krH0K83Oa7MkVQWBN+AXWgcSi
a1qNdFutLsn3AE7nK++UgxeZ0rhoC9EaV35nhsdbKXzloEIWsrBSDNewGL3AAY5ylAL1f8ISvie+
D+MDb/M8egm4GhHzfEjzoTcOiI89Otd31jjnIJGFTHMzT8rV/WhV4twnyEiMpULgSmWAp1E80QcT
1G2nX+ACNYUvzstHD/zLBHOAKIVBQVHSn13BfTOhuFPEzwFAZzrmk2eROn7ndUqz31N3fvqZVxMT
0FA1FYt3L+psohpeYWXi7N22bbTlW/yCkdCz+W9W32KSKjAo0ZA2jI2dulKgn57DXNkDNHsB8qZZ
vX54UTCn+wToEBmXcKV4IR3xJsnqLCSRYqx0bKmduH2rO4nGmKYxBiUvw3xObV4OorvcWqgAXwTk
+YBApPvuTJdXB7rm6zi8ROdf3CsQ8pW97x9dnb18TuHOTNufjmSed1dPUEaG5UgzbIbwzPGm601A
FNmruBA0ow5DGSGmkErL3oW4P2BsMUhvdBDv4prOwd/HqDrAfGigU1srXryPWbZsebYXE+2UziwR
iBJx1dsIF2vp4o641TDoQ1XIkTKUNtQJVbfYNEweR3CSw8mpoFfETMFqMAXgDEV2F9zkv9pnfnmX
34y1nF9598wjC79eYr7zJJ2hhqGk7vjG3n5jauaKI6c9t0jjYic3fW94xBBzExNLl7XyYO8ONAS2
qLGbub6fMXweJJXQ5/NoRJzPpb7mapXvPlbMBSlY813tAbmT/OzhsLii4KgtWBsQGO1B3uLdgcG8
DSBv0rt+ZNaFvoRfW+Hu4hTVPtN15EVvCoY+QfEJJ6HmqTqMEdJfwCqQ8flV15nCH2GzhvXel1jL
gbiJrSjcaBap74e0KoCQuZAJH/mX/yxJzjSaKhcuqnARbrQdr8OwxJyTtkZ4STzj9BzZeCC2ePI9
ysgtQhsexIP3Ki1JDsbOqj24KR6v0j2HQRIpAgRBmtqkwzYJBZ9dnJCSLzGRM4BUdXYtbnzTmbOj
+pk273+QArhIJ8di9dJb9WoTX0i5yHx4rZV822HHfqdDaNzhJQTh8cIoVCDRE4kHEmRtKgdnFVbK
P/Yc5VyxjmxRUgHMZKnyEH+jBcki1ihHHbYGja/GtGwkHE3N8Ngba+6M02uu5Yw5nfXLkv5QkjjF
V+8d7dy5AIWLwIn9lBOlJcpBXcYGDzu6gtuR2eBanOaUED1yRXtwKRINR/GXDirLNIZ9I3QtuVnj
EWoze9BekoTSUmvQAf9nz4xF6APxRCrLtpxa16FnVJt4hnkEUKDhXwf5QHp+Py8p9LDnxukWPz++
dZU8MoTjJY1KIxPdQuA813Kgfei/esKOzYLfIBuzIOV24TLf+4cR32Z4AMOLmTS1SU0TLHenTzYs
Aa1+1enac6IeFm/sM4OybD/dIJFGK7kzzRlp8CB00f29qPI9wmTQLJgxjz9gbzjvgow62+684+dJ
c+xjaSSQAhVLvuGMCCZG0IF3bJ7lQzQ2XFNdy8tE57ZnAZHeLZNRoIjpwunqnTiRBU51HJZkkq7a
V+hL29QHkg5lxFwUEA2yUV7nqrxQRExQSJpfMWwfa3unSw/jKw2XThDbaQ1W2vWxNkr+8lhZ1iqG
DPUgWlxlWnZ8UMBFs4bTJNlecqiv2V4lR68ex0DQpHkjIePtOtj8C+o2agdYl3tuXM1CPDe3gxyG
eSDH4HlvyU2jbhJy4B27EvvIJu1q5Gz+TIc+gb9O69XPJp7I+mYDRhCd19rPw7TyLadlLEHxKJzK
pQo/iQjgs2HC6ofbr3zRB8SA1FJgyo8di//C00MEJTaSp9l+3kATli7Ububxc6mEHihMpf5eCnAP
NnYT8frGY/mZ3Bq+lEtQ2b7vIMRjj4o0QC+wMCeVA2U9/KCOIpxkMXBbQpv4jKwNz4tVKoeDa3M/
HIJUC5M+JHb0oIw1ObeeQY8vvxPcCMWviNL6a3VICLWHZFtLDuIylHot7GuSYH2qM79kfrT4x3Mt
272/XhBGheiuyXN/bT6SFfDq+430kflNRcPmTFSJRcpN348k2PCUHbxRe/OSOS/pLso1QODmddZr
unaFTVh6zqJMduzhuzIhRY54wOXtHEStJIfrv/Lj/eXBhstsQJiI/98+PAiTOeL62bi2wbWJwgMY
RDrIIVzM9G2d1KGAZOeu5nqpmCpOTbzNup6QoQ+h8gyN9YRH4OcljjOm2ENQXPk7w+OD89Tq2kGz
l1ZWG0hhIeYCtWZcnhOUuNXliK0bFI806OeAB0ILjl6xydqeLYWEyLgQMwHqPj0xTzQk66WsNoHm
0qyGs7js713j/dueObkmuhU4/0KoZU1mEIa4ftBTEfQATaa0cNAXfJtsiSTZNuu6lygNeZOyNqmD
9XqM43suPEYCUR21HJxEsJdm7Mu3K5QGeIPI6rRYRoB32yuXIBUoMvpF6nbJOujr9mfIpFYQjJNC
BUIUinpBGPFxj4pvF94k7FUeTvAcwiIoXV9h/4p0qSLVFspA6F18/dXCuBqx+ZbKlXC2QzI5sKzu
DdH8cmkIjc0oLMPavNKiaHweQAjW71QhuAXo9Tx1TdpTdXsY+HHBmavWtVsWnDvP5fKMuWWKtSB0
WD5va86zRRrYHpYsGjCc0UNdquxEOaCJdO5AAdVeRjcBkv/8xPBG7QGiU7oAlNC9UXHRsxVXgAfW
k0OFvxpAVRjeoJMtnVY89xKNVSB2eOlFNuslRRwk1sm6ypwgYUgEuRvOYF1+4/zphg51zdN265nn
pGsRgPfhTWRizo15R2kIh6WBiF6toZWaKqPRY9z23l7GKGhaH0GIC0lJ2FGUU1tNUCvZR7QO2z+H
bK2d8tZA5SPH7uLqwc+raTu1R9odLcDHiBVuza4wJGLOTuATRQm/q8GJh4YjL4OFSEH2mHd0H/ku
x+I1VG79egwD/QySTyRzxb97HMJE31lRJppjv4lcHUwmN3DAWZofEJWmNlvKp5I7ICINHAgIMfVA
5i9C6WZrYuTKzzZuTdox/tbbB3vM8wv5nyYtnXFvn49i319d7dQdLWlXB/7YO4ugnxnblESfHbYm
wzAEDN5KDHoN4uF6g5MN5145FRpLydXRleXNSCvoBL1trJsVHbhgSN4h5Nl0QVGvg42crPPH03iq
BhEF+Oqwm/igTLgxWqbLAs/mLnYKZtnbHvH9k4DI1ee1O6sw7MMqiCiTC+u1NA6X9qXPLYg+L6Nx
Xj6Iz6zgQr5GPovMaEuHxLDt39YV+3YPdwO0rTUvwOKnKJmD/4SYiWXtBxdtsorVtupaQoZnscIp
pDYLEKYo0Rt6189hrzhukyOp+bBBzOFfx7m8KM8HoGH5KpkUqFydX9JLLM9SOwPul4Hx39Q87pRe
cyZ3CuhrQ8JjSA0jlPq0Iktcyi0EaLms0ZwtCs1zrzWnfU1MphmPa8ZvXgGlyGxjWByhauD8e4/b
2A2pC6McRuQYPuZaqiQrWxnEIgEV6dKXljDlV+wtC1crIHQu+V4GkM3nXKE2m7lC272JT6u1vDex
omiEgY5HZoDVNi5mZl1nFKKiTNhiXNKsqCZGnEuF0GuraJ1J1irv42tLDyHaaEt9zZ6nwO3AvnP0
h7CzGWc1OflLqhCSE++zrTNpTx1vLvCDSGNzXRzVGbsXuG4Woj8xmfGFd7Np2pOGV008c1fr9rM7
Of5PWXTHSOa+O353z+ORwWhmxr/tqLym0kHiMkJ1R2PZm8kJ8Rq9DM6b/PsTfH8S4WwSOAPYzJrI
DjnhC4ARkqvSNhcgiRneU+eVhUgtH9WIWwEq1v9TBLcCF7WrB5shEBnp3Lh7/GQpjDJg0nU6kXh6
jMH9IVJAFYm9ogEfQfUuQXWO+uyPYfab4+MBQtOSjQMyUhg9Kz9YUWMAjXbBX2m4YbxssgS8hJah
mDLOmvzqaU+fAdl9NCGnPsYcuORcBtrtyudc7KtR6JARfY74BTV92lSjg3h5QyVx1dFP1V5WdJLv
pN5I6v+VCRgeWBJugBYYF+k0vYhjLjIVRB6yR+uP1vFVZ2ELQZAw4wEml56jaQq08OtlcLONoTJS
T0jfTRGrLvP7c+PgL6cn23NCHuiWBRpoLRLFoeMVDG/y9bQ28aZgBsxS+FyzDXCrrD5gsEabiKJa
2i7TI1jqtZVejW4rVJ645umbb5S/R2t0Ze08Lqi4K/95qv7FFlcxzNEDcpOhyXE8Xsi25kPEO0PM
czsQLIqp9Zsr5JT/jpsehkmqE6IbTd2XXzXuJAGTPe3psVvA0yYRv/ztXbNI2fp8rlIAc5uk5WXL
4+RJLgqINZM/omzyZU2FrO0zPHqbJQBsgIs5ZBDx7O5ei6MNSMdlbns4faO46ZylBdJjWC27LOSM
kBg0D0rKo7KdE5/0Vn31bxVkm+revjMHoN0yQx1szSjpQIEh25cKob59wK2UwVPxQ4Y4Y1851b8F
+qy422fp8zxR0O9WrkXOtqgCOmereiJAujvvxJnDJ8eEeKBm5KjjGOFLuq8xvV/Di1iRnCB47g1n
2LgrD3uUP/6Cum0gPWYIK3oTJfVpfyp6L+ECDm5CFrMCWETLCrixVuQF62/RZWEKOd0acUN+pkD0
bsbSzTT69KrD2Rz2Qr1mFMyH+VNlKEuRSHC1Qs5wHXMwsKEMJWWKA3Zr9xJ58DQvWu9EhrT8NOtP
nroA7w4PbR0WGN9eS+qDOP/OiwxZKFuQdCyun4JF5nLP4Y//4ZLFMsZ22XKamv6WBOWvZ7hemBV8
ZiIG9BGgFD3pHwlBmyPCjBeg0Z6Tko3Uil3Ldg/n0zZKKybh91fxtaziFmIA025vln93by0pqy/1
H5mn7OM3CaJg8PNReZiKs+CNOjGIWA2V8WY0BWGxjNLYLaWw8kIXY2i99ZV5/OyE9mhGvrwdNi4T
PnL27yJMWYv2jrGGcRlKt43sKSXNmWWdSwaOhaqCJBpX4bz3fBoEyoKax8bqX9+GF4cuCBf7EE7Q
woK9RHHrPP8wYho5zO+RV3t/uECcX3Vaj2RVJGR8/oCuNPxFcBL7B0iRVMlIGSBaz1Wdn/JQeuWL
x50mNSwMtm44GUHV5tYuHqgs/+mKuher6s1Lg7TAdtOPwMQRWvVkPZ0i2akDucPNn3YllOocMzsa
BPiXsq6HBDVSAGvid7i0bZMrVPOMgEyRyalZZ2rjik0A0owGwgi+DZNmSJuvrIDmbNI4A4SV/upD
LnU2HMpPEn5BVG6lE2SWjLLZxTm0MxHdxrcZJDMTAUKns7glMepgPE6qA6L/QVKACnlFhKe4REjw
fpAwYolSIYQkdG5ATW93+iVo3k8F1k+j3S3j2yQdnTt1ZZSquxDWYIgNQ5iG83/PcPthaMhrXGjx
Pee1eTrjNjmPZxZqb7XrZroFxNwMNE1Tv7gMa3CqYAxQBuU+dW57ZViCw5QLumNtYmFnoYrpZVTg
XSh3DJvVYQk01mcxqQNO1KrezwXdz3NStxgoLd/jJmwuzWqxT1nk0P/iqzj+8dn8fOtG9/ulDhGp
Wn9/p1Cbl8qjUNkbWPVrfE0LY4AMQaTSk/ZVssMfd1UyVVjPMdgF7MohY7Pyg5L/uJH6+TBEMNRG
XKkuI3qaBFjfTlolFF2QZoDdl80JacVlwPpfHbde/uzgF0fZRqUB9zJfmTXe++wSEmwFnCNIRk15
dINdjGyS5hayfeMtK3T5w2LiZaWLxdX3Iw5+fXupAJkM5lx6RBnoCLa/Hfah6LlxbZblxqNsntXT
3oF6z3sdbLAy+d6cHKWnF01hsLxAHlm90hwHa4RmZ4OjYoso+4VyKoOHMyjIB+CWxuWx4kAU2r+r
rXRijOSZM8Iy9vltJh0R/YqqKWSNCsvYNB1HmFHb5NnulMMP+7q2Nqo2KBY7/SSPoKRJ69x93/Ad
PLNMLMMI1OkeytwtxG2baWcEelccudOGMJ8Z1+j9SbVfbUgSbYjBSr1wl2IeMa8aSNDffBXM3WAq
GZE8ewvk5uJg0+GCtADeKwFEvt75haPcjeeiVAFhW9h6xRuN4z4LOGG3f9PDiflKf0Kj7qdrCP3/
pU4tRtdvQwgYgTLFUI532Tk6COBSrQsZzBr9aP//uKcuzttu8tuxKGDPyD+cucKzUm6EGXCpNntL
x5OqpglbES5JZr8+Di0YwpcLf5CM5uYmnmPfCp8OfmM6J2UcRUoD8I3DNk6lUuhIuKK6EzaK/Fs+
njOcL26SLVkYy57I73Q3TeEDu/IEMrSJLinSpc1zLnu7EsDeRGc1ecm/Fc1rQi1yciEGSugUA9yX
z3gRCOFXR98dznP8NS6Cp5q5olqj0Ha1AWUN8l1wnyjd/A0bgXk7qkNB2JuInG9qMSDpW7wflbc3
RDuURH4MUgb5AsEyTZszPTCsMnbTy3eMDV/Gk94mlLlqBdKWGhqCF+H7+XgPW4uNkYg3ub0PWE/M
7VWHoviqVVBFocgj6OYq5yghZYYB+UB0on9jYMlVthNFTH5BEEfqCq8vtMkKk/tdiI2EiikkWk0Z
CYWEEhwSOD3XnrPIO8v5+tWQ4qkS/hqfHZAMeLNNYNVxaKy3lvaS/AS6hT/DSbQC0U3reC3D1egd
Wf6X/GyakRvAKWCeKoJljaiGrbkk/P/ZaeKCwMf5vBC4i+mDHTEDE8RLefX2qpZPkPK0t3aqN8Cm
hbpJpRXraC+myPJxSAdaWlae31gID7FHSQ4M+aJD9tQ2ZBThChbe050QFeDnNUxxS+1q/seeER92
C8cjJ3jdqDQwrV0WGqo2uwMsgKAg5fAgV6Q4k/c3NyXn2CZmzrd9/WTSNHK6okdj82k/MQ4yzp0t
nKFQaQIs/JEvWNWuq60+P9vFgUJ+NC0NAqsV1x26iiSQ9R+7XxLmwtaQg0m+FGB6cOjxfa/c1ccH
awiHIQqzxFK1FUNqzaBlxiP9t3MG/5G7HvydzLKEBnGeKh2yEKIVuSVgCGmBQ14UkRBXaVaUDU6u
BKemabatnov2j6omZoM6lfQ73bdn003zFm1jGAKRBg/pVMlPLGi0JgZXM8ggwVF80eAU3yWydWgw
6yisJWHf69ck4QmK1uT6Xep8PHJtWlczFdBWKvdlPjpBZZHdJa8myiR6+qurfj49PGUZLPzdMeBi
vcfBVqo8YLIPRBUfSLo/iI4gLQ/ZQjKZetp4pzAh5928IoHtLU80WksBBETxw5hMfBtDWp2yHtM+
YVopb1oTSyxKOiWrqu8F6b8aYiv2INQSIMKfohRp2277fSsXdKiWkXGUlS3oKjaGhfRN8BeVzfTI
IvHIczu7T46WZk8p913cIaYH0kK3ABOrW7uallA3tpqcGh7euPDWg8WbXoevRDGr19+IXCbyThbo
uS70Ndt3uVNO+MAFASoZ2tgQhSOQQLcfIpybb9KY9dH0IP+sDEDQ2IcUrYQUwGxoDScvsXGqE4qw
1pnnUOSi5hFe0QtujSA2shzAL2zElAIVD9TdkO7ASthbp5K7/byF/p5YwAO0fV4hU3jCelJn201A
CNCH/OrVnOCC8L4C32LQbb26VfNOhMlDO5D6ttnLcDOVhCegfbN5Wwqy6F1yn9fYKYfnGpn+SO9S
mEL/0gDkOnbhT+q2g5yxKBtMMrQ/6sr65qwpZuUWOX0Lg/CUBBgNx4daERi2o1KPUVMVvnPuVsPj
yW4MdNacwxklegj10b49+4hI17oi3M2vkgXMUzyE4Vd0uyl6oiKHkGUpGwCYBivgFasVxfDslhde
9Sm1eB6tacqkeI9ZQ5sQj3j4zw9/87OWY3x4BXuwp304QwulRPwJ7VBqZV8GWQDYmQ1AQmu2V6b1
9tbkV0ayvt8s3lKEUxnSRtsIMgqE6UGYS3MJ/4ay9xOtVX4I9yFBXNDWMBrqdpRKpmca6KV3ihkC
GEMkp3felIxqN/EgldvV09sOupvGXH0pAX5KYcQQEZkYTxBYCthExLM27/DDA4lQ+9J5/KdQaYt2
i9toKipcG4STQf6B26ygpCognD4bR64///VBoqb2CCuu62kAN0FWom/Ne2ep7C+oD6SOM8WIEkyk
PUXUg1ZC589PSgIUwJz+5dxCbzV5cdxgXNoCJ9Wofm2aj6kpu377YEC2qbgdxFvEUgScbAi/R8h4
b1JpeKbbA/4LCDdRWZJ225prpFBl49MbQfubihXnXoGsbafDwtx+nNpHqFr/8Nr75+YIioG+1Tjd
nffsWVGGH7fRpeuZjhnZktPJrpvoLEK4hUPpsU1iq53EQ2M7YP4cEmJZC8NqI6aDAYm2XGgS9zja
Jl057zXCNMq0BWMJF6+nD9I9yUaGeui6xnjqr9O4eUcX5jn48IEkwXhSjdMHNNubBO7onTAQT4kV
1KtVH41PbYPOUJW5TlfZk8bCFu6GnSqwGfoHJuTGhzEVjT+cNKmwT5cxYERayOaC1mOqTbUsXfgp
fmURf7s1ugNOnxPu1YYRw9olywF0JOASMAYyDmIl+Y5dgCStD4bAS33Cdzv4lCekDJo2yOBB7fDa
cW6GQ0GovGbCtn3GiKmddhhDVA6QMXuXCP1e+gbr1Fl1Vh00zgVVOTsIN/haao3NqNweW1K8PQCn
YAebYq3kESejMe2X+sRHIOK7vaipTkQVetvI9sNZQFaPSG67/lsWoPx7oqCNg/W1XPFz3LMltfaN
hVXnYRPkRV5tNN0Ivji0db+mZ3/Hc9Jo+zwRqmX3l7mksjF8BWrhDMZ8P+Q5pnuGY8e3/CoLcM7u
4H7WThM3evITMjDT5d8PAxoiuBMYgHhoF5/y0Jr5lY0BW8gg5Tlk10sDvpOfobW1oNP5kLFc4W/P
3bmy2QIZOHrQ1Fws5GgOh+mO2Gyn7xjyVOTnIQoqBE3JSOWQEDYKcj2PpD6ZSrI7zIXqXrYYNFda
EOqeg9FjSYFukDB5fEvAohwfnX8A0WMn90Uu7P93138icWz0JkR0sIGhT0NbuDmiTNmhT6u9MiMe
qzMux18K5zR79HSpHt7qSPCE13b2TcIAJuI+4Dj9/RmTcyne2f8oe05sdAShWArAMsqNlTzAgmJI
gMi6x4NS+quYERM+WSlhPmH+A02GxOUGdPxPd0mJ2DImmYnLe8aEQ3i+sm7oJ/cbnvD0L/NVv0RP
9U7fdKG8+d43UbLF5lH4FvsuLqbI8mlWXayZIfDxLvtgxciIiFGcWx8P339vr0VTS3Z5iGCP7nWs
aje54F3zfDgsTwHgYdubhguZTZ2iBCVEmTU7YN9K5d6UCPctpaRvtdEzg/yL0hBxMT4nu14onEha
Ks5Qp07A/3dB2fvU7RdSB0f6AmiFhCA6PCD6sac5jYCblsxVh6sdv/N5pKPmVhemTjHgv0tdOorY
11a930jkCZ/V/HdewrsXCrksynDac33mK1Lp17HTT8lZ0iawMAHaRg34OtGRSs3moNuNI1ihq8UO
KF9I4du7NuJX+PzLAr6lJo2P7OT8ONG0xhtbo6O3Bt2JafWaJKjcQiRHxdei0kTGc4tTA1t2iRdp
B1ZBPNSVyBC06MOkV8j539qejN3gJiX+Shu2Rfeptt3qtMtwxr7520Znrzev3+GcSLvgGTf4XZH+
XOTUUP1LNZBVeP6AX+IXXvwIVhowY4vuyo9d4NeRUptkHjVb8zLvW9vHYVyzXeouzDgIGrQAUT1l
EyORE0sWlLjqK6jAUq+685Rvf7Y/szCYNYAQevN/hVfXlItVfwB8E/v4HmfabGNUiKL0Jo+4vFiv
kCrTu7TeZtxs9OcP8TIUjjzdaEBRMd9ZpfFbXnLT9c4rum73tDyCY23u5lgHhw1/FYNwhRoehI76
C6XXh4443m0b4iLKnr0CbnC2HDHh6zs+tiQ8H2yqR5Dt/9X6lIBEsNZnB8Bh4e/6eA10JHQNjRhY
II6/QlVbzjS5tqZ2uRxHduD8Q7apvMFGSLpqRiaX1lHvHb7dfT63Ta3ZnkCJpFtagf7ErMBO/IG/
zFtI4YHYF9/j+tjdHD+8EuWqxuwSDE+OtRosJ81g735q9vY5pDKdj+H535OOBoLLR4LUz+dUypOI
mIcT1W30E0KQdS+cY6jtkS0Lj/pbr9kCscisBSRzjIRQYh03CDqkAiwq+ldpiL7J7UWxEYQinXwd
EN5CkEKBR+2uWN0LjhjzGrvSuU8INrPlGTxmv5PbvSp27z5Q2yjOZNYKBOgfZwshdpmg6tGpK4OR
Oxezon1Y67C/gxKeXs2W30tmEpQrslxnrQtbzMxMxwo3kFGOKhX9t6JJ7sq9w7EHE3apAVPyQ7jp
l8Mn33zqJa8mMziNDy1Tm+1vG4Rq+/rtq/Wwpdt+YXMN4zDfFCcDVjejhRdOnEqAl9lssRpQxcfF
eEO8Jh7SWiJN5AjWC80dhCG104uEhxZ17du75dOkB9Cgv876Em7yQML5Xvj4BLtj68GI5Qv7Dxaj
GK8ECECjeYebWGfRTOjtLOWUYDMOkSH05p7r1IQ1bfuDAw13+UyHsAS7yc2T5m37WYHyviNZ4kEG
bsoXfBJa7Wt5HnCL26p9Yr2zvCORPJNF/S9FuT7/0I9hn/l94yjvFZK3lCq9FTZfxqRF+5HOTlAW
AKR9zzEK39gmz0pRtEK2zylB3Jvjm8ack4bS2a+xqEDYnS8Za8CmJiVUQUo9A+LjNYUKaP7vH9Gt
pgr8+mJOJswJhIiSK0kF1oxF5nEz5vgXVIAC9S4tESQjsoLp8iZ3bkYxblaD8ynnIi9IfEGD5nHP
i6HMTYMQ/hwZz8dL8cHHRRJ1RxTapBPhhnu/2NCoC80+Nra6QGjt4MKYeSry3avTIANsNNznra5z
z11gIZ90Q732JOPFF8e8G8qFMn69VrYeDPncfMSPKguwMMrocgTLGrsEu/cvxsK1Xc2/e7nqej7D
bgnGeXssLbVOQZFzvsJx2jGexi1UUr9aU3X+Bof47oquwXK2Tny1IaHEga7daogxaKsczWgwgWhC
V+BNjd/GQrYriFJjKxBY4vStYO/rl/YOP62B72aeldqFU2amytowCdy30EC8RmDlHy1meR+SgID7
2F8sfSB2MKAH03vRuiJLhvC4et+ec7SN3e5LutcwSJM1cgHtkidWw8auAhSWPK3rCkNpMwSOI5nb
nzQx82GSOJdqcbRupk5aF0erudOwHqsZ4m358QTHKnoVHHuI3gMZ6WpwEbaYA4b6OIUAIgbDBDTh
5Ejj5EAUbnl9maKFE2rbBquMRzmPE1BlhQ8rKmXUzpyw4lajg3vkdhZ7+zQk6PLuKmhhMoITG/Ko
UWIdxorBDIy/hMKTI5lnctSAc8MLhITjGEqQiXhn/GmJSMvnifGso+mUGaiMOmgGa39AZw8udFFt
+ZPJOIZCTIRlTggrauWFua9ogNQP4xJNC7bDf+14eLRm14qYE53gv3LBtfat6Xh58E+gi9qXx3Yt
/Yvk6e9iB2oxEWgzO73CgbF5vJ1fWw58x9hwJ3I/LrbFFJM4budW+n3Tk0T5dBqdDcSzr3tlnqVD
Ykv4StR8mIFyvze1HbMNQnZeVKM10vBvvCF31hFkaHuNVrBXQJH0kM6Au2Gjh5THxqaehcGXDd0H
JdxI1GCjF+dwsT3gUFxZ76eUA19f/zoskA605hSCssOUDjiVZzAmaGVL2ozG0FNq+OiPB0rkcw6H
EUgEUu4ApMyDFoGoJS3sNDT05MWu8axUq449M3bqox3YaJ/MjRxZeQEY3KZtZ0DRhP2lpxCL5O1+
aQ7LfvUjRzhziL8tzwAFJNJuF7bzVQyyx9nP5zlp/+DgjVEW4R0kkxbkNLlrmv5wPVB4KxB89YMK
rgy+MX8TN/Rwari7yAflqjB6tCoqAi+UfKJQiGaiw5OcdTBQA6o9Uoknt/HKTp1ARQDksXBVGS6L
+yBKLYVnBUbd+RjaNp1C3CMNr5LmLOqJ0Gy/fTMnq66h0f/gTTJWtiyoCPkV3lYCUqBhHBRzPCBB
9WarEXQFrUI4NFl0M2qeL1oevsz+kGVPmwvHtxNOfGNyuIsxifFZpBIr8BOzZYjRQfqhR6HIeL/5
zZFEZpgbQwjprdrcaykCRTQAQF7Rxmw5sR/pIBYIUringhpuds9pb9nfCOqAgOlp0nkTbCwWOq61
P+tml9bnJnbgZgvpUnu7Ln/IVcYNQgS7xrIodHnF/8TyRT21xHdrZuhCuMRldKTWHXrIx4kd/ktM
9FywQ+/MdBgwGFVTgzjcRuAIT7RTkUTotbbLWXubFZGxlH59COpJXpSd7k10Loha0zTT5eTqA/UD
xxCm+W0A868meNpzl2HzbiV8L6bnAPz46drxscNS3GtNsWfJ665G0YWKk58pcNi5h4JBzxEyTpD6
KOsWMZqFZoNvUB5etAxiO0QcXS7cuP/UHFIaiZ/fs74euKm48DphzRJifF4dkEH2ouReBtnoLjth
o1OUEbnsmC14QixUbXTmdpdT9aRbjDjjZ79fy8+aMpAc9h7njUz7nI1NsnIaPzh4RMdpQMlpVBTD
8DHznDXH69cDlRc3lUpt8WrcEtUO33/oyHnS5KlYMcnBKSXmZG46LW/3U4IIRSlC3lBgxsvCOrLv
J1zmbFfXDGFr2E+68QIaaTjWQE5u6bbOUHjvAreYzyYFkkhEpy4KGhKuv9iTdqPSRHOWdY77/2L8
rYMRjyiZsPna03DLsi0BWXFsW7sHiIoQdLH7LZkDObq3KIj0WQM252nhHVpbhv+ApRqo0vMsgqd2
Bv/4SVpLcJpGe8ZWWV1/ORejZwGhC3doMzywAPtYbjvd9XLSIyl2+gBX1qOpRrahJalVPS4fSeFB
X2QhywrQkC8vK3dnZF7hIQUBAPaN7UkwDPIDyX2/OSlII45ccqqTz/QKnNFdfLEDcrxPrwThwU9F
OzKFko1DJWA0u83h1LFx8T7jGpzPS1rWw8K8hePPX+LJsq9wyRZFhyPrbIle1pjrMlG45Ay9oxft
+Dm8HFdqTeJpYbw9C0Ko2FkifOG0cu8J2cQ+EEOaCEhaiA/nn7RmW7xbt7uFlZk00xiBgJe+qqyH
UcduT7EfLWfQpRBBWbendqjf6soNqrFdusvPJ2XvV5nFBzthO6sV0f9Cn6j0yIJd3miBNJ6g2mGc
I3ku3OHU6eX6oeMNjhg9VgZHOwTe08CQv0CRELCIL71x0GBEfaCSxT2xXaO3mbrMf0ns/2nFDF/P
4ZlI7+/nqXkhXHwGjf32fXRIINJ97ueDLPRt7rvj8/Pa6i6XG/4vM9XBLNp/n/bDqKzngOrwMRAY
VgppGVIZP9J6yBHaoiTaT7BMyLum81q6JqVB7jcFV/zRjyt+OXVcoiRCG+/gt2/8D/hUWELUEJOD
a215fnbveZFUVc/3MFoMip718HXsUyXMYXpGgpY6iUWns6q3NY+76yW0k+SMWdknTaG7PkPqxsn7
g17rwJjza6Qmo4W6X2nZ6HpRS6RicGzX1/xeZdFxSqxkQWmeUfo8kpvv1La05R4oP1qxSf+EeJeQ
j/8RT1cKkewk7uJvK7TM3AE0Om6199twqW9fZrtykhEKUcAMG1X+e+TugW6tv1lysOmTJtXwPasy
4UT+pV7lXGT/qKmkAzsHDg6DMmxBrX4RsnbEGryhBUbWWcFCJ3vspqaTSqkcZWD/UnzNXighk4Qc
vUg0YM7FTh0oK6z3dKJ9BrPhSXwYFM7e2/7xzuyScTM7/RfpZXRHA7uy17LVUlZy+MZq8KHq4fKZ
G30wmB9flCP7dey0qHsyiMxYA+qD+TeKmV9SdFgATu3lBGP1aQiSNWtHppA1eD6+50E++mqzFH1h
m7eua1JSAN1qXKi1YwxSEVxCZQJWUZMBLmoCRIQZ8zSirOS0BzdVeJA7ojOK0Ti/YYhca0DiP4+N
Da4nm0IIZvkJEF7OCIRfz2DICasLP4gz68m13ArRDrpVkw1bGE+RlwjbBBhXB2M22D0Xo84kJiMR
9ZmZuN477GZg6E9oj/7tJktel+6DE8DDc44v4k7Ku6+JHw2gE7WIxJDYtvhKgbH3QFYlbIHhu9fB
bjExvibyjCV2PYtAA+nkl2Mja8c+CF6Hiyd/Ea1uqdDcktqIp3pIQ6AVJMEnqrvzHE4lyMfokkII
e/qpgf3pnphxBZkgL9Tddt4I7aqCRQHKmbaK+E0kMBq6KddsS52iA5aD0skQ7w6ain+Cxqsvu7mZ
59A9aP3HGZQh4eflVS4zYxx7TPlfVi9P0Ub9YRwZ7wS596ybYM05cx8RCDF3Bddc9MtDySuaW7h5
sWkRUjtFKlRkKUdMXHwr3IrEPV7A1Lt4lpgKNpwrsWrrYMmtpBA1fZm/CrlYsLOBWd9I4tZsFtCk
RuTGCtAG8viXdLZXHO/btWIMFrKRrCl8UbLTwcMqHnijZzqt/wuVjRdExkadpTY/gHgT0+5eFuev
ickYJfpovXFK+SM6DUm28hsTa8SEl//5ceeGZZZUgGfU+QCvrszyqVMJNVMdlACLX9LjhjHRuH43
rKjuBzTm0DERDETkHQESFczpJuORTHvUIL8ar16WpWsic3flgCUq2K1DIY29PT0zY3o1nbL5jDzf
pJ3KPiOov7hASeXdACV0D/YQn6qq5iUFKuUSwCXrPO/++uT4lghbUzBvtPRhWOdzWYDUI7p432H8
lXCAIeY3Bf81++V+G1tejbctJ9BMbJiUvWnqTRNf0bvKcjWbDkKURQ3rIL5FIl6rq+u/yY0iYSSm
jr43enHBTRuSh8tymyiS8SYBOuReBIMuYnmkJfEocggCSlSL2i1osiibWvQMpU5WPV5/uKxBlObw
BBM/YlVSdMifYClcAQgKz1ES3M0RxWBxkdAUmnXSD7SIHSG52VrkmzNG/SsQ2LCWx0Uve0KFvZME
xENd7QivN9J1kkI42ZmRQmc++aQos8r9cnVHU+wIw7tLcPG6Yg0N3PrCAToDptq9JYGyblHkUaZW
j2TKV57ar4Bqu6/8URrxQFHvNzDYhHmHEDa97P0K1jaVExr3nZLnPWHQRWYVl9iFBrKi1hHT8xW1
0Op5RPbDppUeTuWCsN8vJhhN4YNzic5cVntlrpj8+88x7qKtgPOZtaHgg5NR0ksFQrv8BVgaY1Um
z3gto9ZpxsSdgP8s2gnYKglly5GS8YT0ysesSu9aFjqeYgZhMKHFTLIQJI5of0YJhrk8bYQJsus8
ksawWc6tx75cIy0s6/ijqSF6yIfNQ1AtXEVtAe8pVUqNDiTO1EPTjX6tZi8WU2kI/9PiZgaQp328
7ou+yWNF5A4nqXr92ExdVu9duTYCTKMch4iULdub/S+EsK8JJmjV1e75EdwD37NRfZ6jCAa540D1
HjkQphRJYFbjw5gvC1Gez/s8TGiAPshvI6KMLWLuWqcpSNrBqWRbATMZkAlD7DjrsSJKuKHzV2Jg
gXERseF6+dKBMDGCeB3GmpilMMzyfExkEkfVMxi21xFkUdXcyfolgKX/iUmhgLqEs4EqHJ4aCH5U
i0uBWNqKIcf26uj3nfVb5mgU1WTVyGoZSfHfgEHqq8eI1TrpOTAteLUcVlYvIMHKr7/p386lHHZ+
1wLgOk9x97pD9cdg5tfyci8oOqsT86o+qdF2dzHzYfxEPOPL7qQJQ3dVnB2fE18BIRf0UhsoaFUL
HB0l+y+H7DyrKS7G/om2dnTLdrOHxHiAuRF4iXfQCXavBJynjjcyQz0tZVxg1D6fT7sSFtQdwDUW
3hp36Tg4mmc8W/d47aedP841a7C0o0YxYSbPkQS8nqphp65z7dBlDpCKf9++U7VMBC5mk73jPcOR
ghfy6rDghggVb4hro3BfsvGBUGqhcMKagnbCWPQ4DpC6ThmbFbl833Z9XKn1Ss1I9TPnZFrouxUA
g9aXNn0UlwMy4IlOniZPyDJChuQNUtDDRhN0DyEZz+obF2MQxT0pylQvYlzdghgnby5fo6EMYbUJ
lHQPnv5F2Oah2FMcJJjQJViTLYMOlZlAxk8e0g24lJ9bvVj1ylA7KSojG+RdlCgqZKp+ip9FQSRh
o5BGvN18+LtIyAa90BE0EVzwI71n8ABRniYSxo3iwNM4Qw6kczu0QsTQOK0/Mz6sKLHhrLS39p9m
bjjGusgFS+IjjaIouPar823EzZ7eca8Muq8ClotjxQHne+KX75X3dnZ6vsr6abX0kFv6+cns3T4E
SxmV+JunKLc6LAg2uLp+w0W8VFEkfpj8AL2grbcbK2vPstWLP4Yfx7Sh173kyOApt0QADiRVYN62
vm0XItFNFLKtJb827IPkIWqowc8EfhNdw3YSc9VIPcHEhnX3iBjoYMuw1wP9QdjkEv3z8haQ399S
btlCSVP8bAqimfgeWV1tZ58uhM94eqT4RGXLkOdjeAP5WOvuGWm+zR1F7iH2e27wrHGNoHszMT/7
Bb0tGR901cMyzGJvENZBz0KcO1Xx4N1ua+iftwW4S24HX/Wq0OB7f7qiuXIv4RnKbDlA8Szo53+h
z8fCtJZGApwwkxPXc09CgrHtz00/W7trgW3UqJf1P15KZig8XCL/OByG3x+jozOC2Zs1wmc9y4yf
vxQ2taj7SP0zhtlT1ZhtpX98oyQsLFJw7HRHpow4mAIIx+uq0ebQftglUr+vU/0BUijgm2nx43O0
OScevrnlTo8KJcwRiiJ7wnNmblD+EtOKZNygpeUyVrJp0x8jfIB/eQZghWaKiiVD8p3WrDeS2WYn
+ATtyo5pMEqtGp2EiCFXduLhS/+1vemZWWvYsmgbz+a+YuQQcISOxCJHV7efmVlMxCppw8Ff4V2a
Ciij4GC5iK3miOdu2H5UK5ADXq2sIbA1eB4TF31fWjyb2QxSyEZ8L9CaeL2WGotYkDnlW9k0A4Rq
3Xk+7ZcpHBe7zDGG/jPBa552p0V1d2I/uRqHKt/bTm837qheue2WJNVXFTQ8IGbOU+j1bE/+9z3o
KkuSBw89Bjzsj7KI04vdygVHzH4Ii5xuSM1XxgH2MqrHjujbnitMD/FSVDfz12sJiv3ntuMNKudu
RSmljqtEK5tHwcTwfHyyIkst8+BeqozKDrQExv7h26NA5g9t02yOW0aMqqnEldlqgCKnPOFCIwGi
Y5dBoU4AKvmnIhHOVw8EhIKzVIy6rhKbD2kLzszLdj3AH+55wtbnwawdjD3d7yHnxwknmWMnU3Ca
ToYqjcoSk0UVcbGjtSsT9EUUHF/n6lRsVMVR4NWVJWcZUmorBazUTw6V5JwMsaXYQ0QCpzDbuHZL
H5sGhJuUCVKg5my/cmUMJ/gQs78pjyzl/qy9L6rysAlbnwNibnMJL2OJr7OncRgJnrNJt0KzoQAO
iUmjhKi/9IxK66W2Gw0TvdunLbMha0MWpODc+dvZKnuXG+/QLFIG3cnmmj/SJ0UyHqDffoMdyvlC
xtSS6hrINrQUSuSW3+pfxpO0M0777Y1IZx4KLhf674PbuBAjiouIJYv28XGFCru80HCVq3D8qh1M
Hed6n+nSJbo8MuvvrTL5w0SYVFvcO1lsZGxwS96H25whUIRvoyZtSNagPqmBL9YbWhmN3EiXZVXO
7nibj7wdDRpAihjpY18iMVdQPX99S2DGPrtOsCqpTmxw/qPgJsdut4Q+p6IN2dIm9uIQqeSp+/B+
WY2x2Pa048/+BcWjyyQuWGUO7TxWuaF0Iwhb5f9muHFHgLRRJGdfXNEulYLqQN/gb1NVq1e0x3C7
FskAK8mhOKfcTtpa/CCTco7uzgBR+7vrasxdCNW8EDWY6BUXZFE2TAunOijzPfJXRRgGdvJXol9B
T7FXBT5ndyXBwn9q1vukFxlr0VBdiigmH01pTLvgDHDIwd0Ie8tWlYetXbKLm84MXBcIHLNg3bR0
HZk+ab/J0/6yED37uSEt8gBgmJMGEn7La5FBgBYKafBvXOBJiXqLtDrlbDG3JGntm01q2HPLgXjj
Lq2M4WZ/l+CGHBq1ODryCwmw1s+up8RaHqZb6+eSCXUkpnuZGLr1e/T3pxXLceD+AbC+FRK7ESw/
Z/sI2OBYoPw3Z9erCedluFemC3zgDcvgqjJsoebpxG1duHPJsT6r94VrAsW0BPAaHRIyFm0Tpa7A
oNjv3u5tD/xkQ8gFCYq99knXxPEu6VhGepgADM7vOr9bcFyNX+vfk7zmKUZcmybMmJ+vAGEzJ4KX
HLWHkAZcT5Rz/uNpEhypK+U40wrln7eIMoC2EccOfeZ7QYdo6uEp/3ltQKPOWZwkwU5gpzyG+YKG
TYffIiGqYhDqKoGUpR93ORgZiCdO/uLPA1JvvXW/wFbKn7EDLAQ4kAY0dDYgfpFf2+CM1VhkWT7p
AQSJ9nc3UPNzNu4VfYNtUgXbah3owF+hUcR1OSe9p9v0Q0DyIanH+kMPNaz+xbqJ/087EEtl2MOj
Z/lLAcc770eiTSpgNYsUOjthtHVXaZycCn2V4MzR7WyrV5QB4aGYsBAtaNtLD3ADlsib9qEOYCWa
swsj1HA1Qt8NOz/SYklV7gMzStPVPr8iFOGP+32RjKmUf2ba464HTsS/ksNnM1vD9ZBqoa+1adaP
JQsejZfcvSxKv+t4L5GDyJt9Qkl0jPNEMb3BeaL1KLRa9vAUMkOck/SYFPSXK/QQ0kQs+hMzXyH9
pyfq0Ox1lJ0Dts34+jjiSAOyOHyH8p0aK158tE5WhWQ77S8SQ4S9mBNDHSfSljnH9KBzcf9GzuzE
WpFrx9QNSPInHjl9MCQ6F9xnJrt1RKKeb7H9tVF5kCPNvDGCzf47Z7DmBYr5PMq4MUO7FuvGcY1X
cOCRYkmwPVqXO4JQESa7SGlkCdZR80KanwGnvH+J9YikbHG8/hgnL+SupkOgUQpPpmOxzOwdEe5l
fRm9UrkHU+7nvKPh8Ej7zm/crr2IOzWf6F9VG3edbhsQhqGJd5FKHeyAW7BmD/jabsCobiSYOwM4
pAhsJDK/Co7RLft+jxx3keLXMQnaeV5/WiS3QsFby4OvuUIguJInaXdkv/rBEmmm454J+VtcmmhO
tpAQXWhHayN0bUpVKdGW5VIZLAyNHWef5f3MCbPluBVPjg8It6KJiYTe6kOfbQ0s53Xj/0ksmHH/
/ZsEXy2rfkPStVNWINgGcgj4G4aWNalTT3ohlfdUnojv2xqO2f1+XxbqPpSssvvpsgCO1fAxBIE/
NnCa4DPkGIAKWgHAU4pod4wwELfV7lJy77XTJUdxguFtPH7QUt5XjrUmP4yOZ7EcbdZZycFQKn9O
hH1i0SOo0TWOKT4yGxtrtFNjYXV9td0DsJQcWjts/tXEoljUiJXqN2lORJX0L+pIhBy7W7NfeYji
G02sz4XJemPKS0kFc/ThtyQMxZK+bYS8xvv/4610qLLJ2qoQ5IxJvH4jBV16dQLNNIzIxfGwbp68
lQ0S6tDVTXgpemFFZPDCe9Ck56db3aqpdaD50t5wxGQmFASvTIbfT5Y7h1j92CxuftdBEIAJxlcH
Lr11TPHtHS3LGF+ZP/LuqfAIY+9u9MwVclJXqwCa+uq+/jh2uFKiaJUyPksXGM4sX0aqh4UwBo03
L8ptTTBhT9nvxCsa7dswOQtzx2Bqn7ZPUNxavuS29qFo5ROW89yYHgskYtpqTeWuZHkluDAvIvra
RegKMtpsgVTi+3doDUeGY+SviEaP9gF6gFOnMEPeuXGJ8A+pnVc4RfzcB/jm9MC8EsMU06MViYQf
xytoyDRZ14MuKYLM3XmaJzlBLskMw/nELmjuxcCvl/QxD0UP08COXGk47LEO5MwrP7eoSqfTkzyi
pDhBQWAVCGquVlhmljCVyMmKd3p5ZnCo+OCUbhgYDLSZ6Rt0Y92bbeN0eOfGrsF25nQMZw3QuYEi
kImhe99to7PpbcTa1INDsS05pU7C0ralNj1eUNs5C9nMK+PNl/iLfU8vtMnEggPe/MsWZIVcXKpI
jYpmsr+53UB+++t2TUO/aIN077oAzuXPeUfX8ZlRycMG08EOcve3XQ/ztBkSgmWKI6KC+J3QHTPy
ero6MSyzhPPJp4c8LIxXjdyJDk1YKb2QCSVkBuX2cFRVGtuvogxeV1nrAfaM16clRfuoVcILiR3r
f5lvXBYKfvi2h9Nmhx43HO8yxBIaLYdpnsgIUD+KW3LXjlNto14FsG+vSiueApb2ghve02MPSkei
QuwCk5Xib2kxXIB5q5FtxKi8xLpqMB/wrEfEMQtUVKhE2uUDSejr4P6g9Gq5MhUPrNp/CNvSBeRv
EVxSTAtmryOHuv7+xXmn5dGTjr20JEwauKymSOBD71cFO7oBCTQaHlbk2HrnfRqlkRQnyvfBvWes
YtFr8cl0VXE3aIN/mlDXi43AU825l3ee404KqKoSvtrMm2Vr8sTYQEKlJCLqxTMAuBWz1rkoSVDf
FkzEUrovQdFYFccEJazBZF2ydAn5Kg6cbGyz/gvXB1GlRPmRi6v0jOaxDohHHyMRV9Keu0Ddk5QM
tcz+S9yrjBrUxVAoN48UAZkoU1NUGM7vJR6prg+zUSaj2XrIF4vWzBKmj6kmXvHvTEVy9FnOSF5P
c5js7U+lBv9ZcKMZVbI5tzInXr6APYqDqZYnmG2M99eakz4Z4ed27snnb/dRaFY35Clq6D+1E3d4
gjv1WswkHsZ4N8Qxw69aiyUcQg9H0sulvFej5N5q8QhHogDwXIRdhsCwuqrysjVzw3gJg8DD1Xpz
TvflsqNWmZAwY6gPxCRTRHJyiC/ssp+6aeNV3Bh/qu58WotuVf+DyZDBd7XJcyxHhSu/k7YZDIU2
8Qev0/gHHjfuTIuLb+vEgpaHrZpVMU4yhwoKvJ57OtSig2fZVlDuykXNb/D/Jx4xkoDIkEfwhJzP
XbUA0qOL7LwZkNtkTJlJ1pwslMdLAnSMSpgbIzA6WeTXFDoZi3dntVgeJyxBKHSsQkiGjR93j44I
AfQvLgNPriG+elNsS9SLPuew7oxqi+GjxackJri7j+M94usfCbut3MR7NduEcnNHM2XW86qyjYii
h9JBjF51YEB6u5YbUHeuFmAY6VCJwQ8oHLLlAaFTsSpJ6myqxDJYTCiGRIDvhQtmC+edQx9i9y7G
f8De5FN1ukw5XUQ2Inq7d8CDX/OCCXUYmsCqGH2pQhGyNgoFeDS/Ajis13bNHrYOy85NoLVctnzT
lRSZmiBrnevhw6+mG9+dQHh6jmDWQV0pvKRy2WgtimYgJXRUeZpN5Xba0w0tROO7WUVLssxBJnAM
Dp9vUP2i9pM8Tzci6KYYrkY/R3aMmWOaMzYV4NYE316OvAgnCxtcxuTmpjDzy6JeeEDDzSsvSuR8
Xsw135op5aKP3/DDfrNgchZghNNMdkNmN3JABqG5OsVQMgNvIFlS384IPaJ7Iaj04b59qJGoICWb
DgFU8/RmJeyNVNwIyLgNPe3X//4HmElpur3X7pVlckKsSnjRE3Agd7bpa2FERrZCpZcyywweMuQu
Inf096u25cAho7kQeaCK8dOiWMuo21ncKw8O9e8uhTqpljy04saec1tB0IldjKYNhandc6rqcNnx
cd+XAYjepRrHcL2JvqzERTYBOKKIhzkTaRfGlxEjgI3AQCYHGEHRDdoQDY1icudYsDAPF+IqU/QM
ocOelONWCvfmHcSdyFXVGjGh5ihQw0D72LdqFizBR/vkBGtmnWin1z9hqAEh8XyK2ADPAs9BPJmO
UJQTpV470gioesDl5LsWbkK20mtgD+Tfooj4sAa7SGppVZRLeKDcVBWoWvewZX3/XhB2vF3SldlS
FO2hD9nqcOis0rWOjbFunssK1nZojomXsnUX0vAxCgSfr608Zjqh57xpbQvYYzpix0IUNw2WvbRH
FHbw3ZsknJuyx2NWnhveaE32RQIvobkr1o0sSloy7vA23VGP0p+xVjvr7ljuROoivAs2rY22Ul3k
mlaXSxbrZBbxoUbYN7OapfsIbASRFh3xgJdhAjzkCzRSAkKir6K6PkRV/WdGzS/N3E9VZ66xO4zm
xVsjEeg5XnO004uNkIE9xZMzNG7QPhhXpeXOuPwPnvcETRa48F+nM3qIbm1p1ATSrg62ZpQz9PoM
LOmKRWYDPe5c0Nmt8l57vPS9I2Mz46XZRaHzsaWpl2YjNzQOsUHcY9am0wwrqvSCn+1EW2Aciv2B
NRYmEchw2nKJOydCCAWzlJFXjbxp+i+n//PLYtnMHviRVgNRGhXcQFssARiynIZxUidBeyAiA7fN
5SWtM6cQjC9qBZQHQjAscjqMTOYC0GdMTMXtttbT2GS22sXYPAycPL6Y3TioezevZ+jwan/9O8ei
y2fTE+RJDhRsy0Ik5A400niGP03tL9AmTuU0ZkHOqTYZVBhLj/5Uw373OO6Zv1YWa90tplBHEt0X
8aiMLfO9DjBiihLr/32aIFu72iqqjSJ0d8cC5DblHUZZQ+ppJDaKuQatyCfodbrKkv6egTVFYENQ
/Kb9g3DOfmuqrBFLURycwuo5KwJJ9bDDdf+SqMmhd2MWdrk8UNGUOQkQ3jGgeWbnxj3bKUlPEnvG
HFGIuRyvC1daKD0WrO5X742C2TeTQ9+1nK5KA7U2UQorcqFhWk7c0Y+LP0VKPzgSskAmmmUU+9C0
7GQMlUW7sQNcwwIFfhASV6VtEtIlpEYlCfJvcfnzUEwLK56LjM1WrgqUlIEzFe4Myf9MF1eJb6rO
JWuygNkpiDuh6zg5k0SWCXbgTHGBB1m/36zI1rzrgB7NhtxzCWku20zZnvNuuY+yrMknbBvIsArk
GlahoeAZ+16q6B3WOMCGT2ubAhgdS70IZ1kysIKMLTi0kS54CKNGSjcTka/uZky+dniOnOZUG/5I
UPcf4eUafmvW5wSnLFs+oqIFq9MXzuSdk9UiasLtMAxG8QIIQoAHPboDVKhpwKbeoLgI/6V3Wj00
TJFsfXrkpPCnQDI3rNHO2VmYLtNqe4PNjGeh002ARpYxGHDyYTSV9sMF4mb32r9I/c7tr5ou8RD4
mMR3zLjwI54Yjj11YucKW9/TV8Al/NOJ8ZBSq9x64XrW4RYWXWplyG+8Ra1UWo0wFCyk18ZgcNkE
GqnGoGYYBudVX/Xb3Hne52nqfiM28OGOOW/pahprnzTjtLSOPgad6BGFvh7xv1N8hFf758ky0Wdn
xXRDLKwfPzMaMPQ6ZiGlpRcNkRVX93zdCq+b44aVogarJJ7GoszjrSalDNrZ3UHpVhNh9qEvz1G/
fgPDYGuVRq+6eXIqftxM/OW1iwEtHo+WMOtuRoXKUacEOlOGKsLGdJyOjnrXJpHvv4m4ZSgK3gmt
nDccArbItL3TdZM8xKwKVDfwVWkPltXu0GBiAvzteqpm1itY0NAwycSdo34s1zNTMwwBCWQg+miK
UabCLChxXJCG8N2WQMwO9vBZnlT05EdPoi5/KTGPw1Q0Xx5lrtOm4qdPhppCujcjXwQ+egFnQZA5
pgJItImUx+E9hF6ABGpAsR1kUSHS1TFdsFksMeFBlywGz5UnHxuohqT8xzM5fJGKS6y2DSQqvrc2
t+59hkpmwz6A70M4BRgFJjeUkvjrSOv1YMJkpX9e45RSpPOnDVAWANTgXGKW9u+0DDuQ9nvrUgsF
HUalUmAUa24DV9SmNErLlRzGH/KhTfioOesJWRO78TJE8+Es0XtGEejRALKnQgZq+NJ/GSFbFA/U
qS6+YGup4LMRR2NLmjUWaykeCWh9LBIyhE7KUJKw/mPJtBvo4pD7zmt1vQZGlMRlzXTd6tLkW50A
gEC2dbwSGQ9dkpCh7cRUSpj9LhazYacuUiVMno/QhlT+QeS/fjOoYS3lz5PBrVMkK2Dlbo5kPe80
deW16wnCxR0xK/uaNNuyOojVGMfxBwF/jdDsfrPf5NZFlv2ZHn7NJWQWqi9Gzs/qVU4qg7MphOua
ueK9l0EDPp34YthemjbYaA1ElAtjldKdW4AIrFyQVYI4xnfGFOxfzCu47srNqhnXj2CQNpb5vVrf
F79ROoYc+/kss7BwWzGzVllaOSPaIvCyKcWEZaPaGjZ0ZUHu8GrBTMKZpm0hnMxNOgrWNquK/3h9
X/01zPi/o3pjQWxfd3xJiU/4zIZ8Whnqj7GdpkDJ48dbxX7xWzozatxk0kLrY11jcugjvRoQq5Z2
OvqZTht62e1qL12jCzUNWo6Vh8A8NBPU8vh0k1L6tsFvDi37h0RQIOZtMQ3Afzw8/rtvrORQNWsK
Q2p5d8K1+1WwD9xrTZfIsfX2Phgh8w+qTyUcvH4UeAOZ1Zc9Wegkd3RS3oP5l8Ec0ZRZqi5esH75
10P+uQGT6575d8lQEZhOo6lFx59uBtv+mkTKibBylFVAuD03y6E2l2n5wcUdxuan29EuJSNJBip9
kLDzI5IpNfoKhyKSftdW9ZHDOmFcItJVh9YWFMgR67cQ9xHF6KhKUKSdnVd2mekX1F+U78pvQWVn
2ymDi0+5+uIUqmsnQMn1tM0spalR1XjPtds/04SXSsGLp0bl5bi1HCcHAEKfsV94417fzP92d1bo
XEfB+xNFXkm6YvNvGsl/axFuujVBuSpZ6eQxyaXCNNuVzf+7uds6M7rjQUcoW2cZOdVs1x5ji97F
rGO1BxxF80pBpBjJKOUi12Aq+Ds65I2tmU+JtR+ftrcHj5Z50IJJ5xGpQk8eBpJIeto/8/YcLBFI
AgwQ20VLvMZz7HLP3xUCshFKKl6oig6I6rcCKZZ+k/YeyhOUGwxPaQlgrZz/pj5A3G0PvnmsH/iH
zSNMrJh/343juOGtqusS65RLkeneH0jNDe233Eh2pIhK6AgXAKVAg9Cm6lb2fHkqe41OIZLTpH/0
u2oyvurk+F5hS/2KsfiRN7/i7XAb8JtetnoTEQsbcIl9FWaJq3OmvDhcREg753IceIjalctvDKA0
onytrCnk0y+d5Up2cJJ/e7CT++vy4gXeMGIiPa49HaC0BC6MG5pE1Lk49LsO5/eN8PiJYN+kwaQK
qx/qy8wWIDzmyFObR70BcPbfo32+NdiaecvfCjxbEfwR/eLlXJn7YWHHC1pBU9wH/5q9FsTBiNcM
nYDLG/B15j8bO9vIiHojCeBBqeVsJ1IVDxABXvbFg67a0jhQ8/zqaH40/1pGXDq+4Q/PF9MZqmM6
OtT9FcVGkf9kdHYmFYSALXK0EiJRBnO+veniQo8Rc6RzSq5FlJHKppbiUBoBInBt/DCUFFm0ynek
4XYjv5t7TUkUvd1wQVyBYn2f7msU6WSJj6zjZVe0M3p0dmGhcBhEa1ZYFuJaQsO0AplzaFehftLs
n4TM5PkFCz9OnxnuN5Hj6r0qTZeBjKXrbVg+VuFCwXR3KHXwKWn9FApze22ylVzsRfKzrXSBx/5D
/mCHfNdiR/WgBwdhF2LDkeIjvyNrZWsv9/fkBq/8FUPKGTBE2/p6+4OsO4Qpg/LWSAbq/WT/29m3
K1OtypRt1UnT/uKEwIaZvJlBVSRLShFOZEfgG/58gZH5LsSO71qvt3VFPuHyiRnq4xrPsSBmSqqb
G9TnQ++5vegTBKRhhKaNEU0iH0NaLEPm5uzACn4oH6UK7KAL0qQL+2U/RoR0AVTnzWJw5vXm6m81
vUEFDLPTHBswxEUXnuDC9SqpRvb+zxcHxQVdtpzhv9ApXiTLvitj240uq6BvQ1cRr3Sj8ar1EbqR
fsIoY6Nc2e3Pcb4/ybbDi94/eL+7iVxDfk4bQuuRdVMhY44fZBj0nupatryT25wG9Co1AKVliG1r
hBcrJ1CXMzmi/kEBPh22PLAqBN/W20JWdRJkERLQ8QFIuwfCnRzRzprs/mmGT5uHdKrAnzC5V94t
pDDNUs9RQwP/fMs/CUEMjA2MRkz+kcKQNLNgVvunCPRkmMyq4HLEZ6T7StleeektTSgnawBXKEu7
4n4B+3U4fO0opQhhrOQZZBAEguAlIf6fGwx7r5ZLi1WWPpEK5zqNcy3pGv70En+6XkKcwOkY1NhP
FqbhUy+y0fXkXHvlNUfyxDGHMSYAIi4xvUTdBys4EL7whs0IfxAPdxH90OxIQiYQAKVWrPnFHhv4
qMXTz22dy0DEFjmqeaAVt5B825oTbZFEOLjT/pCwAEWZvUwX+5sABorUHy0T34jRJjUp/D3vHRzc
0Wiv14bS3IBVSWHo1GUgyJTQjlgilhB0Ba7OxVGHN4rkUvEL8ok/0hMbMQvpe+n+BdjIQmR4fhWC
D+70399q4zpmaAB+3pr+qt/WzIgUVhpIH7xq6Kf1X1cOuKrVX1GDLZtCCIfK+QkVMzgbyv5nTYPX
qaKoDtKsKD6ZPviL8fmzIUrGsAYXKh43vv5pId7wKMQq3Gd3abe39HjxeRoDYxGV3qD35+SvSaX0
YfpGjDgS2ZpJ+v+QCyVnw2rw7YWiryOXDcPGzCuIHwl3PSVK2Z6WZqdGoBuDvrZ+VZ2FoZEEptqN
gH9Nydv30hqE1zdU5fv26wd0exnrPQ2dfSaMR361z6u7IgNplBNdVmpaLAeCg9lqMh5Ojn14ndt+
fNnaATGxL+BEViL1c8cZxsdArC8vHQiORv6RBOkxHBBA4MjN9yhVLiG9agYsNliqnbrBZrDGITDd
248Am/e/2FIDjPKqXxzAK4qPGoE6tT0mB7mG5J5tidHyS6tFzZCpdIGOhwYafhrZuOKTwucQMaFm
+w2OFyv3zOyDuJd80q6gyZDlm111Ym6JuFEk7FBX80kXDbySMUjTatNv/3VEepnreH9unfLUcfe7
Rq3+dp0Hzrkw2XsiV/vctsBlAUieDYUXsrRgt0+OUBnepptjV+gbiOZ/cNN3cwA+DBXuxDPUqtCU
9MF8XCox4rWWq1DNLMk8gdMrOMXA/vog19m6e7XN1efXUuSFpL7d0jxYT923LzFlX/KtMJvIfYhF
L9N5928Nactjxhbc3W2DT8bqccwSecxwxEMcg4TCERVJsBgmHLivG4MWy9+HD30zEDxK4SefG0Sf
FyBeBve9Fz/yJj0eDAhOesNPwohodk/83wTjt2cfNKc1z7bJ26AWDRRInL2ov8d8m7HpU2zQzdyK
wq7VFlSvvbKnKup1O+WzdeS2evdZy0Ai/PDbDGqVHrOsR8fxmaLDX4Rm6qWDnZx7MukXtnwjtkH1
FsXsR6CBEQTpDBUFc4OLNwgq+/x4LUFEJSGdWh2QcItGXdNUNCEGVbZJkdoWE7o1p8h58Mkesuau
t7oPVQtNdQXYZZtsarjvwQD0igIAEz73dSJaCL9wysXelfDz6GXE9BGrKnZyheqJ9aPbRK2a3p9f
FSpZvJZd0/6vtRxRYeQjEzrtOzoqZO6HwpgC5xg8plANJXTIDMpjNiyoDfva/MIRS4G9OEef+V2n
r9NpAMXTTcHjho41XQtGUGZqgEA56gbEQhxawIKb3/niBZW06Yliu4lTdk//RAOylTyYTy5L2bUC
8Q3KfHfkESJ6pHwUfaxQllwxwdY3DW8UYmB2IiaYk22COLt2OdDrBOpHGTuMROCqoacsgb3gBwTY
zSC/N6I6wXsu8r+qL7EN3Jgbul9xMQAt4X6Uzq9WCTVIv7r65M9sxPAq/Cxl7z1toMKNvc07cG4W
psWyPrthgoE5CPBE+JhHiJxB5mMOgPECQxy23AgKZXDH/FmzpuBkn6n/U2XPBRIA7eTj2MgCq+iV
RhyQtLQrI56fFWgxW3GEF0YN9XQk0qfoGm1vxTV3YHxkfI7HASuBqE/6vcNFwyHcsCSGrAfmGs/I
EMFxOfMjZyZ5VNtHV1beHy72djpNFxDqO0DtLKUA10gQPAUMZS762AbjPhDsQsQt7BBNAj5+ilNY
t1f10YAScTmaVBCYFOTQ1oHgLUVioEBxpRNkdPSCx6GbfEtT4/hzq7wIMz/lZCrLYDkMnqp1g6fa
80k/o89z4HS9eUCcsjA4HlfvHKC6FOlC3LQePmHERRrecS4xy2PllYxTNHVfhX7ul5mOMdIi0iH0
0IkNL2/7GtvvZdpykLS/i94zZN04t/mZm6eCpOUn8vzTOj21sOMkubFo8VQrlnnD6WS1gGguSJN2
/ku5rwt3CgVki4cPqHeW6nQeGMbbCT1P/QwBCqs1nqQsBAGKp3UuzhatVl6ig9tTndo4DrxLMXdm
bXoA0Z6S1chrdVBXzqZH4F9TAGFamTa5N1Ia3IBDl9u9i2eCPmfQ+4M3z5iXhTOKs422WpG4wihx
Bc7q5M3BGkp81xL2UP0ZDibA/hBuouR1rf8Tyi5BaQYVCC5dB1qNqtMUBuOWNoQULKnDbehroqgA
dzf2+FoiHbAazJV2s/gcXUQwXvGKNjBN/swXeG3dTPKwMb7l2PSRkIHSqDIJbgfc1ia3WLcM0kkJ
bdDhxw2NNKBFmoMzuB8sqIlbkeUPfiCQP815PUnuFwwTwD0ZzsReheEEK/FD9sopzQ3cRtGI0IXG
oCcUFGzxvCF8khM90ZRR5ZPZbrVGePt2gM8ML/DBR9Jj4C1MclhomjFBK73lZTkv+KxrtkPH60aF
MphcLpKzWaTKEatlPlvB/EvkeydEfb/b34stCfYzjvnlp9+cTRuAjepc7O45b3yBcF8dCXhFshRh
/1vdSc1J6cWWa8nLZs/3iFciUR9qQf5IrsQLala1k0auu6U9vnyPI/4Cd4qRSQ/ETlZCDMoDUAHm
Mi7yCsD8bsMrnqvp/763uzOlja00WnnQ+BcQgFfEMMfS6rBVSDwbvT5h3v5aXI3qlQJzZ4APltWY
hRP/LQUkyAOvQ8/1n72XBUENbk4OaoGOlRRe2U8T37G66EcY1z/ZnHhY/fSwDw4d3owho2RR4LfC
FODwiAtcYmRyj1/fX0vDwAfwq1TxagsdclQ6JF3imAzy71eYQ8UJtWPe+I8Cn0hETqrTkEGbG7hD
MrPhSy+kHpRp9jDOUrgF+CM4PyPKdO0lx8Bw8vn+8xqNGFumZSy4QICQb440qKyGdx9kYOeAgQ20
U3nUwMGd2K59H+8MHQnGeTTmH2R9cTWmN8Oza7AvLEZkHf4ORY+5+Nbdbd3QpEDl3snrVeQaM5O7
qAGK3nJVWAhUYZbGCYUAYWI2kjeH23UGM1DqxfzG4YBWzlo89a9qRTiesTgm9WR4l094hbuMt8wI
KqWOx+UHS9zOqc71K6tgpDDq/s0j3xjEpAXiPeh1YmsoTaAb/hlbptnylUqBRyPNtBJYsDA0Wi2R
KcdJhTQfLOFSi8Oq3jgpGwwapTFP6Gzmf9f5t0430HYA91XcmJCy2vMHukF1XHkEmz9oHpX3N0ca
YtvzA8HMWlvpGwoSaS9qN7KaTNy8rPFEUhwvJDNnWZ60or6I4xzMW0yYHLbK3xl/7Pw9lNQ6TVzV
aTLSpQcz0OuPmUPwqY/MRtSXe0l4Z+GlquKVfPI6Jm3p6h7ZgL2jPnZdj3yjP5LaSk/hv1WJ6fjN
wskIiaxY0+8Eg5BGGuZfBbXxDpgXdm6M7744I+LiiaJhZL3nCUpZjnfGyfO3umZrl8JtHm9tXnuA
VQIMSuwAxHIAdeAg84N85MDHgJzmI8O0UD223uTh/rdkpzzcfsJ8yOv3if6j5Z+A4Mpiz8o6qlZR
CG6pcqd/ua4m4f+hEF3UrE9g6wyQ5Hs919VXXrQRvKusMCYxvht+tVxe7QQ9LRq23ZD783SHl45Y
xGBxMlwAR4BCpwHyldLarOkPLW/F2L+duxoeP/qa0zZgW57rgWQJomHjk+hthYRHN/Nm9vgTmg9g
UrfY7hqmQ9VVxE0Vlwc3JYnEsTb44f7AvZjK+Rm+TEb6ZqtZioi5arjaYVmxvW9XP3dMjSiEG43v
8LmNqztVto62bySISsei0LKGHO6+QaveBOrOkKxFGYOP9CYazLnIAXkPy51lk7bI68xC/a9Z0e7J
O3cf7apkHlF8w8lQmxqbZD8ZuGMzYgPdrs8Tc+g0PlCBwvcz3rRSUNFRRm1rFo0kWJuRzrEdc0nc
k7nA0S0Tvx0E5b7myf4KFtVAmASHQKp+eUWawEgAYsAhL+UCd+GOorMfJZPlViDhaJKlOGwwFFal
S89E8zM6J3Zp4WSzBmNcCbKdKI3whxJLEjwZTSvFGlL9V5QLNyuKDkJWtRpVvY3hE/DtJZgRM3xB
AehXyOeKSiEFWjV948crTcumaGwrY4e6p8TCIMgawSyPMq8Hk/pm0nSZ6LqNoP56XLK7Enpb8HrW
KLAbla7EeQnbIPEZ3b8dkFhaiDOulRK8URKW/DK8Ly5heacEUS6uCkPaMU3WexavYYpt8pQy4WuG
SJ3XB0x5RKxuT3oGvOcSpU8r68j2sdeLCf++N2UsTvSsixbf6C94kz1afvgulTIGqc1rdvrk4iBw
7uwbOlTpoKw5jj7nUUFSjvHZBiZJm4WcDM+e1HtKjKkSp7sN9qTRiFxWxhhMrWnxP9Wv+t6M8Wph
z/rNQBvK1/PKMPOtYAs0twG0IKfsJt0uJtgoj1pYtNvwzRS0OO6FMznR1nT/O6THBRJ8KoU4NZmE
CesGtBCqbU5EGoqHFN9NDSlylpvoAiOxTkww+PVELK7fLaGFPxNmOgGtjGRDyKDw78tCbtgExing
SLP1aS5FMe2iLPrs9udYWQAYvHVGF85uAWItonH8uiuzGPuGyJMnEFQqUEV9Zb7cAH91NgwhdSXN
dnf/7cEhDc4Gi4jABTo+G2+Jo+HBWE9VNej5hCjrz3gaoYSTGUdW2lMo1kBSciOhlTh/V9Mno65W
i9v5e9b9k7v2bm4MVXTwQPgJDyUKgNimiSdaBPgKj/OrY0RXhFLLZ1rmY6KhHF4E6dV2cVdGessV
AppJ5gRNr/ZLv6RpvK0hAuy1+Guzwukt3gJSCiWAZKheIs42oYRKrrQhcbPTsIpY1uyFOYh7tbBT
+M/6XI9li6GZs0ndmC/0jPQi+EOBLGDLrsiUklykSPI07ZOhzH7lVXFvIZLhnM8qpAPOiZ6ruYmG
aEJp4+GTSQ/AnpNuZOp1pK9m0JWNhbGDEQ6h/AqgJj7wTw9jafsKkOmoV4y9dsQvpEnWs2swuBkv
AoNtTbpIeaSAM4Pyj/34GYl3lybFe1jOlVABNLdyJIqgXSQAtH6kf2TFhpiJ9LcjEgR1hToDTpJH
fvIeJQxG1IvfEtRvMUTJ3uo02UjsVolUS/b/woSA+rL181Ne4G0n1nj0fuhbkr24P0dlXwJAUulW
vWqm3E9m+amr6fU/43urlFRk1AImtezEOVv+HphsG+IOQbfolO4+X3KTyYpvl0Blvh9EGyqhPOlD
nYUqA+7EpCIpHfhzTUabVr4NE1sn2936+36iZrXQtmD8kswyt3oHCIlH4q471NVN70jRU4DZ1iU/
/wXgevaTXE2domBhrH1DU4ZSqpasfiNTXMiENQ3bajYqdshWwui6PBtTF/gMoUlJV9lMltLY/V84
E8HQXsTfjY1pQdmx8GoFm5cHfQEgxCy10L1yuWcx68ZjycGC4O1vbXPs2e2b05skx4xeXxVcKY7w
icdArGTxmVCRo66/e9SmRHx2ew93T3wctjk9Y8QCGJ3JLktP1pzXnqwgL9qfRzwDablSIbrwYboc
ZQaoAaJ6vSesBK22XIYd85WCnff9/uTDrrvfqJxvb9Jb7toHYN8CiaJzDZn19JqMuVnzMrfR3vCC
Jy7HXIACOyYnTF+zB6LnVGvAG6PyNKYbnXK2CwBBj99GXpHWG7AllRda1wRGrDLESBMOOSg/f4lX
kXmLS9/r/6F1VXHDraq4AkM/gNUNNDP/dsUmRUeuv8cW81knlvQBqL43o8qeOZogn6C1TFtfg3il
fBrHENAIYxzEI0/5JPhEkPkK1SIKhlMxR7ilDXjccn6FMcfvpVdr0MgSBAPIs2ixTSieFCKXi4JZ
u/Y6W0OSoO3F449GeI7HPyVEtYYfMBb8Mc47BA8mbgIA82C7W057vy5Ggh/Wgws+RG6QncM7CLgE
Q8ajV+gkT4Om7QklYqQ/j13N9rKlalRnwqnkmwd8MfDiZOX1KpnrP+/jRufuggc8HAEmHHKQa9Nq
UmwnB4v+ntXtPELSKFrrvB4AERyGQvcw94ZAkJk6x/bS1NfNVBvmsFx9H/c/MFnmuIDDMn3Hi/TL
dUkAJNbbK0KYJ93kYmvNwbsdBdmd7gDhn/Xgz8HYpGBCbpxMg3sEexe8vkMVnQv9w6bXLnb6L9vh
zGugibfV1IZMu1MQRrj+rdh3b/UQbkRmA7MbOlxEWqkP6roCslXaVvxNLlP50xtPfBSMrxqgLEqQ
1/M0WucVHQ0MgZDfhxFee9V0bXevwbzPAg4XRs152ybqWqIg1G37f2M2ZXxqNXlVSX87ZKtmWM4H
g/BkMPr/+zhkEzuzprWm9Y1+oFxDH0NEpsqW3eGxHVdorbAE81wN3nm78O8C2569NyyfojEby1aI
w1U49PNdQCQblcGJHx3ylTSGjMwu+r4LBaULfTFaPg/+cUgCFM3XObKqt2vIXQ+IQ9xcKFFJWj9M
vQBTkGSpNW1t7gaHz8Q3lOFzwZRVJ5K3auJ9hVDUT46ckCgAnIAh0Xj+O0cg/mWeC+bx/2dNRd31
kXGlm0zI1xiA141FvVt9sAK/9FWB0f/TeoWycXfRhc2XcJTMdXcCESrS5b+cBgP0KfYhycYk7AmE
t3liDQjQ9dqFNvofRa/BPXt2jEIqmmyq8Q/jAahgLFPOf2Te352L9mwF1qiei3Mu9onCw65owpY0
/2tLyUeVPz6KpQzuzraddpWqClIo/+3+fPMHyRqjDN5F3Cj4t60vCVbvjxQFaJsJUS3UspG6I/25
S2zEjIg/g6pgRXnmyxive9MInmA/aMZgB7ofeV//NtaeXNbKvrF+KY/WE9mplkSuK2ybnCkK0LsH
LCMpzkQXoG08EmGafXiY9OJw1PJOpPu8LFL9nkCV8bASkOSw/bgCHSL6deJb3SyBFaBxrp2h9ATp
8MZdF/tFWG0/UaCpEJUKsxjwU7ByOCfwmaVrL82YJQm+3+WGyK8DyLSWZ8rahnKQ8Bf+9f6i5pfw
gglg3RX9KHZh9a0Yx+oSaNifKmqr9ufMY/iuvAkX6LUL3KZwJnIfKyeluPPlJQ+lyBzYVJVH7Ida
3hgmNfoZbDu4eD9gD5IX81j1eZxAz8kLmpvilcGABtqEEQSrviWfasBRr3SU4AGBLWbGu7gTdJmf
JJYTCyJBkUCOix8/kR4P/kYClckRgf5WoNUylXfJJDYRP0i6urDLGeVCwhF2cTgaDBrREHbay29I
Lar9aOm3tjdw9aJiIaX13DBYQTFVvW0Vjg/tV1R491ew8tUOpZNEKkqqlpY13h/fdsUQ541/vAEY
vMZY4TAzffbu5b3IUVNtZIblemmjZPiGzFVhUN2xvfNIhUb5Ku/OPDIYH/kY5OgfwCpASd+Pk3Lv
+pB4fYcTUswGh/Pr1TjaLbdDolKsTj+Y4carmspbrY0KZxujKhlHBLnZDhr5sD7Odpwlk2aX56n8
SrZlPlQcXUjuDjNzi5fKE/CMGXC7rUrrz7kaUo1l9Dog2oK/pcf8OacrSimXwEaQeD2aMU80nv7b
boW1M2d4SU2r4x8X8+TDXbNDllNhZuTfRuTGJMeiplJTELyyHuGoJrpBe7q0d8C24w5zfKKmAVhH
5IYBzjYVAwacRG4svbpYUEL5ZFfm7iDhXjYl2Oc4llABVftJ3ZNAXp12LmcNWury7ZXMfjbM6ACS
Ydj/CbvdQAoU48/qmam0mMNVJg8QHLyx+nzvCbDbmHD24QqX4NfN7/0TB3oZC+2ewqOsYO+fCmRU
AoYy1nGszh9Qq8ALttSPfGgKfs6ZNbgTrm7oh3B08qq8cu1qxxMNPhCDyxlIlSs4VeKF3EnQNQ/3
ICQEl2/yS2B2r6a+iT7/+9KkvRJHbRcy3IO2ufC5wSZJQp0yCctfkygYrVF16v9SGQ7b/LzpMXpb
5OHdLNarLKcUx2lhkpF/NqMtW3o/kp+5Ni8YYOspEDloA6mcEdswb09cYhQiukqGK2rGFdOAFzMo
aISt+BjxNlZ46EF/M/qy2/IE+Lj6UmLjniYHpqy+Bt2DDiqk1XyBBXD4Ut3+tuMMlzdvvX/+43Vl
FmgVH9ah1oAXxx1Cg2HBxhBQOlapYRog9sLmD+w+GxxBhTCWc1KnOa0vYb14GVgXjdSfcxi/abqu
xS6QEtaaimaj0nzFMAKtYKiExxaEAWIZ7koEEmH4llGvrVzI9HUQSvpSZGziU/IXjbM/WLTrdXFM
EXFFCIBHGPDBwlds+put5ZB0xLDecMSpJuPWIYv5Ny523TIIocOKZLzgILAO6ciyCvMAkWAduowj
8w5SCXgUcoBI9J4Lri9WMZ9a/+Haq20nxJ6MpTjWJQXg5TFmysMJ8tSHSLCo5g/UQUIFI5BPJ6RL
zeO/EemMEHeAovc0evxxjIlbULXYK6cu0e87ipBDlw+QwPDAsoEZYz887tttJOS7FN2PIpM+8uRO
QANY2VhrKZZqO0hHYuEbHZb+KRQBTFVaVZqHFywGetR9k+QrUjYjRbuWpl0tKLEpia+2hU40l4JT
Pz5lPWKAO2nk05s9nEjEr76z5DZEs4aZgHexzvoLkawGTb/2s6UsFGse9JrO4BgFFwqyqJz0oM4g
wZEM8wCET83ZRs05WrvDpUq1sWWwHfv5AxVSrUFKD1Iw7zLi7Yefkwa1gVJh3O064i7JZ3JWqpmI
7RLqsUmYWkegEINmsMr021yNtezmi+qYQykaRBO67Wal6fD9fDxQPc0oYoSEk73r/Cndfq5+ro/W
mvNYRY6qYksKMp13h70GXsBXGVq8l+bBP0CCyAxOsHLzmMj4f9g+fz8y5EOP8GyJdDyHE6Lxjru/
QDxvxV/V7fHja9Dpc7LwQ/NMhahg7eStpPSKjTNLyswNolQ9xJ0xvObP2UpSRGH/lyqvOcJ+P5bN
MzQWzVdTECh1vBhiXLOEQMO12n/2nFo+drLTccqSMKI5WtNUkiNgjOMKsqyQLq5myfEb0tZrLOGU
cgm+epFc8V5qnVyr6ozRmGD3YBH3RBEqzc0CuoJf3XfClrecI+RY1QxCZgXgKLiCeYc9xTVvJ+dd
qk5XBkWg3PhG5w1N3DTPYofwR160Ii0801bueXGGqJjmd9KicjhlzbSeH21782AmuPc1UIw18oP0
H3atPDBzeay0nBk1fBfCGCaVN8cKytao1cAB5mBgvawRZ3E61kMrDsNP+vh91eact5eHv63eJSp4
6aYH9VqbiQy0eBAnh0Jj4UoQAxR8UWzkhu7/nIPQDO6hzhCp4TTAhP5TyTnv+Gekts9uG364VYrX
0U4mwuAw9SDP7x5T3LwCJKW/nvbbZXkU4LcKPi9WO2uo3rEZYLpkV/AEcpa1GJZare76wfppMFxr
GY89MlBVOIqgSPmVz6KKDKG9QroGjDNSdR803ljJ39M5KAfPgOdV2hAfpmPwaJP9T+KS7K81y/JE
S6JHCa6EN0rZeQFDlJvaJ2ba//vTvC9V/VQo6tEPtrXCqr3iD8UShEboFsvB2XSp8ot4swGMYM6m
231ctzTWEXaMqmZsBjsUAmEKMy369qBZB2aJEb5GYN5D1MSoRLOjSIweRjJ5u55/jhR7pqTuIKU2
l7HJc2OdoAk0mWMUzNprAuQ12ZvIArhMV0nJOgpAEjyhax2X3TPgI8NqP06GDN4ZO0XGOlMckBnF
5HsXQiSWWTD4N7h9g03jpoU46SbGgUHutX8EaoFSQEfNhdpjRy84nOWfOUPchugyYreZF7JMOiUN
fmYgaU4CMJynsM/DrOXeFvcOx9KFs/ATPK/et00SyXRBKcvUcAQK4LpucUPVUAoPZMmtLlimENiv
wFU/q94r4fEyKfU58ZNGA0m4UoBCE8QENrq5wWXjnUpTfoQrFrI+9llJZ3eS0fN9RbFoGDUQY5/3
aLrO6mGAvQXa9WnADcmBqeTbTsJIpEM2pCpzkkGfoRvv6QHjDjdy+ZaFPbZB7WKgHuzATMfNCWbM
wMB9Ue+fK+qMlMHJUDjHMahhVYEFLKMdUuBrK3YGuI6J7WoY7vO6pv+zAoSiydO+sO+z/DjpvWHQ
jTJexSKlJQbl0fXr34FHzcCFkOjVEbN5cFgpfEVW7fFY1naYLW3S/FzbU7grvgNO+T6aXAuP+SJZ
lN/JH17EzXfetXRIElTLW6Uo3aKJZ6iIfnqyT2WAT631ivpaVI95Cd1kkfbLmjVPdrDTCnX8devz
zRKH0AN+gUrVYRtULdlEWbkyk2GDxIo84oPVyA8J76nShjLOLDiGbMHW8EUz5Ngyja3809fpOye2
Bv3S5Ay0yadqJ53i4hdlmyh2Jev05U/TGF5S+V1gPFI5TUudebz/cSZgF1s+qBkm/dJxdwDrXb9T
ZsshfVEJ1Xyt/OLtTMgUnxdqTLq2vMLPGFPk5f3M2brgl/mIU+DItw7SIkO0Nsxu4eEcjHy1LobF
A1NB5Rr9XqNhcChjgtZXT3ZxYA/By7slKT2ktY8iRI0WsSSQ/TYm3tT9+irwnP/qKG9GYNOPEEb2
Hes9k+8XFIEfr5zZ+iCO5qOKEZqNjO4TpThX1IFqJiEtoTP07UX4XmVtexJRBEW4wxGe0mDL058E
nMZROweaKZ59HqG8P0jgiZ/a7Gm59PPjGFYkEsz2W5OLIjCDycKQzfLdvAETjf5a/zbfK092rPg+
00YrmqfYO0rffvcplVCw1N0F/xDpWy0bQ5v81rz1wNwsn4OaWZQxh3YYE6q4WxPWPKtywQdClGBi
9TuCvUYf1ViSitG4FOgi952/rV7ecBa4VhhMlm9pkr6Dw4WHNwVmC+at4go8KI9MCxCfWy9aDTZt
L5CPfTTDg2tzhMgKLU3cTx4eAmNjL7XdDQ5H/anoalqt0Pd5vt3pte/7lX8EkSDSK9VVYH+H0zDc
B7fgsmtYKarYZ8feGjTEo/ytqw8GQ8vORchboUO619EbtymUJOTvOjdQcS9zpztAF0YoK8WBajD5
3Ql0bS1FRfxiLs1NGLopNcWW9gOwrO28pJ0I7LFQZZxGfcpyBoLvU7LMJfC7FUqvDBNryrynrMT0
mr8CV6IhPJO56myC0vUMbn4HbF5YmfSlDJus9t0CWYR6k+loCFbXfeTwt5smYhCPPMFA2ptV9hXj
wIHNE2XqdgEEgqPL2QJT74HVCQnd+5pc+TXvnQYwty4IrsT6YMBxbhixo6AvAsNqleoOGQ28oGJd
mdPc1NgtIbXb5z74Y77tMrCDNCmVCWP9JzDX1ygmCb7F/bTUGl95FAWmbvfAnxxmrdgrjT4Nm0nG
90bt+bntFGPTGQJlcyxP4VkL1xFcEzb7hg6nMQbiLsDna0BQIBFEUDohIWA/5eccZeSaKboptXA4
N5N2rHcrWvnunCQpMlSEm3ZW0TyrO0skzEAKso+GMqeLKlFi9RLcobdErqeiE7XjkjDri3NDHEUm
s/ywtBhzL9woXRYe42rQEwSsXg62Agg4LdTPOxVfd6nKBkwUbOd6eO7cioQdpXpExXNrKUZbcgPJ
y7pupGUNg6BoUW90Q2mRTYLHO8iOeZpawhV8gdjBmLzeQ+xl6etb4ZPGOZ1U2NgF5fXxwimai5x8
9Y1vPIPhQ88rNK5c/O/pc1wJhQW3V8ysCfcDTjqZ8DfEntaU/iE+J79yHQW+Mt4fQ/w6+OyZb/yZ
308GwViSnftM2FwD0HMSUA0IMOjkoA0EkDtEHTLbb8sKHUTCNjWpxZWJnSTzq5dmHmgQ6wwfxBpI
MxgKDr+55RcC7AxGhxiNaM2zmMwakEzRRbkKgmBZ4MG24G0Y2rX8Fup/3RLEqmgem8bxa2Eqiu5P
E4E38w2sjW0qmF/mrtDupwoOi1i3lJKAcxmy9FSk+cbU1C7GnZChURJJsUeVUk5j1T3D/dMJEPhT
LPuOXyp4Ubvpl/Xggrl+b9JvpOdsapiYcdLNJbO6vjJVRskryytFG3gEktmeQDTjYi1B+gNqiPUT
moCiYyEai4TCEBmEnbLkjEqd7TnxqkqPYRFhi0oVyg38xc1CkkKy2jSb8RtQCdzCKjFfQOsJC5oN
KgDv4QfkFK6r++bzJf3I+qAgURvPFu5IrTTIVr/TLpNWTDg5uOHFa3MIFhXBbofHJwBaKHeoYbGQ
WcD8ZfUNjdsQyaRdavMmrn06lNYjOI+E9NkQthxgeFJfxT28OQo/1sLpXm+Qz11LgvWaHmnoTf/j
McKgRR24SfzcnmU9GKHLTOcbA04kf/f285TBqoNZDY8IZKbDx7c8S8jYqE5XUrfpbXcqyjrLzyfC
Fc1snJMQqfpkXN6K+c6C3UYFj5CebAv5qsfrr/5bu9MnrzKVZdlzxdDBhmhChdMT235UztHF4WaV
Jg1ABFVNsRskACVIFXPJfdIN50wjtQf5pDSbnRLvZsIEZjv5c1n8psz7rGzh0gPDb2xICfQucqGl
Gc86i3QP8ZaEHlykGF72FqgKD4W8jqqzDf0E9cY3fgzk7bHqhNHWC/huaTuwXwiU7Qy4pJkoIvFu
hmKwlidUfICHKbAvSbgiv3WF0mBEmTqSIEQRs8rquXl32OJLP8f0nyVgFskKgCWqVWqXT6PVtGlG
8iefN6+Z17a12feS77doHjFoDYJEi1ZuSQUmJihOWg9n5gzKGwGeZgp3wFAQfqzIY8OMxtTuKvEH
z5qh3mP+49LwRWxVDZhqdsmYJCQbKy7GMBo+S2WbV+KbuihS0S4573tS6+vgxzg3OlX78Cy2bm9m
x5+O9XuMhYgjPZ3gha8GKEJjyzKqAkckgG5FEWO5DEEX1db9+atMAZ/IUBAUhz9OClaNJ/DU88bl
QJZjzCTYCGC9VAFECcUWTQQSM7dxgf1g6YpapcH/50lpn2T0o3ZGpmjbaGQuQwDIb/Lg8ruV0GbL
akjDq7Mg14cFAHnhCbpB8V2dcjqwD1+d/ZOmI2tC2F+iQ35a6rm7jRZoWOdNsbMyVTSCMKi66z0k
dY3tCNOgJEr6jnaYgiv30LJWS3jAIdEdSV4wOFZZvKrtrot5LDVe7G4/W7/5naCJfbd0sJiVqrDL
D2dEVKO1hptxb4eWH4N27HXBQmeHB3Z/D6sHRYZrbhOby9sw+UjcfhGYu73f7LkluFS/f+p1o19L
oGWmEbNgM/Dflwl37zfE+iXwX1Sxmeiav/1YB9Ldzrn59bAbiLN1aQxFtmCiQZZhv2g1nMV1m/2C
0ueconi8SoW4Cr96gzonizQaeIZmCDl5E7nSXx0mJF/uP5y8r+aFJPN3Uj9t4SYkgJijz0UPx0od
Mt19KmhfIc6CXdIwwGB7GKWjOGfT7hAVYdb+77924woTSCLOmftXXEIQe9nmXcmZmLLVOZbL1+Dk
g7dqFka2o4oDzRFHlgQv+nJuH+kwQIzs//L2C+Z6L7aRtTr5KjY5O382Kj204+zo3/lM0zHv+vP9
2m7jeGdp0WQk+ReX/KuNvi01w4kRS7EE/35tkbwoXX8OS17ZFSvJBCwsEm8rzfY1IFDjNGvZxspz
/NW7EbgHN/PYCmoRcDzXHmNk4tbN18ynVaoPICDhT8Eux/xXvE1f2AzfnktFp+Tzarbs0I+L39hu
EMLkxZ6cZs1oLkeQXbVuWhqQ5INQfAALtCPONzVay422UGRmJmqhFAfCG88LoxGx1OIe6wtR2F7l
6c5eNL5e0nfHdWYGmhqGDIj2RajC5X+duwnnxW0T8JDAQwMLPOLghmKpAH+M3ETa/vLwLzzB0OS/
O9oSlYTX4cZPnLnFYREw6Zfa1+r6cmWYRd5o4mmA4yexnjh6gUFhhcPuj6v7OJpHm9A1KzIuhDx1
xRVBagBMjzgyanPZJKOWrig12gf+PwsWPSOvZzFRZu97QyAtqXiIbyZNJwO24vrvS0pWmGS2igtT
4czOouHApdMMZ1DVkYP2n4g1iesUXOD+4fydYHCiZTOJU8/WGnA91ojJ2ahqmj+ab4nRcB93ihn/
rmBqaucf0WgHFkyWgzL2fyNtCH5Y8aCN3TCdDWSy45cns4q/JMFTe/MhLySEwJV+U+Jt8TGUeKUx
80Qs9kbYHllHlPreTwZwndFicDZJxhCJCcBnNX0xx0WULUrd8TeBIoxAmv+qfdsj8ak3PoSL8+qq
gq1av7kgOJM/6516+om8OoX1MPoPofmAK1kEsb+phUeAz9Huify+SgufBujfGsCLEKRqz6uZlyxL
wB8ck9T7waK55YOKmceKi7cnpaTsMsgBbZGjtmVHOMMEpPySqJqMZxXqhQMaiJ1QvVb7loZYSUnr
VJ0YfIXnUMsrxzcmb8kudbkB45GC5Ot+72uefgprx/5qqCHROKeU1stGTptfRv+oRbrhER9pfXed
o8XIDyflOBLBGhouG3a4kvGsq63xa0m4CLImT5d4CBaq4aVj+uQCvJjwC2YyTMakYCyt9oxK6Si3
Eo7vQoJ+nNyHMpW93rXrV+sF0BDcfaJHjLAq2TaCmpDzGF+WKYWb0y20/hk3ZoloM1cCKtmIa/MT
DKRq78yf5eP4+ep+khmzflF84ynJQSlFGG9xNGZ6jR2xqvmtF+nyWpOc3Gqbgt7Pabi7ZzPPL/Dp
+7pCbhf1c8pcUdYXcfQ5oL3j3nBXL4MS0HTA5rthZQPwhNpMAEsx5KrYJulMAB5r324xq0ndBNCC
ZB9OJkgMr1SoNeT9kFXuDxuRzgnmSOtgGwImZR/k+X+BTnvVum1fgX91PnO69HJcX3cE7wFDB6Ld
pbWTpZcX6sp1zh2wPHgDEPRRLe+xzE8f+s+nceD+tuGMv27qdb2S9i7DX4riNwHng7xp+BY9aYAi
4daim6KXnOedkmDXTb8eDP1pFnib/bwENqSCa24ucitUXX+dsI3qeCgbDXKOSicoMWNFiIjv0/qK
Cb8i9M+gzA73hBPCmIbc48uDJ+diYD2hZV/iYCpSodFjLCbRlklpi5hxZZSUxt5o/k3tteuqq8Vw
w8+A8h5jj7eezf2uBgwbblZxDZLauDw8rjUBXb/FT/Ha5L0zWHm/A01u2gHuDdTEf02vuob84lDa
95oVu/WYW0rns9EtJJnpZsCvZrjmF11MDTRKSKmxlLiWaswYkvq8irEIENVBmYXPC7UfVWc9DqLo
d8TjxohJf9lPKQOmkFssVNytYuaTqT8zsjkWUjUFmSWuotX8ZFw8Ibnlt2wkCqTPumKSYKMfqFtD
0f6mjCd8PeW2T5xdlqkLbaIW4WPQlaD29krH8W0PSCtIJTjV90rb6h3nWsv8Bh5rXTasda1U2ksJ
WwE/1r40tFIZbn4l3SwmJLFxQ3NCX3AN8jx0zSJZfYQa6FxICxQMMlXlCyLvCwSZ8HG6OwIwqqtT
HUk/2RPc1CZeWKwrRL6TwGmsDnleNEHOopUm6Qrg05Ce9t1Ik4si87RpRRnBwbukWR2ZroBnV9+x
sUQxJ9felAAJHICAIoEgDME0sE3as7OMUgH7CltkKljI+OmKDsJYMec1EXyTL+bEhCnYELEzMNuV
pKPVmSDzKQaUYvKCUAXrJ1HoRJDx29ck7OtPGgu3qngFELlDhuJFaq7hopum1j36p6Lx60Jnz/8c
QUjtMMQa75wpuT+6Xh3He303KINFBwdt6sjmz7xJFnook2qFBx6SYNbH1SecWG4nEZqNXdqs5baE
Ema9R2IFGL4TcW4EqfcQzoJvf9llWVV5K1LHZf38cwJX/YYKuYMXcsiVCaQofusgVdJ/pqZ6PoJe
CKhDeb7Vrg+YvwboivHd7j4ApfKQMG27p1DJXHBixn/wRaVpsqD61ttykBcJ9v1L2QSRAvKqmTAr
ocrg4fNfqLvgmJwmfH22udGZN2VfMsAeX10WPdQ6+XrsW2Zz5ETC9id2oIh5Lha3p3rYUtbOM9fZ
bMLgYQfQRFE6F18t/JUdokjBoL8kwD0ytfdsiQL0CO4Q5rrWARNd12z9X7cTu8jgmX6xX7EyBs8J
8IkTdPhDPGblixxexuHria+PUVQwb0epwWwSrgkr+QNLxR9k3DLRqhmbOoHrMKgyZtNCR3DZYQlx
y9PlhO9Dx2iW+woquwQxhCnsjbruxicM+cVg0D3CpjSKuk4RY36GQ3aJFdWAG2+lDX81cr73cGw3
vaF+FgvPIJE51pzwNV20NmhauubWjL2yO5aQW1bjj+0XHXADhbOjSeW6RdLzCSFBfQgFWxP9b2+v
rBeSOzB4gAqjcwCSht5U9kOnMJTcek/m2QVnHUq7SE4qBHNFktR41zQQnPiSh0z+A4XQ302+9wa5
h3Ry+Y/7VnKDPpfQY4g+7rT9wr6t53pVbjJ5Xa4fagRnMkZ+smkgHTnHr5sUuff6wIUNylBk6wC4
UZnxBls/qXRueijYTiPD88wbGDBOfMJjVpsRpAeVn550GxauOOP9S/Bkoh49zOrdDTsuIBWLWEcL
tc5DFWNB04JyIOBIYimZZ65GL1KtXiiriPO9wu+Nm22bf5XueyC769hPxniHRfElJd4aMWkrEUGS
Xhs6gOiL9URyzsxbAUNZ/9Hs+nxdAtsxt3D78eo14MFHcWTKRfxZKB2J9UHhe4gF0fU6Yoo3lgyE
3gSSfo3WTDnyKP0ow8hoh7D+Ch7COVRV9NgISXhaawFJo820PYprXNbI03SXWeJItB4XDKQUhzll
zc52LkS1ZkOe6JVQLkgaeFkC1LwyMaqaUcBpWrfK6EgxFJ+WUVr+kGLIO0ZeIlRt8f5NZ8/S6xbz
MGvuTiOGb4HucFAUYNR5wMin5/JvR8kZJHf3BWrQDdEQ7cLQl+84vHw9UdxLwfAtjgS1H1NAilr/
j0fONHE5ATc6c1UGxO0pcjtzUWIT9lbwUVku0uiwQi+ed8zHVm974GrUUCTS66aj1V1lM9cAldyb
GrQV3vc/SNBTcHcJPysxV7ydHCQF/w0Q29gxUIGTTcVFd+FdeM6Khze3KbyGQCGccNV4+KPig4Ev
hmMNJP7zKSfBsq4hbY7XR6etE9BkzVdgeyC78lrHVJb1OmtPzzvk8Pdh20WuDSLbOhiNRxwFY/6I
dE01wPe3xbFvqJl9kWkFOd4vqaIffPs0AjRDOlHo0IKoNDKAJbR9wzcCT4K1N9+bt5pn2gk+p0zF
DJtoZZI5xMUWHRbetCVBPBloR5h3YjDTvVdvRoLvgPvZEvvvIV3dt8334qQKFJ8GcC+aIng4hJPp
2SYEDznH11Vm2XukYf9qk8/4lwg/iur3UBxMQ+bAE6d3gkQY0ByDaxc/+xmzGIuEhsEy/x8smv2r
VaiuQKbhxKRNZxuNxlXOPJ0bpBhKLR08fRH62h8FzXOxRdHp0D3B6ovVU+OA+Q3nYbWDWzfjJRx+
Hljuls9tG31fGlCl1s1q7SDkcqeuhXaaJ4K8iF5E9/ydxdUfjr+NFF/tpNGUKuRcVtKczOkK52WV
g1zF+yzWAx/Y7MxfjkiIkjm+KRlEP7I9ECKQuleuq/Se55sDZsJ1+GmonWG3p3iK/PtjXz6GL+t+
YoR1oskMUXtnHpOTmwlbosBR3EvqIxZQxKtjNnR081kckwFUIYNQ5DNRovW85GZ2uDuzfzJDLG0M
CuStLXy9umJcdXpfv6xX5VovQH64X4aPTZ+R9po4pwP7H4Af1FA7GgeCuqJWnepsJDrRQY1hPYt1
hR9TcH2o0Av9jt6yZYiCrHbq2sv4uuLj9e1/gA2x7TT1XXBud52vAw+vI2+ckQCsoKAMffNoC4E/
WA5PR5WhJHtn+8JxnxpmZMzRjBhS0kHWofcm02zQwb6VQVr6AEpeWeKo8FGyN0/nynlNit27XCWi
iTtQDdI2Sm7FrS2CkkZdBpcjUiVLaXLTsN4xgC+hI6S/2VYwEzP3MT4DpFHcOek4Od/vIju04cJm
t5yLl/j2WltJ2oIhca2MebGs8GVd0ECuQaikaQgjoS+AUm0/IORjm6q+rHgrh+QQZgPx8XcKbjmN
Xpp8o4OhUChxri8CDDs0GP5/6C6BOKe3SAtuFA6XYKTYvMIl31COn9uAzqDXqTEzeCnxqiRo998a
9D0qwQwnxPdkG4bYYFLtRv59VbHLt6+81PHWdF/8LAWWXoEpoHxfDw4JS6Tyf9uTjJyw6FsDpBgR
DW4qy0fFVYamvlYbBUCPN6fcNRAtS/nU9WaTH4Vy2c1XuvSWmOn9boK1Bo40JZBskwBeO3xeLzgD
IPd0/BU2SPJuf5bqm1pMWvasPtkDTLd/WMkXVCWs4ANgm9GKxNSNg3WrcWE1pI9Itfk8WBVsgEHM
Mvt7bOtD9/ASxA9ut+LMmSrXPPuwzNhNvP41Tg6owqqfu7ULz633M6m+TDvvUyOLa61zSGdyRmK6
IE/qxNdzC5aqiUxNvBXLhzyrnVRparhvn0fU0cqdk3O1wgpMJoGVLz+xPZnYvBPYUfp/lTHunkHc
+mHDpreobjR5vXVPt0g08fCJZg9Xs5gOQZNjYsw6a/sKGmU6Bru2meXBBnbGNp/Dkt9yU5JaTm/N
DhfbiJ/uOehNNVv/tJWQsgmdkedIpL7JRANr4mEE+fFqOIEcaI3rgVc4FFhDDW1NFDbfyJm0p6/m
p2PSranp6SSY5arKhCBzUwCAiHwuXPlWksNSxDSiNLDd99A/lOA+s9p6Xed5MgVMgylSV/L/QOYe
/hzKDQw0JmDtucRjjXOF+XvQL58jWb4yO391pwGTbIoMTaxchYH09FRCOwJ9dLyqwQhZKgJDzGYZ
PJbu2pY9A0xP0/dHhh+1asZmlTvPGpBnGkQGPWeNG0SMHxbRIFOFWmp25qsjMa674QwTuiBZGjV6
V8ZTMTOLEyEivJTOjWhw5EYKbRZrXN9J2wYrQyw/pWXi+CRe1WHsP7z4nc7Z5cCbO0/mq8ae9jwD
VMQH6H6kTEQsAxD/iCaFY6JA3dZ9LYlBZmIMs5WpoR4QYpPDWmNskwz4kMw6zyLxqLH+Ym9Zycv/
8amQ+vzEPDmoW+Os8828lrQ0v5pDN2mCnG2jwyNPKrUmC3jU1sf1qIn6mBNtP5iNrZOns7Ri4n/Z
aoKSBmwAxdyiPKhMzzHOsS36vhHskuVbUtQKUos33sodJtK79Va5I5Sdh5PGV2Bh4+o6uVwETyJ2
sj6t9DVii3sCCmQ+f5mcl+yg3HdZXolhbrCgh6a7rs40xGlxPK4fY3N4VvaL+lXpfYs9m9M17IX8
zZv7m8AU4lqrWwbQPpplDEUvz4zjJL5mtp02NLrb15MShj5mPYUtSWy1dF8pDzy6rjNqaljTZewm
nn8flJjpinsIeQ/NBjGlYdhfXkZtKuHE8iU2W45BDbzkAYycbD7OX4gkFBXmU9A8noob1xW1AFsr
NE0PjrwrwoVOeFyehFH4buuZC2IocNYesV9B/a9J0WGvUp9iWo1zcnqkbBD7CY/w4Szjrc+OlN6c
sHCsBTquI7Bm6gPtFQW1lU4SOX0e7ZUCrMH3/OFUW4gvxCLtyYTLMZ251NarFXJYKxlHCxjcQMaN
364F5y/fX1KnXUOndsThpeGvJWEu4BfKqxvMMbyIpZIkzKSiGDxaIEYRwt6uv+nCBUdj2wxVnyn3
HJr4UEOo7KZsU6F6sAhHsSecpp5od+1aR+TzkHwFZtNSsv1qCxrWmhu/k37RvBI/LKWDhJmuSeYs
Em9sSX+LlGjQ7W+qJ5JumYYyTorAvHcsMn0Nd/2EhPcU5jUa1STraabeZE+UIVGQlDO86UMfLnMB
JOdErbwAyY1Y6EaKeMBCAvngKIRqz0e22HgTt0VgSgkRkuZdl5UWqpgQ640GS5PFZUxzbdHAihng
xd72rYPu0Am+0MwYJscnA+IdgW8XY7+EBtQH3EBmDPpK4KTfRKQmj2KvEXHbiFwkwwo+elKtVQMi
KyBuKcZY7VQTQJig9aUE/4VEItq9eGMtHCkG9kSGYMD27+WwrLuSXUQyGt0aBo9WFwgoT8Py9g8c
Mw5GNnGezE28TyIq566HmQo8xHo0L50zrLo7bmA9HDprYOTZYSvXRHUuCwaJODuPTY+L3KRTvoKJ
jhuaE8sLpiCEfYM1rBNWsJDMHLRbM0vpjetLeUU9+AXLRWGGlkFn9N4DUfyFU5KhlutSbxaAaUxO
TzdSBI5yBGiHbx85784QbNS/CR4lOexfT0hQTMDm1/h8Ao1xHzPopHfAorifoe8oP7B7m821FTLO
YR06rKJX2MMNRTLxjL1gGD5FreaxiRm1NCPvGPIJCYcYMCbn1+Vg58eKix5NC+zby66HrUyZfWdK
OXaXJsCy0C5XcMbd6MXyxUUSK4nqIg3dPoEARJULZn5Cc2egUllPyHPCc5THkiioVl1bZoqvro5t
n1TS9Cnt2dfelZZgp6TrRFNQ3/7u1BcZDvMhjM7Vylc8UHhLTsjeDusm3hOrFu37um5LkIFpP9FX
Nj1ADtwQ7x3m2BWHARJQ9eUWZLMzq8uLNL867J/2iCBDewVWY1I21jI12VChA9PMikjRMBYx65/z
f5jQTjD9VOA5SOzSMCARcxHEAkOBXXd9nzwK8vQMDDmtoctC9B++CybSSdgis6dG4fasyEYprIwH
Mmph7byqn6S9z+GmJmFKkBwP8dEZizPyUsQ5Ryqj/ffzYfh9aqKcCEVDgnd7OwutLM2gKj4xC9IS
GZZlAh/f+RAV+A/iGVQ9dJofxsaAuZ0Kub2//hRJbwVHoZ9BWdA/NE7OgTvnJLQiCCfEJ6B6lh4M
cD5FSl/hNiZbPG8GvoNhQFbHb/T7OedKMH3uPjNYXlAj7VX9qNb8iRQl28Snu1fiYiz9lxaFVYXm
tAmPTYUaV/zRX9h24Ic/MYbdKuiJms1CooSp09LCtEgiaF/8qvLkCEvW4xyOVPUOQ7lLqf7nv3uZ
sduDMMjXzYMDicGnJZkMXuCrwMDENMV4CFRq+Blhae06ijNuI8q/V8Qjj9c41EUqkzJOUgcRPsCT
rXNoMXrx6uCdjVxpP6wrKIWMqlLuU2Oi6Cg++4yMl5zs3qJ7TlzZYu8ra342KqasN7+wMJrduzTM
/rZlIz7+zmNOgRWYJOo2rkE8CzVesZqSLQQQFXvH+qKhJoEsUXCwnjUvwgGYbQ4JkoDTn09Iz1Yc
B2FBosza9aJmjO+MoqO79717/N2BqrYSc83/1cFhsks/iZJoIUt3ywajgoTwh5rZNwF86KzPQOvF
af+7Wft9T1YXwW2ZeVvkZClbBqD5ATH4l5Xm8KLOyYaIYolwT0t/+0sQhc6gNEK14hxQsEwExPms
3A7ULpg7cBuPT1jsTjN6FAcSagXRjEOP5behz7I58aMN99aU43Dr6mg1GMEqNuZqz0+TYulV/BbI
IA+zYO8k5YrSSxWB+Xkq3sS1RA9r1p39WFO3a7n98ElyYE9QChdpMRpY611JwQru+2bfrOdRV1I6
ThCfadEqDrt8OqXaoBNrmhCGvbVqJN7nM93Qpv5iE/zsTDoU2BgLWRv/YVLOq6W4QtnWRYam5otR
x5XVjA+MKmgOz3/5k6AyJbSeVGp5lKZnzvuLt6afmfvizVCsByn/yO/KQroYq11v9bAngY4XTyhF
9nY7697RGaAKtUetub/hpg7vazyYSZEKiogBrJ9qKHT3e4AfkUx+v265efRJLMrJVGkDL/iJIcHQ
5mmX+oH+IMgh6ut7p6S7BF2PuXkFGTS1als/CgIVD1th6h4kH69EqJ5QgLUDKaF9qF3v47CwYbNf
Pcn96eTQQi7xR4bejqoNG41LHEEm8ZaKDU19QAsOToZIMaz/hID4A2fG5zFMBKy6wb/qQugZRCjB
8wpQxmw1Gi8JGapqKJSsNxVtg4+LLKq1IjF7V+Rc7H+bjlw54k1OKwyCeRqDdrFZHl2r4ffZymy5
TMCHRS0rwZE2HcNQ+hduquDMTn+BEpilerAQTwpeupxUnQaFfixo4bXpBcxra1yo8i+IrSCXSGSB
d+6a6/ZJBPHqQeh/P0n/uj2LGENJYepVkiSGaPFNDvB5yK5QzMJQz/4hNOJemDC/+w3ZOYZm50el
kzRJn1sjqLlya7hQQNj76VpYZ3CIcveC0inAxiSaCvIlBUajMMwQysOk2Hr5UbWMDjB8+2TDSGVK
b2VOhHCwb9ZM4XulslHdi14IukLmV+TECyNbU4Z/3/n/l25Vcnb7j15VtzmtE7EWBw3HF7DhNZhZ
RaT6TE8vUeUKwFcHFyyIh+GjSRXKPSlFMzmMgvdt/1+lojflq/TlrjI2DLJ+thWm5r5TqjdlYkDV
fzqGhAuDthVR07UCQqf9VylO1JoVYk9hvQtTfflRlybeEPqOwdQuzS9vzmJaknbyrYAfYWaoq1hI
Zih0OGmjNqSL7hGtCa8uTAY3shRaCbuCUGOvMscShMraZCqHqqr0bIpj2/4uLQkb56gUh+YLMXZ9
q14PvNkK5nCWGCEAJR08v9cmOph38ETsUycpge39aicIjkZMZFnAlfM5nH1+EYQomnIuXHcRcoBC
SkCZXSg7eu2oqcY6NwN6IRGvg+9x2r/+fSO58iyTCn5IvG/HvHj1DRtIO0ie+c0Ml2fSuLPkkVi2
UbM6/rxHLPjMFUYKPB57LLMBc7YaK9rpc5yyuVJIbOfwW7+mr4jg8xhmOJniLS5iRwrVWRYpKtDk
zzbMaKH9SREr4wQGipo0gSYXbJ0ulIYv4AOtPvZPYyKmZ1ZiedAedgiohL4SnRZqmZYJxrwcY/2k
4u5mNLsxInBE+ElEXtDOTuJm7VCOaS9zDIrAasLFQ6HCHRuwpwWdxR0otde0PY9WgNZseOZdKO6B
b5jPm+eFASiVHsijElqIBYYZcjRWcvWJcNL1Ss2mKG8HKrYKdKQWqcd+hhbpxby/QmQIlrU/Zt2p
dxORIOPj4M3Esh34ucV6W7CI1drSYCNwmnSNJ5k6yU/ygC36p6UmUy0zXQoNrbXEp4x638463ZZh
nASaYxx2upc/OmfSHRhQzAPddeZJK+/R904OaggPRQQT4+tyN3bVFfdGHb1IndWui0WxqyzPs5W9
sBV4UdRxNVtWkntHELOqciH5ugx8k6ktR9V0tLyXNZDMpjCVnBkhE67K4gZ+wpEu/0Pk04TzIJdm
R8Xn1kSNPyaTD5/CBGA4Tcp5czMvs0eQAsDF6M9dBQxSqKjiqbmI8RAQCyDuifvWMIerRCaZ1nX9
49oZLset4J7igpmbe/HtG3gfe8qulR8ZVf8YZlGTRbcjSs5cAdLGi87ATTexTv/6BgUrc9Qtqidn
ksYpkz2ZTx4elF+3nH+n4txISFmvkHAnjBCoAJgUqFRNVxxxlEZD8dzUM4qlKkArnLcpxYT1gOPv
SdhvFF//513teFyGx7Y/nEIBR+5CYZxfMvdZf8XjZzqR/AV5zLNffH5KPTc+O0RURZzZCeeak2KY
StZ9RBLwCTjulxPoP+/+Jexhq96KWLMHCQsCktyBkC5V3KndQYgEaR9Mw8h83k8DZm0CHwF143H4
ZH5BYs/J/MWEmleUMJx2+/XVZW/rA59K3KZPBuvJ9Xa3nNNTbWL5BuMSHppna70ctaB3hXIrkphx
jS80QFwfLkffak5+qJz9uqI+e4X04mfeDY3efjc+sKw2jWYsbDFy4Hnb4P8k0ZR33vFb1Sl3OR4U
PSw6SwsGHQ4hbqVavlPxVfym4rvl3x1TRBYyrMZKHSV6L7q0msDIGuEJtdDGzQ3g01wm7A1hJ9/R
oX0Gwt9lc9Zxqhlmsnngmpltm+hveroBZ2jEbQwQvSfTXRiEMK/PMJsIJy4+WCX2MGFxDhqwvNJn
3fBIXIryINd5MRhwZmm56xgj4bturq4Et0UoR2ng4JnUdNjzp5RhmTZoOx91z3uwI3kxARcEVM7f
3d1vui7lCMQleyTp71WiOkieBhXqkVWIFspxm/kiGWfJuhTor8w+carNNTb1u3Y9Yb/NiFEoxhss
n+frkhV1WZsP4cTLQ25anEXaJF/ACzQWa/JBJg/373BykQCHcJ/WF3omnC2XY5Gs9VZXrM/NdFg6
cEdKgLwl8Mu90uXR+vgUeiTjrj25Ei9TFVQOpo8TMLW2+c/g+XNYV8+q8ax3itifMqxh19U9Rcmt
M1uPdj4kbaSM7Z7E8WVeIz0NWLguf5cGYMN/wHgWimy5aCYrOf2Rwo6i1OJS47ama/Sx/J/m2S0T
Q1AtEdEwrFr/hZ8Uk9mDOZuHfnBkOHoR/psPkQnWNRwDMwuSoHPtxWRoBUacco0ocuZ9E5M1z8Bm
zMzTqtqWWmU+RMj7QpAQDaHF7rEpI9Kwmk6I0+DI6/H8ZXzYyrJ6SNtdkVGEgx3MJejuWYkaaF2w
Jvs99+XMd9KBcabGLuECP+Aw9/yKj47wZZrNuTs/66wcSmAYyd6MkXMJEYVw5SAvKMsjchKCeU2j
1ZSUz8QDuOj3LwN1GeNpxyVILDkNBjCpIf4jyOb1AkD4JF0pTG8C+lizvoYeYmoUJIaPzFmplUb4
MAimIMmp2vWuoxaMxeOZzYqTSMxS+SD+llcbVhqF2511Fh3HDXAWb+b7LIzTXg7CEbzk7h/COrI9
ql44ZwIhk3ORPp6QQDTklN/fcPG5supN1LXXkL4qId7rxKM5NP3WBGG7jqqQJC/IpRTo4Yf801HC
SzemO4zR6IzhwAYw9rKX20OEwTPb5gWfrPb1sGhPi8FXwkwAeIHufdrU6UKiv7fUg56HZk9MRqSJ
fgUlPgjXOyvHRJVtAu49j+MinkXHyZgZGL9siTKNW4Tvecwqh2maOZwLHai9E4eDkdzie4lfIZB5
+uMqnhWjaI10cGcRhmK/2w+6UKRs/E0M7BZxd240vRF6XcQpgQRIf7uYGxGFg/goec5UhNmseDc8
5Xx8C44XA3GCtTCjieru93zvfA3jmemI4vuMup5tAMOd7uqSpRhTFsu3V0u88OZVamJuDCJ7r2Mq
Nd2UBlEGrFGeBJxC3Lo4kLs6W4j7uwBJ+34NnN6hZCyPZSZrgHIw7jSIh7LjcnKleVWNJSFFtTHV
ocizkiFYazjeGdyLLmJtCfzLuwLv9c/5jieXW//SLAf0EGdwWKjAyAs97MM=

`protect end_protected
