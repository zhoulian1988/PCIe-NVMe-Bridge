`protect begin_protected
`protect version=1
`protect encrypt_agent="FMSH Encrypt Tool"
`protect encrypt_agent_info="FMSH Encrypt Version 1.0"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2017_05", key_method="rsa"
`protect key_block
Fe+tViTRi2EVqh/wUAvtwV18wAFQgpfvABMlQvE5VeAqlIo0s2udfdDZfS2CSJCroSp3nj3vFU7s
GIPirwFFTsxZWDcB5l9riIQNL1xdGkJD95N/bVb315KLXS+Gh0IHdlnSM18GgfEiJk6PNi0n7gIq
hGn+H6a4Occ78CSXiFj8yfrTPcPq48fg7Zc1ZdVWpqcNTpu8lrWeNnI992uyNFIrASspTHqR9H3q
0Ceu94T/sJzdTo5tdO05dFFsW8tgbmRuLWo+AQ08ztq//7WMjOJlQQK6O6+/ZIlDd4Kl6q7Q4Jvp
Djh9YzjtD3QYSSdXFwBLA2CB8Fp/0AuntdTW6A==

`protect data_method="aes256-cbc"
`protect encoding=(enctype="base64", line_length=76, bytes=295632)
`protect data_block
feGcSM8E+bzqQMWerQBPnK669rybny8a81d8xRMDAlAB4RbOdHSzqZjSjfLb9KGEi5lIUjwhB2Oh
1x6z39nNZrP3Sr9U/tnKKGbbMkuyZg3jL9cgaUsfFS04lT20VAYb2e/ik10dZPFpKePg1TZgWnF7
esbLGRyxOpFOBLmOcdDIc1tQ0i/YXDJvtmTDtPokXylS21FPsJCmGZqcdlqY9d3T638kPY8HEPIv
8ygV9tWOorj5vgP47xU94WAL2ihHFTZNmbafCGHaaRGX8cQpCOAWew2S8tKXOnSsByXne+8R3cPm
QeKvm43/A9GCpDzUURJNUtm9cQlMvKfUH646Rg1uye7xaiq2CQQ7UwJz/MgmaNOTHPqkhkYUaSk/
UDv/X1vtxqEXdjHo5vqcuAONorKvPDemjtrYMwZXS3PGnRWMaeUW5HvsXJpvuycM6MubY/4TJra8
g9tGwgN7h3Timnl730HI2xxPoImzaPQIE3WW1a8TVV1KJOg6YyJd2IGihN26XfvFqnv4WOhQawBK
dYqgxeRn9lOmu3CiMM3uMmYIPdz/XEULsHmfbDf08HufBXUUN/eKNSWtTTBS/4PYs7fTJAgvuG+C
QV6fRSw2IGywNJQ5D9AeBvk1VlfOCTLB9XOhz2OFPqlaxHJzXkOMNss5QfadmdCwGnr1NPhNIT3F
nQTcqOLPtlbGEb8Be27peelZDsXxbOjg1IHMjBsp3+iqsDgZDK2W/JpvRdswhl5zyWgOdxCEHzkd
33049Wv7bE0r4yNbbygesWdQXaUPXrG+zwIJ175GLYm/MM6ke9iCihyV5ci2a4uHw+lZmS+yjdWL
R7AUm1FjTBr3gBljzJ5bANvVbTg7bSrI7PZsskKEEnmAAIoTfVMJXCSiQVG67R+En9vH+6U8zpPG
rpVIScMcJX78X07w6zN3eCHdGnltUN+t53cT5jIM4WIBO/efzwKnhaqF8dUmKyjgJb0Gk7HqX65B
45ZRKUKbg+C/tm1UruKB8pHtbDC/JcUi5trdCrMx5eUOhJ/t43ZoO33YmjdslCiqdPVxnEfCP8Ds
5+yrZwFLkgC2tLw252PxPWuyLQonuf7dygY6fgiUsCG9Lxz2SBYIk8XIrQolfDD5wvNRd7E5H9R2
voMCdBL6lc3F242vHN3gnPusRRMtkPz5DA7sLnURTxJ7dl7HlxjqSdtGvdJaf4Lk4N1j7L7p6D65
U12VivQYiHwjKDUsz92lpbJjc5G6VlGtvFn9t6wIyPLUzY6ADxlLnF5yY2qX1qMFm16p0NjdL9Tw
yadAKSJ2NxWLp+PSgeAR2gybKEHW6DXOuww9tnR02+m1cBaCNGJJPjtkBFeS8+Akhr838BF5U9bt
dEwVkM0NPcG4AV+VVXQ/KMrKdFwJ77xLIw/SWTZAlKmdjErIOGKSIF91BfHpxSmoJfhqCMsfmUcb
x41m0ElHG+AuZ2qcu601h9jJD5xj6idjAhRMKgP2NcxNwp4xLIm6xj76fYVnDTpbWB24aA+rEx01
q1F4I+vcQfrusTtYsA3w2crMk9q8uRjzaniazf1Pv6g8KbVBDF6X3tCwuq5HEoei29juBrOpq3cJ
ZQJVbloWKwuOPvcp3jAupdF9bATeDwiEQYTgRjWIDDRKUuck0Du/puHT9vOy2mFiaj4WQurjA6KR
yPTXEfM6P+uZocLJxiPxJM4vbn8caekCsjY0lIiHggxvBu3vFvhJYP9bqGLjYisVpmDctCIGZt+o
FxTx72wbKYVF2IYuveWZ6/GEdSvPLOfYFX32UfLzY0RNTuaj1zrJ8gHPjOA7K7lkQCqm8loe60CJ
5IMPdqeqiy3RASAJXjwo32YV6N/j8gj243ihNwSgWHM8FufcxoeOT/VYlFxDQYTm70HsyFQ5ZcVQ
mR1H0TVJEMcR0xPTGWn4qOaMOfP8ASYWSQtpz7jwoP6iTVatNWEJyVb7TNPxXMQSlHAolyo16enZ
unUENuZlvZgDeGFJZOhMIyG4vdMCUcFO8LvtWqXa3Rbm72oV7OyOMVxrGMbTl4ERemwOsGGivJJ4
Z7p6RQDCWqt4SPbhrPaIVg2j5Lyn3bD8LYCqgRv+VKcZeH/092ukruUNpa6HSKOkReY78Ao5bQRq
nMBrAS9OL8Pzs7ogao24d8VxNKflVf9dJ3hLe7rt8gp2FAalYOWyI8+bHXDFqB7ERLKAqA8crwL4
87pFlsRC5JMRV6TBhqipw0HjsBpb/8MU6t0nt8/XdZBOs8tqM8rpTGGbQ13i1aG3USMS2vaBxS9E
e4aAzc8uU+qHfEeqCUyb+W5aqSzdx6f2ehNzkRIvUvjHEGbL4Kpt5T7wgxH3XkZaFqFBc+pdXViw
teNWmmUbrX10fLywYU5Z1w08LvNYyflQtxwrUlw/K9iBlNSdSPlLzOKwxW7WqCOsT3chC57IHUZC
s9pkOirErLMkkF1KnplxyLo4+MGkMje1UUG8HItJHWS/a+G3Zv0r5wh+Q4/u/mvtbcT44DA86Lex
qs3uWRgv7jz7I4pwMPKdC1dH7GU9sBtY9/wRI8gHtLAFDaZNYVomMdlvZTxavB1Af3Uxx+y0juhC
3WY1Q9sjqRbsdyQNU2eDbXl1/xGZAfliiSbkGVUDLo8BG3bL1mqtLia0cmp17PsNw2QqXfqnWr9v
leb1iNeibc/2tyGuIUyJJzfNcxZYAciAJzAZ4pH1BaVafX6zanqWFc+NjEtgsQkkQRnaoRGLqI3t
IX4RcaRoyywnrNAfbx9UWNTdNuR0JUqTQtXmlHK7l7EhQAGTBepT2PX0qrdV3mooYk4ka8rVY7Bk
3Uq+e3SoZAHYmzh4WyY2am6bep2xNaBpyqofSDGOioNEtUWpaDCefTY/Z4ov0FV64HHr3YH/0ej9
Hc69Lrz9+nyxoi1eYtKwag2kqonbME0u5R7IVecPV9V52JawCN+gZAomAjegRoCXLbRqvjBNd/bt
V11efKHNH4XLGgWeTI43eDb3KsKI+4fg5Kqx3Fg07MbLceu22dcPH80pAPOHuidtCf/gpm0MHArZ
e88M/R0bvKfeEdOzL2VUeQRV5gg1zvVKVe3t8KXYMyKnamn+6zs4kPNWKIh7epq/SyfqaMlUrmSf
CASjyn/AD4oRe0zqQx4vmLg4HqcMaDHQ/2Wij8yk3I3oiPVOLRpfnvlzAUBEq0LZ7/O55O4xGmDz
UHRGPk9MFIi1JT7WjAkrS/laHMeYxsyoIB7UFdQJqjSMVA2cjWd6bVekNWATqJFwuXkQ9mfwuOcK
6JyPny8MVv8Sq4Mr49mcfEbG2Iro9sADJjMgNNjE8N1K9rK8Vnt5aejsN4ZMUf+O3sB1Nd8ALvJD
cQcGBQolaGrUFX1hB617+/54Oy1z0ggRRSb1VpaKs9ZdoDyLIOYAoysmKk9tV0qpVGLhFr1+2TIy
G7kWJndf4CXwq0bn2LK/8W7iOixdCpqyBFRtcwAm4ic0oKnW9MIO1IoQkTl+5YTYjkLdyKu/+o7y
49CU0I3dC3u4aQwguUsb3a0yScUaCyj+EEPLKrSJpE+6UC7IVppfVACSxTLNm2YDIQa0+wJNizia
giDuYIpjsczutN3uE+P88f/lw0HEqy1xn/0kSI8PsT63w0Pc8bJj6RvAEcfyWidYEtqMbGc6+IYv
ocZjoCQmgT0jDc/x6CZic3H5u5WDwU5L9GM4GwBZOfcDALbYE+9iq+lGGHscd3dlOHKol3O0wVfl
lJ6OzgNAGVoKnxqeoQAKg2dI6zUPu12OdAbR0xzrtcnoSiItauxe1lXPxHc5sLTwyuD7cueBzU6S
54lSUREt8L64cIGiR5CUhah5d/sA/ef6W+1q6RC3PYxAAQa3zmSx0P8X+l94dr/4je9wz3hmHA4L
suLH/UBYxt9aaCQ5nf2XSgemmb5uUMmfljRW1OwvYZ3pbCKd6UeGso5/hilbknHdCc+z93Dw6prN
6Ho/bPa4fr7Yi/253p7H/CgZkHe7L7k6nGHmaUiAxclD+62TXLMO/ehNwPZEM7FaqfZhqMkttMGC
R2VQOaRgbiOQzUzCjy85zijtCHqg89tn641PmCYTjJGynMr2UeoLxgJ2TlOnC1RTy8ljw/gFGz2p
Mv86coRUTaBQSB0K1wr3K2gWvQDiSrHv1HYE76aH8pfmIYFmIULHo8yhX+2xpysjmLSjyagHpUzS
R0zY5q5nQf2Z3hy8jycf5zkSjXqpVEzs46DiIecuMNux5pugyeCifOO5m22vNw9g9hm6Oo8jTKSg
Un3ArtpgXO+VhVKK4tmox7yClU5cvhBfXepSdlL4bbGPuxKkruehm5KV+XSEJ75qeuUlnA+pBl/f
uw5KHu8P2KGEDqmQYmsOIq/QZc1PYAPW3wYMKLacdRbSOw9GJzjf9wG6Rbc1ZTqv5FV2YkhWEZ//
9rQ2DRDvOkgV1cDUaY+zrlInzW9kn9XdgGyo9lQKTV5P+pbm87cdxSigqFHMay7giKT1h/bBKfDb
19Fz5hbZMcXN6GeUMqcObHyACxfQy1B2etsGpkZtRwyYFHGnm68I8ccvEKk71D5L5XNmVD1osn1I
iwBysyyY3IqXMakyyvQU6bpYosYAppu0m3cnNROcsTbpX+hlK5uup3cJqj7ZmTTfSX/9isFbvfU4
MbHBlIndwlV8cYsGi714qBNiZNm3kiLgvbP24x9vfcvGw4E6zUp8oDct4/7Rf7QDg+SB1DEEr35x
J0wbCRo8/SUMABiYaD/OKVJMgSp3jLMTSMD8fHbG/Nd92HZ47I00WGQ5wz8W27HGuQxOU25tw3vU
0uFE8D+/oa7IT3OAJbCnb7234mzIUcYRUPZTxv1km/V09UXEM5133CkufTbvVhJTiRxT2D96wGo6
noypFdH2OouXhRApL5yv1i+djCTv36qG0zlwUG9xgKT1pWXlD1e5h3igVA63limuqhCYJPqtIIJY
VKhP71nc+bL6VRI3lj4QXhrM2SezJR3eAXh8TEncOr5XNq8EPmnKGnls7HSFuA661wKix8ti4VOI
xBPTHWn26IB7bXH/lxDUHUgDUUaOCE6lhdn5trmZOkxUpmRG5j0OWJcal36sMHI+U+K4/YXX0o7s
tskk2VTMcnatCY2AZhljPIOeAisb1agSOSj828i5Y6xSiPf7f6zI7CffEZ22e57H6UAIIZpJc4YZ
uyfpP/n8xpw2FwY4++/SPXVpEM+BEptEuhPUxjQKGHQFkW+cJJSSo9/M7NpGjiJE1SWZLbMMT1Tr
NDovMmWi8CbfWZcN7APvT1fZZniyB9aZOANneo/Q6zjftyDEyktciqixeucKpOjxfyHRiKkPhRqT
mX7Ynixa+kuZiQxjHw2hR4ab7Mt4v7GOtnhh7/y/QFQTSHkVJjKP+eNnRt/V8y0wlC7r8D3QiZQw
iBQiLOaiEoDP3oW6lJPfwIgjToMkf3O/SG0FDsB/u7mhgbdKLLRHUGQTR6hmliwhHyEWJUY1r4wA
t8GzslmzyN4lviR33hQIS3uqbPGEjMxOXtlcqk38ThZygyb+CaujfurzCOZl88/tzDFqEq/EV1nz
JQ3JSj3No8EIN6It03yD3Zbyf6wZqQlpKGjRsDXDcJ2kVK0JgtgC2mFBs0W7u74ql6Mxgrh70YlR
kmk5K5rB/syIgyhPhWNeifDpg89YEq7dWD6OxkuKiXhEKXzdtEJzImppTe2WmVQuXtUrMDcTvK4X
8zM5U9JyFbmdq+yKRs7P224p1A0vkYh5D2XAo0XnjyIeikJHc2oqxbChdmaqfEirUBJqhs6tHSbW
p5skCu8c92yGE9mKwy1K+2NAaN3lCYxxPnDOX7cCvEb4zecMYbTzI31X4pcW4juQi7PcACSlOa6L
7mDZgesav3uLxA5BkEHNLCkJqdXZ1OyGOn4zIsNlc38tL6yPt4FBKNgDTzjZsX+QycMz6X9ThAQC
DiFGYxOKl2PTjDgzr1OtuapjtgIecMzFUQoyHJrmpmQC/gnE/8YSO9WVh9VNPr0sWGGNvEc8REWg
CY4JFny4WGbX9HbyNTspChkur0IIzSPUTF62HaeAhlnwGEUqwc+6gEPJoKYi3U16XwyL9CEDlzxD
Lbhn33zKpWrSKU7QjR0wEkma3YCp1xqIUcpf03NHtxRjeE0x2vZShz/mkl00BgzXm0raCPStGWI5
Ww2C3SEmvxCbmU+1IgUx3AseCKm9LpcB9HBzqnsST+nJ35Y9DTYSC4UNczzw2QClTwM4GeM3MFIC
s8g8gxbiL12PQlNpk0I7gt7GIrjXdQbf/dz/wL3wPfmQZgXzE29o/CDK1ohzO2qwMA72ebsa45mB
1oJrZYZH40JHOioRxoIqhJMaOq0UUN92mCQyTCFhHDA5YpsZSU/cCnMBYHr+DyFLmh7u+95iBaJv
285dT0fHbNGHoCpW8lc/pORgQp5KG19MHdgUIWn1mNyCR++bW6/OdXLvGbb/KzHJlik8TJuVpGaP
UmlG3CY3Z7uVKsH2Qk9upBlJDabFIHsoh3+W/OErsEk2BvP+bvB9n0Or8nM2DiKEgcaQnUQAojwj
4yB4X1g01SxQod36QSbKznmOwRdP9SGIZDrpGDVJiT4YxduJUQrfPD+hl5sw9hVSeBV2bRbjDCr2
OID3DhDHRhTDHUNk9J94SNlbY57PbZ2fLo3u1t5PaAOqrfxHLuQ0+QfopIAzL937rk7DW7gxqEAA
y8iw71QnWWLSPjDNDDh8SGdnQqjRn3iIOZa0XZ2K5tvA0qrzGPOGWERXj1cHn5sDvQFreuM2bfwf
5wyer4fnmHhR4x+8wDL6hd4+ptHZQdIuKp+xRYX++xc+TocWPIxyBUEz683CdeqN1dexLUvsJ0ij
KFi5r8O/N9cRpQ3byD8JPtPU6nMs92fv3u63kGObPleIYMyhoaqdznJCQFa0ewoIc1C7EEak1aLm
xfr7bK5wZbvnQhs7rt7hkPLUGxzRFLalvPVXA1ibAFZELJDkLw6OzunF3yh1jG/TlJqpn95eQTIe
RH6hohaPwHr/KWw7MUi5bC5keHvnsq7GrlamGVTLtgBPFXge+Sv3N+rOQkeDTEyihUqjVaBvlQWB
O2MTPnquqxMep9aun22gbGpxEYhcfvVnWbwTZsYgJasooW1IOLPLQIn3kDWPXodPx6/3FiEGvfaX
UzcejbFO77dhj2t1NX2+EDb8z+RnA42/5NEQwCHIYyBBeRv/iVohHxHvNYF5ZiY7UjiTHuQ3EzHV
O58gRClHwduMRG1l414xZAtEwH6uBz0hQf97abVuP4mWLJycfGNNjwwy+C3PYulUtQa29VrI7R39
NYsBfJNwMBW42+D7vkXA26hD40ZrznxYzRzSPRtak2cmhP7AeikORG1B08ONh8xRDqcm9ZiSbsDe
w2h9MfvDt9D9zTNHxNDkg5cEF+gzT3UwayzCZ7mE0P7LcXTAOgEg+pfg9XjbVpoY4EVgGLBjXjZg
PsB/P81AI2PlC1DcOdxtaS/b/66RpowehvpwKOTBRAztDjX1vXPvVW/tIOnv6JB167ZXJnvwdvUE
tkNwYx0o72I7t1WzeEqLN+A2X4W4cZnd3EJlkdnRG/VQFUR8bC8GN35YWT9Q7zFXYsMZFr6relPU
YG+z5XyMz0AVYr00xnUlmo7NRz0Q2/9m+nayVhb3g8iZtxXm/baNZPMyq9i+sMszHJsoF0JKKhre
BcYIp2zQezQvWaOktcG+XiHSEP/iF1muwSuhTYO7DUcnuDl6fwcPNqLBolJw8W5YIriW2wEcsKXi
v/lCmUvW5HFS4RSQqKEuqKaMBBwEcNOLqHkc3hwbvRwbhTlWDigfMPNGXRvUAuMq1/4WRmZrJVbI
hkPqO7kSxuN6T/GoEtD/Fa17h7UKZ3nsKifgcwqnxUigJN9CcU4fyIAVI/VVo+vM3K5MH2wcqQmk
m7t4+tynOcjmzxVBOfWRkIgXgXqGnSEsfsHBxF/R6nzWVZ02i4esL1GmLvjh/HNTjwujWNeFD62f
RdDlX4Vo3eYLTsvnTlXEEDASPFZ/y94tjqCupQW06fvULP6zceTQ+7pH7aakJwytRr/aDf58D5nR
weJ7SadfhuLJTPzoUCMAZOyeFiEcRa386twmxmApeh+15/2f+b9Lim+9TQf8NU5PJFaQ0nMoyBBX
jh7Cks27akJh3ES1zFAvRwDHSIlot2ZSKvaedVLenX6UPXmLHQbXEylCVnjOSuI+P6jVvKIHZtj1
hmFXzg8xkClWErmRtNXoVI1s0atksae1B9Io2nrfJTswL9onUPse3AugN/Y8oF10rcKPshtI3zII
FWnNu0i3bRISv5DHn1R3BRdNSbU2xJmm+5EaJMYeRKlDYM0RFh4xRrJaziMCG7mmPAQgkZe8v3Av
ReNZn6Xg9vpfvBObgXOW7rDJS4n1EIB80ai/P3dqMX8+Y4CfZ8vkBAEF9MFnDiLr7TXX7Vesm3uB
Q5xzsGez4vMeVH9Yu1EsQ7GWxGKrlcpvj+a931cZjdeiPhNndAMqlXWJiE+QgAaicyflvu4CyY2k
ljEYQJH1LDdRtl/4IXJrqu+nWkm/e/REol3znnPS5/y4pljsIKT7zi2GXgMgF6pTlqXKJyP3J3t6
/DfN0vnMPFG6oHhN+XR83kGVyJLcI+ZoszlcNVyU6eS/4lgo+1CE1SiAQVy6EVQe587ko36GiX/A
pPCjfItrEhPSbds8h2ZkVYXqWd9AkowTqE6SELpzh94EExtb65kUeK5KUljm5zdjxkUEpgMgeUjp
WluSggdj9x7vHm9u+67SDh68vY2LRm5nhXupTCHEKb7A4AzRZ71k6F9YlwDvN95+7GP7wa4rw8aT
og4ejcYmGENw36ssrfqyWJa+iwolS+h8SZee36c4d0IjZu1/G97Qvm+y/5wgeLmqZC8iUn/qR7ZQ
SEjfJ/ytW6LfW2ItfFU/u/Ix5bc5KOUrkv3hdIG24CCQ5rYAoT963ekfa19lm4v/fqT3SsI7J8fh
+Mk5w8sD+1L/DsSUiNy+8adR19QjvOCw/EoehxfuGB/yqdfaCNpeCQL3s7cdswDc4WkDvE43f+Bf
Y/U+RhHlZj4uZ3W8C6zU+iM/MqY/xSLZYU1rGyH6smrsgWXbm1dDgNveh6XzSAJks/t6w8T/E9Hj
dMElmnMRWM8L/83pWwvZWFPwyJqFXGskouC1yyWqNS/UtmTPoZYFtRn8+rV9ZX2gyhY5M6O5GEwZ
JIbdRAooC3faoGY8MPFRQ50vOX8gso/Ygnxj5WTYXAFfC/RCz4IvrerqW3Va1d19dOWTI1Eiy32l
pi5G1jlMQ4LhSLgSqgJ1u49pyEYG8dmJyAFEOzZemr5Mk1LPmt0xK9/RLzNq5uTNG4tA7fas+TsS
ocuwiQ2sqRRjbeS6n9HJq2UiGBDYK2SJQ1ZWgh2KQfxrHqfKFRVsuT4StRLwj9h9bQeIVPpdS6BT
sifOh6MoBBKRcL2PiscEKunuOgUCRZWeI36xtFaCgai/6pD3iWU8QGaw6aGa8JnK9TySAvLYAzCn
Qb9M4wpHnk+fak5lxPkh7Up14WJRxeYr9CSpa99cyEMnxoyHR7Y8rg9LK09y252N8zC2PrDW6yZi
WPlNFWj7rinhaO7y7skpo4TbA7jDspkyNsZhNymUi29gdEbMkgKBJzbnbPdL5o1GYe/8b4f+Zy2k
67SpCyzu7cEEUlfFTYwUAisgzQpQIQCq9O2svTGBUzQj9qBDLOJge7SCPIzbiYnhlzSZGUwn3aNj
gSjwi+NdA1aoi3cqiORdORuglqimpdyUhsTgjvFK2j8iMHH+eBKN3oxBi+vDlSTnm8b0L+1R+F8M
ERTlOxjsKJMgSeV7lfGa89ylkqu3xYl+eGZxOwFnluFKR3V4lvY1VSj3KMhytPkCipPlcro3jy/W
0YG3usC89yYyqC6clcsuaOBLBlNGP4xrzWEsvo4Lq5eVDRPSk03faNK1JHR00vhQuk8LacKGv1LJ
Jge1yL7qUfeOWC0twk2uoKQeDXdGuELE769c9qtPkNbYLQifwgFSoIwZR4GOb0sGFyj2Mu/Ks8Vp
N4bipaTAelmqJIETglKZi8j9mAf0qvr/biuoQAeeWWPsMgYlXPzfx/qjsiWwvGL5ELUDnvZU9LgQ
Ihp8yHTOHiHW6ap+0nNMkZ+qW4/RhB29o6BseWOgG4CsqfMVfYLOMOgDhSRy0+CcfsSMc2+2sYBm
xBFv3TQ6jDiui4sSQdSCNdsVS/znBNijCS97vtrpKB5phBn4N+iLlhhDoUsRkI3fnWMfZvjLqHlJ
LsICpYCqbzLDmMJV5sdLsIJRFX4xSFFXE54cgttxygNV4nwnGH1oCW5VdpTS1Z8jJv8+gFAvCYBd
DhtZPGeXxlr2sR5l8FgxPr5r4WfDclLyV+1jerH0WsK81DgJQEua/ealX/P/rUb8Xke+E++kxF8X
M7lopTZjccK6lSu3FZSLuAzUwDkMdZAfkm3EA8jpymy4sC9B013DEKEJDH8V+HEenKv4lczHfgr3
nXtJ0Ct1oHIorm9zSl6AhlnGlpGb7qQtvxqSkQodWs+BPpyXmIqz53mFp/88GwjSvfpfA5/Pd+jS
DwNiqQE4jnp0T1eQklxz+znTzvy7v1ToHe7N7+WSZsS9ntF2gsphyF1Mt/XdHYWMS559xYT3Fq97
RegHc7anSX2BQ5M9Eb27VssEJvdYc+7LgRP5vdxBmcVuGJ1ijBQ8f92gb6Aodjw1cg2LB9Jvw9We
cPQSjgcQpF8ydIEdfvNRy1XXlizuuP8N/+JojAi67LKqksB8mng+Wb5fEZeuzpVfDwXaZHyN9/xA
AC0o1kQ5I9W+EZS3abHg+PFck81QZnLmWyL8IzwDBCMI0znkBqeW2XxVRl3zfA6a2y+YogbATXGw
BEKx+GINqJgolYqBhnq1sp4aX96wZK9ZX9lSLcsXUagFJflhAQv5bPFRyyU9rxRJ8mnR24K4pLZk
hfk8R6kQxTQ30/TSAwPfTdpF/1qjAZhedopugkUvd3qiivYmgUsEBNH6ToC0zU4coV3UWvCGO+kF
8UCXJgbLhQtGJ+UxbM06iHyj5lck/9G+A3VXr45JXX7B+jWeRp3pdMDit5i7i7RocQ4GWbxYkLoQ
2ruOFaoNfkaspTpszMQv75wpvYwxxyR8Zq4uE/Zc5yEZhO3n9V7BVlFZoOLDm6c6DcBbcxnipp+v
S9xizGii7GRv92i74gbqWT/0VTJJuULC1pK3bTiAPSMBQk4q6fkImAgSIyus7iAWDoaKBpgm1GQD
AgQiC6gs6tvUc6CgrW2VmGM0mDGdEpeA5c2U39EYPiiuBZYC096wTmhzD4hw1c/wZniZRmp/ngV5
RmGa9IQpdDlOKHaN2pCUwoqsSd7yt22am2Ze4oIoLkz2SbV2kmCXTKqtzRyoEiKTtpsK1PAzKB1Y
EeSLHbqHG0T75MF8+85rDk/wyisvJ9sxXVkhhI0gIPXo/mqcFR5Q4K2IOOAFg2WHhUoJvlMLVrTU
zl+0rwGqLKvry2aTjmobSVjnDltMZRFQ5rlqOA1F+/j3XFya814ZINvpCxC6KPtIcIKm0pxPAqfg
uA4AHj8aAQpmDouwuiYWNdyVK5WcAfFj8QebzvnRLVm3ihAIOMXxVAdecR0+M17uvM31gO0Sj6Iy
yMVcEmbxWjjPTQHgEnSkZVrLPNBtxfQ1ypTRI22mywH+Rgqx3qCDSLAmkzl9Mc3fnhdji6TKP5Cb
EHh9byaBjSwQRAq8VEpVAjx6cUvrHqzT41Y2e0lm5+saRL/hzGWK3U6m94MwOB2cR1HohEbOSABa
CcYB8YU5jLKU+EpNyqoIkGZijBRN2DNMDX71fJ6Xv67GFH6BJqzOpd6VYqxohVYFtla8vF0r2VWV
TUYWv1OytLKYaDRLlng7AaPXjRL+lBYUwYgb5Lw2Gf1IngwhsohpZ1NW8inbc3gBYBisoj/An5kk
lz+nTZSc99Q+V0kRrcExwmYA36fbuH5gGXigX8f7ktwHjte9Pju/SGD/+9rxSzfn/BKhQzhEbAHw
Tt6GNOHY9HmpAQPBFUVDKHUUoCvzgluk6SeOSuVoKXN3Q9Q6wQ9Ochi0tCsjN8gyKUGyAPyAGxNe
nXSKCiVxzjXQQW6/Q6cM1Nnc2Igq26D04IhML0iX33jsEl6G+Khy6NZIVKnUvDhlHU5YMXQg7+qL
iGv01u+PGfnnlZoB0KBzcSba1WHrSjEg2uymReaF4TWHcM4YFBIQ0RAzBavCLgK9Att0T8sOaZnv
iWZBadnNrFYu8UoLOHUlHf7f8OvGyBMKhp1odTgydrakugHvQaFgXDk85ZgGF1GfPKJ02ty0n/Q4
EUuKSkaIDEmLFIYW9e1vZWwtMR1eicW9KIrvS2LSJusSCf7Tv82ZR4Tv1N/arATJKLBFJAOKf6TE
qXjKQbmkOS9oS8qwMxjQ20apSQrZeXf3+D5b/mJHfJ2I5DbV+38orkM6UvTF3L+VfEqhEcij4qIO
RYbu5tUsgLRPZnYv/plSr1RSjDGn3SOAmy8FMmUjztHeoxkmlmkR8twp4VBNoHClGUUV4YoUr8m0
w5m4dAaQ5GnflT8Q5/Hi71lQutN0TRfXLrXXp2wiDThKR80Bpvg1AheFaqQqmSi3YaycbWk7rjZs
uQskSAVMio7jtNgnQV31+p1FxgdxYydOdm92wnmvIIDa8mGJ01zTfHW1HkAKcU7DCTIbew+v4oxk
j/dcYjcgdIXErYYtHZ59VaDIzD08v94DmkjcdPS8SeHBF3lAC5Srv34iaRMHVttVN+s5ysJCppY8
T95PQlS6DTggGggPTDwLHR4jCmKnKg6ayon6qA04eq9f8Y1WojYMuQQ/t1qEgjBPz+FRVAyE9Tor
naj33P7EI0G8G5jSiIoVKw8vhY3QWAKpga5xmLO8LT8mZ8GEGKwKYyZbYTJRXwHKaVi/aeUr2KCz
SB/JB1caSHQHEPIFwVyfM3KzLA5YpLbbhzpl+5KnDwqmjwsNlGgDt/43UDhEawZ/+Yp5pwS3/JVT
duUMO9FmWqA+OrdGZ2GgmGQ3cjdttZ3iGJwOAwngrpk6fXFm7esM1GbL42TGWRop/GNw1uzXk69x
ksRBzqqOyDP4W+L/p5QakNo9EEeE1pc/LZq6VEBMZ4PkaS+3EGvncNUZAh37SPjwKH8L2lymt14O
bQYNit7z9fYtIxlYeE+jd0NA1bQ1+u7VH4cFxavPGfIlLYNMvxxbnzCNm8uQfPQJCrwi3g6OnrBK
UHx+2z+pdtzjE2A2mmEY9xfoS/yjlry4QEE9Mw9wQw9ikcptpqrqXgEjJ5mJBVlkLcIrO+4k5HRw
u7uNdecv1frLZvH+HkrlPoF65EPxDTfLc2QpWdRed8sODn4zdKjOg9LzF78RQJefQpKUHjfvkEzA
vfZspO5gwHXqdTvbU4wl/auiOL6ANfXDfeVLbbphUWRKwWPO8TRU5Vm7wQxN6FuxuH6twauoY9O6
zgLSVlh6va2Jmd5XNe5CP+sZHum7iw2Ff+oGkOJAaX9Fz+MV35kCm1HpURqbPElFggjav2NDs9dF
q+7Eafa0xCITCM2hgmiXAhRvQC9o9sT99ua8eFYNwXFAwhuGXqrzynnqat/x/ECMPDFvwPR4wy5c
v9muLGSC77uG4ksWkuGcbWBehCT6wtLavmca03IAm2C0fQWaX0DgV42RB9TIDkgwmjyR3v97ksIg
fuixqbRAS7b7iO5k/2e6t9Rk2Dp2SRHMl6/mStCknuONWkPIGgGQVUjfSs2JI4Mizeh6eOpgoVWW
nclTR4LKnagMPlloqmDDPJlzrByzd/BjB27DKTScV4fI2kEoH45XCWIJ+5Dyxzv9TQL1r/i9wYHK
a7PfaRUHAW0gXrgYtKOV28sYeGm3HjXImIzgGz93ki2Nlw2BTtAEWBngFqQ/5rMs5Q7G/85xAKLp
Zp5afBd0CP8YI3OXIjPOSuuvKSSjMed3CxrtrkcZYwE1U1u9Blp9Ay//BDqC6sPUEtkq2dzims/i
hF/qORLUbqef/ejlHId8Gk3kCAQDeN/AUIZnXmv3uEX9DdFIzQounEyv7Kn0FBatTXoGo2owvrm4
+pKWSFlMfCsupeNM648bzUg9Z2V7cMoqlxLBzjCySlwpcjeIj2YogF1ieEz0qHvpiCqXeqmrHIuf
8Q50h2/wML2CPutBl4xuOGhDWM6pCtzTpfy3GUyAHXmZuUVWv6qnDSX9p3w1J9tCLbCiiYd1PhOI
PRMJHnskRJh1h/moXMb3/wVQsxTSxFVhCFfxV4hq3ccoWnQzofh1QEWjabc62WRuJ71sCOCA0Xl1
KiWiaDQ36ze96SSTG2oDwXtktPMFmiQrH6YR7MbmRORRbZMYHoBMkrBq6948PizaaGPyvn/Vwxw4
ZNGGYdoNv9ZfiMXEW8LHOlhN5hVlQzTKmV7WlE7VfKxW/nD3KELrHZZZrxYMns/AV7AIFlJv6NDY
uGGmfXYAUKVwbEB9Y1ShdEcp2E+jW2hQ2DO13trdZbu7muPpm1L3pjXsSWlzqFB35HTXG0TmCdQH
G2UzEID1dP8PijCbVKMQhxZJItU62OL7ms1ZjlngoDddndTASVfpR/hSp58Exn2XNPDNLPSixI5T
LJlztK9INRsyx7k5q+leVgncFDGDApICfYBkcj0FHv+JhiiIixHUWSz/8AdQh8QKEXz4A67PtxAP
XrD1Q4U+io3qJT6xID+x7BwYm/g+9/uCa6ndPclGfap7CeqT6nN+GnkB9yu6lKAjCiDx75VvlVhI
jgJoZWxBUsovTIJO694CDYkq3tegRXTnVZzOMB13EmvS+A+c3ACOVJr1GgL67xAHKMnC943q4sXo
sUiBZVGVGZ5qAlUAgyn0T7jCi2z+6rPZGweuwMbnKXCD+H7XtU+mme0je35Auc6fbkOfNnpP6Bd9
e1zcv+WaS7MNP5Moi2J/IebQGV5hDf8j5h0QRpAjMxTqHk2a4LIZMd/aNBZX8FO4iimvxyp0PrEf
Wx7tMXX17qyGRggWRNjcUpOfmx8WLX3VD82pkwCrHjtPr9tzs//TtawBjkoG82vVKicgrTW17l+J
HDWhiQRT+an6LrRc1ERNFcsYnxcNTlExrXw79RW3NLXsq0I6ykv+REcmg8rEuj06soR4k9lo5hKX
u5p5fuRz3frKvrQk6XEoVFurV0JBhoGEA//Wj7tK0ZNynyPfAh2RTgv0OJrMOnJxCcYoeHlm/HN3
Q6z8u6iuKERYdEJsB2960D+W4unopy8OWLNtQm4JFBBDRkbE13qWODiRDXnzlb57zIQyrZxtYKb9
fslRDes2FgLcPNY/1UQJHugsOQ3lOOHni0Q08tIdxkLG2K1cTP8avUleMGpNGL4WHYRNKKQ5tzhS
fctJormAmnySnMdi5ul/LCJMwYyfTPuS6vvioiEi6V8SFJKbMpbDyUZ8XboVD3ZcEnzlN1SJZ8Tc
oJSRfANB0ThwPIhxJp9eNfDQ8Aza0bdiWXnXSIB/On5kYyjm2aiE3EIBm8Anod8pMBV8bEuw/T+h
rLuSvkdlAEQMV5c9TkWo/1bQ5khLg/QR4KfruVDvS+6UiAc+997z65wghnN6j3SHE/6NKtUEkBV0
LDWmPANHkPNjWUYu/GzQ9kitD67YfvHH4DYJsndv3NDDUcs3jNqXEYjPJkt9AFneSM00y5GFLE4m
Ni8Don3KgMZxLhxH9mAmzifPO8b4W4LngWZKVBpiNhuxQ2nd4LfqG1dr3JSWOY75QROBmfrySkkr
Zrkf26iPkIcA1AAGfB+Fhrb1VBV4FOzbuc4D8uCgLu/BOKyGco/DAy2tg8Xyw7ja+o1lzau2391s
5XyTjYgaJBPeNHOebPayLU6Dtd9uyXrXetDFCY/wwLQeSAqTVTyVD1oufiq8iUtc/2vgv/u8Rhg1
QjBs+kEqln1veiRweNNl4os47S7m/zJHVstu3z1rKolD98htiiJ2u0izPh5fv6mM8UZqAT79Z32s
n1UJcjDb0i+9KNOlM2MNNLWSfODVvDueB5rzGqyFIv+zMKHk/Za4D4s+qGRx2YqIGoT5B3sqkzEm
0NolF4zPxm7/IwwJQ2Rqlo+7bnQbvXU+byuC8EiQXp1WEUl6iFsu4T2HDDweQdl+w81z1JlBnyPF
9sq6SjOnww1ebTxA3ydVMMgFIJhgjE0TwQqXhH7KaUCFnA6ncdvGO/YNOMdt3de3AkNLKNZXpHNa
YC8Hdg+TY2aJs5Ll3FAe4V0Gp88JtqxG3PW+ieokeuTqQ8vAyKs52NiJdCPAMttpMPjO7V57f6Z3
IQke2U1f8Sv8cX+jdmo24Wv0PeK4udz/j0R8N9fy3idsiCiV/3JeiWw1t5njbJ8iAZqe+ncSm3f4
inegcxmTshM6XB7mN9x46A5ay6PP6cw2OXYVmeZ9gAhrDckM32/sdRCx3H4pqnOPCJnfIjioI3e/
KWp5tiYfqoa7B2yeuFVr3hlHbqYSJ9qkicLIx3aRfM7w7w5RHxZR0XK7vHX1Ce4N6+fzLg9t0WoP
HF6t2ZG+pwr2GGU2CnJI70QgnaVYDPWylG475qd0U741JtJuMyW+bXxYjXAMIVZ3i5q3DjXKPrcm
fFygtBMI5lmkXS/eAW1CKgs0IlqCgk+BreIfBj4tvwkemaeR8ymNk5yRVgOdoz2q7eBYre6ezK6P
fXz8MjkqtWM/jviTVpx3ihv1Kt40pEnPjXVkAP/6+nxMJWli28+LhtUFbIA+ZDI8q+dD2GskfokB
b6gRGLYSFRr+NWlIiLCD6stbLatdKYQVXPUp9ed5GgMK8WKIl2CZvo4BfMsk0pT8+l8RTFaPZBru
tZsMsUVzOIzZNs4I4QdoKcSumxTQesR5JukJSvVEvm3DpAQWKYocojyNmeAT45eazygUrDKT5C8t
eKoc1zi5zxQslwllKuCdGuMqaLr6hPgf3G3Bc1nuQkfkiPFtd9IddX0ywWnuXsaNiqrn7fqBTwv+
tQmdfV17Lr1B7PshGGYE3WpVOHGXK0oIk8rwJmicZWLVYc7oH/x49esvbAv1TAjIxSyYlgyESEyo
oR+sMFp1LBLINCml00y6qyRNrDy9JQUdddEUvQL67xlX9xUO1rt9rf30dweo7UjDf9jF/niaJy8Z
KDSRsV5GXUYrR+iwjLjACyoWgCXoZ1V1blBkeiCjrPcGKEueySGOwYcTuSJt6/VuKWBouJ0a7Ory
9VdY09VYqlARBz2tNxKGDvN5eSlXLFEDdF8WnNMS8A61MePATCvhSn5f+5BDx3Ko4cyRBPAoWMVr
QpAbTRobdEeBRhInKq1624MC1TfnyDjch152L0KhwnZoYhfQr3p8NznhzFHd8k/Vtu5encNFcdIo
M1bhVTEbkbGoMlAeazYsg71VF3YuwXQ5MumL1bVc1l1LqTlKrJPxmZM1iWrWmq4UuC/FHH8ewFKg
pzN/XCLdvzGxa2HJa7c/YkLacsDPDVZm7jsiAJ7nNBugntqDKENP4oUghvbDOaw+vuKYM7EPLZ1V
fqASJdyoiJ4wDie0zZiKCq+m1pBrFZMmk4A0InLIatsfJX8xOfg90WGib08Py0QDzhRIvLrsjFJ4
nn54PCLy/yfJF6SARyQ+2TcSf8ZdAKM8pIyCmSj1nRAYwXkN29w1EWe7XD+pT4BPX4VOtzmUIAVs
JWpF9nZNs9Yv/ORhtYNOgAdfu19QNKX89TmS4Oxhw3eWVxV/wbpLhz78n9oPfBl9CD9+5mW6sc6K
JA3f1s/fmmKeeBIUOFYp0SljeMPIcWIr3Z0gulwvRRAPrCiDtZYJ30Ihe/s7DEf2kKySYwPIPEXY
ECkNMTRvbZHxYKjsn6tOkoFQuXzyrghfEI+qA5hpfoy23Bsk/gQkGCV6cRHqOiDp0jXwMz9MwjVO
vDfCDcpcxdw6wXO1eYXK8k8CtF5xd8SKdtnlSHxyktts2rx8fkisO9rWBxE1U7agRwUUdvIFcIbW
111KQfMF75iukFGY+MXvxzyACclOLQP4wFrTdrjVpITt5oCx48v2c3Au6C1o8daSfwIfij8hayMq
1R+dT9ZYz8XkNkUELHOCtQAy8XJ5ya/pJPCwo5DKn2R6Kz3OZ2mOXew2QTeljKtTvax2mTi1c9sP
FCxJUIBhRsWUOd7l5DKrRz9pmSB+1oKN43AFS5CmH2WNCU8n6jl8KQvcvhlkt9vWgWqvMNTwuR1A
LE4sswaDRJEA6ZSEDy3MiBvoy+SiMvV/JipmChjW4VRZ/Z0YX8ZJRcXUsysiF2vmwPBmfIXF8wGz
eGm0/3KsSu7dyB2hlNu7EZ84VArnJGo+zV+dTwaIINAa0FlnSZ8b9daTzvhhkaNBiuu8hpeC+m+A
wge+oT7WoWEBsWLcToWs+9zHkSkk1/3we6TPpxPjosLRSgk893DqAWaPLRrwJjyHG6CowW2GQsMj
LLAHh+4t/JUPh/CbxjBiPI3FfinmMOJXTgPsi3nzF7lKAEGLsHdHTm52Yu5/V0CyYQuZjgq+Hqxx
eiSOkHJgH8e9tmz8DQpsbG2ijufnXk9XWx6Dt2j3fzOCKoSTxxL0rnb50nhVLulewA37bolLFyS4
HiyrnjTygBsjYG5Sa5T4Gdodq98ASzP/uzOmdgQf6WZoJMyj8lbH+CdcBsITFuU12fU7PifE9SJA
0tPYB592izxg7jhV0wLFXqWp95dFGgAeu5qFYLxYCbmhYqvMqXdE083ZYvn7xoGHCHadAMwTaQzf
6YMa6/CMluF/Pg9jTI8B/iP4BeLCQY7tJaQdspw2I2csbRL+8F35/vtl1nXiaDmua3j8aMrEH9UQ
taAlJtyxtpflGvNzTbd8Wef7zFcTR9Vc/Vga+uobjW/IOCaa/8Kqp1R99hOUHs+Ku4XAGGoWceLd
bHRo/2KHV+G394OFiMjJRCqTBSyHmsRrqloNbFk506LijB2Jow9YKsKjJo+RiQKnuYBG6GsKM0fH
YzxJwvawGFyRBew0GvmfPhMS22xu1Yn/yDSsf5jEmiFuvrlfIxtB7rBJx7bMplkdqK3mnRcn2ttM
ccb7j4kIWpErXHduE5Wl7GJ8s+wdjN2hcixixkpYqRrKFgG6Idy5gT1e+L1lpLtKLUCG0QCPFgQZ
CPzyF5qpKfEJRun4HNz3YND+P3x+FyDsqQXsjStHkrGLQAUDzswLdeiYd9FGaUP6/8vEB2UxGE2+
O9D/53bMMvg5wAWi+sXSOzZb3ifOmLPdM5hz2s/jvF728KrsMPs4E6HWnWHIC3GZbqDrvGgA+bUR
3tIWc5ZHZhG2WdwlVeifpwzAvF0KSB8iOlj5OPfQSkKgqjKGgS+DkPMQL8DEMb4mOwzpasewWFmN
lhfbBEgU2x6wosZunWPLOdzVmPBkXnKPvljcIfh4K+g49Ab4ABtyZ5ZcD04Rx11zRVwaJK3LucLg
RSxOzqpvmXz2Ob1U0jbBnY2qp9qTWW5nmbDs42ZbqiH0ovBYorSRfaxUYpbof6bMrPr003OIuROR
YGn8jQ9yaS1Kv69o87xCz0U7YLL0G+8ReB4t3zMBFYb+jg0GB4QKjjne1ErXllRdncrsqlvyJ5Bh
73UbJIJWOu1DVe4u0S/dj4KOdGl/N45yjUTfUDkG8OM77Uxr/GxynwKtL8E/9f/bfNf3Yyap9kqO
BN5WFnNOq3UBpw/0G3J4srMuH4e0DngYLWHFdg0dRYz8vpuOgzF0uj7Nwgf8/CmH0NAV3cLKD/sS
U0rDn9CrcM4IqNCDPL70NW4kAWm2Kqg+vfb37cjgQHwsFUy8yS2Vc8zytV91r3a3sPNosHzLf0Kp
5jf+T2b9P82d4S4t0+2RHzraC9fWQUumgxzD8NYUKH8Esn9pCW7USaiHx4cEFCIpyTq2opc+J2Jy
/In146BzvQB0sO/YdnCDwhEc7h6l9X/zRtYczuTMCvDF9BBk2F4+je9BfBS388a88tWecDMdA6UN
pUlfKYaLB9lTv/Se3yKyuumpKS3tDhLUdgvW5gW5fhiOBjDmlAXkwX1JqlXNUCCp3qBs57/9gd99
psZuOEC0TbuOjVFFbSaPPYWdBcykJGZDtRSBXAkl3AVG+YibiV0u9h5qjgPNZ0n6VJ10ZMTEs7Lo
VETKLWPSnNYJeg64TGBHAnNARUAOR78jNSHvu8qTlHUVwwa4w7Wv6RenI6xdUfU1ZCTwJ8QlRtt9
SMO7xnPiBv7qmCqeAmMltDom5aQn9rY0lI37unTlxJKVQ8N+04Nf9dDLUntSTuJzaawE1kQZYbUM
A0oKqGeybQsgQ86kEjifwQiBGwJdT7k6TwEAAO2sjiKQI5OQ6/QZsfEe0Xlue/9wMAFef4bO5s9l
8uh8ALaAj/PS66jc1/9sSyGhf4GosvRq/HfSZBXFhDQK1NjITQG3sVT+T7s+kjCaQRVMMq3KqmfO
+gQnZoglWVfoxrjMWtwaryZMNiJh5IyWrwQk9qSVH2ElAQouG1XAc4Trua1khjUY9aIb+MCvdRtP
D/hZeBBZ41YKiBxwSp7SLcT6xvrH+7q6ohgC60V6ybQ96hjh872fw1XNTHHKjIbxaP+q3ptoAiRt
xM2qlYdyZMjjkzunHz9RaPzdxdLVS9YjPcw+CBT87Y1l6Y8jz3zHNK6WPP8AMwC9LKRjotwzBiph
JPNkQHVVSs5p7vfnIH8jhnTbwgrFpGaJs4WW/cLKRTRQX5mlu5cYYgT/8YdqicOQgg3kcO7uvCnd
vr8nanJX2aN67EO2Hkr4INq+rCpbxcbeupp/FDXAsoXpZYY9/Q9f7SdtiyF4sS48WS9Rrh0HLcl5
1e8VP17y1ZMQ2vYJ5ou/XJGCGA2dPl6K6xnEzmODk9t3jhOB/U2UKqGKgp/acHbnP3drYpJohE9Q
6RxD+cQWGIuwCXBDO5E1YkqLiVzkyeJ/gz2oSjAPzjCiVxrHiFE1VK0Wu8/EggRPUybh7w2CqqiV
m+MFPvlm2Fc532gYcCATD7MhTlWeVUrcV+MUO05c6SepFDvr2UvgQsAppfV6NIXjr+borh8Wc++A
+prm/r58QXYDcxWiHutaQQaUFdPRrTQENEYscvZLeEwuZ1x7rgD2yujxX96JtVrGcgKRYFumOoSg
D7FwubEe+HG37JpdusiMVVO9BldpyVN7ehLemQ2EvI7qFPEiey1wrXmN8CqA71pQoapxwjK5Bzpb
26dHnq36U85nShOoAjoBbR9PzTfASj7/aNG8Cp5I3Q2ovnk5GDiuO9konQ2kZM0Z8yLF1wxC4Jo3
lDQpKVPIaNfFRdiEURNNf+74pZ5aUy4pRS8XcUEfD0UpuR5Z5hoCBqOHh7asp/QvcbTFr4q7JLFA
uGgY5XXzSQ0/NCfCoony4NmeS+YefrDHVzN6CMAAiPPfv7YwF7rxyQgavkAMkpWx/KFoiMbZm6bO
9pCqt0D58p/Cd3juW9NVZT1mujVInStKkN+Pdlehz+GoFcDh9jZ3irhJ1wMgI79T7V2j1cC4seLs
gzOMfO7dteRavrKqDjplR1nwCq6yzuPUdqI5E+X/R9ZhTOE6A+gkn9hrS9uFTDOe7Dx6xNUackHT
KzlIS6H41r+BVhwH8zwq2jekaiBBTaR5Kh1N/dQUFuQzcoQxqLbgek7qDrVkZBkNh0AlV0B5wkVk
RZmQQqQjcqGslgDd54VaamFMJX9+Wx/ODMCvTjfgz/33q8EwV0uIvLwlF0EXH1iLqNCjU5oM1uzS
mODuf7lbKqSY+us46/vbBC+Zp/pamE9XyXeDg7Kl2pwwNRJSg8BTxdB8mcrXDukE+l1I0GmRQZFy
eUERK6c0/TlopYGOAs2kcKKFzkHosPOOY29d4eSTxUn8daDqww5pJmAhox2LSliVSRaWCpv+SKTN
Tbkmu2PWLNQp4xDesHmyMWVi7VVXjLoJuQwMRnC3DIN+DQzEFXdQLUZ1GCgS5ec3QMGc7qAk+LOG
CRvt65K61C6RSwFmA7qGaB1+sRfPHyZA+5SkRa1jkkM1hyk4e0/dr2x/NUat8223I64riQ1PWMeu
lb/hrW0kv/rZJK4MwbgJBwvVE3kNYHeu+wNHGes1sndTPEAmlhVTpSHucwLYXkD3WLg/jQRtJBlS
vZfQHIwnHsyKIAP41Oa5hK/F1+AlSqy0O2mtQwH9Ug4J7dIz785fxL7dRkrbVLzZ1oHZl4YQLj+1
eXZwwHj1mYtzoR9mBAxj0a1xd8BHh9y+Wvi/4q75nmpKatjEHjCI6hfT45ImjpweyHQbXqKVw9DV
vOGjG6c09FLjAQJzOdQDXmt0yunM2exaDN1A7h0MmAiaW7uhKOHRtkfqt+BfP1H0Vh4oebe7faI+
uIHfNgiDWd1grnoGH/FEV/vCt9qQNh1l2NYjBVxtdYAefLzOynBga4MObb8oPn7gzENLewl+bFC0
U7Anppm4m3KCikH3IyS7ozYzOZyItETnNT6VCH5EoI/TUhmHjwOJGZHcTX97FvMrbNQs95C48Ivg
Rj3+EKRUVQsX2zb0UdTXwyr9PvUfKwECsSS0r9pO5s/AOgN1U5ArT5spZJPPDu0UvQxxWuWmLybU
Pr/JSHymPiB0lCu4PD6GcnYUO6+ErMNMV7MC3SQcq+ba6N7vbqD2oGX1TVGrxyDwG324HVmLezvs
3KLRXnv1p81WHdvL5XyDjnvuKZguRwmoH1TwiF+TclnT9hBOb39EJkA/wfDzSmCdV293Weqw6y/j
1QrwWxzq/Sd9FKpln1lI4z5OfnjCpB3B/CeuoHJszf3WuhfM5EwVOWcy4m9y7UiwElWxBUOXuWc2
gUq9a4gCP39e9PYPColUJTJBv55KUx48CKgiPHC1Ab9GNUNqYfmK7CAqfiJeRLyVZdelKxxF1xI3
17syaMcZXAqTuDyXzgt1q93Kz+FdTzDMCj5kUmwv76OZTFcWImEVy0fzd6ISikodR20HL9uj0K6X
2M6swTXl4msP3yCKjs109B3YVC4/+gyAlw0TymE0GcoWQXTktrfrFpQhP070frUIkZ1wmSZ5VFrI
BVIJPVmVnigTx9SHXL1RPhtso4h7loKA6aiSonEC7Cw7o+ms3RPMZTTo04zETbW6iBfIfvYp6GRm
CmjL6DpD4NILD4pMwz/b2ewUgA+hFvaGBejcqqLlfYQEbtC78B1uL64DtR/lB/3TXTWWndGE1a4N
0QUsJRaq5yDld5G2oH3NUvdcFrAg90Y2NH6CO9MifcgMPbcjeYG8P6TzGhNN9juwwcIJ0aiImXJh
ZBo4upCRq8x+zrX3OHR53I7HLtUcy4U8MjL7wqE6uP4sTB1NMJpRoMa5TcGjK0MpJtbNCsqa72p4
KoNppXEScMw3HitrQAOo+Wcl7aLDFyqVqha+eI9qU1oqPqllVDZEn9Vxp1Joqd+zUTnz3z8Xm8do
aosGAoKsGJkjpfWkLxTbDcJ1/ZPumN34W/vHOhQG87r1V5/HAuORUKcsRVZoI7jiy/rRbWHo0XfE
X32AQtBc8YqQTaFvcbXgACpPtVMJZ3eAo8I9G6eZwUBbATqpJILh7Yw/A2wiHLSwtXLQ6lQvkg1A
TLLsAaHbPd/0bxee4wyh/ttqHzgei287iugzGnVen1Ux/le0eGkoeOGHi0l3JL0255cRbZqa6Ufz
q2/5j8h9Uy9IO22aWc3LzjVD4paGlJj0MDXsc5A/EqjzZaciYvk2EbWVFybQilvpVqhTbObqXWh6
J2JNvUJKo1CL1WTFL4P4cfxsQPsIUtShi5KJAkKGbyGfX+g3jhVv6mRymmQuYHhFte6aOhtcZNen
fBN3LrTWLxS8ld2koNMS1oqzlEQA/H8e0KA5EnoR7rhDsVnG+VFbPLzCavq7yIFyJmydP6N1GU48
4MgB6JRydMBW0+O57IQjdhsjaEAPBC2k30CrgemEdjWSzsP5i2NpRpy4uZtQzD+mGnSNTPb6xsVD
qqliX6bieNOnn2/QTjIeTeJUZRplPz7A79lHtgljKEpqb1Nea1BhG372Upd2WCLRlWv8PCAsb6Dk
SRvj0I1lr+CwAbqqMDmTVMUkZC+RW9Bs844RtxR/rLGJOhD1yqyaZ9ToWLy5udSzNIVq1ibFLcsI
cmX2znRwVW/ERolWhWTayH8UZ29aNlvbVfyizO2HvOd1Q8sjPmipogeDUJgrjNuDf1e8+eu3Q//B
Q/okZmhvQOK9Iz8wJWHevsv9rTGphHP3bqnylITlPs6n7PeHBDqUMD0RhDaRrbBN8hxm5gbCjff9
YX96vIgDiv5IkFbCJSiyrq729I+Uc+B3rQh4wUYqOlqg7hjFfEEITZ4ceoRgTAHD3L1fxKBjm6bJ
kFr/V75AzZUqx+xOG/jgOR1BIoDCKi71N6xAo37X/+0Fy4FGKP0WX8a6V/2wYWXNYXUip1/6HcFf
1/Dng/asnQci6njYrHTaHDCamhTAJa55XpPJMTJJv8fxwdUFOJY7Za122gmHtme7Flsg7hUOx1ix
Q9Dwdgx3i/MiDwHVOvXyaa2M+sBOsRtJ5t3+0uuPZqu1vgAYr0wn1Smm/8v7CewpFvmuT7OWmcMP
AuskF80aCrutFZY7q6k9afSDQTFMuh1mvQzSN6yEiqrDuPLYrunA0zJ0BSuYTJvFdRu7BdxH01NL
mAaVrTaRHHESrGEvYIrB/cJrSnfNqeJL3HUbanh5a0G3r1HnJhR6EvaSyshSE+1K8ykCHRv0eY33
5ylPS8MZQWoN/q0SnAawh4JCUj7uo0u2LMvUao6xxrY8KRttKynOQkDhVdErXWMjUXGT3xtWtaHt
7rz3eEoaCM+Wys4goHr3aQHqjSc6GtnN568IVf7fqZt+tGRah1oaGdo3WnRrhcOtXCqoj8qYhM7W
JwUXk/8fn5HyOSQeePojz+vana7FhmTBMuj129Hzhw3ay2sGLZMwKJm1bSMoeqwcuixtIduG8luI
eSOp3t09TEavgGLp4I7Dz6XY8DgeGrKHi4SZkgYbk4WbKkMUJRcxdzb16uiFBuCHnUplJPea7HQa
vGaup5B3+b3g2tBP4tMrWA5782tR7jYzBs3/gzx+50R/KQulQ3aKarmyXSjS+X7CmXOoSqtBO7uP
sFHBYh0R4+8Wz+cHKq6sgpm2UBRU6gAxEvr7F7bl2U5goCgUg6FPdJ8e3cWtkt402jTE4jCTX7pE
KU9vdPvzj4w6fWazJi5Fq4aCH3BLvov8KNeqr6vj0OpsChjzEeiUeWKbYzUhdGeDxBulBkI69sLD
Fes6xInNZAEhDr4f1qVqE/wWnlCZf+UXn5Njh7EA+7a79UuIU5qLmHZafrb21KmTM+mFQbo3Ztsl
BdJfbx/BNA6Jd0JIBXAHFvdIgwtLhLqDEjcfaFkYYOhk6dAAp2YRCKAmoTvjGTLDPabJfqKoZkT/
osdCL0ddXzl4HTOdl8aTiIUSc4pbOcLGRmA1BlqDvuBIJeM4HvDTEM3RZ8cdh73hcNy3J+ovRlcG
ixSShx7OQoIoQojx8JkEnM5jDA+6Yf8S+AEjFSI6RdHiR2/eVRREUK9Q1qyPl6bjO6+9Q+aucUTv
zTzZGzy54aGyaY5wyW/vy7fKXNLOxTFCIvCZvZoaRx8x1lNXvAZ+Yj7N08m/k7Xk0Ddhk64uzcw4
puxYhyXutaT8rsu3CtFPgYbwH/IpFmv42plhpKkHAA8mbduBIlRMXz1sz2XKRrZATO9U8Px2POAJ
1/Mz2TUHA6YjVK5ZlMk5yli4u6DeTtZuOD6sTLcNEJkcPsuDXyaNp+VkHC6QLYD0v0VQE4lAT+XB
IvvRE6d0muK0EMoDwr3eMVd48m675TepCeRYOw791JKgHcEtmkpLOi4PNP5/i87+rWmDMcfyRuze
NAoPO/0NL57BigmAqTakKAGolMKUloNCiSi9YfRuabq7+xyDLKTFxGQw0hGZmeDbVsaf8fhdqykE
Rg7VqAT/VayAYiqr6t5WUYdehg3kUqhOQx+Hvrvu7OeZmGaAeuFJvBeFGcxb969lk61Vy9A+GHNm
0wIrA4/ieDqUKNshwzTbCs9F6cPCgjBPsdOt4vC2dy292uHxfxJfdN25uRVS0uZpGY4pRY6iNoNw
LbFPheOmAuBBIq2Fd2aamMYZMc9xedsDmbSnAezlNsc8WrIZP3a2NWshNrvldVJfmBhbZDU3IOSc
UxsXLu3cAoLO6fEOQtUBTwC7oUjcVHulrZLVd5gMciX22xlfevzFLuMa5fIB8YQU68iZX+HtOp5S
c8Tc95jzDiPvxYtDADGOQelNsO1w7pTZ3hxDu+GIFyUzef9iGQ3ksbgQMAGTZEhRPDADGY4mRfPe
/m1940bY/WZE4cu1B6efDHojY+znA0/GbTynbk6b9ld31v9wa20kWQVSAeczld/qSl+IFB2l1kuK
ShLe2NFMtleZukaJ+jdOSRsjrtXbII1xAaDuqh2Us2FINZ7ZIezeNuMzR6RC4sy3gjUzVJvajwwy
BJ7OjeQsbZIJsoqELpMtW4QZezNIdpFdeaAoOT9Mu+UK3fCW9RrIF4LIne++9C71RFT9wZrktpd+
Q7bl3wGTHfjBKzljr58ysnSxI+7rI7fVslljF4JwE94+PfNqdCE774lTB7K6r/bnJ3zGQrXMO0Uo
G8w79fVey2hcIN3LR9qo12dHtukrLsB/aougtra0/UeMARpbbuUSwkSpMZkbnqgY/xANMeD1VWz0
4JaqsytzmeyWiMpsztP+OG6lk0ZdV0fUU6/cr2PHXk56tYK9PQyCZrA3WF6cYJAF4ajkduTnprRz
WgE6oUkMZqBCPC+o82fYtdMZWqJSTuiKCd+MpPmvhDIZ+Lqpb5dP8XMKyisbzAn/yw9BMXbqTdCj
BYY9aguvsYU2UFeJGA+AF2lTE8zbMlvVWABpkDwehqSg5vkOfa1La0gs/eMWyBh5TOrMC99lzxK8
xxKLIrRpAUWzBBz9oeB8NFZrkG15Vlml1uRoDufpAgheg/fG5Jv2p/l6T/YI0mwMhNuzwFxJ9bA4
ekilIj9u/n6iNTSt/xLtrH8QGWJgfTv0zLA8k5yvbWs1ujb539QW8vUtswIb9nJuH1O6HHH7T2tm
A48NgLKJ1j6E7dD/LFl1HfARJzAJw/PxspNCfoUSTFzLb7lfjg9GRkeoWmBFyGoBjB4KKMEj/4re
vv8+rZi3QFuST5CiVPFv9JPiD5La5Ezxa89EF6nwUnEZ4tYCKxM+lmvOlrAayVJOAErm7J4MTRDh
hNSLxfflXYUJabKMZUGYDzF/0xxVodkt5vAgKdpdhDPT6lGX/X+aO+iDhm4XFC4ZvSYRlZx7xusm
htL7lwJ3qxaMeFxy2iIHSmlOOzDRJYUceWkwO6L/I76Aaom6MpRKrRCqTBtd+lbRAS07lrYMd6tl
v4ZcQnChbM9+99ailnH1vWTfqLlrvtxVEHORdwdWFIHZrfuJ48TjpMeZvVgcCp8I2GhOJhN4YsUj
H67XJFN+nHy1bPErTTcusf9inQ+dfJ9/nZNGUly4J6GVsDN2DovuTULam8KfZBX7fgbCJpv/LLnd
BXEiqkYpPo1pr8BSkmt0i9CadAcWqa+BdN+lVmUep4IuKcNiEnK9HT3Jlyft5OI/eXSiFYdx8dL6
ksYdnc/bjzVp1etopHr6h5bH4jksTaxoBhGgjpjvff6mFDb/z+GL4jveroyhTx/sfQ5HPW+VPJVp
o2OuAYdVGDpwYyp0NXNUlx8XzEmMYrK7NE1fXpy6Tql154t1E/bwSNwERhegqFXoxKOHFVrxfKgv
kfrCsuDuHBObpf3voBzn/HjdiWL75JfUK306NeP11oxJ+Nw5jVWAmx+vAFWZQbCq9QXtj5wUMC2Z
cxArcyCsgld6gtzo/WDCFDDLFr3670V843OdOORBpEkvImpxRl9Sv9wLpIh4rXfyyOMYc9Jo1S95
YwlA7FQ6K8T0opR9wUJfdGCVBYKmfCs7zyyTxV4nlx/kn5nsXdKYjT2HxlL7ih0B1GAPaHJkgoY6
ArPK8qjG1jFRQJISqlOXuyvwzsyv5E8mIpW4U7nKi4y/b1JavZH5arO3FMWF2fvUlVx5mWxDNjG5
8ZJpYT6GV7TXdjpgCVA3lSvHWMv+K784NrXdG0k+jQvVCMcSc6jzJNqM0wifzylzS/I2qLWxyCdF
4vmGtVDLX+O0ooy/Q65KUtX9HuxVxwXPa2H4uX81zO62WdgZdgtsIQ7N1o2P0WemPwL5WX3jKiOZ
svheOVLbh7qaVibv98SMevxkKkbbxvMCyMARVLraV/MMlsxjiiq8XAC5Bjvh/2yzt5UfZfiHgVtH
l53nqxl+jx+XWhYYRiNuVMwTQJvyfE4dxa4PNJkQwGcf3rhHSpVH/bUTlSE5LZDDKwDambKDW9lw
iKwaNoKGbn/DhAKyFJvCdLPn/0mDsC0zZKkeDEquP5YAB96rI+lBFtuaEBQzoNMMy7hv6bY2bYiZ
WmZUL7Jd9US+UADaa0gLsolIRWCn4s0EY/EKl+SKucZfQZNLtfPwUo9AZgoKNzKcS1ssvzUR4RUy
TJHbq3q+e2JIw7tb3CTmFizQkEE6fhnOufdHxWw9N8zGjZAxCQ2P8pkmVB78buXZYaejp/mp6Y0Z
ABDfIJMiHdHXSKcIsZrK77MsZtwPBmCMq/OZf5WA1wvcqJiSQYdHRFwk3FUFqt7DEDLkRoliWKX/
IySela2+xsd17L9PLseQXiu2mEuIxnAzVxuQFqVHNAYBswlbNx7MNwkqQv86CRRAXXMdxRewKJZH
ahPTCUoH0vazU3TeAhJI4WU8DdJTNDxjhd0aTUk01eKJ3wXB8CIegzmpopceUrjibeQnZSWFUaP/
eNpLRoHvT8o0akAdYsfO8e0JC2lQmV6LKLR8kLVJ5U+gyhTcp0gVHzq3B+Yhv87xpFbDfHTrfEMf
Euln6PSkdQPuN+ftHO+j6BxofRmb8X7F+GagxCYLJkIMWQnE4AgVtY72l60DCWRVeP5pmWOE5iqi
336Z9UlNXmFve9ym4s8o7E49mkOC65g+6Ps0N8Av/O89c1EAvx+V1u3jWwx2FIQbybzvwx8umNPo
ii/MpQrLkb9/oTlI3KHk/AxNAMPhVYe6MwXzUW8/TxoPIZK26i5v3iEgUyeOJPQvsD0qJviAXFQf
2cU5q6QUrmR+7PMIvB7NRCRry2Qi6B9l3iDkcEnHL1WBiirY7gzd0GVjWiTy7/Br+uyZ8pBv4m+p
qqCIK1BiX8d9L0n71LMnC/wLKT833GkVtKS9OuLjbPZYGdQmLsYWEo0OsQrv/SgvJif27qYTu5Ze
hZ1L9MmLZMKCXYCai52kn4Bl6IG2evoNrImty9HWaIIYtkjany9qrHXXlWRIdAdrVC0mcmVpmmEh
EN2BU5UQ3V3H7ObvCrsHeeHKq0SvuJVK05bQp6gBahQXXc5Pg5fyykjDKBUwNeqAfzF/E98wdxnH
/xYgS5WhkUCqefBJzRx288NZB1CkyrCztDgOVYJH4TSeSkZ8qf5FQmRNteK+TDJVzaFAONz+s8bL
VlqZD6jYqYmvpJVeSX0kqp0Ucj3ujdyxD/eEHAyhBqz2n3UWGb5vvpolQqwMv/xAl+VRCGk02dq9
WQEQYP/TU54XxnUeTy/u8jODkjAWs2IYo7QqYlTzqZe1o1ySFo72kxBjT1QateeC9IZKfB5t2yMv
H+xwnWHhQA+T78R2FaAfu9vxEHYAgHPQxm+46ENrEIcWMT2tQQNNvyrwP+yLDpq/5FHgFKncDka7
O2GZVm09djA09hHbgixx/UAewYwOu+rpoAIktSixpTw4NgRL5LMoiPNrxFkr4gIOTubDceqb+Kyb
BMib6/xk35QLfX3/X3liPSGunkBCSaYwfbv48FshDjZrVrRUpaj0pr9vLXR9Qycc5Cm7hUbg5Oe+
PbMx8jys5Q02ejGu39tXjATL12FkPjUwJZc1otqH6gg5+I140kSmMNvPyxIwmNRvGao2tjQZPqDo
2ED/NzTn31u+Po5xxnAekxENG2NH7W6sYthZUpO1P9Eigfw2QtcHZGTQh/WCjYpNbNt5+ktZbWNO
vpxFvbgeXnaWDrHkgMefB+Vd7hCI+B6HpIWa6BPd7gR5srQgrcm+72RZW/m4TgC6qvPBY47Lz9nS
UbboDs8V8mUBYTSu0azVetYsQBF22NbBCTtN3sbNg+E5vsRB41/glqvVCyVdsjAmEXMQPR9qqn+a
driwi4PpLhIKzXWpgghax5V0O3/7lhIK4sONSEB49HcM1VsYYlgA9/JEl8/tFq2sA5Miuc1RUzgi
63yD/4wqhLHSj2RGjVCqMnCMokoYcxB3mShzDZr1DXvlbrQezw76cDNhzQCfufQkQ8LiVU84mNT7
eZW2jKtLW1AmCirniIlHuml9HfXAmGp6rqqXdNB2CAS8deQIS+3S3jnW0O2K4cuAolP7nXVb2bPX
8vXhqqqkstuYkDOJxVHCscPwfZhZggnvN+8WcYmPgGa5E2OSkZsHSdyT8HjXicrlNUH2gac9DoM5
yEK5bLL2pcO1e/gOz7byY4yKWgL9s59P1zFr2fQ4KEe3qQZDum3l/VkiyZP6c5XvKgp0dAbBJNck
gsBn0O+YXzCeBWkHAHabI1HoSPaBeHWznOiqaOtZHk13tRcfbODKSNZJhqc0WYbDKvAlf/yeiIKN
g8bnj9B/qNw2jRwyNa8UoCToFL+H4MniU+AQJrQhy25FtJCandQDZhntQo+6aXqYFLc1Hxp19yHf
jb0SEq69OaPzr947A7BuwgahUiX40uTC7oOU6qI13lZvjRhvhPMJi8v/jBL++e6dSrY8pJzJq2h/
4WsVj80VGt5ToQIsFakG6s2J9U/NxqqqPYS1F4WSiUgF5+kHtwrtS9qefpr1rxQfI8/kTfzSdF1c
hzxawpnl06dMhYfBhdRJmWAThYcu+cj3k/JB0i6GtWvATnD4H0yjfR4JpeSY84Rgtd+FOn8FyyLP
MDkNh3ZvVr1pzvXJDadIy1EZuTQLJvUwUlrrn3+AfMP25aC3E+PQdHFxmArXJTGluJVpAzAsaEJq
vgM64L9DzttfChN3/rS5uQ04mBcZgpBQXPS21Twbz8z+nYHd2wZa7Tph3Zf5upF0OxCh22kOVSm6
EuhQ5EpUYDyjvi2Pp/FZy67AUCOJGr4f+n5aDz1uQhRHY4fy9x6cbfJjUukzGHXCOZm4hxKY9MJ1
evZzZqAJTSpZxm+I9D4zJp6p/cD7a21M0UA++xNBpqloxK110herGE6Uz94rDeGqysCMTTMGu9Kb
+lgNmtmGDU4e80uo4nSqxmTKB/trqRvW2WDJJOc7O9qY8FaeZ9pB8SYf/8bQL84gb4Fe3hcn+Htd
C15UruwsnME0BCR8+DwkBinSz4/ra4J46+x8BPDtzrqCvAqPNWSldbHIHrFtyF3XDGkNcvvZZ18O
ohcsOb0Shy3iIgBmO26BX8AuBSW3fybnhZadT7YGl4TW1X7xm5/8foLpXI3UVm7YMxaQCmWvCEQG
eEuSS7XFC1raC2MLnKewkkVpiQ0uX9QL0HY1Low9odm/MVwiqmNXabBXeZYFnq3YxGOt+SMbFyBy
mkpa6jrnsg2SaKPMtTZ/5ClVTP4cIIDIb94FcQaUrG6XWFyx+8xNUjAlspjVHVqn73AvyifJJvYG
hRB2MUKXS1+GbdIUqW3EjrbLpb1y6DTEyCHGcYoAVDQkgHexGO0wmt+WC0/gkKPfY6tjSfNeZCE9
2uPHqdmyITRsJCVZkCNcnER4pPvO8BSjg3TuvjjApY/Y4Egg58dEU2047yIwN7O5od69ZPUoi6Gk
SeJnKynn9fkYD216HYeDQrtZVlbaWbLd5qYcf1PrVdEFtKgyPrhHSblDinbflJfxNcIgqnhVn5vF
RsVOLmCbRLyLH5eMkKufdFcgpTXUcRLbh79OaSH3A7HEWG/BPuZ5skkVSnIzhA3JcPtnpe88LAv6
X3WFrYTQlOhICXwqN+lzLxhTMgfLROmZ73lvJA3ie6sM9VmktiZq9jrKIwVk30BIbVeCCuSdm1w6
1EKkKU+8zYgXv5YuQZ0KcXnvc8fQcwOqO0ugPZE8OkwEyHticyKY266NLA0ZFTN7RhlE5jWrx99x
Q/evdbfH2dbZYRXrqbVhoYmC6mMlKmP7KDeewHAVWlijTjiPnhIm4K6ZycQy65LH/oLCQXdmqPwB
zMS+qF550CfH3bBC1ew1NJrCSuz9VQXdwU1cCTVFQRT9legFLSsSzGrjs933rserKgofnd+6T27/
sEyzxCWKSzqQHWA4abvNttBYYvq7k87uYeH+KLcWhy5mEVDiduTtlXkH2oziQSJnJA+1fKQs4W/N
SF72cZSCZMJnG/DIph2N3ecQMm7GwGfKNHlsBJIuoytvTDIaBMXBoXU2KcQ+cumvtrtTJeVz0Att
UTuFiMlRNJ3FirLlGScecs6MwQpFxnXIkcwSGq7yUrWsZfSy3Vzv0knX6QZQmng60cVknavFTPML
wgD4aj0QX/Kpn6tEqBzcDHVTjCqKqiWre3QQOMLy5N+YoMhCkOZQ/KeKBu9ahYow17eT0lf+R/Ec
9HaMjE04S8IAcY7nZy7UtfKw+SV5OT+lNCUsOOT+2ybpgoMMOfsRxGm8SwZM3xDFSfEQHypuoDiL
eeZtTnj7iztP4/H1EQEVQLVxOU2YsAMokJ749NjIqTID+WqP5F1pSmRD4ToWEXynenrHSOH2rTxi
+AAx7/bkCG4hVqSm/mZYNVEjdT3mQqFCY7+5DRv/0sPLCimbvT/0y7m2KicC5d7LUchpuJP9+Lny
OG5nm1aVhjQRmWdeou8344lUe/ZQt3e7RQKZg0zBGGBqBcL8h9F02z4M8D/BcLoupJU8cb+r/gse
ZGCWyJ8f95LuI7U+PDduZdDtZEWDq1CBGM9Y+WRvYt8Ago/3XsWRHTTeS+NLet7vu69gJGL9oaCp
sqE4u/UG7WKcHKsLrkjF+/cK13fZj7cMRGUKuAU9a89snx3uoM4QwyK8r6EOJLatkrpHTL7jMLjj
XrxYVuTLgW8hldGJuPsLSUsgsILG8kHYL1rt6IWufACC6gpk6ktwbmZouOJDVlER2gV+l0UCqy5G
CAoujzTal0KQuosrHC8IY0MCADff46nB7SYvdqQpQFWmBpJhHUuu4XXOex2vbEzwlm82GTRBu3ZY
Fb6NhdC8eJV/TjG6DiaTsCb82v0KgOLNcWx+mYI3r+qhkOFLLur+zykRytIXo7xStqVU5hl8z3St
4QbYUJ7znObiUlSBdTtQbBsm1dKUtl1Y9Ge5oEpG2XIAiPKgH3orzppzcP9GBh//JqOOMsn1DrP6
LIp9l60n6bb4i5rwJrvau68v3JEGz9aPA9Vc5QN2HJg7vgFu12yEkrTfhEVRuk5+a85Ip2tXqXww
3Z+XJG1JjHJ9DThiqylYJtsTl3P6j7ESMRnkhmS2er7A4DpI3y7J77Pvtxx8aQbErjmLuKfIReih
/CG59Sbmlvfwyq4N1VTN5wH3+hWjzWHffUoHWv6KhU4s2YzrK3sCYbtpUsYpTlY8AVQ/ckcLtt2m
FsIRDnoFxsKxJwg5bM6yJ5UKkTSEc2/J2zgNONREk6OL5U2//1SZM6S1LyhgHnfXpLjXIdRs9Dt5
9cAdJYmsRYMuUa4fz76q+874BPfqnpOgdPF1QiXQyDv1ALWsvWDbWkPnq89rsNwjXfKY13PmwLMe
cWJ+4AxregL3hZ22H+10gkkrGNbhdodpC1O75WoLatTuUmihMyufJZohVwiE/wjeMZC54myqRP9l
HK9NYUTmn5ALmmxWwySjEPwZcpgVAt3ZY4uGzOWB/7NHjgtPqeA2a2gnykExusNdusYdFgSesnDk
/91/wsNl30s22/uSoQ/lS7QS9NINfM2nVI9Y36Ba52amHN6H8LdFxP9tKcAuxEo889UG6aB2bpqo
jK2X8UNBuf+8X3M2uFyXnqP1NjjwG89KRMQKTObjb/EYtYqQA9dU3j5if/LPSkHjePMFnBgL/PH1
STdHZke1I7VS25nG0tiOHDT6caOsEJSX76zzpdFFapg9shAtBLWmw5m6WIs12uq5L/gAmLiHBIyP
/ndWAaE2LRv3sxgiG1Bdka4ouXheIe1nfIPXgmtXRioSOD5xyfR3pmObHb3a+ow9WIjjHwRh+ULM
nqeu9L6qoOujuGLUAfbxoTI+6FMGZlEeRavYAp8BfUU+ov55Itldv8UwU9zkfHS5N0uV8ijX6piA
54KIdAtV8Obxa4D/TjKrYIgp76adWfVEwK1F5cGqEaHph3s3zFUOr8vW3IS8pIqpspmAl9YsC1aE
XZ47Dom6HVVIqeGoIMxPZI6oycGbEL+UCgETR6yjWqkqFTleM4GyJuUS1IhzSdCxz77+Lqg5oo0T
m9TKKmjgpYQgZW0oPZRmgoZ/gL1wmAbu81jA5LFNPA1GLWQbVwtNTW0Yl8NFSLXDO7hdLh20hbyA
uPG16pN+aP/x0D89sgsVaXekl7Oxnjt6YWTutLn9dOjshgI1EC/9vD3xDYLlbHkqNc99KmwBCcta
AmFj5vqRzajEwUvRbWMvgsQ5dHL7AtTpogIG5iuCcNbm8MyFRASZEUTP/Wn333dtfdZ0v/pn6fQj
s2IkA0Y1i9EtFwqq77+qTBeYiDJSpsUqYem6Xs6ma6gQHc8rvLYi8Qy52W6KKJfHZnFz7TXlA2VD
bOz2wbgs7P/JLMA7Efr2l+V6TG12Jj3j29uNd3cCyrdqrZbZv8PCP/P9dq+T7kiycKLUMLZDD+HR
KO5JYBHuMp4/a6faC6nY9aw7/PcTBbXWdO7DUwSVqgoEQlEl25mf+E/k7efCusIM8Du+3/ldBWVm
n9UNXx3cpbNDFvP9vi6ivIHXXf46kocFpMh8z7Q6E+F60ZPAE2S2tPh3yhwXeK2bRnAktvfapKRN
5a5dnSMfzQ2bTQPc4AE2+05yJ2Y1M49mGwFyKBqg6SrUQOgrm8h7qzgrSPzMKNaIAqaNGE44qzjX
HOHFG4Z7BUhEmom840fDKfuvxa2GISrvAfZ1E/DNKnRA9wEnsL2i5EXYeOfhbLs7Nm5l7AHhZ1v/
5q8P5BcU8QCldPvyeK0z0/CLUY4GnzUJvln6IgiZBjIndT1uAdXEu5EDJxQoCFfWHbq19C/jIems
u220BuglCRPwoL1vMKjH0EYL0qCLFt3skDF+HB0CVKZADLkZWawhOUnsbB4O13pUX6eldvKcdWil
eik1Sbh0KLtpZ8Qhs648+1d2sTxIaFjJDULUDHmEf2v/1NM1H2P7eFklJ3cJXjfmWTn4Y7emIPSc
DCDevg+QjRVlrOr6PuMj0mZd8kHLV5QInEuaMh1rfXWdZL2RS9g+xPdxFVI4Ze97uu64+7QvZBuX
eeJR2EPPMuXiYqTXfgv3AF0s2ks2qc9L3+tTIGj0W1WJQ1ULciIzZ40q8SLwep4IG4qLPvF4XRmT
Z/2knN8S1iyLNY3Yj6924t3TH0QTDr3KSWOE8n3FSO2f4woZzX5juKkazK4TM+BxfOs48CufKkaP
yyvO+AGZu3mg/xoko4eCBielbDG4v52zIOXqIXarFmyNfJox1HPOriXKMOHoDn6vXhR3xylU3dr8
WZm0IDkqanph6AvyCTq3vIQuiyA0GI3ywHeD/AC2ngpLUMv9xrk6zz53s55B1mth0M+/QX58uVef
Hsq44YfRgyezL8ECqQFdKmL1xenHNk6Mxz3eV8MdDLE11CwsY+2FxNj8KfcFOBpm0JM9PUvywq0/
9nqfYaTzRhbeXujPi9ih8gJkD/LYaX7EBghtVrxyjq9WeklkK69qIv82fDlSUOWFye8m1qYo//FS
rsE1+85BVzRHS63J3bHKwndMxHjY9vYXloP6pTt9Rwn2E4mMTPGdY9DxqsWrcNaNnT8+sZ4PRyO8
XBVaJIDUgqodrAgle+6arv0rZBFdOIzinh7HqvwGKVv4BViLaPtXrSec7Pq9ICaAaN6YzOZDrO35
65ZRzo8df6CbFznY71pTuDNXBI1XP/uM4TzdYfrszJvbuh0C9BDFvtveLEIdG2BCOT/Gg8Pqji35
grt8PzfFn6S7D/vThBcDl38aFTLsHxKeaE8BSabXRto08+719hORpz7B6Qi3wDZogyFP+ckpbnmh
/ySvNjLflrF13P5kN0l/Z9NBrwFHMDSRxrYKEQ1qYgZf5lCx8hiD6elir+XF7eavMbmKXAbGA/L9
YxtXEzQCWJuNrFs5KOQRX1UFwzAxxvGKqUn0+8uNI2ZLCR8NstXG6p24IJ8ZkHjsjsuH2wxlj1OW
4MJzCSubPYtl1px0PQUY97BIm5uJ5l+c2P8X3qrPM+GEJuwENrHDcQ80LQ2Pnh7MMD2G0gatW27V
kJMBYp5pG4ZiQjB1/2y/DHZODlz+wqLHoBPW2p+iQkz5adXADluV6IQLk56RQjXDQBm7AYcRA3m4
eQf7CO37ad7R4Tyl0O1AiEDuEl4bKTcsv5VQS6tunk/Jyb12VcdtdfHCpw9rYrn6rbOLVvpiktqk
kz9Naw1k//qBgSZB061qIYa9+JkU6JM5O7iBgSHIHvijwRkRldGb3P6W3vIs7H/6ZOgaqSlFJHha
B/uEcWKMzXmWPqtGSmcRCzgZguVuRtYtXqhHzj+xfv8SFkdP9vlvjADKlAHZ6X95fNr/mFKn4dKS
taSUH3GzWUIP6yKdpSZ66sgx60OG1mb3HKabo0YRwX+J/NWdsEytogIqZrwQl9A4gpelsqL/U/CH
7wpRJ78pLw0sUG3s0Jyq43DRoaCArqsL8209nun7OVMWKgQs9oMu9gfSg8wY/BrmU8OeQPicC/NU
bqYG0b1Q/TngpAiJswcb0T/0RZ8MOpXTrFWAvk21/021zRFdLDliGa1Rh/uCQQ1R6tZukEoLVM4K
Bul8Vw/34BbR+ZJY/NAMiuHlN+NQ6riO3SPXSWcESdKH4UM2nXIvbt2xMntz/ycUJ1XjIUSSr1ps
VbDkH6NQi68P7UuB4H2Am45sSj49aNGDafg/VSzWXt03hwKz1K4mLX0Nm44VdgWuwRkbtfTtnVY7
ZRTeF5FoQ2ThH56Nm5Oc0BLx595+o7Fc5e3jMJNQACq2saftJ6EBFYSV38ycUpQuMSjYkyAjVsk+
1NrTuUOquVswqQqT1Mh5XEVG9BiORVyl+6/ceQ6/dSMCE2bbDJt8HjOPsGgAUKYllFyVTSAW084f
Y4RI+dGDsbNlG8RZrQL5lbfywTiiHquCouRuqSJRp0NZHOetaBw4a6wtkTPi/Ersolfq0ZUcQHvx
y5mD8vPnH8h/7UWrEH9mZRnJgBz/QbW0eLlZuAOLrGGh5N27yqtjLVtpCBfTy8aaj4adqOROt39M
C+i+AkG8DZz686NqYNfdi7fWXtuQJct23XIgqurprNaacmSvBBpMJT3Na/fQEuuSUptKY9m/2VH2
0sngTMv+Ta7/U292tGeW+Z43+e7/DI+Kr6lvYjOh0VW1tYWVH2cBaQxWn81Ccuj4IFltlC6QJm+u
7Eu2c+p/wRzeyWCJouzPyy+D23br6CvJlplxkTUtK8k/2QfLXe3cdI2HtlE5WpN+jlZd1ERGo1Zc
mWjItFeZThL5lszTvvrtUlZ6Ol6kZe9aOKt0NxcVjpT9NaQ+H3kw37ApBBzeDXE7ZrY82lL9ZGn6
SHM1AUye/4Mv9stbLdriKZ9YUdV/J05vTWZk6Un/kjPoNWNQm9/yhrV76xA+eLF7dUBIoIGlKyb5
ptuoxG/PW/HhuOEzZeeEF4k178pEPElPhJDonAOdp7q5MYJZkyhBJpk6fRxeQB5atC36vuEqhHrh
BmwG+lLLac6wXWVgWTmos+wUGc28NBXm41l7sE3L5um5Y6K04KLelJYpEukrckgLCNAL0usY/RAr
/IPlkgfjA6WSq4v8/uOmjwSQFBniRQ72srXR7LItvL3pMc9VcpUWqC57nAJj3mN8Tvws6NVxzwE9
vfY90HxIq78zbFIbE3V/t+jfTccqsQD7vzxSGFcB+cociBnpg6IPtFIaF5QtZAEMBMpEQYpHAJaA
GKZacrVLZTt16t0NGeXZYksYgeKo6PLPhTwFB/nGRRL098RjzXbMGv5UuCaKz6oajJhig6ztyUCg
4Tq1rcDKTiWsAsFqcFjS8UI6PQrd7Lfc000p2oTgDyyr7WDrciXP9CKy1bbW2NkfBNp+I1CL4F+o
Ccz+ilpT5D9VLypAwrDZ6ziI9/zFebOCqpGtTVPyn0Lyh//8aokoOD96n5NRG9iBspxR7W5rTMNF
aMElLVfrhZSLaolXb15/zspHHhjw1ZyDCpZlNLrxBN9Uq/THRxMS9LNxYGJfVuZdf11LWNlf9iEe
6LkYG3QOIxd+OnzVZ8IPOzkORWin5DXPsvg4qN7hETd6Z+fURtaY228xw6UrC28DYzlVfXU/D3jA
BI5/0DlXITyvMu/Do/EknfraVUMfMgCwusVLIY47MYNh311EOz4Uj3d6nCY0wPUPOi8oqzZctaab
qCeTysHi4dSq9SaR/b4v07yoWqe282LV9wfvH2rgqIygRe4naD5psp7LLEpbDaggYnVff7+aO597
eXM9d/T//dSC1kRpA1n1Yj2N2Q8yb4US4V12CzLa79sCcFeSurFBK5ZfTZBOSVW5XUnBGv+mNeVO
r+TJpncnjGwgY4TxhZSsf5o2w5lKzZj1YJFLvMB2mZYg58Zidal392xJjLtkUeQEQFQT+jQGwsxg
GZ2FlOuziw3ZwjQCDqI06SjMwRvmc0U1hEcJNRrM89mTuyUqfukX+UJ8TiCEjfWGu/AOd6fVO0x4
XWFNBJrM/YGMEI6iw+YojLd2y61EH2dTMaC1biwODKcus7KmiNohcvXdw9aIz3l0Vx8Oh81R/p/0
+C9gJbRd7jmYqv6kXQl57XePnNY7r4GQfiJu09jhKupg7i1hFPdSp/hd/cwg3w8Q3j1PuUiZdPLW
xrxSOxWFlB69z1CeOT5jJRrr7JmUTCkSwKBYckAhzvl/Vw1T8ynS3DKkANqW3vxtdRnxV2MiCKg/
cO79PHGOAHDaI9YzUdMR5Lc0ZG5BejHbTG/cOQPi6NF5lNXrTWelsb1BJEOWwx1MTH68ajRJ/Jtz
0QheZd8usSxp+y0MiOMMLZdoUacx6mGfCdsEJdlRY0RFOSdi/HzD5Tj7AN3Khhh4nNHuSwb8sUkk
3Yw6dT+yTqqaE5GHx4DNQ2ATWxYSmgFiBffIZDbyDh9i/+ws2DydtDUcwd+HX8WbBN+wOq8hCA/3
LotaNP3Eo6wMvrveorx6dvhcT9lx6wH0y+EeR1Ng2mtEOjxUtyfcRPhhu02OflG4CUgScfEJiX5G
jXZ3Z/BYZsdUknjZwfpJo8Omf5YjQct7ZZUG0zO2yGW4amg14IHuLYE44sRofYsw3Q9o1fsRwjw6
OBDop29LKWoRJ1Xmh3S4WH7dAMsRXIGJUVXH21PiP7ZFfAEhdHFigMJdpuXKXWv01qZXiumoMpv4
wQdA9DV0EDfZfqPG0V3GEvGqKsgZE4c1MzlZe0bktNt5Vcmj82rr/dR1RSi158hocpkXlZQkxud+
oURYYOve915erHorh3TFtUQ6qEPelXNvmKszfU6ig3433pIr7PIEk1F6VpoQKvIq66Kmr5ibp7do
w/De/ADgpllxG2gmrQgTQC+qgWZ1zhjlP9POCq47lGVTIM4fk3sZakbYHe4P/IfG+1E6nWQJPiy4
pkm1EynQhjyr2yXgARS8lh73yt8QN8+aXGTzBDokL6cd1ordK/O68vStvT4u3TvS6itfVwBlU19D
Nek7W0TeCgluwsPifhm/w425HCsScpgUgBtv7pOPArFji7C6JuF0qOAf6KI+iI+AYLepFw2hpp4H
gZPCghrQphqEXu81Z7VDRId71J25ZowBRM2RmGYoHG/sWR0VhouT/0o/gAFi4rVMG7k8uHEvVDgo
GNOXoUVaNBfipBTSGOlj3kMUdh8kcyaj8VLN9mDGIGuvY9nUR0NOjI+BR52VTJciC1c9Hb7PZU+i
3XeeSxvLKVDc7l0eqTVcqjadzrf6CHJdlDnIBOU4FthkwrJvY6b/A8VppGmExsrf+wGFVy84EShN
CtjohSc3lz9OF7a5UultAKubtzY0xTEeB9Qitb9HT4lv4pxshYpBwj3zguwM0/2nFbLmF1i/sVfb
IdR0OWbdtUAovIBUGInBaK+JvCrtD1WQzBEHnHvk4kUFxct+n7Rdxe1txsS9LLEB6lZwp8g8P7q2
+Xf2VTjEfJQsAIQiYnHvm5GUourB8fRAQkloNTnLU61DIjln+YPG4TbtRuF6xPx2Qy43oIxLvMB4
c09govWAk49jjYJQvVFV/MvAX6/T7MigcG79BniZqi9dzDQQBZJt/CrnQcLeOtWHKsUTl+bhgNuR
TKLwR06C+JFzFILZs9mcy2LHdFq4rUj8GYbX2tTBxB8DwdrzhlzR2a7gm2k7NCuZn+Ifsj/gZvmx
HQ+7rQgzz9SMyJbF+qyZwCFJxQa9VYtAv8We12qCbZpAstWU2ZL/sKNBRQO15/sRJAQNUVZr3bOT
+kzLZ4YYhxxc9StMmMkZMuTpzY8lKdSgK6fwNxDWSofGSVeuPbZIczm+uJTJO1CLXoUP9evsxig/
DqXvSGHL9YOcx3i4GfLvB5ESI5W1DbO4A1Gvr1SYiv8/rgkZwhDlzjJ7nU9FSnbieesRAExSKPof
pKN1iob8ccNJBOioz9ZsOfwFjMuweKqF+lM4ikAAV3AZ+pfE9Oa5X0LOWQU60PngzZjVhnKrDs0q
B0RWQR76JeWBprb00aDVHESnkBtyDQsaqdXqyL5rmMTMTWwS+BR0qFc3qnwdjRfynaqzRmRM7c5Y
Ypemmp9/LJMFY/CBm19g+ZIq7tP3whbE6IQVR5JFaFkIvsZ2jsVhxvgKu9wIa65fajF2rv0el3Nu
9bF+TduAa4aJcs+nwQbi1ZaxVVwbl1jL/fOOfJN5arliWrf8keI6SKrgB8IolhWUi+E9nWqMsNgH
BxtwokzwO4Cqqo11vmwlPF1+8N/49Z6mbjmFJ4apVgKpVO1BoLbLqQelA00YO+QPzaGwp7TjAr7o
BLlPDU/ra2DvwpxtD4eHYRWcOXHFxaS/lHLiAl7y71SukT6zVumalqMvPkt0XfyESDqfhSKFB8mS
XT/D2n4qdblBqtXmzPDSygyZBTmuyCAiw58EVJjzorzk3zsj1A+YfeKrzjuZDcBUTz7l2m3aaz/k
0sD/KrH8rK1Yywmw1fGBVSLVNUTTDLEuqxH2P/BTzfycs844OQoXAdkX7Hfvnk65BIcau6cgR59o
K9oiJaXjnflBoboTnCl7WrWeB2byT079V3oKMcmgW+m6R/JKQPlW7/Y5M409qJAd1g+/itzww8Jd
ZbHfvjSa313qSyH1yYDhl5OJr17fFNZZsPsAt4rt3PLVj8YNnchuE+Mu0l9us8ushJ55582/TLU1
CN7QWA2VBMHj6d0BYPAGEYsdRbvxvTdXieegJ32M8cUo9ms56cdNN8WLWxoMxmfY3JvgefvNWM0y
tcfI25Av0pAYAf4a5uy8gG4eijF7Bhsf1xrXMyxhmrnHBlhPR8RwRGByZp40+ZCLGt4m4SFpY8h/
Fo9rOGxxgqt8CcgsZ476LDJ/RMZ8C97yzW79KinA/uEFlai8gla03XB79gR3PwWloPCRww2ciqTd
SQzUNqmHZE6Fl3KbhuN/cb3id1iXPzowbO7tMHA3NgZLN0AgxI1KZlDZN7DYTQ7ecmaQbsboIZdq
znqXaunF3ERtUty/G9/oHmP39CBqBqORmS0kB7xaz099hEFM3EklpuO7xPYCsgSQkZ3GARnmZ9BE
J+NR5skUyASHrPsCS3r5JjizcSUxpVnt7+uH1zok5LoPHysLFO9X6k6+gklxq2bxjglkZOnJ5Pbv
XTKIuI2wEmaiyXSRxln9MeQaN4XJG8NT5ibRoVCKIqqwy4Qm2Y3JIFWsUCyd9JbKE7QCjsu21Kfu
6V+Q9AdljNKJkfWaNubutSNsr11gJ6qAf+hUmUdW6hjUQNmHnGk1VNycA15URDwPY1QxWv6j36OK
zWQc7VdF3RieRiN9vn1DonP4A07E1VsN5O45ou970JHQNKcS9qzQIIo8/55uMTuKd0lAfCmvnJQ7
dPIm5Q5VMUaO2Vope+rQYMuYw0hIVlcpR6b5oLklrsxtj6e3tj/jTmdLRdsSSbHU/4gDiW0/7nnT
Zleii7/pXTQH7bU6sbHnTrEMEPM1iZ0F0iCVxyXnoXlrHRnsFwkneCb4xN2jGrE4GX+euwyY1IXe
H6k+zLET7pEZJAB5g3OpsSWZuC2CdqZglXe70cVA2KIXKy0Y16ojo+1eNbByaPrtuVnEn2mqGcnf
+i7wfyYpvsz208eV3b57nvroSrLAVTG177gp56AVcj3guG6clNepN06ylUPDexFbPOCqFd3dB7Yu
gmtAm+HApgPXOTNuMZmxvtS0yIIPcmdVtmnYMgDM0x4XPfOa+7oYb/6h8C0dfbXGTaWvgTj+op6f
MKBOVlmv+fuuPrYPgiiJ92o+a2UKNTYTZFOqfLmXUk6tEQx+mYjkhmTQQpOOFO3+2aeG44Z58Q1j
nZJtZZBLzkAFvbG98U5ZkzvQU4yVDLY+114adqjfjeWtafU4KwAJHSD7AfGaoYfqnEsXeT8IvtcI
hzDS3wjdR4JgKEe6KWTLqVr5Lj/xjvBHFt+Akvw859bqg3mRJ2IK3P0bUZ7rgkWHDEGW6btvFjNQ
pO6LPssUeomiUIwpU+cOXiLUPB7wG7RF1iFUM00oiYIdYMpXtq7nhHMsqr5pbsvP4AMpF7qQlVv/
WURZ41F5RaM2JpoWDZ9DsXJgdAVi2cKAWrH/RKIigH4fWNZIRXkj/FotFUURx9TFo7DU6EhM2668
IjEtLm465qxlSEwC1o26TN01xWgOpypKZsr+hZgiMR7GVhxdL9C8QDvPwkC6Y49KHRXlSz85/flG
mpcfqq1HtD8zFNnyBwmSGxcFR8bWqjnFUs3uz43JQGp4Wmj92v7FpH1yqd0o3yv47k8bGS9w3e+q
zkUa9QjF3ga0TVj1OxiADEq0G/oj7Uh9bb0xHkj3m0sPdQBnFb6LaMQ1IV4IPxq0jly9jh8SjgwC
s6iyURcfn4+33WR7g1EHyqH/IhIRG4u6Rk4L3CsYm7xNDOm6X9KogWBop1hoVPiBwNh9l+UrSPkq
oC/1YUGmzSnTZtarYboDGLtTIbV55B32plbJ+LBbG5PB5r39uR5NzZGq5AI7XG/hx6/fIqZFS+GN
o20rD//upVrtNNYilreJtVHDisj09QzYM46YnOw/NqHb4nYCRzNo7b67dJRVeHnd4dPdRwGLGqfR
oCF58A+QeLPaYgAcMe3Sd9qUnis3O2QDVWvve0pGIMbDe4OJzj2hp0haY47r/ogBAl2LWQFzH8Yg
ve5WmxA8jW2mOas2b/HsbCjO9ojJ7++/vvzzx7DERw7XnqGGdsnEiRtu1jA+pQLUPsNPi6b4ly7g
eD/Yz3YaKE4QJzlTI0FV2vKxgCy7NCrcUttdroZdvfxC6uVmo1p4td/vHW+K7FttlhQsGzCG9O1Y
kKpxPvASmkUlVrG/Pe7G5gCgM8eT1iY+yqqzyn4GuHjkODTzmFE5Ijp9FN/Vss+YmlUGjfGBezho
vnrE1sS8G0ES8+/mdJgmNkXtqlefOII3l1plZSBo0HsxemoWvLEVtJCMJfzDV2Lh7FanQ700LvfM
Xvfynjifb1yxXmsnFyU1mUgBgK3iMyp2ErEdFcm9T9wmR3uORUvwac0/dJmrIjsuaR3I9PiMHfwR
qIHqCjFER91BvG0HeJPOh505sz+bal8K8i1jssALpBYY3aBiXk8oVx6ywLBxZ0KIfkZ901mF7ABq
oYF72YvS1qQvZsQwmlFc1Bm14WNuhe9Yh2xeWkVSlqldrlDqMPfESbiFRrHdbAjvxNUj4oYnUyT9
Wv2D/GR/do+kQ1pM37xtlkHfcCOM95cNG2+Uv6aj96FZtjcjFwTy0t6/hZLQ+6TqXlKZiuOKChM3
pPQuAhI196mE8tnU2JNx6tHE2Te0kYJTG5OtMsc4tyUOta1LkzTj5XeI3ipeix9EB4VM9/FfQsdU
WG2dDF7vofYjrolxG7Sw2DEmFyAtbeckLOavizRDt8c7BbjxwMM8dJjaoRxviseWWX/kcDVOYrV1
BtS5iR9ImVpPZrGk77r7gYvSauh5oORE55dy7vd3Ywuy7etFDa+pKrJmlYJ3AtK+HtdHxSjQH3QZ
TAgjYgeXN3N2YZm1WvN3W1k8kA/uDNA6KDPJW0JqPv+qi+f/60yQdV/hMhy0mcs3lbEqhmwui970
nwR3DPy337/kEW4arP6/sAaH5CyryEr6+9m/u0hB4dNwi2oBfkVdusX3HXjtrw5UJhmEk/pNnyDG
+AxtSRtN3/PCJM3beFXaESB3dXlKdips8dYqhL3x6dZpcDc/M65+4RYHPskPpptW/1iGLC9WlX3O
lHZzoZvdqfrIVmOEvUxQiwoGe792zdGPzwT++/x32l/ZvG8aaTnaBmrT/FIezkk89SckpMpu2odX
+eP2w0+fjTJs+IFhrtHgZgJtGJiWsK6KZ+Qyg9I9aymrXDj3p4EWlqA84WA9bXCe8yEayC+62WXC
kPV7/9UY3VQ70NEDoVRirAP/Gm1HlBJWfRo0L9eIErEXMG3HGX1SLtqCVd1dJxSA/zp6BDs5xcc9
dhVsmyOpohsP1RUpNiO4SHXvcCA0zP5VYT3tRD+M2lpXWLJ3iwlTBKlgYyAZH77ME7PYKIxhd8xO
jg+sYMmlpodKKtcIhkNYTUrG3QbUX5GY0dMGBsQ6/FP1e01NjEARzRhdDYr9RGBaFsCmKTAShaXs
rUyDSVBfP2BxMEsk77USrB9DOx6SM7QZPYqrV/GqrNLwxturJ2JnKv5a/qxlwa4MYtqYcxbpH3EN
qfd2MNnQp16JN1y7mRUuNS2JmngA71TKVXgh2ZuqcQ+NheA7SlbNsji2Cu2XvijRjTIqw3KyAKm2
VuGmbw5psph6QGtFtMxdr9b/SwT0P9QO5QD5F3pouaXBdGPHM624Fkvx5g9WQt8xO8a3ZdVY22d+
Eff/JbDhS9AlI96Fe8MkCGkI4BIXqJ7Xk0Ubo5nKdtoVx+Jm0cI5aah49qNr00krz45MxITxdr2R
/8/nddon6n870KCr5ct2QDX8F4PhFZCV8bZ62KsqBVnfcqchDhphNUOjwK5N4WK0jayU2hKpx6cC
mH7JRO1fr1FKDIjDoDjbbZKX1nHMadDVIW8al/9ot9Gsby0qR3xnOrIc+4uYmOodF9hOi2RxF5Do
hRaDIP6i+QtDbV/TugYalXqOGwPceGKOXA4/zztoLPTCZYTfCHO8/DWyPu2X8Eqq2G/pa+oZmodo
kJ8BpdRHdPOZKPqIfXdlJsLOnq8devFZSZJ+TjerUmqYHSuDsRskJM/KO9Hdhq6R1xcNTR8lTsDy
nYzVKDzgIvRPfiHbQRsymLkZ8fndRYIk5gIaa82j15Sni8nkMsO14PNxERgzUZaoROIIYP4ek7fw
RZgtULZbZ5ZIoK/Bo6A+QM+FmOrKCGifvsZnIOFoiwKA8JCEoyGyemMXRi+hUgXexBsDjGaSAxDv
IjM0bOhRtLfaCpkOV58afE9KrsyPeVEcfi0/5bkyMaxi7M8qwyTbswg67oFVZ/EGFRS7Uzsu1Jfs
m8kKP4Vilqi0w49fsbwxDvDUoqP+6jXvPsj4nHteHgNYOI2+IHNtnKC1hhxlT526rQtpC6BEE23U
SI5I/liq/IdEbljpDtvQlwPCVAjrCkH+CIaImMnLnjTM10PgaWzz4H9PxqAQvvIhjjwBV8wwWEVm
gvPDr8ediCASxEWX/ZixOP+vbEH+kWqmskymF2rco0snA65x6dhFHJVtwmjxhj/Qj8rzO2igt5/U
H6Ao7O4KoHP09tzysooKN0he4NMSBME6MfS3YIXS3OPrDq2KcEuzSXIm+kaBBxV+Mvv+N7/dcF5q
kwnrqLCQEMmZMbkB9oeBm28xEYJhOklTZ6bwiNtAIFsqOPCmf0PvW9eNQzdN2mkaZlHKWLX2txjS
r5KniekznJASTkiPU2Sa/CYiEDtnbRutHQ/zOVLeZXbv3h4fl0/dYLPqGFRp6sqVqfptuPmPpR8P
aJ21KRLdShvm1tcqLuLgMnwlBzuqhZgCW3jxFCJvY7fXfzfl8U9W3YAnlv25kxBUtulZSn1QZuAt
8p2L0yRVM1bYi7fRJUO9OBNe3AyxrzaziTlnRGkc3vp/SBF4Qx9Qa8VsrWlj6A4QhIFIDow/eSlC
G6JyF/eefolfSECzuE2iMjCEaMVaz+QKPGhU/nzTGKSq/54eHOtHsbAD+G8MLGkOP4dmuIP1ZydI
iYd+kJp+jsPZPfjSK2lTYRhxeAh1kuDIqq2H9gywKM2qeX4r+J7ZsSNEgf2CuElpf7JeaCbCNK56
hebCQ0w4M/BzGeTgo7OqeBuKQE1LMwVbuNwIOC79y0WfWKB/QWgoaoz5YLKcjhf2xziym65IWU9j
GzmqNlJd+/9EaXMHI98TIORRgWqXpDKth0+mOah3E51Udhqo58aGORCqb6MUx8Yt3/lbtCzHs8JX
CFeEdZe4A8/dSkfYwoRJG7AOBDyE5v9uWUFoLBlnuqPTemPDNW5PiLus9c2HEHOWTo0r2i/7iAFa
0SA/HX9RfwcWIQufx6XEktcBd3wRaE9C8QvskcnAb6pqN7GQCU6MxiXICfu3IvG6kujf7IV8YMVg
Fmt/eitkC56D/SQKAKDMm97ird4B1ERa8f2CBqoPbUpT0wt2CbzuNYijZlLnSnFWLhE8I6rqHwij
hv8mb8W4XRJqDSQc0+RTE30vIW++jF2AWWgLyMwBemNDoam96F7o6NlFKtyV8RWNIFQicTCsLSrP
QTHnRF8v6fFKOFpq63hHE6Z9zmFdAEsw9wxEIYBPg4+I0atHnLEJR9SBrtgtR52U1tMfBgDehAD5
OndbAKsAkRZ8hmLNMcxzVMEwTisQLXKVxVk06AoYML94/wPmtadNKEAR2ZoVmfSoL9vgmL0xQbMO
g/updNSMS/hCkHMeBVsqlJL7LGQ38dt6htF2OX6Yh4RgCl9D4JZ7R76AkqJr9z/vd8s0Q5w0UFrz
mgkZ1gZpcAfFrSkZjCEcTAuAzLdmlXTA1aqpxSGhrYwxdpLzP3dtkqIRajEtbErKfLAw0yJerFCa
MSecAH8TPB0rAnVy+/HQOAp66SofNhE39ydU2uedDMraCm9oeQsxhyM9Be2/V+Fe/J0CPb1oNXol
Ca6T6WIrMNMqaoOajbVWHi2XJ/ynLVhKk4j3ZbSTBYAGS/lgJp1bAas1G1VknGk5h6zDrWascLv/
7Gmvh9owZU2p+jpK3mBSkhayI0aGqHGDkwukHPzeK0c7FW3cIsBk8agHXnjA4NS8ixoZTO0EHRTm
YUdCwQj7lHIpGBYWqwVIFTs6q/M8xpHywQltK5DoS/XKFaFMNEivhKvbDaW2mJyb0cLv7q5vHRCs
3q5f4k5Unryo1qQUY9e1MGhvyyQ51HyNYhoKqbmekCylvNDKs19C7OZR1E8TyvH1TtNOl14r3MiJ
9Npsqc2RVthrK+aviheC35ZLXllVhzuHCaL/owQWI+Vsk9zeN963ZGWb0v+Ft8s5O9MO2rF4rpxS
UzP8sJr4INDJEbG62fJ2/zLJwmPl3qUcBFkA3/xNSF4LSU0uLRngk6x933s7z0O4L/oKr58lYTDs
tIHdjOS6KZl/By+G1ep7r7M8DoHj0I3ZKE6LePjNY3DX0RZ6L96qOa/6p/3FLASwwOFpvfpOZr/F
QyuG27XpOHcTXV8mh1tB+/7L0eH/YbiOcxA73JHJU3whLy+SbevP3gqtNiRC4YBIOtdx1GP/XW3S
qQmVarNdW0fZDBv9d14rGcvMVit5PBYbuMWWt3gguBbpLu7j86SehNXhfOcYNFmtKNvlf9u66LkV
kKpQ03018A2H506Uf/8d4JYyjqGHYE9dOXjHjfxWBLA+KVqaImwb56B/3uetiG5A5bkPHyUNt4K/
A8Oif1B3ZafjWjy1qWadbJvIUabW2VCwVK5r7zX9AeymHAJtodfFPWZUeNnVWTiEKfd9hHHh1udf
MVUlhlYefVP160rKEe4ZDaF2pFfv9cn6iKXnNAgzPjKJ8rX0KjSasmvWlNKy9iqivR8SY6Rru52c
MwCknkmit2T273O6+fYpr5NxSZ590JJHG3boU+Ja7joTFE2/6CbYWBW2op/Gd/urMFidpscnD4yK
ud2jvboafSPEsvrypDHRZGVVuOb1iE3OMyeYNTEtmZSvxYcBqLP3pi6aaOEVZa5kLy4ugmpPrvwz
QSZF+qHVIjDd0KlXY8Ia7olabZu0r9gxNjr3aJ4rpsFnO9C75tl5Cla/mLyY/o3Vo/E/rSFISVUM
QEPP4q8u3XF0oetliT7kzeGVv1ZYueC9euf22wLqau3a7vAUtIvtD0OT329P8aFNHtEXUKgSZgtk
K8BMrWO8HQJQ1wzb/5MQU7BQ773TSc5nU2ebPSwrq/WBW31ofKf7DYQNd2p70KCH0OIaibJMnID1
jlxraO6ooiUTBWap9SuKT8QKGNHkjllUCXYoUv0t4xGByIhvfaFev1IJCrRBaAOlRJpArwQKQB0G
wRefrSOfcJNVIyxnp51yY+kAeHZ38ef+dx/CG4m/QENbw63SDc/ypb+Q1WzOsQlPp9OzC3OKy5Ln
9UEMC5omVTGKVWWbUoqIW03Z6yvhW/Oep5FOMTa1VQp3HVUoJQ5FRxEXXkzMyBMS6twB73Pjl3SW
6my7Tya0LOPunRSr/S38HSM91df8R1IAlUjyVjsrXIQQZqCcxEGsv7lZwQnsJ6lep/+Rf/LqA2m/
FE+jSKGdOI0/c92Cthjm78XMV6UCPuzLlpj3BAeyicrjCKTZYjVsncVDddvCHXqCwqcFAkU4uLD/
HqFpSYxfd1Byf0uQrsPxK7/lWzWm+p7kEB901/9tLKz+zQdwUaND3EhoSb4D+BNFK7lnLz8Oj+gm
slnzP9RLK1eOS0GOBbKHwTeR+up/2lHmG32E2aGJpCeX1cGMnO9b25J7W7n6+UIv27PKFVBrrU7Y
JvRO8iwVYxPZzBAJzP5PqRECEIefyehCwgNlTSB+d5MqV9opk34C/2m9ICS4F2/FallZhMW5VO0E
fFx2N+Ms7L6kGncEZpYOd/Vg5+mqGJ3X/Za7BP5tSZ/FXEXPPT5nNLXuIXybCGVaRgYlB6uO44xD
YTbgDlizzgjBtHgo1LSdrAspyaNHEC14lo/G3DYiyl3Dxr1rdb8ZoRTIeQo6Puis5ymnyskF2I6W
6sgEfgGIKarf02VcwjBpy1iI+pvnI1sAG88/pluaCmuD56iWo+cX+vKdKUeJduCFV6A39al4Fqe3
a5CrJco6LjLoawL2Nr5D/3SPzzDSg/LdvCYrVowyYQgEQwEgQLHQgWIWefsABG8b90Rs86sWtwyD
o6qK6WqjlVMVEQgS2TNpVZ+W2LD/SA62jAQeBYaStSOeJSnybHbETUhx+ChjfbrPPOiL50Zo6Vgu
IngUTF+x3XdR1W3D1tzJJ9fMBydP0r32mE0ao+jJ/6Rw4hkxeXpNVWnEYE0zXIVhsiyVTWI8m2gQ
9eNj1Ta9OQZ1bYMfjfZGgH3wInQ3gi1K4RYkRaX6SudhoXooR53O08uzwPFMg1HFdIQEeDeSgaUP
xyoXH+OGGDTqTRPH9kXSAcPlywf3voPTG9TSCgY6fxN4rEk5I+1hewLw9v1P87CkZlkp62wRJB8B
F1w+AtdC6nLSglWif6pLA6WpZkyxI1IlFsBbZPit9aPCCR2WT9t0QLVEgFYHby5hu/QqVJHY5JGf
i7zUZf0JuJaigJAoS1bEyFVaJiJGVJMn3h6D9zmr5LjTZMil5G9rgBSz/Fnr7wJE6p0SYg51AQ5n
vLvhNaTnLk9bZlwxhL4+3O9b2wmGbAXrHcgzFMJoKeHD9w5sMalG1FGb16VlgeXFf2CaXGUGmCbp
ywty3JCoInxZIId3UVlShmkytOclmDVGrK05UxO8qOCBJ73X089KcN+7ZBuGhRJBvWrEReYA2lhr
OpYLeGVl+vJzFIL/H7rABCbNUyYrJhxqLapjfVWxtj08H4ABidyNZfUlbXSVHuqHoT6L8P2a+Oml
HA/nw8ZqsM37rDuqLaMWmDnvuZceTsp58WbwYlmzCdVm2ULX/ljzkZ0qiSo5k5NGrBLu/PeDHbWK
Afuot1E6mS3Dau1NBpFCsSFCVsFLR3DLnQgXwuWosgz2LfjZB0IHF9Nm9MA7e662tgcXxXFhwxjR
7LhuQSSKiFe59p14+n8caq4B3k/o9H8Etf97VNkdpaJo25vRpKnsXGjJZ9s1PL38f2C88Sq0k8Ka
a3Rk8loBaYgqXq3tWTQJYhhIocrD5mPxriu46InREs+Q2LVVPo2RGif3hEEZ+2/lyvWFenOfuOfO
dpOdTOt0qoXDGuVwJLZaXX/Ez21DkG7dZktxnvB8d9Su0cbIp5Hs/HWiusXQxE3+B5RfNtTQmyhZ
A1dHYOFiuht+brriHVwQEf6QuT1KT3lNcR05EAGrUQMFyIaOk4ht20oERqnRqDcFjuvAIiuXUxPD
hQmx5CAiQcPBmTi4k3ytDlPBP6Tkhz+pjZrVqINtwObumYjXws8/whph35XOmlvli4hlvEuPt6U8
t3Q5Ms1A3oLE9N3gmXxeiVeVYaVQjf0gzuiSSMFJz8OnItbiZ502ytzoYXhRgiBcYswqP8nqJEFo
mJotUyuYgYdbOewaUHWMq47L1Nv0hAl6naD5m6cGwLtgcLgJunSp8Ext77C+5e5b64tfdIusV5PW
sASx2yDavTYJXMyYv5vU4QeFzB7i6NyWQFItRV7kjOjHcfFPpR7l8yCPurTzhqT48d/hctm1hnjk
mVTQFHtXaAodALswHjGRcvwGQ2MPB01nDH5sAKhWVFcDdGzH8NsVDrb/QhDv1PNqvJmSuvu9dwKn
4ocnGe1jI4dniknVgpGppZANZJ12H4oft9kwbD2dOxLGob2teJrJEtN6gnjXxTbfoBZ2QMnA6ygg
7BU2wGr5im43uPlpU4Um3Jyk1U56u6OpU6XvAjeG+qC+snpG/H7xbEYbNIUuJksYwVChXxoPkUba
41vHwbl4jcnb9PS0PlqiyOe+hOXBa1w5882DniDKrjmm3DImG5n4rcpg2ydhyPpfjpgpWCxVM6up
tef7AU81O900jksPZyQT9UQoMGr3/cRCOrnJ0iQVLy3U7g4fW/w7TEXk/Rm5M56KzjWdXXyLgnmJ
155J4oni4SlVaX7F3Ed0WFqzoKIfsL4GbwZ6ke9vq7ahXEjvOk0lxTWs+qq/tOOiKOc39C07s24S
Df/aX4x0pbnfdUaRqERZ5/ubwoRbYmYrJ57PhSQdFvPyMR+1b6mQwDbGcN53/3grKVoLA0UVKR4W
3ubShI/8Uq/GylcSj69WUUjB5sbBn9LHnIXCjwL4uUtBPEAaL//mqC2nYuSsp69sp1GM0ZDByMjD
iE9bJ0xoBsw/+QgBfjjLIv/SGWvPy+zKegykK7XPg0g3m85Jj5yuI0ZCOgAk77DxbGIgRVDBFHYB
caAAl2admLjM88gSbZFz3tZLLi26fNTKP2gegPQG9xy+tlV7033gKL0Sygeb3Islo6xTDPeQc+2U
yYgq7T7fFd1IM9chgrppWTJFs5+bJUdKDUW7XyTMdYFVtbNId4XqXa/VbPrwOOWhYdkqCdLCny6B
fypc1RN0EhjZRbkf6k3ZyS9OfSNlKRcUNj2t33u0+hcSqPj6GkslB+Y3eJnaipAxbD24Ol0gspib
zt9KyCeZgHqOpB+uJmXgnYq9edpm5YNmQX8GmI/LAokU8Lal7fD1LDhOfH8n203cyI9pfLdGL1SC
omjkEUgU0BHUmhpGF9L0rOthrtzNpnYZRkHcTHfOF91fCnfRCOBdHX+9FQQdFtWKU5kMghJsj7/J
GS90ZKlSnty/UyhXjTwzXoxKgU3eFb9cJPDjQ0rVO8OfzpKPnd8XQvp5DIXVWcyZi+HVqT8NZTqv
JoqeoymkNIxxglVqHo8k0maDJHIEz0YCkPl+22TfC3+mdpXc750x5e6NnmuKyB6iJAa9DzDGKI/L
u3HFCVk/BOqSTpxuG215qjTnO2PjOBAHoPP/YkEiInp9RIkvB9vEzYjSSbVsVAaNYOEkEKv4MBtb
Ucmu4g7tAUPmL0u+TpcUOZIBeSp2lWS2KvIghy88sbFSIE4fZT/u76sl6Y8u5ncV81FRwjmz4pC3
QwaaFv9ilxcUWRzn1lrtQ1z/hO4f62vtchRaIF7Hx05vgxw9Iiwb/N7LCFAB2+UsPlhFCqGMLUid
zpdDo59xSPJ68NmJdrlwLvWra6XQAU+bkqB/gwTXrDps8XyZF+9YegWcam08OoZOpjPhm/NaXEFQ
xFe2LdY5VzLjCjBdK/v44MsjD5Jt47Hd3CTEhOkatzkOJWksteu55FKnua9iNC/8gByluGWULZJH
BWXgytkrNxieE1XIoRLeguKwMPjPj/Ew1A+Q3HgLymjEb65Cs5dAUePKz7ZVk+jafov8CwqgXcxV
NTpA0ysap2IgG+cq//l7XX2Wd6XNCukZTSfp/z4Bl5ohxCKIqIVaI6R30RFy0Fw7PMFX0Nl9B8UQ
kvritvrCMppg6wQV0kt4eiAU3bI3gRqiIIPHxBGyOuSIY6+ydhuAcCC3lVF/4wrtCnwPHlW4BgY6
yqMdg7V3R2G0mCKJYeT0Tx0YLXdgviJl5g9WanbF5eboG4vLodPgetSiZHkB2tbT7dB1w+sUiavo
HY6JfiucfYLzuW+sfSUAiITLyTnvZPVyA1xvydlBBqHFmhxz5jk7IA4rBAF0ScFN8XQ2Ey73xciV
CUCzHCoYb9BO7iy1tajtOH+Rc9gPGuejNBKtybWGGaPeH3ps6t9aPyTaWwo9KGpw5NtRiCUcUO0p
/2mSZ7IBAKezyhNZvNrGzSpncGjW3q+xCnSSMP1b6WhSwYE2fgcTlyh6aVN5O76w7whwFduEi38b
eRSThqAbe0uqis8mzhGOw7OoA669PjRIBtEzaS3L/ozJPpm6zNLkdNf6txOSbsXlUuIGQgZiU+tt
AW6EB8Orh7i9Ml3/J1nV8hS2RRg0GLfnl5n4vrBokZ6XxhLiyzmpSYZiv7VTMeASz1vYUCD4A+6u
a50D5K6+F6Ukn+ZdpQYKmrPAeBw/qkST05LcS9h2Pk3xxbi0Tp4HVzhP6JrLaJ/buEi1nSzSrOrn
0Ln5u8B3mATeOgOa7LugE3w0pJJnY2uuWGW4XegDUO+2n7oMvdpiGkeCg+PMmctBfTSV8TqOzRdY
9VJN+MbQqpkGt+Qbr8lNLQenxhRyOIjiocaWsVhH1IsZ3LG8YMbkX0BGbCYVRQXEfOpfEjmmWHAU
P2OXq1M5di/HqiL2Y6H+9NOEVzNgHdwtNCM2HBRcwtrM1mED6Ou0yQH2logYYUQ2srtWOxL/a5B6
tqwQ+8g0AqlBn8macMFHDlBa8/Vku3eFNPfoXPjV8U8EUnYOhWM4Mg7vCdhHMXlwj/AdDVlLiinH
NBv6AfGBDJCuHNJWxYupTLuGK1GVuwmv0lAObvlJEDdtCTgAzefUlkX71PcaxosH0G/srMFvbfaS
80fIUqozRNEcccaTw33MInDNWc/TscD/LHK3f8n5k1Xcdl90Fu/1t4oB5wiOOeb3TaV8eZorqGaL
+RAaoRpTzNbG+Hliz1k4krLTIgcsttW5TtT/aB2gZAF5YjbJft1flLJhKzvNrglHZP9f4jaci48s
a5sigNRK+ySzvKDRau+klDOgTStotCdYyWBv74ev6y7UkD+tvdq/l9nzGhmqz3lhhN0zhJ86JnKh
lbgBmInE6j+imCt24wEbpsruHUfUpnFhFQ88QbHt/WVFoA2iT01L4yVwD2Qfz9N9waYI04tfKbqI
O2Bw47uOpP8GodwCciPhhvMf4zQPc4ePnODbCnTNOvT0+K12cVA141tiYIEGSF7YKPFA1zLZsw3m
uQC49E/SeocCtxZm4Y+Kty397o/ZYnu4Jh/mdhlfDLAfa63ut6PnwBckcxL/gGbGkEblnyyDr5sD
svk8bg9GgN0hVlrrvgRUqPx31AA5/1kUc9GJnUMGgNoJStdjdwWFf7vOjwsFkJb67Qy7CGT4ZazP
PHWe2lsg63AcEoUTub1Y9vELzRxMfnAdboFlVi9+J/bqg1lsVyIX6SLK9an88/04MdA0sdBbJD3o
yozXPDPduWBUW3xmg8ryftkd3TGe1bR+iL98wIPXovBiW1AqJm4v9UGUWe7To1iOMolK9BuTnGxJ
1DwVpaijNzOgEodO8HiWo6G/mYjInmUAVlO7MjhkpuTW9RlyfyLyOf5aqYWyZO02l0oJwaPGs2Bn
JAD9LIHuO+KZbsblPIvYndUFAzo6lD3JW+oTZVg/e5RoqmiU8hMRF/dQN6CHco2oT1r2FqDIACtg
Ym6Ws9uIDQYGSrsFtz2a1coc6wkQ644AoPjVXqtI3/ZRMytCQJevGTO41hoHTuKOCELgoqmAsrsJ
yLPTN952dfCKSlGm9XPvyJ+vX6Xu3Bi5th9HgwUeXBt/+3s/g1Rj7DO0bEVyjknEqyVlVetQ0YBP
SxV4JGoojASh527Jdw6gXFoiKF18QWs6PYC5MCMmjtPlKN7AQTihDaW40KGa+wqOLCUmgOAeweEK
GXyqNfSUIxd0i95zIvS57cU/kOk0J6bOUE4ATKue6H5jyg9F7R6kO8ZZ3kOVecglltem8gJFnhi5
D0wguYkByUvQ0OZG/WgeO8MCr6/NF6o1v36KRbsqHrlmXbYgNnQbhHK/vQeYu3lQ5zoFJ8yMH9o/
gZWsG5AIbjptrDJ05wYtNXyey7iwSJZ2AYx65MpAkceHnFycO7wlXHuVrFZIPSprcxX2A5e6waUQ
K9vP+bztEUjoxMYYMrkBOIVxY4Xc+nQudetTCONUMp4Foh7wnyo40bz+55ePhbK93owai4O5RUZh
XvYXapEWeX414Xb/nsHyRdAHL9G3yKDCSm5Vx6/fdcR/a78e5d1dNzAQAPiewZlkk3gk7U8CHV2M
GjSDrhh6CE9KPwZVezBwdOKGO7zBksi3e79MEyeN3tpRb5nHRetaguIyT87AjffFy9rmkH8FL/du
YrFgC9V8tZZcso633U0O+yfUw1gz+pSbuCKYPXKM8vBUAWnXg0XTzJO48gqgtFsqqz4+5mezl4zU
3l409EQ513I3J6NhLEBkUuap6CoEVIkRKl3whQGcKY9UskwNdzOeKChOjikDQPFZvzBiLwFtx/U0
oA9m5HcVIdhkshMeIQpmgYFM1SEUVlhApXEmE8y7V5ECNsbxqQLjxeW2rqrl+r7Ptrn8b5i4DRPa
uGPa7MQDXuy3A/MIqTzWfClc8S14jb3HVaPEYCjOXBsqyaI486115ygxV0SfrVGbn0wAnq52hkjp
Hx8jvoS6urglG08syuy/W7nuTpWCsZly/cbNel3c9zjdcTpJPvrmBgwRylswEiS6jL+8r9VofW9F
OX0U9+LaG4bdQicw5SgxhR4L259YfR3COEHtyZEnoHl+k6KoVmYkhkrNAsytQcQgInwc83Q4LD3y
y7h6XBd+fzSbfIWivmZY0yjxDsOzim6uo8wsu6PfJyhfgc01kimVsTUVmnsoOVO83ohff9BP4jle
qZM7txy0+v0e/QWTd+mOsX1uN+mVm5V0XyA6vsz98n+BeuT3YZEUavqcbBq2BzL0tW5qSTZMpUzx
mB64XHRv6K2UdKIKA1zuic2I8iAGu6ZY1dBIcgcpQJtMJTU4eZtCU43spAlbsk+ZrBqzjdm+C63j
X9Wp3sAema6ogWco+/6RbK6oaizymEq20/lS8hjVeRwWd932hHqDRikMoM4t7YD70Epvi7tVKKiM
OwLlNhLdjyDi+zCRdEXgMvfw233OkJJ78ambEAozJAjiuIqCNenBbYL7vYlvjT8wMOXkOB3zotZN
cgi82iUb9jzYJLsmDcmFkgY2PttXVRvTtAZ936FiJLJ6fVUOW93rUr6V3rPQQaWlkVa8cy5ZuNbW
igRUmvzDq6qpyKFYzZPZWi9jVsvzc2dVn+ewUkpvUdhjkMVPE+egsJSjb8wlQoPeDaCMIEXih+TU
ZoLLCGZvw7PBUbY/wovMAiOwijzNgB6jiI9lrko/QA8TUebVf0C2PpL5I40+krh16GzzAAEhR3J6
VCnbLgPDMXOfPrPMW1fGJUqAxHf17s+TBU262XuRInadVvKOJeqon9zR+0lLlha/KS0V+E78VazM
UmxIeEowNYZHcYlZvTgvKwHgnj6f/lVFjQzwRDc2Cdzzn+mxt70DtM9QBRmdYHh3u1py9MS5DKse
sc6u7HdqUhjsXmI8wR5oQCTNRaKgWtalJjEMgn0UobXaGkA/T/cxTUPodZYs08Jnge9cvIIdgihZ
vM4Ej51c4DrXkN8d64dKeY69JrBV1TaVi823m2Fm/0OPsrDHSHDy6Vx+rSduJe7kAxpPxwUzfk8j
2lsmX3t/2+uH0sXDTk0vKJvUBdO/rysxEeOVVx7qMoZbezK8giIf2BWVx/0SrrIhEDHdSX4G76xF
BCK6JED+pRERRtelmVp/OB+1r2sGMO1O3FWIj2B4aVJFfkdoddh0Ud6q49sGe2VKL6meG+3I0rXH
GLNXlCNDRLenaKuw6HvItA3+AGHbr02xdc60QGOi8Y2naWhKOP8vPYVK7cF0FKYV4fXbrWdVPRVL
/h42eCNtQ74EF8qK5J7RFyk5T3AAagRA/VtcW1WzeK7QOFGYS1ftXIZYq4XumlBU/VFK9WOs2fJ2
UjBhZxXCiQbhJK1jvj4eKbYHhKzYdTA3mxD5r50tM4AKyXvLYO7OLzdKblmGe+71LHWuV5mfzhWO
GnKZR6YCct6tTXNwnMEucJnC8AM7y4BhZfJqFHHXsJhXFBjGGiWC2GALKwq3+OXbfeSwU6NlWLDx
d6kdiZiguEVBgXmOtzvsF9kATopAVkS2qPO0MQwdSqrO174laW7wKqLskWJw9ItO9HZP819sHxvn
a26olSjbXncuR8wYkibq9RGwJq5UQSkPt+WNubgV6ifkebqbkXdQPlJ7PXh8BD0TDBHvDjRYLUru
cKPstaO7J+m4CPu1k/FavdorFWnnS8aTRXkr8Hzv/Z4BT68LsW8+ouNdjXfMNspli5n+GoOQL/iy
G0mYRQ3CTM9zbczsPo6fA13PRwfpEaU1DDZtNs+nCRHW+k0Fb3O6WzePaZ/niCN1Xmri0h9zOjaA
qEI1sakrYCkVWhHgWDLW7fNkj2o76PB2vBrt28c3TK7xKAhw8js6uTIWtwCFjWrKXMK4UtecgSXd
dz9RpNXHiV7X/cNW7J0Vh+CqGVMsPXDdyeX/knzlCmS4YJuX7N5qGMdFgxiLK4aN5cB1z460LoSP
C+wPD9tB9Ov9E8ycfbVGFLSR9K7vR9ox2xrD8V2zU1GA0XCeFETIFTkidhLDCXOGat5OfXR8zA9N
ExizQRVfnbLRCuRM6WBSfQhtVH+zN4FEAAPX/X8h5xABZQEFBG32VpZW79mlt6mb+s5t/bLom8Kg
+d/jgYk8XjurRTljOmsWVYlSvDnqIiHgIprKmyqgQMJ43OvH4pK2A+zaVRgn0I1iCtbKHczZwSLF
Qxb6L+WC4WzB0JuU0fs849fFljoeeHeW7Xg1j4a/lqNrSBWP5c4wsCnvYKNcHLJ7XwdA757xxjGC
r9pYkM8lAskmSN9kSE3OvhGkE9xJvQ/R5kAE/Ky8TLZotj4o8kFKaYIrXNUJ2SK/DhH0NKTAXKNE
cvL8TpYmG3dnmNVitZXvFPwjhRTuAR3nknYTPREaVY57HVI5gB3O0BdoRwNPV+9LNGJp2QfCTfM8
zmva607yZLXeVhelcvdOJ2xX20k4U6u2Mty87OHSnhy7PrkPsg0ne1tI6FqPacHedSb4p/QZEJyY
HnEXz8+4A7mvxOnfHzSJkho15WT/1yKQxYBHrYUB36MlaBDa8OIlGDV4xBVJSUrnuIR+W4H5eiup
bSP0QzS27afvHCkL01Y+7gFklpD0NewEk2Nc7aTEt8e0we7IYxC1c43sd7n8WeJvWBRh24Vlm8WR
6ES7ak3nJO48HwsMgqTbQHf3mQ+KfBOeJ4HCNHJA7DReAlCPWtD9jk1ygBcHI/J1+be/klGvkvZx
uVzcgDizlWMEex+V9Xq2TcVhh7qFniJCxFRfuzdr7q7sxl0VlNeborcII7fMH7tohTpk8iX3aitZ
yQhU4WlRBae3YnWQVw1weNA+1uy0ot2JA+Kz26iUZfRA7ilj6v/AJBdXapmENapnhs0AU8RPgvq+
/iUS5FJyU+iX9y45efTf8XA28SGHAHMUqa6jcinqDBV5M+/ip3Qr76yWUturM5mWr4x/Cpn6Btn5
i/RzSMAZARotFXSbrrFPdIdR1jA5vsnn6pUV8RTjG7y2nYmY9riPTWTEcXdJ0sMx1T1jthUu6p4+
w5ixvnMa030pI8dWHKSIYVY6Hh5H1RBrFmo8rB5tfcsmCAwYYCKbBpCUecumnlqPf9wnN/LQl2ds
/P6sjWEAxa0l5M2qVOApMw3Z+P8LkbcjSXBnNKb52VSEniSgeAy8WlHNmu8s+KFZbxF0OeYMKh/x
EP9GDInXethX2NCZlcOSXmSFwoTNxTtAtF0hz3fUJagndDI9FcbjGJwF4gPrV5L9yCaWudjdVzeS
xGEZFtNOs7Cg8Zf9tbmqzo4Jx+/rgzBEqtjkVq1Nb7QTP9hkyvbBxmKuEpIILiVS0LMh+rgvlw3Q
eObb/U6jfeszVVduYtbdwuFQQap5WHy53+FqJ3ly8OARuWLssdcKpd+wdFHvSIb2KCaFROMkzXIE
GjxyyQU43N4qG+XbzFGwuWNwqztibQQVRo6HWrdWMW0OiqBq4ssLsjr0TDGf8Kg7X1+uQhUqP5mD
T8SOuP/o4RqeGUzSyYckpm/ia3PQzjjqKAEWhrqz5p14PVtMVUYFnObqEahIrXCr3o5dpG7mxUqJ
b5GtSSiAle55pXcDyS6RONcqkfxaBvgPN6FfWWXXcmEqDR4RBgjNpD1Zei6qviwTzHXMI4gYFc1h
cE7aTZ1vbvzbUoIcyLkpzMauGKmKt3lRTSAOfTUqO1v2ozKT0JR0h8ne8qMUyIVSkASid2hyIKLH
x99XXOfrwaBQgaBbISJY1IzsYwDtZRPFPUbBHaTdS86XEsBtmwIkW9am2697D8qt2+GCtToTNEyW
EZhUrJnSQFazhCwGtq7mG1ySEfaACxmHgYUxy7SIbWpZMQ2a01Fd9yIRs+c6HOvt50Dw8JyYMkUi
peRJl7aGEvA4cyavW28AJAaVDQVrBBUUqMi3Wzpg6NyATtOb3QRmbdoFzALZuT60KwN3zKGqNIMm
ts2JYV9D6RF2yTj9hJOW7SSvepQPjcK/G3WdzFhTzRPVnJB94lA2+EUKwH/+rTJ+gl+qkHuIHe49
zNHTIPEL8iz7fEoYmyuLsVyjV1MMd2+zgZOjouTGMNTkqgDaV33TL8FTDb8uDVN+DOga04RaliZs
tVjr/w/1faoj9cVvzPy5CHLIalFZSM1g9xuJXJW0x7zFXYm666M6DIIpCoBz7opQDrlIRxMeVjns
l3IMizTTDOvYGG2Xf3XcP53xg1CdE8xB7ZRbfsSE6/zRrxJVe13lwEYFY/YD4j4tDlB0A3jWKWW1
WCPNwYxj3H8EHvvkJZOvxfl3M6gNmCMxQOQL1BknHztMrEdYtsCgKAIWFmiZIC1KLRENo2x0B8JP
AiABBrHsQokatPgW7Ix2KAbaoYCBvgM4nnNAYzkeZUeL4Jn/sps+lB2ujcC4Yh1nuOew+Bu/9UAh
cVrX1h3LDPm9mf3SxpZacbZasl7g9qKMBK5r8KaIWocmisvG133FNrUJIDgU/Q5btYc6TxhNQoY6
WFF3/Ixn88WOEfk+weGXQFKw8SP5Ey0K3jPYYecPypgxrpKgb1ThOMi4/d74Qg3PHqT6VYJayfdv
C+6H+/bFwnKKIBxi/5YKlSIMI8/gJGj0eQ7fsIdIGLyEfNrBwPUXou5CUteawNkt4v+YAgZHIJ+y
+hbGGLa37zlRdUeYmBQwPWAPp5EnpnRecW19cAIuuXGXkOBwSXL/OgTN0h29A3oc8fERhx+RwnHK
qiOs7grOx1lMXEH7J4NJJhJAnUBH+vm10jVcgAYdKB51+hD1unde80iGf/rJU+2LcEEoXGcQwN37
u4o3XMpc5/iSI2OtcWa3j0kwlsz3X13HJXfYFXtENwcJ1Wk0q3dtuDecXVO3Bf87nKVTyjBGz8OS
cRrOpfCUX0vVVdipj7JhIJL2ER0BIQ4BMhwH6R248Cbj/IXGyVSbmxiYjvGlxfKQqeBLsS4NqFL8
f2cRlUhzDvkG405Vk45izBIWwZ1NjU890C3aUmuGbd8k09Ce/P/xYPOLTOwqsSwAF21jc05gV8Lg
imDlTMgaiM+hTHX1Lij6hm2Wa3KaRbo2GM4LZv+jpBE6yVCQChjreKXvqutm4WzVzJwu7p5xOOCH
CS21CL9OF1D/ZZIS+afOIVUR916lVeBW7yWzd/0qFHlHNkybk0TS6M6HI+Utxe/XBfL7SbXIshib
ytZUFs0h7Kj6YgeDQeUHIwlxAy5Wqmp4NqAzro3IlWQwJkQ8VYvwNHdJBN1VM/GiykKtt04wO37y
dgPcf+Hu1OdkeH56Iy4vDXGMsuiSQp4zwHVmvoXBsUnYNq5N5xH2FgjKAuaVwlcfVIhwFjynlA4w
z+dFeTurFFSM65z4JaOQ09aY7U71CI3SJldVIV6b4yZnJVwybnYNrRwdoFtgbDze8POPB7HHtrLP
obRrB4F4taHYR5TlaoEeJH9IxW6bmHaVt1dfwTTEUviifzp1RonsbMaAM0qYxVIBGllTDLTsUAPM
1Jq1wwhVLVYp0qT8fCqrCeqRHCRjPKg2uAsJZOJb9fthkDf0k7c7deWokulxqLZ5XAUOegfSMY9p
+G+cBDoNdH4IIkH3F/D+JLSCV/5tGhOoNHN4n80JGTxkRwauStvBbNzObdpU6rEQAPXsaqWWxIqe
3DNMumTETv1waKENS+LPvEpyQFGvy1qOhrMja664Yyo1LbVmvlT2vjww+DXpj+Szv01BuJVF6Jl+
uFjdhROgjPHkV+JTpcxws4O8Sz3WJK54D4k6amWxb0XiCOrsJt1if/55RNRMhGAeWvUf2W90K3sx
saEnkgznG6hUVAwoV3UVz8U6l9mZy01r3jyGV0kD1bh9uI2cbSg/MgY+I+Hq6DqmGBJG5FAgoEaH
k2Snxb2dd2lZlDZ0mZMLUSabzSsAS8DH34684sXD3R04H/APmsm79JSrmiXXg53ZXu6VV0DhSpK7
TNLsAScw++3oINpJ/Uh4QN4uUK4kjGcYdArevoHVsxOBOKnbWBE4K1BU0kwL7x5FWm4qrddQwni6
WaSzAKa5CPvgo2yx7x143UAz7BRgmBUlJGK4jr6Gcm7vQWNuUfWjM1OmYSyrZip5s9QIMSPklTLG
uoAGdbpdXmkdRSB3VSdVJaLEDv+ZtijipnqZ88foAiri1djI733Lu/RjZu7G7fZuSw4x6CPnFRvH
0+OMkhZiktY3P83PeSDWR+sCxMqpz4JfjpqnSkxxnQ5jd6cedXKEAg/FvIzI6dDdrpklnRJav9Xf
kxvkpP26jMTyMF1tFup5OwfBUaYNla8e8RqF/jycl+3jEnlNldU5v0n+oHW0weo+9d7GTJFsv6r9
mpNRGEQHj/lZUuwG4N5vyCezJaHXw331Sa3IsZqkofglmYBEJFTYN5SkxGQs8giTeRo8VYri61T3
oWT6KgNuvpHlAd38VVHNd4aCfK/2rahANJEJFiqdiK7qmNPBCFnOjSMGEmn7zvGakGLUsiq9pTej
oEY1AZo95MceevrA7hblWacsZEY8Eemm72FX0/mP0p+8gKdRQQpy+2LLFPVes8n4hPfvrFxHj+th
Abp6O6S5+3FOC53pbsqxJvNsr5cSdM791RKbPyLsHzLPQIJt9YKG56+kp5NcM/PrWvzSwwtU8y3J
28PbuvaGD0YUXt7RVyjHEgbH/hjJzJb4pk9QSE1AwQzcJ5T/N9h78Yw5t62pGCAGrhdDTl1s/fpW
m9raLWkdUyZoeK+PCX1SQmt+k9bjhFXf1THedvmPUvjrTSk0a7KfwMpQ0a/TfJRt+Zs5x8hI0qC8
hyUR3Nn2McdhVNx0ir+CW6TFvKRR2TKhwrL1QCjSRJ8j/snhGmBYTC0GQOHozmztfxj2CutUCrgv
rCryyufbD7oHjvOc+6UOnIQK6SSNfj/W552680PhvYPkJXC07XdrFhDgDwwK+wMIBx+Qstvur4OJ
60lQjzK7qtGKOpOSqoUIMZf/1Hm+MFMbdUKLvbWM04DVCYohsu3OTp+iY1StiVXiDO+WXcmkGqcH
BEAFDydWqPfZULOiByg0Acy1VWDPau5t6w4Bks59Ho71izB0cOw8cK2vBmE6u7r5vcaEAScjOctj
v5Q17KUlNuBH9VOlipSRNJswF2c9tE8isL9dkCmPkZfJ7ijw204qrmyni1REw6iOdvo0JQPFQO7I
PqJgJn3SsJYOW17l4R1WjLfLR3o3C+ak/jViBa3Z95m8vRBD3JjIga0dI4ZXWN26TrbADQUq8GRk
JMIBPN6hw5V81W8ialphAaSNgKKXBavxzWB/qQ6UqbDst3MsxhE5JP3mTS+iQDus2j/z9pqoGMaU
x+J/o36IduF3tRXosEGwfnuBIVZ+zb/YlcrWRT4d6+vtS43yk5eRugcUswGIggB+ZxjCOQqPGKPt
WmmRWskqeoEPeRpCm/QKWfBmjFTHrP/NFWcuqqnL7v1MTa1ThvTxAJV++scjwQPMrBWskH3NjoQE
kqR+oocFrNv0I8y+EnfP5viqZUUce34TYTIRPNfqNtezmUsVN27bP0/EeIqrJ4QX0roEG+2M8g6J
dbxfVsUh6G6f/Zetpsie79UiQCV3iHeUGTeygF2c/6ltY7VA0xHuuZD4bZ3IMa4HglSNO3XgcWNq
uuEouJvQg1iVh3LQJwKfIElOmAElsl/J9YhUHQRurBQRjK9JNMYI2J45APb6Fof+Na3ITajFL1ka
9Owf90DIynpHsGOxNfETknp7JmBy1EC3MEAEIB2gzJ0VKWnKD2ifPnKpiFlHbEpbL+C1OKadu7l/
Df+rBLp6Oa7zoXBIDX6NtsuhjXwPUF+WJxulHiAFzFHiB/Dv4m99bHhEKqZbkwp/hZmzj9q1lop9
d4QPKsqMfXYx16XXmukhWOj47Js499flRjTT9OD/H2qB5R77R3zcJQaSFIpP0AUfKOKI2+NbP2O1
FGOY7DcnLWZRgLj/oTi3FKr9YhkuZTjzXC4OGv1oD/1J17miS95lcUmX6dBzG0ucQTsSN/F6Vl5h
eSSZ+xPnRtAnBh77NVnEsQJQWp0r8PJF/g+pMBLVWj4QXz4KhvRsoU6DASs7O9vBJQFsAiyyJfZT
J/sZAqUuMmZjMQpwa553wSBVsSGHOv9BMTX7C4YbjU5ku12Yzc0it/qYSU1ReLsOvatH7uyraL2m
siaGAIhhAiWRo3uK0bRFXbru7VYl7kac3P/vEm4Dxn6Jsc76I5h9lEn6pcROoXaVmwU2xEjrzUT/
kqdMPbx8WYrIHpgImSKvbw+azpeGPxJaVvwGL09BlWFn5/t/sqlQCBW7HrhsLMS0c4X8ownE/80U
zHZ0dbfN84We13suH8bLv18eqsWSPfCBPtgkKCVvtMWehcwkC5U4Fs5O6nvhVTWonQPsh5zqIVpp
FaEOafwxT2zlAwOAIgTAWnYW5XEB75CJc/TnaENPOj5GKkSlD+T/1Y98uunsGaq8QGWL51r0GJ44
zejzESOo2BFcfYtCI5g8CQGoXlODOvYgDycsvn0Ewj7yW4xbl/vebDoLELRbQpDHtQ6usbuGEDrN
Cf7r3tiww8L/njvf2Ag9XNW4HQCjKF7cWpwXNg0TVEEV0XZSMjXswQiq0n+5oViOjpu3tTVz0RVQ
ZP5ncS6vgPZvL8aOQ5kZ2vr9grWUVpwflQeVkrIHrlsQt1Z5NFLnpUbVs5u6VgCcC7bzVL41FyC0
7R6IrKFsHqa0PUZch7+kqqkMAdO8pN0SZlazvVlNyGQVkJGdGciWi8j/Z1Qt+ZfTM+dhCUMQ4OzL
8BDtusRABv8xeRzJVH9xQ9X2GftCdXN6e0NYeJoCZhmuMIPwZZ3zcGTYnJ5mcqXLifatF1QSFpzf
8GJgPNIX64g+EOZWtp0bkmwjFOmcn7qgABVhvCOfCdHpQGrkJcoRjXviHR/YhuJAxGPzRkGezQU7
ZvUAZL2BLo42R4CIdOUOmoVTxFtDYhJJnwrkxhJBwxFJSCFDUHE+wPBWv+VTRfsQmpy5AY4I5lPa
qD9JfczIjpUja88LkhCZjP0Lq6B0/Ot6uzlzGzmj2s/T9FjPrtBjBDXznfQwhcyd00PYjpqI4O9q
xaHt9vQuPRXFAplZ0ftUIhl8XWaEHPA2+cS1qbGDbX9lV6sss2OavdAMv2s5oM6GMrv0VOsUBh0d
390lQVZecMpHOfElzxxnDv3LM0lztGm/A2/koFpEE1qkYJyHFVBeRvpV5VwCPvTsNBUyeyHfEGVV
SG275QlOXZjCHdKLqVuvLfTgHa/T3R+dd6WVGSbSynon5CBsJiYJrBmiER5ZrxG1ojVF6zDTdADh
W5XIfo7dXXguZBjduGoDRO9rrz+n0JYKf2F1x1kHeU5QHOJ6U+dfwjHSvD6l4KDTfDdPRALvIXcc
OSMb4jR/Uh8OXpaNe4GgzlO1A7teIRzZ0Ifzr1d07WF1bkVuOGLCHMCNJed99T/iZQBoMMXJzrYj
Bq/muvR0gmn90DiazedZYxN45OxzClDd/eNdxQ9HTIVvQf6ugOEav/V6p9p//Fs1AtLpCKb+/oyw
zk0ojio2zwDaxg29m8z2O/GIbzsnpQ1fV+RuqAemKCS5RdnHUydYB4JijkKkqost5VsLSasLoonE
HtVyqRjBAaWcQvpy78NlwGeLGLAXQ2BUZRqQNPKJJYuGOPHiWYAMPJycueB+nhD6CCcz35GvBlFY
7tg3P8mWHt6wWTVJLnj9xHzx7RuwDq7a+1ccq+yqUHuD/1Q2WVyPSsZjNZlg3YDn6+SSqzpVjUR3
+aSUDSOcUOmewum7yE9CF2hxKeTlzYyK/JzmTP98URQm9vnFwCzfpgXXD0UYF6T4uWan/Q071zfb
R7MYHn7LjHNCuYnU7jnFMU6Ym4zweZXOZTEwhLbeOpYhi8BWOGXoRzexbI6LHqK0VBBPD1EbaSAQ
zFSA8hHd0ZcwSk7qLtG1LHkYMbd5auqQAn3PADxnKzsi9pYxFwn89sWpxOgGHD6Yig5MSONyD15k
7u4NVRsAZC/Eh7MXjCEfcc2IKmmzBwJMELvscnrqwuyw8k3NbknMmCSL2ivokjqLgchvkb297A/2
D2Ae4Pr50v7fdsPcrpCosUkusN6v6iK39xDTCz9QpJLZWe08Ua2x/N+7r9l/PCE1+1MqvfsLu7AB
nFSe9MoNhog5XFtBQP5ypesydIGc5gxgnKqUa6zdr4udHXourCkzaXrwyoRJNdUvOWpQRONa+YTT
ClzQPMtb7b5Dbkhy9ekcjohAYvsFEES1x2dTfeglQUCDsFcLtHssVfSQauUl3vquWYFEa1Wk6BZN
5m5eg6zZyjTNsepmeylRoiGBTHWs+97tQO65Ln+Uyexc1qdxRhjiZZfMIDYx4veZFV2srAfIP81a
0vy+mVAZLHbWbt8kVkAvmB+0F1WDG1Fk7bNl8Lpd9Bh0Q+AWVKNq8tby8NtUZ0MImQZbhGrbnr+2
HMN4ZWIE59qRTzDCvqB00sih76bgHjLkA2KicKOUTfza3HBGBIx2azVAhfV4/Vv7gduw4B67TO0J
Df3Ivm4kxA+UJGGtzH8Up1lCFRwokjd6yg/69Fw5nfyiTUYSCQsv8Bi7VeC8N067tr2OM1O4LjPC
BsFPtmPCXzaIj/fAbA6Er/dmtKVUDV60uzqlGYR8oE5ToyRPjqoy3TK7HlzXygPhoAGjZMaOemWJ
D1rH++lYIj0a8JgN6W3N5I3SCqvvTe4TJarxjCiI0lRUjudXCwkJ7A7wKDEh8jzXEfDrNs6PBtrr
KB8qr+BLFJu0Xi1Y0PASMOygb7/F8/rJ+ZZ2o+qLpM41yOTzgHNhxfIodyDoZHu/uB2AOdDEklNE
6NBF61tAjLjnoBpEj0/5+lk5cj5QIPdBgPt69qNJ6OKE+CY3XEyFF+M7CelElLB77DtlE2E8sTjB
IFM2xBEt0ykLx8GxJRpiMJn1Z5gYC19KO/y0NPF90QZRAIZNsYXpv72foJjjpwC22Q3/Gzi4SrDC
MVGSImGRji8HYVULLHEH+del4LdpCJXEEQgEKiJqA29LSn43TsFdKJT18Y3pxbl5/ZMdYV0okjya
8EfnhFBjJCTKudZNRSOq7polILzWT97Qr3Jy3LQcyPwLnpFVW5TbB8glNnZG0W6uS/xCpI99TyPH
drUGX/k6NV0LApwx53/fB3vpmX/4sVWJBNT2xpgm/jbtqHBvrBf5C8wvGFtFi5weH5ogfAabejRT
n/y/UIiGfjHk/6C44mgodBqH+zDM0heWQ9YtOzPDghZB8jbrLk7kv5jxn91dyUwwVCvEWW/BySKk
3g/oMt5KZDpFAu7YU99eLFxuFUah91zoHAPWgzq5x6TKVF8tz+s+CY8aHy2DzQo34hW8krsivAE0
rCm3dIJsqvQ3CXvAhSQVG2wAWd2/yLmvnK3jRkhui+rkM4oy/aOgVs0nvCq1w3rk6YiFccKFcR6A
d8//0HIXkorIo0bqkF+++j+UIhdpW6Lllwxeo923RTRzZbpOnAs03G/yohs2nrt6+NrNvIZ9Hld5
QO8sbY0a5mR8UBYRm/Sp39AIxs6NQJ1Fwr+NPdNw8BQKsjO60Eox4rbS1G/0aM8rGwZVB3dOw5JC
zBj3R2gu+YCkw9ZOYbfzbpwRYqQba5/ehoIu08TF7n7JXIO8fAqCGiR4xfMQD/ElxIAqHd/VV1X9
vInn6eYBjQM3iLpXaiEQzcuiSexh8oKFEFVZv8bAG9j/+ALTh9PQNvmHc2ekn3j5QZ/fYv6JomDi
bsFiQIMbb+egwHiSwKz+1CWrAbSysjdBnBCQP/NMBTT/VHSeaelRo7DwxGOsqILOUQ1wowzkeckC
cKeqvW+18jM3E8ug2XemrhV/fFzNFQi82JzPxuDYB+KOMUtoGNIEOGaZCdfQD+u0jO/pt+DSaJ4V
wx5Dn492TTsjMdI2145PWlj/B0azSgWJAjoJLFXAHvezr3afKiVX+QZpVRvHs+rseTbRLCuUa6mw
djbBg17c6EeEDxPnfkyhfsl/FQJzujC8mUcGzhxAjroDtLgAvU1Xb5lqawg3oRt3ip3y/Wx3xXl5
A86Y6NVBpQBVG6I77lGqzEMerFi8ucNTgwBx/ZbbD93cSXzM0Ytwd/f5aNC3ryp/H/PwYbodL9vi
Y6TW69956eYd4i3wjEX+Q7cBKmOWbYZAYh0yAkmx+QS4+6pQvWid0i5zwA38sw5O7Mk02JSbBEr/
hbbQRmyfz+e4CFlJzmPB36zIjXIaLoG3je8jlbiDQaq4zJ7szuFe15vAxYASdAKWnTlEWrQsCihX
lVkwM1W0RavsbKRQiXnpQ2A/rUi8sjsCqf1ONwyzF4enRoqivQUv3KVNWwlnNmXAdYtrY7KS5v6Q
DZEnx2HPwO2JYIcJrWMIBjTW8+1+QIbksm6K5b7aL4BGzX3I/Y2N5p/2NksHyMEvq+NNm3YdxeMl
2FEF5tfCr50QhwafsQby8ozwWU+be6GYfrtItR3EIuQypgnyEeJZvBkT4PQOX4kgnKvw3xYkIGke
uQOVztKTsdmZCH7cQm71+CCFFTfcUX7Ug+KOHfwurkG/Ka1r0G9Y37ilfCzFwfeYmCGXZ2nc4g+4
3c6Q5glOYYteRJvHoly5zY9vLXpihl5m7qy2Ya78YS8E6d9lZPV3uZL3ep+V9R5Uh72tJkDV2BFq
yyFQAX4ZId0OitUaAcwjxvrjX0xHA5XiRfHxa9lSPYRuiE4bRJcs267XKxzef4OFsi0LBFqHF2A4
gFFFNP5JhvIiaoaVBRIN7ryaqitzIC51NSXt+ebW0L9buH+JyC0HAGxbfKanidJUpAJwhpJjAwkc
guVQtvYd32GilZe6fmhQwOkrZwesF8q4NQbxqkuKdHe1luMD/TVQ2SAuN2UTR0Y3+CSyalwYLPO7
QAB3irjDgwR4/KGkQ15LC1qnsRDvPOVlZDn7VJjA4btMU0ATqS7qGfQPwVCtxIbnYwY2MeAnguzF
VQKAbz0Nw+JYLYQ+B9MyeWGmYaAPdjVJnozCQ4Dd8iZ3QT/y4ZsQrrTioJgXVe/RRY9M2Wkbiq2c
EQzoPUDkbNu9R4he1+ySYouttg5lYyVaSyewUTXWCs5Fe0AvUPvLRliHEpienv84F0VKhAXq21nu
5Fd17nF3XZu6pQTKXgPBQUvRCWBa4/aXSOmgvZqilZueoHisxBmEADB9hIE3O6huIuDW9mPsVUxD
MfJ/HbvJGlhh7P7wKLK9txK1wOOwQOkHr+sYHXJEIHYwvuWpQ7qiSRxLuMTBnT85cu/rdVmsM5Sy
qTf1bUzbGv88A1fSAtd8jbpMz7w3Uz0K0G4gDvHwZUNVCjr6CL+8M/ZybEVseF0J3uikznqGk5m1
pHpftGW6asxL/rpVhTYDNVXje4ErLbjpGODZ9U8Z+QWqYIN0ijOcNtmJEfso/KKObUzcPE/at4rX
uN7yo1m8/xOfU9BkGTouQRZbMO9Lgr9I8za5361q80yFJOSmXfB31e6tYk1bIwDgm4g4M3XEVhWz
VNr/c1oNb6PpAwU2pw+ilRwYi1s6X/rO8qgXmtqll/MoEJhMGTUQm0q6RGZd8nw5nk7wl0QpLMll
Z8WbW2zhCOywzMiSbZBLJEF8SKirk+na2yrZB+nwU7WblFUe7cDSI3sND7gt7dJgPiJ86o6eUier
dZ5EW8rdMRan7+EM8RBJIfoAWrQWKOxMaMZywmDcU/6iACmLwvKKOTR5tyVkTma4kiAqPaXZH5NQ
gg9dE8EdUyTOclsZT4QakjWvjS00uQJ5L6QJCfhX6zdlYjb1y3SXDxVeZC38IoW21PMMZvUvm0Pk
mwpxtAE4X1k/xsBiMUAuzAzDxqatHcd3QZAJhH5L+hJ0SLVARUHb/BZlazdQbGL+mhDUzVTepXjT
eqSj2RgMSQFFMi3tK6hluhzeFGnJTchv4N40zm0ErU2f59EWmGllaQHXxvbZuX+e+Yq+TcpACYSD
wifViEX787KI+3JP/7N5ym4hZeZn/lU8N98K3lDizR3aGfV8IKOSud/PIdUGydM9JKodhaOIHMmL
d2jC+FWSqSAj8PgyOYNRR0KqATtAF3Mmi5R7a3fBoocQDKAbZKXGCAODBfJEBzRywiy0X4KrmVwj
ZIcRSTbHw8KHNUChkwGSuFu7UEmUIe5uKSD1jTPSoc7bkD2j0fLWa3oGI1vOZy2fxHOqrSztGQi6
CtrboMgAzLLbueKXzLuFn1xFS4DZFnL1Q1DpoBTTnTu7sHphOMjUbTZTXEeXizz7zGtR3Ez6imds
JukpwiTDJlp+dMgHscCnEP3MnmR0B/LXC2pb+ASPLMirOmRNf7jhpMzgYpnh5QX4zTo46g0jyz8e
kvwCFl7gcPnExDHdr8HKEkAirzevJVd8xwx6U6UIqIXMNLGxkWdO4ya0wVZ+hpV24mdM6DLDGv7p
jepFYhXMApBPEC6bDcSpps8sFoVIQ6m51oDuZqezDixbwiFHu5U61/XK0t1JxPXVzuOn9KjMsOVG
hYoaDU5ssgwHBHxTbWOC5z9Bzdjkxe9T6Ips1cDLTxkiDibwuVhnR/Bs4DfGAMRlsZvgIdxIFDlW
jJBlSX2bKQGgTKZDNN/pbEvXcqmt9h0xx9n+DqBoV5Ij5O4Ct6iJnguVTuJIJHIYy5ATsCtLBu0j
hMUwtLmJJoizepCDECbT/YHo/JePK7rfqk4s99Smc5aUCWv5aDh3S7lFEJ5e4TSg5U4H/f+FQSKy
lgDVXmn6MazpV6IfKZX4A3EcNKJvZCe0FgRjfyVqDfyVEAho2g6ublx0w40f/XSrmXr+lIGu1al0
A4EYlQ2NFVCUjBWy0NcSP16obWcmxoN9+f/wj75ZI3eGz4O+sTuVMfQHIsGdCt04HuMET70WO1Do
jWVKz+tR0IDA52vxCZJdLPvNxGIeokn3V0ABcc7clzRmkMgiDX9QI7jyb/HzOtzwgCyjGm0rQnIr
IwTx7MIVaKee49bIbPRXnN3aZsrOpsCGQHHguxB3lz3dhURombe/Lk4W3rWzeVBCsAxZg0w6igXZ
qtYQH1IxJ0d7bsbgR0oMXHwT7dvCa/c7kGoP8YDfHP2ZI+v4i2dV2TEpwmzS3Up0fb3FkEI45ldR
x7JlkdMb3y5/1sqC0obE358CVI61XkSWKJAnmSROd3pwEOUusO+qLVEWhqup0p3mhukNJlghn2mA
asR2Jyx2d9THrYAKWO701XYOXL/7Tc0OdlX4pdjuDyCUdAIqIzYB5vxTap/claETxJ4AdmNKRf6m
MhR+YwmE0YviJL9L4sbSsAy9GVXFED9DD4XVh4T5UaC0kTyTcVnlxv6Co0jZ1fGdUqBiAPPRK9LR
uVfDeEdDeY+UYmxLgIVsVJAYtQGK2IoZ86q6bOQJAA+UlNELh+JUY3/2geTBC1M1xEleMh03OGN+
46k+Rfl1wA81GD0/psQywfnKxIZD/J62DWWeZsTwkOsfZVJtPZfcIRPx1yPV8fTU3ZLwY0cNH4FR
jJ3duirWQMqpTzhRoLR5WGS/c37bzUtdU8+8HRIAqob4U1yo3GBjANz5d4uG5hQWs84e7rnVpDoH
/uJsm6FK0Oejv4ZGsrJdGvIyw9nOC+SLjD6XyM9EJfhphgreMhAo5dlXFhkijlS0rDRX6i46opk1
pYmaGxN8Ovyp6CLnBR8dvf9fA67NNnaAyYtWCfRSu09zRe3YfmU6BcvfIXE6VSbjYXqFdVlpzoLO
RRXvgTBTalslEYP6tkxkyU7Io+IVZT+qZIbSqYg0Vb8I4x215GaG3N9UqhNfCBIlVRLzpYzRq4Js
oub1m8qVaSB+ZLHFJH8bHFghQkq2spw1jCGzwrKBkqk6hbW8uwGZaO0szWnFDkmAaB6tZJCgd8qw
JtBPSOkyKjWUt9GGYMHDX6dGZtJM2cF+D8nc2pigQzEoxys8zniEgFokKoCRF85xKytxf4+SPBx4
7r39sqxVH0yL3qv8EAHSkA7ou6cAva05Vxiiy/3bD6EV0Wt654g6ywH2hWBz0wWYarVKqESAdGSk
cPMeFlKqC7ffAhE+ao8dqy+WMPD/Z5fgqvQ79iZDZQrRzC/4Vx7DadfNYoBT02mIqyL+MeFoOiR8
KJCacF3u0JymEQkyNUDCiQp7HG3KJUItOW3ebT+kj76GlPJCJp70vWyRpMkmGbX3kH3Faxl9ytED
jsingc/etIq+33CN5JWKzxSipFu2JTx57piUz5CYgg6LVxM/dkUZGtOD4mOBbl/3ZOwLitsvJ2ew
Nc7Z1CNzbcIaUgKB2Q1f77oteua9G2fZlHoGMDpxD2NqrlfO6tBEBWDvASa2G+qH+jbKs9V0Ywin
K/2V8hxLu+1Dle3RiW4MvVNOS0MlSUrEif71CDn7mlXIJ8iy3bI1J2x2pG9m4wQ6lEDXykW9Hb3s
7ZwTXV7Tt6XrDXoek4FDlDmxyHB+qUCc8qEGimhZYXSR+Q92NBiI3Eh8XP7DRo1dusQzm35siIiE
bZt3R1PWdNc40dy3y28vu0ErqB43qpzJ5xaA5Q/9hT8P1NtsfCOcpi+tj8DyoHdphEkspl2FtD0q
J5wC+kKi0XwPvhcbdWiBrjgeq+9S4UvXqAcV4Awymr5LSj2grs/wYCgSxyMGv5G5fxMUNRS1qJjx
Ak8hOIQIQVxjHRsDb3yvsPcfN1G+xGmWKVlb8XNo0SgK72DCbA9FJ7MZuXmZu1aE8GkgWQYI1zra
Blz85/Wj2wsz1Ckx65fT47R2zgEDcZKuHcJ9qCqFSUJqXPQhWyKeVTrr8xwlR/UnE6N6jr/gminy
xricHU/Gu+E9HnxOAF0ScxE35YEuMOGOtrgO4Rcy4eVFy6Y9uE54FfvlLuxL8prvBX6ccrJ3Vrik
UZ33vuadoDtIEFB1IoAZzE+/HQloy/El0ZdDzOL5vKfeD5Dp5uJeXq4PMyb5GifIUuGYaPWiQ7A9
0t9tkePmrQkT7hGIj4+UESdxv8B9hTkJubhNkA9+kt4fzSpVVS8i/8cgjBEVC8gl4QjdZub1FDS0
lsQ7IMRMI/5HkPhUk6XNIHe2XtawZ3sjDFLgWZQTauhXkIm6REMK8hZCp3Ex+4oReKP/zrFE4VaL
84FVOKGXuBoNvXT+e3Hz3DTX8i3Vpb3quBgb4o/583USydhwL/jDF1wUBuZoeqIDBfibE/XUyBki
oWDoMBmaiZMmBBxP40gMIA9/ZhfFoMCeT89Dk25g0QebVeorymfJ89CxK7NTG/pyrTLTbl/nzbj2
dlh4euVEo4ZvVckZ/ddYTV7IYucbtyjAR1Pk75S095hvSRf3BnQAhPelJ6IY4+mrrbUlx0hU3olL
YyCKVy3LJAMPojBojtCCe182jp3ZajolQ9kNGIP1Fn5S95bfis6/EUr1bcrDXY29UvbtFVRvDMqY
OoXMWe4JDLGhUlJbNsjWxT2Q/dcp+EaR7/2mc9SG7pPYRKD3C55PLKACgz3gAWqwFog91SwRk/Of
S9LfYOmpTjpBWfF/foQs3ijTFAyAh7vvnj21lNMaV/36pPu7MCm7z7hSidzuUQQnCua++CcpfFPz
RKlGJZeUjJtJrwlyeuVuSYWTXyUVz+IZg3q4D+gpcTD5nrmnPg8rO2rtI8rvbHbIGG0nvSOLUHml
EdvcZsd4RUxiD/jmcmom0qS6cVaCxlDRQmWBr1dbGfbW47B/aReUjTG41wAEHYBkbZRTOPQnBS8P
N3UHsfpeMAgNpOblU3u2ZL+A4K1KTqcqDI/PaaWHf7B0nLmj+bvRV8+A8MdsoXttfXZ7LXWLeZxY
MOzaNWPBNeebI35EABFP3plFElxu06J1d+lssNaKmFzs7bxwdYJcD4HvrWmg9QzcUEtb2Be+ne+d
yIM/WdaPmCGxSvqBlca51ZZuaag0gZbpe4gUZQC1VgZ1NUBWIFhqz9c8YWvtkYobAA4VNNDYF+zD
v2o0ent/FydN/zBA3ZnIOms6aD68tSIXDI0/7SpIUxu2hTz1MRMs9Q2OPJrOlvNoCIwx+KQX93i5
b214LQ/qbjbzlSa61+ki7XVFP5fX73nlf1JM4wsJYbM2oIFCOHy9HYXNrBxcj8tqAlTxZWoRy+Bb
FduaezdiO6oGr62ZiEDC4mffaDM0vKYmprSUWRmI8X6UhAV14rw+SAO6Zw9dTFCjGiTNR8AvEAfd
IQsUjjfPkkeZHozmOSEAfYkL8Kog6lIQU9E6aScXzCaHilKMGi2Z81drNko/IoeNJfWlG+A7UzGr
nY+mq+oS/iGH1zMCGZ+f6EHuuWdF3Xp4t8z+j7bd6uD1rMc4D9cDdZLWG2mjvK1KWTBkWbqRFvxT
c2BCytYPjqrx64RGDLAUipbTEPRZjFHZ4uO2Obik95eoKBi01F5JU1Khb2gbcIOHSi77lNN+Kou3
ImREIGpbqMsActWWzmnQGfpsK54WwQZmueEUTVj1DA/Wgwb1c/Bx0aQNNVHYX2MZa5yRn/yxaT25
FcpFl7GPLoHHJb0NMGw6qGO0t9EkccuUguw0d9+c/AXe/Wog75zbN8bLXui8lVkjVueJU7KpV1Ta
YxJoN74SBVZCfenpy27MBOD/Zwln70aRYwOQIw/uexuEDzlG6CP+Bpl/0oY3Dww4QvnB738zzTgq
Jep1Bko0wJ1NDBPdvbucRjBNI78jPhMU59ihF8Hscbc5xiu6mV0dLBmHvmhSGrRx5t2aDl05QIun
0TT4HSbVYroJTtLTw+VY8sRoXSJpZLVfhzU2nFsxYfwMtHNgQkh+2DLUuGBfF9uuBO3fhs1qcFiz
kH4B8+NlhZoAwd6SNYxD6RuhjbfU7/wDVANVW92BvAcaMogbqJh0Qs2yhQXk6gjV4po43+Xk/+6N
LUT08j+732iRANf00eP8x88nXEC2I0XtxKvXy7p/F8QdF7sFotD9bvv4F1Cg0Z7oFRB11ZCogByn
XkQDPpeby1hKjfBcj9TEOKtKGA+WcD6VTeAWsRcGUapA7ZJlzr1LhMq2IOD1zg0LFc0Mu3r5czj+
Uwd2GqribxFMB3yCI5YL0Oj3xigCBmRafEIxw325+wf9smLvJmNrUJnNAMqru535CSFBf1vgbars
kJDrKH38SuykkLBA1YGe8gUgHjDPFTpi8kcRNJKQlZdqNgML2kHUoTJDjVRcp/iecNs+a8fBh3ji
ZKxlQy5xnAr4JI6R7YABzxmSx7kfjBBq1EuWNGjwoz3D8HE3Xp9pSJMKYo1vGavF8RaUrX84wpBa
iqicMV5AVIRMAQr7W2gVr1ZHl7fnbnKKNtI8h2quWlg+cKI4Tqw68ONscFDSDof7YNvcZ+vmtwjq
rsrtyQvdYH+XVPqjEf+7G7W2SvGqPH8zSOhWnUX+NNME6D4AKxzYqc+hqltZs5yi2tNWyMOTffl7
1Ps1CH6YdCI/0Yoe7bto3UVF3HWPEDnjEybk72MGhLaGeR3ptVo4Qsr7Adary2ZmFIEyTwcMMlvx
xnx1IOWaPg/0QOHOD+iJ/vEWLqWZ3mAG8GkDP1yitktSUH42ENyK0u277XhBDPrLGBH3RyVJoVzx
B95n8M2neU4zdDX8n+lwq+W9ONm4tKD1xpV+z56ACcJ+rLWoWG9AQwgBcRlGDYWs5S8S7v/3SGhF
KEQ6yKPOax4+bxZJgnNqNzfZ0KKb/pXB3PIUwJnN5S0ViU6Z2I1o1je0027oYAx96x92ZlfhHbox
CKsB2cR3jENTqn1HObAGY+woSiO1dQCE7P+6V5hGdgv62T4NKzGTvIYoOf5UWNSy6fsQ6YE/n6SK
tqa8u1a0H9KFnXdiv5aD6WIYnOszSkgPHyqsIrsThP4QU370Tni31jM6IF2zQHtPQjZaEjBvJ9CN
mgkDZD6qWZSuDKeqhJiTZmOAMOO4nusuET95gsyKHTxgZPthRHVMbnPVCgX7y+euhGmKBoaMkzzc
NwNqqYRnIXs2LPpMSefKiIGZ18+vRMWIU271TS8I9dGMw/dldQpcbbUboJGV9qx0Ptc+P8K1ybQD
ZrkMk/NOkRm7B9bzZjuz9RwULL8lTq8H83zmapZXAGQexL+D6VktQrzgqBwpb0NoSdKw0WAayFt2
xMY1ewdD9Rg+9f59gnLnkz7t9pVUZkNbzzjMt+NUi/XWVP1ZOzNxCEq1KQYzZZuLUxMYiLk0Or3l
rU4F95iZMtOhtlIeUII/ufJ05UpNdpLhBepz9szivTTUvvbg7XBPrqyA5u/G15U/XG+EsVaLvopS
aAq84yQQcMDmWUS/D2Jq9uYsRDuw4MHRd4CjjobSWi+SjwmIhDdV69WKvIfTVf0z8qal/7jytiVg
MkvLqo4p4tzDJQVKT5YQRBc6QrzL1DVAI03kuThMCkfwpXLZv9V5Efhwsx9XvS7OR1P16ESx5XJ3
VibwWEzwtm1gFKYe7Dt4uZYgY73M6JtKHkdHu3zY/opx3q3LAwe68t3+dFBRPJ2JcrjPocXr0/Sh
Pslf8EyPfIHq3mQq1XpwVJLo1Znuwb80jc5vbHSU05I8veK2aHeFSONGBhdUzS1yPY4uiIG3KVsE
RHHaLM9hMnu9xhf2k2HeOnV37/WfCb/BVLsonJ7pGf4maESkchYXItA9APDbS1gTzn+z22dZcMNd
Bt1l50BHumEfelBfBUPMk6IwmM7WVH6Mm2QabDDeKRkmSOnkBf7/9k/CPGBzkTWmubd+fOmS+HGT
dHDSmSqRBDjOyne2nN5aT4xCA44YTWr+SKbl7191IRIFBl1Wk+sd2el+BmyovnwYNr+Rjf/bVYa6
imUQS4fcJqbmQkbF3eAPNkqO/NKBl8wnGNuSgx5RFZueJ4+zQFrIc3pIHgsC4jqg3OhFmG8Tj/6N
F9Ka5nQzwKWsQfpxh/sXuBUnZdTL5orA5X1+D5fBRdqyCIjEw6wnWgV7chByxJOEoWkO6jks/yOY
FA173zJQ97pUoSwPdITCc3RMmaozBEFziEBJSPBYdWU/N1Ghox6rrCGat8jC0iSzPzUb8d9eBQjE
A/BqVM16lYfoMsuJjsbQs/3zqhLVWoG2mhZfLZSrM95QA563bad+nE+fHDuQ1bHxKjGOAhnKJsbg
t+o7ByQeWkb3bwjdb3UznLjFTuMUl2MoNIwgp8Gpfh3HBKaV8t7RV8v3RXN4uFF+8SF68WS+xgy1
BGZO35f7PSgCdDEDFnO7UkiAQNe/7YHdTr2IaYKs8fvbpbCqAghiPqvmcJvqQfjPA6cv62+IeAG3
PDGeuBuCzVrPNFQZgLXujXrxVY9jgDf/UvAXjoRi3L9/UkkSi1lB6HGiokTzL4WgqDXN2tnmZXui
md/0qIjx+2sHiKYgh4soVP3JIbNrOn4R/TxfymFrJvlsxXoqsFuBbJQWmI49Waq25PspZfHuKppo
OrhKDnS2LLSr0QpkosG7yH3JArIosazQoNBUGkq7298S7bmbrSll1qoiZb2YaWmq80lGN1gLUQPG
mS9EssoHEGywOn8mFdaQ0a1YTZNBc8N/8fxBVXWGSiezMRWqraGiQxvyFrq5RR/kfjXRny+L1lTJ
OhP3OtTsPm8qGERK2OovJZSfHUTsWcBiQKhXef4uGvNkyTx+MvqiJmP7k7xlEiTRa06YFibMysh3
9h/VN8QdFpfCYsNRLKB155aD1WiWUcO5UfXBCM2aMVyB5n827XFIUSLBT4LBDWkY0C1lUGn9zdI+
0a3sAdv1LIYlZq4klBBLBUq61Kt+7RI0QdHU+NKt0gnHWyahDIojRIZa5iw63ZwCDJmr8PwwElrU
ymV9tiETqSXbdko5xK7r4MZ8PUbIRk8kmbDSaXRK0qrNOQzFIl84AbXNjLzSVdRXrzzYD/2KWn+c
TGVveiiHsEiciOUCL4kMfVkwu8QwS4eHvx+BZ6v33wnsDhZgbmW+PC/MaZM0Gqkir/jzeB4AxUL0
llKXkppUOnA3QnOlyOkYOSEYfM5+bmeVl9Wsm2D+/VjgCNjONvpXI0Uj+NaXeUJ1hLCbPYtcOVMW
zUzUb4E6vB64r3tFTNfIsGixj3EaweT2714Wzf6vLplkaAJBccZe5Qprxpsk4tORg0vjxGqCFuTM
LY+wzwlSnQooPC9ew3Yscg1IBIcwWMXpnRKNBR3TRGGk7ZYbdJu10+FIwpdG8tilYE06UVMKwV3f
gIALQWNJqke+CMX5Nn0CwM0sz9/WDnxvDfbzc5a0Dj/gRq7T06xSAecLJadhkDjK3BQlp2r3x6SL
4zuXK78yqc4K1PohXhTkR6HlfNE/2HJ0rYtnCchPNdQ/ZQ7WokcW7FQx+hOm7u80S+aPGMe/Kulq
MEj1+Z5PUvqqI6LcpQHm1t1ovhNogdbTWQp3ne0QGZAxbSxdTpdNx7ZKSwbAFytnqXQQ57AOoHc+
e6ynwSyep6b8t0zooV45Kw46vzN1p3056lb0EL4FPQZJFiMRhYZdfQqTLCkJhl0Ld0tkRUZ9HH0T
z6g8f1yEiyBjvtfks7Q7Z6HctqGpa2Y9S6jsWJsz6tV4jl3aL0VweUnz9O0KS0QzyXPT0yxTJfgi
F9VpazxG1xhq4S57TFpOXRg94K2o0wiyW/4xLfPle5S0qn4g6/HaHWt4QGWcumYkYOgKGjRU+c/d
QMvZRlImXn5LwqVi4MMa0SCDfEoRZrnWk1ioKf/xDpzOqzWil+EqLYM+bcq38O8QdQXXzJCMbIY2
qlhE/jaDY46/fmkRonBo6HT/PWaPkXPanBKpmJL4SwieBIyzKOqtjyqKHfutIHcGfHVQJCXxE3bD
GroYhSwnc9OB0fpIPrec8YdsH2r0ZZTvkApATuwy0QXMlioA6dl1itwqDWbb/1tqjGpDeRRmJDH4
+NT0qVO4tzzhNU1KOuKW3y7+tudkHhexUGdbal/W1DRSjyvBnSwW9rYALplHZvWtrGb/EMl3B/qk
T6jM5vNOtsBAt/s930FQBBqc2DOUe034H7NcZSpQ04mljKSVdR88xZEcmxtzYugxrk1U9CgkWwPv
FuupIabpmaojupYUjuBonG1FywTsI9oxkC1ICE9R/njRLfwxvF/dc9qVuASndPs50fkEM/kP5qEb
j6k7AFqrcs2IAfFyNaqPmMwlVCI2vQkEI1mkAnJ/Y+1qRdV079QnzPP/q8I1qUccB6kMfGNq50C/
TTrOGbkc6n4fsl3ZqzIcUApXotDixQ9X4GVXMbjIBJWKQltkOJjFEs5X3XmeZ7MOhuyWTEFpDpDG
KmI0qaGacocRYJbYUdhveYgHzVOIV+h+qO8IZU6Ts1I7MabNOpBEM9ghxIzyhnLDyAdUK1/0F17q
Mk0UWdjSWMYn5ZW3+OoxA0EdazaH4wuaZChbCiHepM4A54G9HSMOd6FHmdG1NRIaRnRMS6KaUzsq
NY/xO6F8v3xU+B8WvgYHhp0kSggbKUQTLpWEdUTMivVh7xigP9AUnEFZrBr70qhMDMfSDNHLBON1
Elzgom6dJ4FiXVjW2yqAQSFD27U7q/NdUCKhsjg7S6RnBSKavAW9bw0mAtJiTZBujJu/7x6NiveJ
NTd4yKRZ5i23k3LpfQVbCulV1KCMUQIS5XhKh6ndjQhHKRYHdVFEaOP11uzGlDnMSiyDbXUNv2DH
a56jcsURVQgaKEQHryinIlYDEroxApRZlu2X9KcNbv+VbAjmQ5sLWAkUq2RhuZJg6eloII5HBseK
R4pev2goEus1mKAGLpsEn7GgAClgnXOIqFUeRfnYmF6A/5riZnJa0ZAJsZwwxvNFaMpWYT+T4Z9L
1+tUce7h7ExUyr/FTO+KQQVUDaxEHp9j16RYgeDTxjwUwc9oxlIR8stKZ2nZMSB7CAowLyk+bLEZ
SfVANCQFaq/Jo444nG9e232ANFIFcZkaPHP+LWMcHXH5J3HaleFkhcL3dGSx7LNKqGQiW5FzRmEh
SBhBYUTTdrzSXx3ubf3ppz18bKOveqsSrLq+mVGEBH2PMvTQVBW2hMk73kRVJb1VXWmA325InnRO
bEqSlvPEaXuUFeyvDo9L8ZGncZRm8YxySZEGv+0kcO0xbmJYPfvrJn4R+odTeIPRlLr+sWntpfq1
+IGqUIb2+B9zChmfVrMUk26zxzKsdkqQtACPTxnCZ6oowRiL8t2aZlMADYk5gSHwFypIar46fwnd
T1yPTIkkwr67ABQ6YkVKZc5ppwGWgvJJ7eQ48wPw9a1h+Bga5k/E5iDTEj/FhNsPAGRur1PXeKaE
3ShiKz0klxrpXIMM0MQqlHfwA8JBZuJ08wXrQ0hWdejdAHMOAZ9mxnX4L/5qqJbppyl3bPdiUeG2
QzpeUizR/GAlc6X6N+PKDuhrMRW7dj6JFTMNnJK4j5D4cZU6a/yGvcleXrBvOVIIgMm3FFD05g/H
YguyZ1TV6VEu8ywtniZFN8avl0r2QUfd5CpbYtTwYEyg4T7kjLmObRy7hBNz7JALTNbgbvGvY+wU
oziZcaWbwvjz95Q2pUWienMkwCuikpGU2JLWKw85z2Qyg+bjNAG1WHo7bARk246Cch9d6jfOsf1I
fd7AMGDW7EJJOr6soRm1veD97pQEmPvWPkktSWkv3oDTq7zB/4P6QIlFGNMQT1/KWkrEear4jMqp
qSNZfxc1908t9T1AjS6tiQ+GUEuTBrGRXuLafDdOJz03JIX307BfYRVpmprRP+WoIr2b3nZ+luWX
WxhK9a907FS1bUHSFySX/ht4cW79tA1MLbassgeHJcMKueGqsuelmofapo/ENDwMXWc8R0zMevOF
WWDQllAJbAil9/7egEXI17tP8hXSpCQGJEL6ZFEJvU5aOIXBiHIruCkjMU6axQ9Q3YhLb9k1TZW3
7IYHJi0ls3x623ceKYtfA80ur/40LVZbAw2nLpMgOLwqLUaYSaodeOW9V1lJ6wvEaA4x5rwjuGQy
20prw/F+vyoFXMrl0jPyTTcI9bhoj1iuwZFmFo8TDijhb263Xf13gFVdXVS7ojkIRSyXioZkQanW
dmxCZVaQKKIieyVyCPiP/vouD+GUMcwZvCOW2UacSrR4WRTxDmTm5+CrP7WfcAg6XEqZn+DUbJph
YNSVTK7BfE2onnhxQpE9wezZy33zqv0J8mCcaMHo87coLVx3jSi7nOykNelTRpc5vQG2hZiqLCWM
rbvt7TgZr+Ls9fGeZq0uamwlaXhjbhc2zwm8DCA8YMZi+XsiQ3CN47XCPFXYVgfzz8ZThjAEO561
DSNSrbKmn8K11f2M8Jv+bgtIaZoDKXFdSW/u8+ECEaHjwzGvZjbHPWrBj626dArEYO2v/sl0nhxW
Pr/FdwzwVYN7a/bbRoXVpxyYqbjbkzlvFkQVhEvzwyDqoOaAgWfZCE+XN6oE/KwsjEpe8GbD2SKb
9w0vHlhu5c0tKx4eQCwZOLfBFiHoIdbSGNHypLIbO0E59cWosg9L3E/QgxdTTP00w4joBSnSFN5G
2hvhqL79ESe+Z0qLGBKiVpRugIo1Buc0BPKCtIhqWRC10OgMRXtrhb5bagdW+ilQSM2y7Fu2bBYB
DQ4ciu2h6vjpNckNDLdMeQK5wXrACaVGMV8wlE/cfwXW/0hNy1XU9Cc7dsHLv7LdsofisOTsAPQr
6g/4cWVzoUHDFubshyP0PRSoM1mp4RDI9agg8VFTOF1brUA37M9ITgv12rrRwAq0FmdYZuRSoEOW
rfJZJ8Bk4TRXTac02mM3kp8DsfgRTS35dQUUIL62qsCOmWdNcAEzbU0ZHZUuEENKVoe+Ve8Cbwi4
WI1w9bwd6rYuhqJIcd00seWF4ENsXeb9M2FVPB2bOA5M2sCdZOKDZwDi8M/BgQnIIrdWaqB7nVdw
E3v/fk1kxQ6SbFpP2Ru33nZk2UbKZc+bQWWCrb0B7xXJB/lR6tr+K6E6OYocmcu0G9P/LXxV4XUD
hQ6NqVUcsn5reJ15PM3WKttfGNM6aT8+qUUpuJaTEE8+wbGUesyQoqHZiqRdvTXDWn/QVF4sx7AG
f1+18Ezecu/jFlTAHv1KhVkoN1rKdePUnZaGHzT6qdwg7oZ4KAyc1wYMVr3iKlzNKzzlgUF8y6JT
MqkiHVAEzGTrV8tghU84muHWiMb4MiBZxdd/8CxnkBkJyIL92uiwH7fzZ0I2jpLJYTUaRueK35FE
CUuCQhLXgC5MBDUz5BWT8qu2Mg20XuJsPhrdiLjdhM7kSHF48wjSPE830doOsLRZPjAYmXVGORwe
rhMFpPBciTE1eL4SoTrgeE46Aj7miRKSPJ0h1VTljhxMQet/RtqJDTOUqLHoPJ95vMY3rg11IjYl
yiI6AQ8YvINorfU+ii6CDCPMbYU3tLr9qtiIkjbASUXpwCUl1NgwgTq6Q5yd6Ud5qnpXxlDOF50y
bmQiGboUMgUXxzxi79knoBQB9zN1AWjg0btriAawTowt30IRVgpLcUYNGViUYcWhr4WkCaC2U5o9
B15M+1mvI/OYf2IBtRckTcm0FovNCzZ4LL4LCgpo2eQkQeWB/I6IE1gyqOpnyMh+yZMuIZHRmV98
KR35lsibT2iTC+XkfQOBgIq/7VSi+lC1RpbhxuD76k04Om19dr9RUA8v9lOo9sxS6Gt+hxL38vv1
nWKEC2AzMdoq41dGllUvgzAaCXUv+b4amWnF1QshWBWGL85CCnIYweertl2Er/aL5a2zq3AQLHVY
rqKlg4p5dPuOL/W+cKNtf0HA3/h1T8wOtB+KqklHR1QSUQqxTMajQa8476Lx0p7qJVMln+XyWDy3
NjINZM0NgVhJHplQqLIA8xRAAoT1xq5aI1tpGBxr89kiwOVV2WF+rSN6rF5rVjfTwnyW77QzvgCJ
E9LZtX/+O8NRawrc0Lhlt++L9vFiGezBHjgqzzbBfndNVx8tbVjZ1mm0r0CNqvUhtPOHXeEnW8Qo
HzFF3gyX/Lzyr6uTZkvOecBFfI41Do5AZNM4O+3NG3+uJCTaJMEu3e9jzh+vigFzOaLMio45TSBR
FwuSGqcYXQYfsZATjz//y3TYCF0pqCiCtlSJX6O2mlI2xQFRwpolic9w4hWMK6EHLZoZHbA8NlhY
goEQUOkxFRK1bXtFWTqyCRrP+CHtNCDel0Z4kVoHSwO9LNv8xQOU1luoiknX4gJogTi8T2iw/1dC
f7H738DKS4qTC1M5Vq/7xRRgfwO/3UdH7JjxFzBqDxgqNv+b+Ubsuid7kl6j4Klcu8UiroQUsStt
F8JYteUVgiFZa6ha0m1GiXYHaYLO3JEwCNOv2Dh9c7Sf0qPzPmyxUTdtRAkrkR1utzGBKE4A9nmY
/o4ZV5J9UTZ51IfIjGpM5POl2/Gg9g5MP7vVCs01nJ2/AayBlaN4/iCR4omabWmBjeF3fKYzfwXi
eJ2avPEiB8dX6aHAXoJ3guWxIVqOV+bQrh0JWv8hRjB2c6Igl+AJuHMKmE9clHzxLHSuNMpHRiXz
AHIv+7QNhDauqJz9SMVojzND+g3FlV+c2NysGE5cr0S132jc+tfiUmIxGgVycvnnKb3VGjbY+Pto
bInCSNBOAHtc6ZwmyzfvAmCMg8nfbP/ILR8mczr9nj45lSZH2w7AF2urSyjTL7+vfqE9LBil8gqX
U/VYHUum/+o2e74dgmQbRIWA1D0hEqe9QEfS7hkILxXlu4PZuqZsrJzI76CBS8QRsdVs0H0/XuC1
j+bWorBN19hF1J+Aw4+m/ePunILk3QdtMM9iBa5Xzm3PXjOowr8WAApwn575nl216R3G/xO+IzjF
p9KJCoef4e7DzLAf5y21starx5i5cEjxgdWQJKfZZRTm+CJ+YMzBRL/SX1csvhSK2TnWNGEJuGe7
A61E4W5m3oGiNYA1sbJzywDH6cU9hGdwom9YCBN0yH+ClzxnxG2ns+KVDHnrrNNW2LCHCy2rXuPJ
6TTj2z1yLFNYDH3TSTIzJXfLt5lJGSNYrFY4ze6FoJiY/ecJdDqr7qDlZ3ZQrx7lemqxOta4SpHv
N85eUnV5PurajmYdSiPoFd8cmqRYkC87pykgIC5QKVdtZfdB+fuFzq+UJOvtdVICq7kypwGp9yii
sHFd8OLUv7dC/RmS61ILk9uP8FLi8oJIWpj8bohvfR8aSB1P3HCdkNi8CcNrQ5Eu4Tg1PoUQTdm6
UNhjUa3rRkR9CMM+dQyxCNfobKmL3TeauM49mugEPq7sOXzhwomISIyk8J1gN1K/B4ghDRU5Mtox
caWZkre7RBCWk6wdo/Xk4QopCm7fCfMkkxddNNH3S0GoD8Y1yXdd9cBDb7h7bDuFf0bt62784Gaw
0geFqqhnW1h84E7d9mr6Ho3B0kQ9caZU7VmFRBo4KSxYl1FIMoSq/LoAABaSqgKj8K+2pwvnvSPJ
F+C/0eqUKYposDjGfNT7jNjmm0QO7SFJLnRJOlxNCmyE0Q1hV5RtZk0kQ7TCitbX+WWs5U3eee0z
JMhrQ6OtSxNmoOsXnK+9tGJbviO7ySXY25d/1bkEFoatNGIMfLvvQ71U+pX8JvrRZQSZ7piBVdQP
LJtesgFGIDjsbr0PNiVVQktbApqRWp9qcR+BOm5pleHhIudWttTCHWRWk+g0gPxNbQ8XazD+A8FF
x8vr77FhzkRcrRqTD1yFU/j3tOrbHLJax/9V2PB/MuVGyfoXui2qXQ1rQ3HleJkkEFVIlrNjbp1I
PGCUmoeBA1zoZpw0JC/+0LFkGmUhfb2EEnY/ku4YKySSgRX284Tci/UYD4D3Z7aD8ISGN9jYi1w2
tEZXOBlHsJC4xomcn2h6PFR36tv7IJjxEOyoL+L7ClkyN6VRezQ3MHIqAcCoUrLsE+s1Li79RK08
2ZEHEQtVqTgLIcXgcVskge8hsJo9JlQiETM1FhX+HwTqckTF2lFGSbdI2ASwsKHmLY3DG7B7LDUs
EF9FGPC6sHYQWUMS4WolqUgX4ZI4sHQyVfHJKQmmNZRthrmHqKBsPsikQdBDDOZz1xqDy2BzjOk2
9GGDDki98EOAskWzZu1qBNq079AP4xgEWlUDzc4XVprpdhVFj1sP8wJjLnauHuU32GsIj/0iiAwP
4JSPabcBENj0xd1hOyy9SZZLz9x5oTA1SfwjJP46gzKqzWlJPaBhXOmzVE5iohtKSN6AcPXlWyZ0
BkKO9cAH9Lg8GH95ovYjd7ygItjghlTCENfcABM9HaWuWDXsKbseUhn6uQaL+hchr2Yb6m1KvA69
/swecvjPeTWxBTIvIcbNTxi6q82sggBfCll5YsYuCQ+gp3afUmhastEtpjRqRsiWp7oWIS8wRhan
CglPz1jpWK4gyjld88N20DQ7Dm6TQ978tmTC/ZFxznNrQBv216WbUTdm7dkJfOAsRnlLd5kQiAGY
aCKKc5Yn2tDcu8o2BlLXORm3mnwMOZ5SLm6zILgKg5PeensZYqIBczGOPRQAVUUGVYeIj/CPq0MS
DABL0/ZYGJ9BfWRJTO9Rhpwty2pr/NNZN5QEJh+d1xstIPvZszWChU68V7kJqYR+ED19Fshvq8FA
ziuWrk41UqsDhlPMlUkGauP+2zXxIlWpH1+otOkgJb1fBAaUUtJg1HuVT/ZIIDXguuCpKtBZw7dN
SZBz8n71Z/aTYo9Bsyd7ajJT7tpE7WnTsEHRIjH9MsU5333KQZE+b91lm5wA7BdtuDydUt9v4wOn
mH0+PXLnCCaaMnoH+GPMsCufdOfDkoW7wWQSfK4MVXtu5jJWUVf3VoU3N6fMEOz95gODTDN4L1+E
brto2W7d8jaKKSvXWvbJlACbGRrO7yogCPmuOgAx7UzNCKabO+bYHCxWnnw4pNnpAjSC2IqA5kod
4aQRIuzzAAUXdo6U5BOl1ImrIcllzo1/lMDL1Jvg0FVC1odgwajKlGfMtSjD5/bCBmIwQhw0HZpk
4WmZvxhUVUMr0/ye9YapmRiTK8Z2hIUuvyDCAdAnqool+S9biX8D7bEiXZ7G0z1M8sh8PFvNGIPi
NPgAfTHJJ6QzXPAixRNvoNfY1Gx+ylUwAvtMxRKIwJFKa08Wegj6jsWgwM5JjEDX6RMjAvZUJjUS
uiJBWevkd+ngFgWwlQdx2xnfHGMqVv3QAR3Q1Cjudbz29YWHmydadZw/Mpk/4+OrWYf6JwbgK/B8
uORs1b7CNJGQEbSzNPubReKd0cC6ip0MKkzIXaWisRLTWaa82EAbGylC2GiRBzQ39K/3Wj+uaWHx
3gUiu7KsJPXPhLzKLYjBe2X45+QoPAU/kksYO1LFAMIl60zWLvQ39nAvANlFC8bo+CM0QG+7QnY7
78JqzTmPZjgDTe3Q7muB2cL7KlxxS7TiZMlQdi+VJskKIKluRUDWTRt0csjnfctiOzx02TmAL4lw
/9d6feIczNNBC/I9bdXKWTtHhv/8vOe7cyEapleHfNTUwwgMX8AO/99OQtEfWmRDzfO5SSVRrshY
2KhlzX+dSWj4020kt9mLF3NKae6oq5O9Gsky/USt7eRAsECzaIeOO029eGq0zg4Wg58wbqc1r7nB
sNwwh0oww+gUojARj1ewsklEo9kxWuxrdNj1szAUhjKAvLccme76Y1xTXJ1rJxadYQROy6L7GdVc
0xGxHqlWw6Xurcwu/vAlm06tF1IqnJ9TPHqRfXx7KHofj0krX5LpnykEpmLYw4SgE56OmuuXkvQi
X48EXZaQcNuWV6+iYHjp2lP3J9n8x+kE02ZWeNS/oI4ePK6s5GtSbjSWyy2ej7UdJ8VXYFJ7N19A
OCOwp+Fvl0A0qr8LYqyOpbronkqLuzJpEQPnmB9pATf95COYXyXCZYOmTPUvpSlWCRZTSyQJ7n9w
ZyaH2XhENkKEgApYio6FAYyBtLvw5boY7PWwgm+qoqXItdQ5ckCrRr9tewhlFHEHdwVN0sHDllko
luv/iBYa6PA49QvzsevryNQv6gqgDczYZVmruvW0NePg/JMuXCs3P6SxUacMyyPqUrexZGCpMXt4
/MoRQsJv0E4eHCHdapz1h1NulnnbwQzs1v5Vrt5L+KxLLcJpBR1x1fZUfueKH6sCF4XIH3HJcTFo
Fxlc589UqOdNvvQFv2Xj1XUttM740PFAlCjCjboiYWBhKPGUtvzT9ye8ZxYRSZS4VtpuWWUudYXY
jMN7O+redRNH3jKKyuzULLwF7U6Fda29fW57khNj9TsFo+cEvf/EreXpNuS1cGeE/TL35PaA3ZUm
PuYRllvgGv0kswI/E4ttrSHD7eYrDNI1HWA3ch3+clyNesEJgws2HC+ucgPaiS2aJQ5fwCk36fX4
0b/R82Y4/DwpDmFhR8yr9ds86EsNGaih0+jMCmzOTmnG34sLn1kVpRCFAqyQ9divj2KYdrkr5GCP
gNY8OswzxGzuKu/cZlXajRfAjDFZbtlTN2IpuRCUXXC47vLqVALBCa3+NNvitbGsyzyuYE11Xav6
pctdAusfaJbhE3ZUvMp/MKXKewpxKm2nrREA5OIXm+1jtZMcZoUN2b9KPybybPbbsp7BXQq9G03H
sZs7mCQzvSXrMCZi9+3UErzgao8/HDCWvOUOXOhjBQuyiM4ZbyyBGr456Z5/iYweldmv5KlTrO8q
DA7vziBeXAhj8Rj3ebLflf/oTDwh1DSk7cyRr6JQS3CeWMLkF4/2ZeUDZNy3dqaZVCtuKtGM8i2x
Vuv49MS8oVyyUj2/PXrV/z6Uxr6vxyDsJMM29/zkns4ygSVzGohcsJ4fViT23OBw3/ZBM2HObDpQ
I4n9fnMW7Z0vwptdjcQ8r+lAN9vZz6uxu9D4oCrWtYADwASXu+AMQzlinc3HjBa4q147SWSMHNeN
tXbKTDS1uIM1L9Vrvoo+R9n5EQ5cBo27fgri/qOt9fLBCSVebDOrkazXwwlrl0VIsuwkytuRIwJY
XNQzevp+Qi2i3okJBcTQppH83VmfCWtXP44rKCo/0s/HfYRWtkPtVMCxetCNxCXBsJQLk9NF30F9
KJOCE8r3GW6DNptypPWNXZx6b4mGtmlOIpEHnPex3E+329gqrRrqF0RbNOGiYN/OoK6cfGAJ6lqQ
tQAv6n+b0hnTkphfYatE5VIn1JA1X4SLYVF7gvIm+eTrtUCXk1oClx5Za0hYm/pGm71EAFdQLRKq
85cvssQZ2DtzORYLzxdPF669smFrFuObaHEDM80loEHe6zkgH29in70whKQp82E2XK6u0vc23wVn
ml3oDjI2b0mifVrges83/n9idEPaHpKDkDi5k1oAU7ucRXJ3gSQKdg2MyYlU2sQDdJdc9qSIhzAn
oulaGqiU465wMgWIGUo51iBrh3apBuK4kYriWAcohdGdh2AI4BqG1e70dn45FCpslwby0vu+SPgN
KGLFG7g9godfEeymkiuEueEP9LaajM6unCW38ZevlFDLSTc7jj2v7O8B3b9eKUOtWzehT4kcQRS3
rNuS4WR+/7ro1JNFIxrPNOpC1AGbh96gDdEJESKTScNwWNL9FclgSDgXm2NFvB9aJH8fXB3W43Ym
dM/IhAfAGKsbjuf3IrtVQZ2jpprHVa/4JNizxLqOmqVj88ar9g2Ht4ZMIv/QzQLZ8C0lGIDO0euQ
uNH0NIKcZEpPcW6VQaYwsfuQwg7UANps2JbaXFgvUrlICt9XV0VUoRaK0B0O9EwcFDziYRX1oCJj
OsTsVV6L8/BYzvrD5W8S9fIyQPRkB5THqfsm9hbiZ874R60/rSzn42MZQgmD32gFbpsnLUuxsKtO
E86VJzLBIdJrU4xND8OzADBNrktPlzxEp3M1EgkeVemQqPlDB4OYTky7zjXhdgElWCiAda2rrDKx
HxjlevLoxuR/DdE/xC3r6WXbsH1vDKXBviJ5JqbbX+WYAi8ttzyhuV6FgetDwil5wwsjjM4bzke0
yu6zdmf4IVfGsMy9ZY8lKQiFnKUuPtYEPmHY6Rr4qI6a+CxO79jaLKnc5ecvQioy54IEiRK/ygb+
SIRajO3eOQKEiMsHrBTvU3mXwc8y1W/b9d4LdL6gmRMdXoDCV3Q6pWDImJ3o/lcgAZGF57R/e6U7
rqZPCpkoQU9Wb+tJjYhKH8u55VoJjq1KfXDnp7s/cMO0aoDzlyu/ie2AF1KZWvzSRecx877ribSf
0ePzZ5LYap8bjfwWXNgAV0MBIIvGwqbZzhbGk8agG0tWshzqPpbD7s3W0MB4q1BMPrIWAJ3w4F9g
3Y40dVjfnYfHPyhvnTMdpQXh8EXkstt2vJ7tAfC6RGe6Q4PPGAY/URWYQcjHX7VUoN1aqkibCGZ/
CheN7GU6cVZ99CZeR/wU5ZI4VVEgUOCHh4i3XLlCqbfDPpLWR8qfJM+b/d+Gf1xheOy6fatMoHzc
BGf/YOT2egcVgfhTgswvZ2CjOGAdQcToG/MfoM60G9YkcAQBBIlY7m8yFTFfYSJZM54t8qrl7TnD
8iVnA3ycsLtsfNnGeG4imuRv8+sGJV0PPYj/Bj/kp0/MW6NwB2sa1KiB1jIa2rpF54/oEyfISt+h
xhil46jqCfAj1y5jnwgoRhDZlG8mvYzmscTh0rwcVAh/uPKMzAeE+7l92e5/wL01YunUX/UQs5Ip
DaVDMiIsMXT7uxgBtOvafpraM9pgvRM4nRpKo3uX8YyOhC9SghxNLwmuYVcuQBBIqr6vRYiGPIVo
4nvFQKx/CBbYMCSIQBKyn0nT9WV+GX8bKQnqyiDA4h4HgvhO8rI9TVZphf4RFQA1iV1mLCg7X+UN
ExFXcjl81xufm91UtJbtSoNqPKONlWgEv2db6LgePvtGdeJ/L3qWz0H19xoHM3F0AYnRZjlKW+Ah
wlMJ8DilqcQK1p01l1N4t6Dx4ywlkklvt0awHZNfetGXXOKsGAOVmAZD2zPcCOZxinGg5bs6TNPl
5OUsUq/3qYLMx0hAooefIg3W0aUdH4GzryntopnYYGwHb0ljnQrx0a4yImppgjX2GOLtu82MQAPf
91hmoIdw3+h6+a0uvEwCZYhnfQnW5DUZrFqZUTUbxqroR72dG20WApA9rSEZlYGAPbyaDHZWowwj
ou58PRZ+tOuP/7YxSDGTqoqnsxNJO/l2Lq4tTuST0eK0SRbM0UonoS8ciCgvlEIMdSRxBHuBuMRM
ShZbE+l/WDjwLPq2007rY/YWYnQmotylfaxwVovsCEDoorPuH7JtIa9z7bqXxiBCsMTQXBFP6s+d
FL19M7llEUhcEqhhO7Igb9oMN7xHbMOoNo+1spqcAhWnKX06QcdxrF2zx+qG81ant1R9ovp0svUR
jBeqNQIa5+9dVcgKAJYROSvwt4B7u4T7pFUmaJ/9QQ0h+VGIT2v6iF+pbjxa5L11N8ZCH/fY4Onc
BIOSw2LcSylO0xZUafl9Rdj9V0+Nn2GnIefN7tCjg/dH5UmIp5CkA3CiKT9q9ReNEBrRm+Fm+ZSn
yAuJqN5kucX6W28MhBKbc18Cs2Oun5L+lVOnulWh3d9yjKic6eEoPJ6dLk+agdBIQNjFtXpkDzWx
lctDWrlz6/SWezHbc7cHeEI89sXR9GX2THBQ9P6DFPG3bOpVXKkR264PMwq5wSkMJihiXRwyU/IN
lY3MgKtQx0WmJra27nsIpQ0z2oFwQOAe32jC/ZKVIF32epzVoAUys228oo66d8/T1UWqmDR5CQMO
+1cOeGvYmOHRTvAZpU766nAdYRkPfSOwq0CFjvspQir1mxj8yDzk9iSvpFiB/PVbKreSquPfqbPK
gCLH56LbsVTTqKGzZvo15ZuSM9FZKSxfpguxpgbbiJTPsk86IzvQaH3KiOOqwA415I959VCNKFJ7
Tq4IYh3B5gIt7AbZ96tUXM0IbjAR8h8t86H6FIUUSBjU1JEUPGAWBXMqIU3qZvZdp29R1dl5IOe3
9yEW6+6e1Z4cIpsXc5HjbI76tCLDDVnlqY4lnfFs8dT3CQh6Mc2BsXBIeCSUVTkc3z9PQkHI3gLr
BaVTP+N++K9ntxfX5a7BIaejWbRBsJ+pdl7u/8g3LxxNXg0KZRRJ20l8C5vWLobH4zxIJV49esul
1CCXZj/seyNXSbyYEx7lI1Eog3y2fpk16mIEztMQGzdHCM5BfEco3SCk+5Fo6Y6lbFVxRITQZP3k
cmw1Tav098MKHJhyvTAIBh++ru8DP94ZwwL2LWNzHf23WCcS+w8BNRFb6EDzKSRjU9ZQXB7v9lwd
bRLiiizEXplHWmjD5b/2l9XuXO0YpIo01UXnmMvXexP3pg4fj9iqczueRDcnzvNwGzIWFsQvGc4l
OF9//21ivzUOA3NmdFq3i/YrEfHkOkPSx8ppWiWcPC5BK7usvcvAUzPrr1BO+UbjtDOv6SEYUBg0
c1N1rXosj1VZSSZP2dsQAuV6YrJmEysF1uHeEpCb+PUHFY6yXWIf+Rna2mHfZN2Nd8X+3VdiUD3W
GpK4V2OXgwjZcRW6HAzAkw4fiyg3PA67a7AmF1heC1CF3kyc2hhQ9iwV653PPw7iscLZtcQRb67C
UMhT8I+T/NMU5wNIFy3N4/v3+GRPozZINnk15DWMj9zDg1gQloQEo8CeTAbQXo9bXY6BfT+nHv0w
UY5zjX7QvYHhstIjxBPnTYNVOMCV4uU5qikQfzRX9clyMpf9iSXkulkJMSyzy9evwnjZRTIxQaDq
NVN/3QYCXygCl3GzSYG0d6QMwZKOCaiIhjZJACScsAhosi2bwKJE+wAeOAosScuoeTo3x9otEwFT
gmhTu3a/SaPIkhoEcLdTonyVvoY4cBNoa++UgUGYk/qlb4bCEP0BL0U7+ZKFM3ZWxbIDw48nlSr9
4EWrexc4YP70ufrrQcb1WiOjEY7FA794YU0CndawMfwmFvItIi6kYQ8OxU/mr8RIiwJSYcdfJtXD
US8A9o6xNdDKiVtfqSF37Vm/LIAWX4otEcNQlbXAUeZECMQ7dlkosGA69DvR0wfSYJeowRq7uyPV
yyf4gXXj4sMzB6OjTmLzvpNahz2J2ipqrQxCoVkfnwwxGPTOB9NtC/C8vgpcdmN+uwEAdM2y0FLn
UfQA5+QxeLKxBQTbSxhc0+iMLITovY4l1CvC8SDU3K3qP3b+KdGRmTxwzlmGTUUYoHulh/S9xbr7
VRxYVxqlvtZmKLYWtUYzigDro8jfTF7EWvJOLyMsZqF+raoeeLP/bqmjoxbRyEfob6cgrq4GRk3D
hS1Ayl0puu5uDENoUgRZ2x/I4SA3CrQjAjQcQbHPb0IyFSd4srW2HUUsL5KJ/Tcx8iONWM2wF+E8
qupkcj46hEECA9HTcB2FIiJYSCB3vBr/Tdy1J6Sh1sxaJNRAgUVXC+a4WSMbNZRwYBYHk5x8gNa3
DeqZmN1GuEXy7IjxI5rRSmmZSq9S4l5aAe+yBl6amwQkBfo6OI9cmN259M7QTM7nw9+aCRe8lBtn
5NIGKwxpxiRbe09N09Fjv2dvz9zaXCS/8W5BJLklGPwHIa3LLVR6sfSa5d953KED6oLLskynayJT
rPIx7Q0eRdM33m+fWiwgrFT0UO05hETNNst/N9uarh/ERYkDygUOWAAFZ2YqkMBfTVfyzz/sjoOC
EHM6s/5D/B6J9vlS1kI+Fxx70LVYU4mtthpDFgrTsub2Kb9/oxKAE5blGgZqu+U/XOOa931UY0mT
kx8w72INUAYXznNbZQLVBUIN15G6PQPG4OE68H1jeUkn7OEUACARY5uJAHs+y346xgiHmGpMA49B
BkWTzVnY/vyT8l29N3vDOYmENbyTlUXsjuetvrZQ51CeJ1hqNYGkHcwysXmUL8XjBfNCd+aUDnnz
nrAwHYdmLXTOGkGYqWr7tgGPUpaXpCCSqPEmCS4u18/eZCP68aDsVYgGH/jiRfqCB1cyWKQZNNB9
KFWG3XFX44Yj/BQPGDvN4AhcPZ/L1zG6gzPC2+2gnXmxvAc+FPz8jU4K4Ak0xBV2juyWo+zsW+NW
Hv5ISbcLMaX4orYkyndqUb/qjJFvMi0pJ3yhpWKA810evTEpJnC/JR9YKuGHMzTgKFAwv0cQ3pJT
tLPxKcW36WP/Yz5YET0Z4gn0Cs2rluRm/hk2P54ftFlhE8oAv/R5cTrUCtoLEEjLh7jDTDO8gC9X
bvIo+/dtbNOq8z1MF7xkysGZr+vfuvtW/9qt3OFJ/wV7N16B4mtxKPhBPT8gXxHJVK7yhmKdp7My
yCGL6ZmulLR9VN6k2ANU+j7juMgI2Vaq0RmwuVtswlUCWcQz+64Y1lZ5VIb7Jc9FNJ6UVkyMXSEX
vMx5Q7bnmehKmpGA/LNV6pDOAB5oac+nLSgLWOYTgZCpdtoQWC83UUUgYaprK/SSceQVEU+tqCo3
u9pB6VsjSmekplnCHcjNG8uwdb8qcVEd+QICfsHLQPDTqTpDCKFr1kRfNE1EB8kZcynoYfO0RV9g
gELR9IqrIjy6znxErR5aZnXzBVpcIbHD1PF1I6g/XaFQIGAQVbvA2jO13AMiFxqrfkgVUKKRajjz
09sdKDJ8+76PPSTYAC8dNtynoV/8VTbYMavnMi/ECtXm/UFwlMonEbXkq74ezoHZ0CusqswKmOKS
SnXJbv4o0zH9zjLiL0AsLe8aYuHtWlIfNBWNQGWrAmeDvOoH95isb3yuLyNSyqL6b/P4boztNLKO
5SOFAQqQwHTJsBwzftcW+SqNk/9Q1yPp6GwI9zX9yk6hK+14Bp/IGSpZaYjuX16w5t5QaxIGBl3q
iYnRRnJY4e0puh4RVPaJuazZkpThyLS7fwwy7miD/okWsPEnPF96Gco067SgBd/6yqh1DTpuhfui
Drh51MeU1snkAXs4/0oIa0pQYDhO3d69ahtUTfot5jILxPdst8MCslLuVWBFVUqE/PsocmuPFb1z
qRt1ks5l3Gvcz/gfnCvEwLbTAkDMZSvb0yNH/FY8e4GYpuqvXAKx/4PCymtRXY46+j6Sks8dwO9N
afAoq38BwDiuJfWZEeLLhxcfElCroxD73WLojwZHvuIRBGnRjVZpWZxOi3C4hhsVzWsuhwSuU9Fi
z1xU15TkRzxME1kEV5TA1GGBzVocgxHlQ5D8NMqvkvxE/0g6S28YO4V/pn5zQfXB/SVNg49PFojM
uneyNbcHagtENgxksEqZtC97Uup7DZilLQ7OAMngqKoT4H4dvOdifUZYK1DbtzXMahPQEATNWj7v
xjO+VGLx+AUkJEXfOJt6MR5u13x9tC16FmuPI8aVg95WoEQVvWBUPx9aKOW7gjClY1WzSbgeKi2+
qXyFkm9scvKppu7EoSYPkMM3QfmzkCwfNNNdTRXYJZY6T6vK186MCfpyL1hlI1IFXk8E3DKlo+Q+
neI1ENL7Ve2bI/IBD4CiFe50ikLk5ne2qfcEOLqd1RNp1uDGUxPqzNPfVlotmsmNah4HPGX/OL5V
SrqWtCeOwq4XkkLqCikJKtubB+yzBHUf7KsWKF0xPbxMCipzFRpgWYD0jYO4x1ofWUu9AUaTItas
3xaUfcCtQ6IKRntBCo6ZLPQ1eeFrUYiwWlzbI8yUBw8Afqmvj7lRHh8ZqQPZcUHpyzjGnufpK8Bt
FzSuGzTI6ALxH7mhmGesUd+hFTA/wdBTFbdgUlrDfK/NgB8tArxkP0yWhPUa2lb/tIUN2/qw9vj6
plY3gH+txDBTK0+wni/MS0hiJUvTNDaZ3796z/rPa6TRCDKPPn1R2YzG+tLuzpaPD8PtIjih7Bpo
/O+yFF5n+OZIlsbESe+DqQQuxRd3pLKDcsQDDhbnaD1dNWCA81Y3dAbVny60ghGOyzMnI5amQ58P
Uqh6Qgzfj2bz32qBEg2DmKLx3qMzpQ9MuaAu+E4JZxRVeJZrq+bHhZCyMGI5y/w8EN9DXKiKXtbE
WY21dV0R4EtRgK/wrTgzaiS18+D148C3PO3y2CJtA9rsfnUcpMH0COPnp7FoerdiA2YmSGYlsxZh
pfZTWc9ewCcDGUfNZpOJkAjADMRmV2PSnGLjXAILfPNQPHXFJndPaChJE/httenY9d03YlDl9JHb
jUnWQ9Lt7xL5WMDmgYdS74y4e4aLePbeYiwNcUusAGNELvCimW/S6PQIF+xbzYfDQ3a+ugCsnDPw
vkoxRQ1LO2RRPyVGZAfyoj4tkK7+Vf7kEes5ooCCimF3ovI9ReJ/7RX0Bj03o/z/EgEhSKNxH6M4
caRMJmBblYThvwf3Fuld8w08rLlsDLQeHgDhlyKWn4j6eEO2JVn6HFwb70BE4/VvafcFkphJKYBy
OvbxM+9oauJKnW4bevGXVPLCJap+/kPDIoYpBcKP6eB/utqVmAur5Va7LHQXkrMf6iNS8vL0Od8/
gytQzFMJP8LNBXi0vg1jWuW4Snzd/HSXJE6f4AL0V0/c14yUt5tM8uWkekSHSVw86CVbH3Fd+mRC
LimFtb2b95+5c6wPNEAZX2uvPhERqGSGLqyFMvBrcK9hESELdqWjLRb7kF43OZlXPmt0DkPmValf
3uugOViNjBVTmWbaT+s9lmqBMxUkkcaza9SwUpQ3eVqy8p66ESEFrPZ03Dk8CYoEsGkZfhqZkolP
1T+VPJZbFcorwOILkgWukOtNYnDZxNtr8kvzgtRRnm/ApFEZi+ZwUdmMca45DO06rLC4D/93VWSa
1mjiXmmKSdymOqTEWPnBO1aCxtcu4djXTTFcnr5iUcAeOWJy9oAPSHb+++9Mk8xRF0d8k98Eajuf
DtB7zokkCbD+6gOQLqW7lGS2evF9EHJW4mCAhbS4TwnxKgnhhLEMM+BnIerdparTS+M/3fIpXW9o
N0JVBx9YIaqhepllWKw61uZ1DqZe59oLfUUb8JpawCwa0aWvxlvDWkJKzaQObeV5O75hSqE4oqKp
ZsMP5OJvAxWQROaFGZczD34hCsFJXPk9wlETHIjT6RDUwsBsaJZiihxISqxlbJxSHawfbKTu3SOq
sbGhNwPkTD+Ua564WuPldHKIYZhcBLKUQP39FS9yn7UDz2NAMCenYeINiNP/2B3GwyRlIxtIx7Yx
SHfnUgLeDiIOa9NdAsnoUbNDgI03QhZ1r/UFX00f+3OgqtelQ1jkHxnB8z3Ehx5GnMNPdob7Md/Q
fhajzqsrlYP1ISxThyBDVIsCsmIzcQLhuvGWEQgofUNwzody8dcPPmZMi9tWMKC2MAKkjwia8OC5
9zUIGS/6ilQdM+g5OqexPiLqJHnYQ6UhguDFagjoBZlulQ/Gg6gQsBqlybBKKRCZTTup3MOVLaOb
X2c/ziB4Rvxkg8S3Y+M5P3Rq+zqoKPzZpP8Sg4YrUH5wcGmyOkfDBUn2MeEMmDrvT/nINqdLlucb
4kjF2MAQrHAllfgJ+8FBFE7PWn2+EA4YtmuiZy0hCY1+k4WDX2R8Bv1crw2PRMM7S+jeErIdm1eg
jdst+G6X5I4Yh7CGtVbb+UpcpicGf8V+seg3jQThLLIu7gygWmUJMqakz0pLbn4zpdOHoQxW+usV
YyAlPJhCyEv4YUJvZW5foVNFeEnsRidGTfThiP8+O3jxIi3H2IOwRA+lh2A13+Eoy9ZT1KSAW5/k
JNje6hG+yuVlhBK1bkpoFuJRNtur1S5nfBjQfzLfGrG/6Kb4Zy4QEHOVjq8xMYEy9fJn1vgqOh92
n1HiDxBgLEQowl58TPTuYUFu30MStYsuaJF6O7l6wAVtpLy/DRK6fZ9xLo+BqaqS/RNOgCadoYh+
wxFs6JM+lHcNrl79F7GA+/zDI1lKKACF2G6Raxw86B8nhmn6j+mueyZHWku7u1iky/VtZa6KCKU3
2RctK38EWqlhAUdKhCDjskKOzIWC7eU3Dm6Kn2OhMP37iAMV7vFuurcRDRUbBfXMLwjHgec8/Nfn
777S0IIVSaBl92Z7QEEEk2ur3HOsRceEUWPHcEwS2TMfPj6BxXntAEtHi9z1y//3g7lmCtEId6/Q
oQSm0u5YuP65AqanogkeXoRibSvg4A3fX6J6yuPl2sl+elJX9YxYGePUTWOYY7kEyIsJAWbHubuV
Htx7y6pVqQ+KxEMWKKF3DbvktWbsgNo6DOFncCsYFW6eLdUPkR3qdY9HgHBt3mQPfzs+/i1RCvs/
iepiDs+ourw82Ox8H2oB+f7JxU4NiUjARnnRmy8QY+sKFB3XSPFHwc6wkoGRCUKjIfJKPEnIloCJ
kYuSsJ/1AVcDSSKagCmNe2kdus3PhLoZ8odxmu616lxrxg4pAlqgimnsnw5RYgatvpvBh7107dMJ
cP+R4YWqIXCZLI7HcbDe3/4mkSpVroMVAeL/onSn1mvs21lJ3epTRXIgtEO9CnGHyL2r5Y/CLqWN
E+EscYDBvZW6z5i0218gnB6uCgl1zy4ahg3kx7eiaAYP1zQQfnIInSivi/OJz5qtpM8u+GTm73lO
Wl0WLs4utz+jAjRTjLPNy6uWpulKIVeqkNDFBo8HODCsN/5cR0RLZqa8WF5Q7FCXX23/D3UKrpYu
nBKE+WX5Zz5jqS4zSuMBmEY1XFtm+caLwEVt/odESJWsNbJuLBPapQJ1MrMT7daB5wsaYqT2tfKc
qRVZGevnuXV8FAwtkKrbiUcP/e4+B9O2uUIPgcvGfGGZqBuMpgLCZfakFsj1lX8u3ZA0LfooFf+k
juVKCe5BK79PRcXAx9jZNhQLDNISKaK6UuvFXFRfz765Vuk4gsNiLW1PeKzPdxZ+tfU6xgn3PPKQ
RSTkAgQUmmDqB+xdKsSz2K0VXP1dOVCshCE1zJPUK5JiUH6cDQLmMwCuTiGYiic50hqDxrMYomgb
mDAJRgpWAJ78F03Pd//NWkCK7Af6EIjXqsyzDpAQiBdzq8TWAOjkxhsH6Y+3XTRFonFEpErWCcwk
Hn48P++wpNsfRHABJZsJV3RR3sKrGTnoiGbSrAxWEtbLooLf4NaKPpNs4vrDNYgD6DwYLOWZX4w3
ms5/0o02s59X+rlwjPsTyr92qinpbfNjR0b4iImykSc7GdmlR/9JoVXNJfukwV+7hzvcmd6MgwhR
8wXcRDbK9tcSXfT7rpXIrr/3Rqwx2MJZ/mS3XeCeucDQ9hO7NVsQoCuZkW6ilXCDUKggbxGGAiIL
mxvgzNDAnXEGtDGkP9iTRWoxHm+2jqxThZMEDhoDESSkS3yeyEvwuJXIsr9d8BdAihQEYs/uDl/J
7G2x3GWmgX0WwtvBDkMWWW8AFFnE/iAL5nzw4nnLvaspye4R2aP7pPmHp+jLz6TImjlYXGded7FY
2cQUkOFowVmo2MO2Tr1asaryCWBF7khnWGUZuoOBNsZ60Evx8K1/juxk3jCItUCKpNt5gDDwdYNi
QdX0BxjfL0hUtyEGZFQq8gdWSh8LRcgVFhoILFXXmla0FnoUQCbVzERWETOV1M710ELBm/LX5wT+
kbqULKiqmmgpUlo8ZakC6O1a/L3MT2X0MLw9Zak8J7hhAhLCUAfL7OqdkhdsOxlDua1Q10VrCGXi
vBmBD6Q8Z9IQxZ633iaz8rfCl0OvgyeomQjoBxGTC7VbCdIppTWSfRRnp8eDMzaJ2PnOkN0vuQlJ
8GDzf8lhOslTNR6DZBQxXtdUbAURZNw7a4EI/XZX9CVNDLinuKkiLyd7xI8Zg5AQaSv/95HG6BM2
zR409Rd5yHIrTuag4kD6ZppbbB+Qs2k7YGOLVS0jny57GJ1yMtOvFJ09baeIGpqQ93SRlBbH9U8m
RIcyCJA4VLaXHJhl02Bj6uUajKmJ3GFjdvYcagc2ydtaEGefZaU5aiT50XG7ENqvLqdjfMEr3K0h
jB3b+L91CZwvK/hsytbzMP959uaGSs1Y7lNXAyQAxaHZ2+Mi6T7oDkMfegL308mU3ZAzPXDC23JK
I2140p5LlLgy0Wi/QTf13FiJ2LaMms/Ina0bEVg40EQ6Mzy39wWXZ7P7Im+eWL0cqb1nts8z2RI0
K8RfDBnTWKGzPp7E4RBqzrxtCANgKDuiPbB7avvipfy1GNpe+jov4kLkVRRG9wMzvYLwNMl0fKLq
qykxpJRzbZV/Bf3/GFn2UcRqQihjOxVoV3K32HW8U7W6OT09/I2WOWzLAFb4ZQ6Wu8DD5P6Z8osu
ToCkcIfzqvzi4ckIhPskNfV5uRD+FAwo9d8ng3X4PRsTrE2Fp+Ct5S1D0kRydl8QJU4WvCUlxZT+
9srYvre8OA8R/wtiuw/DAIz6BBjpg78AOZi05HB2ZCePBjD3F5ZoZNOj18acxoQDxOUCZPqnhGt5
UpxwiFXpXFiPdAVDb4rlPjbJkjDrRyN2rIQimeSaDFlVllcW/1Q6vLKNuxSg3r7fwVF+i0VmqCgc
hcB2xeiC0Abhl6i07ioJ0bsMXZzycVHSMo6+FoRCe3Ua5fAzHDe0pVJTdCnQz9Q4vpisJOwk+twY
ZjE5hgL2Kuhpnk5hlo6wLWh+XiXwwRlHBZ51mdaMVs1K3d4xz36BkzikOzEFsNgilPJ179/z16Th
wPS//fOMXJ44rmZD80YWHCEv2ZcAkEjBRNMSYU94t6pnL44JEXWT5nUQhhgOTXwgEas/SnguOtJE
QOwg5DmXB8bPf/x/GnxtxV6sq8wfcj6WLTScfrrP06FIeXjPcixZPkdLalFIfk6BMKPZ4pZJBbn1
1O6ODrvxgv9/jQ5pO7ttrieiJEPYoDUtrXTAEuG7tu28v940AhQrld/erNtnDc3JB8yRcRs6ZNeC
63qPO2QtsOD3EZWa8+BEdwok9tQVylxapzFnXomWrKxrryz8TOGMc5yAjZafd5m/coH/YWUpte/b
Z58AYtgP1ZxwWkLvRmlEVQU6ibxptiy2TWO+V/Rfjl1+UqX7kGiuRZiYzAXXWoKEyHdwEMwMvrA+
eZYmoqyFnlJvSsdnrf6X1PwuQV9q3YBnBDCw2LhAarNPdrX5dhvCbgScYdF8bffukWGjvqha8ZFj
YfUfGOsz5Hw6D44i+z1dV/Bsa7tR++0v1QFWkl8bGHnUR5UwV5JqjbHOwcsMJ7KGAwkR7DpVwfBc
AnbAgPHL3NUPtM2IISEjHaDjtS+neo7HvR3kdO5J7lUd9VWm6th+3TTecITb4g4V1MykpFpQ71uu
Yfz+lriPgnAkzqse/CEP2QVn7teRTGoBnM7w8n41B+nKEJBViUGrvqhW1TqLgfAe5FSQgccZWnz0
tHwUGiNjXTVCrqeyJSNX+r3Fa2sGp2j6I3dzMz75PnXMXoGeVfqzAPzVu30hFC+YhU8nf4xMiJt2
H/MlOH0dK+Ds4+GF/gmzAUs3RAsswQlGDPMGyU3gjDGcYWILera9ZrtlFxFFhUcv+ovondxTh9nc
6AXNkYip+nBXx/Oz5wQy9WmLeLmGOqdIc2wBSZpPUjvV1wQ726iHqvkk83VId9+NqN8ux/eBjm3W
WsVuU+ZoQMjqO741KQHThgGk7KIYDzykyzCbgvqoKk9G/aH2r9O36tJCSwHh8mw86yewLb6XBXs+
R8rJ3gZoz0pZG89pXgZIpbxtRhSZUTZtfKfqovHpgLVlbnAk0MrxgFmhavYLHmgSps1i4mBH9Fsr
8cxVeUkpQnAMzo7hXryjwXBVFIyjC3pZ6EKRpe9ZfclfwLSWr5FyhfSVZMgCdy2YS1ph52sJJdYb
I+SDhbVnlkXU9DDrJuKz+pWtGrTX7xuDS596Lyo0RNSKDkoVwlz3NUxGUn2t943KdmJuQIbEjyzP
UakVcLxasTC43ayexhflBzGiwYd9e7/vWXFMoyv0ZpRPBud2h+O4qTUKYVyN+kWIFO0Ql6Oc+NfA
OHuKXLwz9SRzPdSbTqbuHvEXjNtpr7ao8KXnAlPGvQQKEOAPmiGNxYopz6qlnXoGh9kgXrF5T6AY
j7Cb5jC1aSwF1XgPSrf7NsCPntuv6c5poNYZKE3Tw4btOGnRO09NZhpKnlpQDTbbRQkAf2mEl72/
xCuZQVyXnog7f9nNUNOG7ddRUbd7dLmza5lqI5DOBbyTIhcWUYIYA73obfksM4ouN69RN9M0ZBQb
k4I3bmHPe82WjzUXH0o3LNONHUY9q9DKE67gyZrHowiF92Yh2H3mqTVgItQxt2YwBb/mmEMLcwc/
d4omiXY1JpbRIKTLdWx5UBVg16lazQ06nDbPIS0BbIa7TDeGhHa7XiU2KpZ/IAwtm2DbFTCKO6kG
1xwDlCfJZoirP2tfG37sGBqWkuOuse7r1EI634coQBjs2lnZl1tgKNu5hsASl9kbmbh/ohpdUTHI
9P4ZNLplprmEy5vHDAhSxkazeuu/d1FZ4y2/UOdJTPNHVYmSqN5jSYEVH5v4BkTQY2rCRWJlK8KU
HO/VRjCPk4GjbeLwFG4YIKLTbUIJjR+nX5RgJ/4ltRGYWLoAGqug/BGbP3ZyQPy+Y6sHFcwnQI8h
2Bz4Lz+BjwaHR+nFiaWaIEJ1XJniBaOW1eaFS9cX8YG0vUy0MKHVYbv73f/n5SoxXq9gpGssuWPG
JrapBmC/U8O48QvbLMqGGQgcmyWn5H6vSW/5d4sy9Hzv3nxsSl5aoPmy3/xQ2C67woRkpR7JS0fP
2ny62wNzDGo6d3ObJ03EwuQMV31GMK8Gu9YgTQJBAaWic1pICVKprAm+ErJNwKNqIHgl4Ugcyqi1
978hkJRQlyUMKATTlam7XAgktWbD5VYB6NvSQU2xsNlOpNMf1JaQ9h8EzcyT8n0byzGmKIeqTNX/
PCxLSZWfFd5+azhEDC1UhSbPJwM8qerKPNbFuIADSLnOY7Iajq9dMPS89/mIjiB+BuS00wfR9+ky
4c+KsSqjyIkk2gkCnwuvHPVuYRPA5sOJ78kE5YCyUsXcMvDijIbEP+o+jkHeTsaq+0E9olxCKLRO
W3W0mWp1nmCb+FKlX8gdiKWVM2Nz+E+eOp4LJHo1ueRNbS8crdbfH/S+jcd6NXEMspjnsQV4BGDJ
/4hbCedjLl0AtW33luCru4ZGz/LhIM6JhuNebuOJEVPlm9tmm1BrQh7SK1YJ/Ke5TXSuYJpvejFS
g2nUth+I1h6UmCd40ie0wEOPoxoeODyfXPu1xbDhbHZsV4Fgy+bX+vKmHq6qMz8lQs/Kq/ArHIFG
NQKLLdkgc5nAy1c5vyQ7YqfQ18rbNkXaC58V8LDoH/FSMwgHjwzWhY1Rs+F/GQrwqaXrpYe/L+LD
fmECmEH2RV5lsS2F2ZLIZZcqnna3CRkXTlSet4f14J6VpP/ad3BTiZWzvur+Al36mvrljJTVtGFD
YLRi6dZ1+6HuDxsuGOvc2ykhb19x8oGvxBwxvqhveADmpwMAo9apJUJYBKcE7ViZOQol+9OSb1dr
PXbhk5yBUoWP3qJ4+8INN6x2Rjx8LRZ0/gVBGp94kUjGXYJ6KdRAxj6TvSm4FnwCfzM42Bh/4DL1
aCOSXIW9CebGwhWZTSEnv+9GmMxPS4rZ8Qp2W9wZRg6ge3JS0E7UttMZk5FaRsTti0L5mwjFxGFn
YuGTNDdHRh8I0Vn0z+N4wY1cYfTQNBFo/NDTrLsmdxe7Jk0eTDB+1GCWBSfNM9LPaG3QtrYnV4Pg
4fsIAfHAZa1nZoxWQd/1tcAUrLDbIzgIQYf1Pce8tfS1mkAQvuRjkrKQbfAXhpZezdNEuILvoiu/
H+16F2j/kSvSiilRZ7DQvuOlOoK49016mJAq8a2qxX/9NPLPj27x5EGYfESUIK45YuL0rD9nNic1
ogYYoBfYYwSqSn2BzILiKoHbWxRZHugdYfApCyCIRpjyfDYKp5/02sDuWTw9TsszmI3mGZHSwXMM
Jp9WgJ3AqLVPj4mgred8iPY/aAcYemZvjHkNTqlsICQntC6VmfvgiOyWu28ewasvMBbH5tdOA0nO
tL7KIOY6xGGlJLi15z5Wrg2XJ4f9E2ZfQuavlmVoc+MAyT+42BR1n3ea+CL2M3pMajw7XtFpsodS
mnfbUmk/7e/sW7BFwky0+WTBk/x8TQU9XMOUPpTbbtTI6HrR6qkLBJcBxBTqdGsV0B1ROiG6Nk7/
59LqDOcv1fSGN8u4h506z8k9o4iEga8qa3t/WbUsSH8+4MJqhCJ8hfds+LPIosiuxMc8mrpLyv1X
GTDun6asQ3DOa0rDy+REGgneCd1vFS3Nlx06XtNltb6eAklqigrpQvI1v35mnWsmlLHulBhJU35V
KhmudHfZehgzH0JdH3IGup9J9F4sY+sy76+sJWoU7y1BX3oJQ1OJsA7ETCpt95lR97CpHTMtgIvD
Y7vbaGl1uTuXTLq01OY9eFcKcyqeDbShFkugq1uhRqj3OonbA2V4EZ7G0jvPfeioMuyNfpUCxaok
4qCGskHKqxTyAdg3AnSh4x6kXTKOm8Ek305EyHA5+c71CMQ2fPYDQNH1KHqgIHq06OOYCEnRxC0Z
duTfTa7X4r0B7ujYe7rPVMLSD05gg9Pi6NbgLVkRLdk5SSoptHCZN31EJMZJhIVVwnA/eCryFFAe
DGHqVLjFTJagoLPTC5Vl9An/KpeKyRBL+/atSFJgWW4kH8BlgK73Cd604bossdwTPfgnmN16GT5g
UkXieovJScdpMSnTVwZtmJVaK3uW9vj+7QNIj7oKp67+gsTbVx52cwXoH6inZFcUxh8Nn30b0bkZ
jx3gTV/rc38w4N0zkU9vKSYeDvsPtfkCVorRvMzV3IDSPiXcPI6jNp5qlo8QYfrt12VC1XcYGQru
wT9WgnL85deB6vSowuSi1SaLoe6LgdB5bgqzkGvpIeQ5gTBicYSl9ndkwIwjclgRRXTn49MZhOP/
wgIJ9QqF3GoY9z6tArLoVVQ3e5ILZR0uZxdomPV6HdNedG+t/nvTzuzT/o5S0srZ6Tb/s/GgQNpI
pCs8aCOiIU6mOrZeBA03XIBS3qc2GnJBHEPHY0Ynv3Sd8GwdmhKQKC0Ic5AhJlHK87ruxtoy35z9
W3Fl0Kt1d0uvuqXiD/9ffwZH9EjcVCceGdVW3KUt1H41j9gpsj+uA+YJIDQuKBrPrLyB04EBm1WP
PhLSal2J/FmowEMyVuiumDLqDg7vTQpJHccRCqLP8z4GN528iva1RwVccsqjyLvSTN7Y0YXlpFbC
YkXvwvXp0MxrxsJ6uq/0AEV3bEmPS9IYZnWkeVrfZ52m6fA1Ojl+0byvDBCVtC0tazeizBUCbOU0
pBl0KgGPTw+P/wBWeXMVVEo+Wr+7koJUewc6xAkehdLmJeoe52auPRHQ1yMumIKv1kD314Ndn9Tp
yhxVzzHRY2bNCIjRUcOX4ZtlrZRre6LsmsDMJXpzNzMLVZ+fKPPnPc1gTOZEYOIHwSD1ckZKCaUS
mxjGr9k+2lBthhzyRlfG55QmB+rQ22l36v8am9qNeIeD1Hubk3IWV/LMeY22U0Ivu+ANH3N51NSL
TrotG1q3lEBfJVykjY04P5lvtTiIZXfpgjjlksILKgrXbyDXZpRf/4HDFjpfKLP0ubBNhamtHHmz
5X5QUaEcyYEpDtbDOxeW9VSQ5EATmLlVc1b2FKIt+Y6Pk1EMC7ExA1eMZFJALb3Y5TaksN8D8RJv
cVpE/Mbcf7K9BYek0s2kXkped35OClHF2wsQjWYgqYoAHXvrNCZO47nZW/vGKRsiBPQEa2ukX/hS
xYu5TYKNZrwUdieR9/p1o78o5+UGVNN2IRiS+XIHrcvqSv8iSXjrx2lVoXzgPspk6LRnK782y96w
jBl7RKMTBBLCHuZRxOnJHie/lKlsMQ37dwq1UQJ1lA1xK1HMyPp5KNwVHMC5QMJAzHL2c5jLyjhe
vZloJL40HRtO/wAL5o2tU6OP2Ej5v2Y47T35mnynkwyl+irOWYkbRKXi/4GAKvGchSL6g4ZUDlCY
ZXLkmi/dZy4n/D5GRbvha7RBI/bFaqTxoUtsxLr1RmNWb6QQJL9fQvaC/WgY1uTE1Yus3YWFKU1r
3wfMpGMSup6B9At1y6KjwR1NIkHg+ncxYVcq1ZjMYRA1ykCVCG59nL7GjURHXvk45b8w0C4i7+Fk
wZsR6m4xryS1SwsZDSyfXZYdpmBGz705eODZ6/xU2GOv1pwa0V8KLELhCaPyKJ14jOblsdaXJYa5
MRi6zHrd+HhqN38DNudm/sRCDfDgqw7wkIcoJj30vcrS48fSIH8qSgwQEqYZCGCDhccly8vnUe0o
j3REWbf8h/yXOdT5pSlXe/VfDYKLLctb9SFRpDpnMX5g/MRys+/i7aSl2BEX46aYAwyfrxlsAGdJ
6DuHt7AiN1lRmHedw9RgG6sT8caxpN5qBPohs7JDLpMeQ32h/6hObyMune2MtMkANQJoXyENog3J
nIyRRQgk6Udve0kAaGZ3egiOAsnhy7fGMcTr9KUBFDDojjYZ1belqrAiOLeJrPH7JBgbKso7YHNH
CFPQYWMxE8Ia86uLsaFNGCgK7Dzh8iqqMttu6YrhZoAPui9IEK0SlaHpg8ZXzHkkV0/4/WvAW1FE
vUhFIGZ+SHKnfUzkbL6z5pVzxyICHC4r7gWDkZo64EEyu0rJTFmotrjlaHiVHnfaQjGziAOcHZkh
Kk4sCtY1NvNTw2HggHaoyyO8ZHvGHWgVMQuNwToXa5iW/K5z8DNPkOmead6/V2uM9BuBECME/vTY
6VPl78iCn5pGtBMvx2J4Vn8FkUb5CpqHXELZu/ZlWEuIeCgIDC58PBxQnQoUjLn3MULpvWK7zH4A
qTx99uik/IQ/HNORUPJf/D9IklYxOLhyZLD0jY0oAamAN1/TP2mHpbXkemPjN7GDjYvdZVkXiVaI
wrdndemnOVH3pdAOeN99hyWRaZAMcL1+y9NeDYxo00OiNcDHYrch71wRa+r/ssEzm7tf/yG3d5oH
mGDi3vtu+OcanxH54TYVDileTUMX0+bc1UDbdeEZtsb+JLX1Th7bJcXHl61dEYDmUuXyGhg/6Nb5
QOESHJNIryXY2dF9pZC8AMxRkbMHc3NHgdsQjqW+GZ665Pv6wPi5MD5ludwKz6TRQLtdCOpX9biY
IdJ/AvIHA3HOtHy3tfnvDUx+DUVy8pxdSLXZdH/jAuK0Dzw9qQvZ1cgNrwFEKhuM3GnndySJbnJV
Nh5JrtMzlQmodrg5tlZeK0MZoIuORm3dMidXLjg8HPlmOmIcUEr2MF4U92OgbnrheoaHd5TXzy2h
Y416lG37S/0snO/WNVDYyxLIXmHbXLRAxPtN5vykor/kgxUYhfwUVB0wEqSBC5T9QoasvBvTuUmC
kixPNqHv2YrX114lHsYeNcYVBa78+kbwFy2s9gtZOcob+WdjfZQsd+P4UGxKvduHVT+zKh/KYQja
mWvRhpH7N2Bd8ntqd4pzZA16T/S9WH96EtAvb3c9ziRNhULFsJ9P9z27a5EJcl/dr8d//E01uCmi
UIVNLCq04S6Zq/TogtQGJ4JUFgy+xPsCgCfaF9tqNgKawZ6n0aZilcxksj+xugZUCkXqJFFWrylI
4zwvhC0RR750bCXs0NfFufrXBsCEzEeSz7CyZAEEt3T8SgAkzX4Os+ygu7sjH9ZjOEvfd6Dwc3tP
9Ii4JuqBM9cNUA8YOMySZJqWngYFGxu3+Zq+40tTV316DPfdsccl+bb9u57pxTvxEaP6/YHMz9SQ
Tn3RQuR0ej/CtykUbXVtEm+tflrO0wS+nWRuyN7p2wwDc2YAne1Y9T2QGyCzaDLLpkeMSJfwrsrK
Jp68sXJAMBBt4+jsQWhUlV1W07rSeh+JdrU3B/mKiGL83tQzaVd+kyjl2CRzCTaQpbpUJ3c/X9hZ
e/21pgbyu5sEIYpP2wk3Bhu00ekx34Vi8Hs+kL3VuCT11UTI3FQxPS5F+LecgsgI18VkMMtwKnSv
4l7SDHBLko0Q7+NdAeBhFA1pORFaZwBaUBT4rGyS5UaggalTDW6c55Y6iAyM+xBIPDWQaqfnsOKb
v4I1b2eZ0jyV8JejT1VIJ7uteOdS/lli7gOk8CNzsCZMv1iC5+9h7hCmfewykCynhMA4+ZfwR9wy
NhKa3qY+FYi07rpJt+oxgqPq7eadtWLu6rx356zVl1kWFwHy9xr66Sc3BS7bxuOKCD/P+ytAZNKu
RrrQOvTqFfYwL2lP6WQkfFMkplEI0PL5KHI7bZgjP7FW3x38Y0b3PrpY6TpUn+zuNQb+kHrDrR9E
r6hSWzlAJnzhyDw1KTsPsUPsEKVMf1lF5E7INQ5gAiquh+FGqSpa/f7Nhq+i13yuAFlmlpFePUf8
iUonHTxANbuRhOJRaPP0CQB8t90EjvLBBHbYWBuryWA0hav/dgbapYzl2wDiQRWuiCtrb/rXoXbw
DbVccCAlDJ7iHJ4tlgloAHLn3AdgAwwAFfgVzpPc8DKwdD/aKQ1lyfb1KhZHULsSI5mAPSls0ASe
ekJ+VKQ49rc6o0WgSfvwzndusZR5Q7Aeu8NQQhnWPtTGJ+GfR7rEApYLxznc44w5jEkDiTjw1ttG
bO/Gjl+TOXoqryfzrXU0AGTQi+DYUMJZYUET5AUXXms2thE9cm/Mmx8z0eZe2OkS82sr/6aO56do
5hon8Nl+XCAk5hJMoyzb1Xng24ZdxCsmUXHf6iF0UgDMz2jNJaGMAhBW2wwCylE/wjHxz1Wgs74d
AAU+PsbJ5dW6rGDMr8dIl+hL0qh+74Q3r46bU47yZucZYdM1pdlcX7P+oHqWxCW/7yUkfubUeF3e
KWXnL5GaM4zE3ZHrpiWCqkb/m+5pB5jvwD196qE0XbXegI8k1UlF/jraxhayeIH0wMgBw+i4SQZJ
HG1C9KdjApPnzt0ZaVL46ABYirSd8+g0pKju9Vl0tdoSaCroxOQb8qzSR85aT0LXW9tdpEWreV2j
+3Vfca1aFaM4t6V6/vkT5mo3KTCDGkS1UFEu5GSCopuABwrxIIO0TFIK4/JXZGx5DyYJd7VLiBYU
lWNizF9eVl2go93qZJ/5cz06/LexX6JP27OwA461dFPCsdAHpmJmcRrWPSl+LkA9KXXRNTdnU5f7
gCR3EK3NzoqMX1bqVJx/JMso8bE2kyLXlACUOJ+Bl/HlGoK0m5wjSGbMIdQyQwFwzEjYJG7R87Fx
p1swzuQr5O786mhv03FMMKIcWyiJjoFiVgTUjeL/p2cQmki/gWZWAocWD437QOECBEgZqdP4m10N
MXpgp6pey89fB2MabXMmN4m56JKOeZguXfQtg8TxapI4wUiOko9zPcmqscwNJX+UH+GbOCfQvSXM
jI+Ox+ahsiwFL0qp46BIimPvP8F2qganNL17agit7bRPQzEg9YlzQQxx1b3xwysr/Q38sYR+RPZE
XkUvQKW1va7e4d6cG1IUTMNS8ZghyT1O+ZdGfXOC3gmA2UJHmFFDlXtpbhWrcCS1RTzA0L7dqeRV
J+aXGH3/T9cZyP+Txybht0RZPcFQggt52Z/TRkrtgv/GN/52XZMRskvdNeOGSd2LELSS65Wb1+Ed
Nk1yhJzriZJFyjR65N+hUYmIxNrdFJQINOHXtry/51cO+YWpQe2Lf6Rt35TRWm+4YqGeRFFqJ3IS
6tt+9vEBPAyLc2SKC4SuT+rwz3C8/9SlKRAq0pCxO6C4oq0xdxbOPcmVm8ZYe180C+BIA4E8wcOg
BYK/lBMXhXG+nCuKtoKn3w0tkOt41qYQoW9P82sjV1T/Vcsm8eoaDQeFwv1HkyX/rB342qi+toJd
j9LpzWkrpJPCfvc8kZulu0v6Nf1asP6yx8gicyc2f6n4RJaVWlWZixKGfxMHbDF8BX6M0YGlqJq6
5FR2Qm0PGbOoKIDhYpCX36+nIs3h8X/twnBD/WuReHcdJmDVU8WnBos6SByZPkCbIQ5t2u1Xf3xe
kyl8E5vpd4Cwg3i6qvWJ35vBFoC/+F5ON0RfAkrssrrhOzge9nMSGOVpnAMOQwTeSUjwmSjPU0Eq
izsgCQOu5vVo6GGO7BKso194t8hxNY1ImXMAyra5yV0voihtq+w3q6Rc8ZBsd9dF/E9I8YyloYTm
yGitzLdTUxuCr7uXa/3iEj2h2R96CQyCguHl3hksAa2y84NJgaCCi4RCJGkLMQ9lLGKvXMZYVvx0
hiTKiKQAGutbhCRvgQlgVXnz9t9RkjxxUzDKZsUdv+4vowLVYHSt4QJZ2ID14bNFc8OMWKeLHMgw
VpBGI1iBZtD0aORmJt8q8VTcFRcBjhb1ZSdabw8V350K67X1nVwgvV8yUyVv9tzGT5FcDLkKxueq
z/BYmFwBINsGupZWJLR463OiBeiSCOMqOI4zqH0stERL8iFCDCEPOEFcUTJrHVsUBlcJc2khWQMi
IihjC3lI6GQamM2DVg1S+4kcgYrtD2oVF2T/yZkWGuJbDb7dXojpitTF00pzN4c6DEHdf4Tknko4
RdaOWMIuLynUREoEUYQAZgFvlqJ+iR7HjS8U1sBpKa65YCxz3RjbNoA4Wc7IRpkMvks2zyjra3sZ
QpG4G4IeM7YtHJy8VA0ascHq9jr1fRdQSZ41I4F+3mdxT1JU2h05tqi2hR9YmjiGsP90KKLJSQtf
L3gibH7tZrkTsOmDIvsGi5mJv1C3AYlUswiz3AJBvR5WOvrQ4BS1Cw5tIhMKgL7J6eFfJEOR/1qB
3URPJYW+L0h3VNB8a4YScU4TXr84FL+vWEQNXcpHFSo0dW1wo0m7o9V6jZX1Bwo/GrfUf/7h2+j/
LhQnTJB9qpUHWvAJYcSVWSiYzaGlTWwXACQkmCn9p0dPBRlt3t7zDEteXABhaZ1qf9xEDj9QQPz0
tcYq73IU0vLBlLqJZjKP66541MaNsFQ+x7zUKGhnH6fImRdBcbjeq5Ir2J6RvEAvS6XeTYpf5CGP
F+2oqzajs4qBszE7FBhhL3z4MiegDprjOC9fli7rnC+rOQ6zNFcWRL5GuFKFvyT1H2Oo88dGhfW8
PEsqfMO1e/XHQD4Gy2jxfsGDrbN0dT4zIS6KBGl48R+kFNSqPN80ePKBj7uBNC6UD5bEOoOWA7ia
02EJ4Vm3xHnqqOmgi3v2e7pIUzdF1MvtQdq7SqjLrDtwiHsUhyrOUS28LmrygELq6Pj85+ZtXGxm
wyR/7CZrV1hjFbdkQCnI+TK/T41wfRGL60BFgdQvlCKeFaq6nfvpKaK4ICE6PZd+T7aYN1YfZmUD
F4nrScwyA4Lcd/NDLohmaD4aoqHHHfvF/KgTVsEPiopvF5eAH9n0hhFu9iKsBiUv/zwBnRTwEscg
+SWIIxBdqo/xx0mnkbU+DNOdDEiuBeQtAosX6uZ3wM64s+JoyyrP+ADOG1o6EgIxIISVjyzG25W/
RrA5nfGKaK9UbyKs72K9xuW4gYJN8nN+yMBCjSc+feJ32CEIJ2cwjXzGTSIxYdfqECsEVfVSBIFA
4TvQqY2Crv0TnTtQ70ddAjXVL5LEpiGEMXJkiihPqh0G232YTdBc4se9/ZlVWqt9wpf7/SjsObD1
SAaTBdnDQbu2MNZveSeUOCrcms5M+oytKuIh8rEkHnJsJbTNn6KN8fWGKnHAwbVQK7a0CWK+Smjl
AGw1kq61Ly7/oYmDq0FiKNz94SavMiDtBMmf0gNH7pYWrf+gF/fg86YKKSHQ8L0ukwda+2eVmUc4
8kmOQnO04gduvTfDXTJAWdJE//XnoQMRlz1vWUgjVLK23juOnbJ02NrUXu5U3kJNGHWjOyom6Bhy
CS31KvBbMQgNDfp8BXlomOlE/b6/BbgkMEpUxYTNRGPm0CyxKA/n4byZUJIv+M7WI/ER5LLrC6RP
H+cLNB6JYX25oIuNL0193q+5PAyef45vSCnhVlzfczw4ueD1/bLWIBlxpIvdsv3o4goDsgBHg52J
IQctTw9e4BmKbcEL6u3SskRYEXytGMifukrI8/bY8eJiZggUoMamiAMHp3nG0kMoHVUIX1jYv9WZ
0WOSJ1hzma0YtSl5n0hx5fqJ+Ik+SJOjj7duUp1FkpIWVY7dMwO6qfhxPKdRWBAVNxx5bCHvIYOL
ahDgeOXRJw6w353CsmehRq1CJmTMIunxyFJcRZ7hNHaZKNbJmdR9XuNv5Pi5xK6Uc7YR4xIdB82J
QAA2rVAjKECfftWL5i7CX3WDKnJT60BSmUIp5vVKYpqa0O5np1JO7zMlwviJx6Ldc2DMY4OL4eUe
64K09NDqJ5VnjLGHHilnCdAtOtLftiiCJX8SN83HTjl7wk08wZIH6MTv8eqmOOkTYMcwtPHOQHHD
K72cfIk4gFCBN/hIm2uZalXkbcjolvJrzE7gxygT2wMLnoQd1KRW2EwpmnL3X5Fva7n3yIItVRnp
tLQF2r4os0VmlMJCdDgBICg0DDFvkRg7wmzKbB2IaAFSN/t8ySfoOfjqynWuN15JU5tphFSt3RoR
03igl5XQ5hJZP1Y1A0ruMqGkUOB3qBN3jc61s4e4aTJsUy7tv459PXJfxjRove56xqpE9nM6EhVW
R4Tw0Zznn7aO0xwWwA+V22Whwc7QV/bDmjQfvDkxFJvhPQP8ZoJL6RlaRHlsr8NZ2EKgykUGONgM
4XKhH2J4OaRgLLGaEAYIJWUivropK/YuBHoz7d4iA9O4ktJo3HIltdhJBZb1slCG3TPxlfJvcaIi
eNVH4JNafPl95hsmHPnmk+v9VrqJkW0V7vWBGoTLutP/oeZwB1T47rhHfQajKiYvLsP8tTMO8Ga/
Yu6xgbD2Fbl/6J12MPVB8z/CuYiBwWLnPqkclsJb3ylZ40dRolIal8gcUYMIEFOmoF3bW9SMTUru
Tro9H5oDHHOQ2DXd0Ek3K6iqSPt+S9ouDou+Ce64hrw7b4fyweIGvWI+z7XzVhSbDCySW7Jdvem7
CsdQ7ttX2BDJzGCu5qdfUyVHpqP3WWaOoTZz4YPt+Uupu3Z3pEuPDfEJfjCTepelC8+eY4BVjnyz
ZAbEZ5+JIS6C7odwVTDWob06LBKsA+8+J07PznsbjIWclAqY41aarYEjgzDRTX3Ou5hTDxQ/ay9C
rcKXX657lFIW7HO6WBJ3MfSl6srHE8byyfxcwPJTgW8i0DRq54gQCn44Yv0uWlPHlBQ5Mfr4mMMP
FQkuDs7hFUZ+YcwBaOPn2suQ+wMuOKOBWpSq64wUay7xLHpe0e4b0k49bKYxoyU8rXX0vQOD/BeK
dF1ENmrEkZtLlrxQrpklNC2d5sCtfe8YeZHTo4/XXl2WNQ6bqZY/Zrmub0uX1viZMoPlrczvF4R+
wRb/xFQsrAi9+XAKNkhyDpvH9Y+Q5OpZPYiXVi0c1Qfg0hGKCj2B+XWWyaPNXCWmHWGlcK0V8SW3
FATtv2z398rYJWoJdpOT7ciH50Njh/TgHU9prBuIlTfM/xOG3t7SfL1G4xlsjh9Ky7tm/EjWzt0s
bouPiAgMIPeBiz9evhDwGuch9Kk20UCTY3d4mrLdl9No7Xl+uDKph0p8sESGbacO+pGpQ8HPZbYO
8RCy3EjhiBurIj3VvxCAth7mDBTnrsE+OR6GJgKl8yesQgF6pr76w6AP7jXitIViXnf7FqyQ5fbC
536U6GlnwrjTQQfN9osvw8Z+oS8bFR8mFEtmL7jKdMG71bVQJXo6xRCj+y6nd7P0R28XJZH2Dh1U
Jhy6XispX16mzAmrA9ZC/V/umP3tcOm29OdKWKQoR1Bkyn/zu/RhvceWa/XigkLZVGIHouqSEcSv
U97Ghr7DQtwX9CUkgo+jpe2N6mBXoV9TKY8RNRuxu+g0MqPn89uYK7BeVF6LzWGaC4ZAGdn2QlN8
rSmd2d1H/HTiTSk4sNYuCSHKnbNDqnr9bCSNnsAf9IHHBjw4vqCKxNgXLi7fxC3hHPOH4YrJ4sKg
uKFHAdJbi6MQOUaW1ig/E+U3q0rO/53pce8QT8neuH5JIDMAftlZLl5HM43wZDLC78RSkR9i4s+T
eqMhEqD0up3zeRcU0Mm++JKOZAT31wLFTP0t2/XgvwUy8tfU7jEgEx7gmThiyK1UBtJo67Wi/6Qo
nFMbMxOEinBUM2E9ztGQEAPHaw9XnzlD4fWJrDTkZYbb4aDXYQvWfOcA+rA1ZWrP3Q/Pl8cCCJK0
QhLS8shdwpeOhkaYBzcMdR+kE7u1uNf9Lf/8Zbw6f1yCAjfh+GUOwhzZFWurPttMd9TKEi0v8iTW
nwTshE2t4bGQ92/9VlSOnWl3qII7gJ/cKfYuoZDVukFDnU49pBgXodsNOIowbLYWQoImDrPP4A1S
s/omZu0abdCkmT+8EQ15sDJJqfkU+w0t8zJxMSc48uDYUQxx4q5I9YFLIEN6Wbkz9sh++en7Tgs7
Ab/JaVoXtfk9JWdixAhrvT6P/8hmqYyywQEeVv5DBInXVxeTcJMu5neQHnZpKeyl/mPL5TumF+BV
+ym3YwzRrJzWz0d2wPOwgL7YA9dgwOqXf8MhRmg3a6BTSBKkfdiE4piKOOluimKACGCPW9dfy38/
YrszqakKdt0erlBP+Ez7U76YJDXOhqxLQk4ZUh3XPLEHYCfOqpKXn4zTLyjZyZd0790pJVfz9PIl
kfZFZeEKeFt0Fczs/GWm2OtnV/idTjYcpRK/2ITfo+6qHffbYIX9aSFOLj7UyDt28nuND5p1qto+
R+vhtYzb309kpwjwLNusfiesir/kqJq/OvuYFLLeVr5ucd2C0NFTxcIEL5AoBZ4Jj3Qw2BQpXoTC
HBaaBhMRMvt+zcbaSI+R07wgoIDsI1m7sKmFCBoVGuXpezL+FY0vujcOmWlbuHw7r9RBK9x0UlYb
IlXgBDAm39pK13FtIP50cWSZpfgABI6472OQZ/3kXwtuMIb3W0mcwf+XU2qLzEiPnmN6bUn6G38i
VUYVrUhOOE3ylaheGDfctjhCJ4w6rA2tG6tJ023y3tnMQmUse2mdJmirtnflcfR7Rt5LITtGRJ/F
cFqLCAVnzAnr7V7UrRjZPvK6Sikuij8xxRGGgDZjZT70NsB0oVlmgBtV6S2WsqLrnGLsnxzUT38J
7bDIDPqARyPLftYEUUFqrNDhEGe4hwX1QHDL4V41SV+QNiDXC+nsd9lFX+GSib0LX4AbuDc4tpL1
9TyaOhQis4/o4uPWIXNWdTis2+F1p++xHBm4YfYgr0qRImzZ7DdgFrr51babVfLfKT7YhDsPDQrK
TKaWy/mb0UGHMwfi0XfdZA6l1M3BmaGiCTT9S8dAPONbfBSDYqTbaTgfxLbSYc/3i0cnx9ShIKlH
ebPOurpgLRREVEt97Mbl2tnI2ZkRSoe+K1MaiFdIHZ7lplxzeT69hA9h01RRJVA0wppKQJfGS9mo
ReQCl+yX+t5swzt9CeufwFJDB4zChAmr41QXvrZ3aOAK3gJNMKgMzvDEK38UboUkGB9fXG4VMN+W
3YSj4lhwn6XzGwEaslTPyQq78C11jD6hbBBE6zNUBOJt8Xkv4376IZMWPKecDNKkLBCspktg7Br6
pkLfmJYoBojppMRRdqxG9vsiWUYozjYfpNsU+ZaAiOYNZuE9C2fzxM4qVqT1HKSvREgQXeTLXO0g
DFUCBAR0cvsGmEjfZD2ZdTc/Nd61L50fWOoqjXP7SOB4a0NR42fBwLpB7n3hq4ko/WFaGScDaaIo
LD5LjYMAghY9famf6aJMv28OQnN3Avvc02su0t0AoOB2Iu0DPA8oRYJIE17F4GGP4dz/M0KNINTB
f4I4x2ztj+6G5QAYW7RaAK0+BUaM+96w1q1x4Ph1wujQ+ILIm7CmSE9rE+fiUIbKsxk6cVpRHCyr
oAhHBn1V3nA3wDDjHJd8eTMQwHiUxDRQSXIDwJcym4f8Om6i799mueA4+xx68CxiVxGt+kwlpRXu
pYZ0sYLJwQ6aO5KxemhImV4OzlhGblfwQYeWVJWlXmLmIXxc/HipwqqCulXazJKr8HLGYjiaBpuc
xRvpia2Gsg4Ak0WyIiJ8IL3smLwVjtbutwLuZwt//ranV9llV+89jze3FURE06jeOzAlbrUaaj/Z
V5MFFJrRfTcxXPkHgxlGWqFGPxoLcSM2KitTscOziWCpKCyIbaFA8Ulvzhuhv2Q4xZ1eCHNlr8tC
VIrffRFKlQa/UfCk/O3rBAp/15NNJQSXJWLvoZ3ooFpJ97np4pB3kL6pl2cGSGdKYdyJy3XqdVGi
vdC7CnVVT1GaMv8qmTKXsgh+byHreMzEATGvZ/RD9nkZmprH0gjBBpwJwxZL6JWXrM+WytxiG3Gl
X9ymiM3LlomsN7nHezfa7UjYQQ8rqIhhDjTiC5XGOZmfoduiAZXgbP3duiPHGO13oSCQnKj/ZPuE
8CtGZVilkHBP1l4p4H/mCs7dxdY1cnuLigfyYP50UnbmemYfMUEDILBIAHt7/l9ov84qxGrb+r9w
t0C1jZcuPrwBOFvLzvtr1GYnUOKgWVmLCX6aEYSR/yVyeQVl+3DLgG6+3/2ztavZeV2ru+1osWEe
27JXHoOs/tnkBlGVqITuHwu05vvNd0X67njWpIc5otPZwVR3Giz5qZjBL2Q4jh6dmV+uElnlFSzQ
o1VZmAC/go0hXsOLu1TBQba1tvUv2DDT5erG2GRCAIVzf/SJ5bKEKMOO/t/x0byYf0ptsOzF65NU
37Wb0nU0614pZZx5y8rBWob1/Zpd0TxbEtf8bBhuFL4YW6aGN4zZ4N9f4khuCvnr+Qy2THqoevuW
SVH/nj5oeMC9B+Sqha58guV6a9+e5QMd4sxfQroLJAAYdaTkJeHy4N89f3J8lIpB+X8iZfiPG1wM
qBd0AteiR/2G3epX2xX1O17dwmOylMBx2oBpv+Sfcq1qBdKhGu9K2gHPsGRZGyo6+8GpEaRNOfOb
bJoniwOHPJIiN3S7YmgyqD7NRdnOOBuc6gx0D5PF7gDgIwwy0Ine2nVK8sgwFXkOchGlQviJcyd6
HKY2TOS/c0qJ0kIaLSX/zcNHhtlVZTurowtBnM1Mlatg34r07VHrvoBhzRpEpaC/a6GRJIcMip+e
IOepUnLN872wqFZtd+4QAmjmUXAUBvrmX8vKjnJNTolL+LINTLy7zTxSqX4E/sA1FLghPZjLJgRi
z3/eSOUniKoCuh2/9TyPUCgnOwcK1pQfcttekdAn7Tz0VBvYQgyKNwnfRcBEmWSxlWov7KdfJGAZ
9+yE6ljJN/kfmXX1fKQbv8qlh23kO0llIJC/hitGb+T56jJppPbz4SlqfLJhIF5V804TXJ4kedS3
XKxum/HzHBZfLoCze0dbxl0yeoWG1mVFnirTNeLvmkxZaGcXKYNf/0wn34nXNFsdzangLJss0PEV
g7M38pk2SunVSZlOGbJZlVbQy/M3knpOt33eE2c9oy0TnjU9zauXcW/A6YXSJNo3jZJ/dMTutik9
6oUP/DwxuHu/DXLp5cAyycJZu0WyTP73XvhJ6Drfn+Gbhq/knLHf6DcUarTpqVm93Bnm2WwhkqvN
UGNWQWipwtT0J/MjvRerWH3ENb+QwVfQjGETfzbuW1aEAN62L272gDxuq6xJqTusUpUNq1mQqdfl
VICZdrecQyLkh34Icl2ybWfBGvPx08Pydv680oy3dkyctmtImq3JoEogF0GR0kUqjykDW7FKyFKU
Y+stvwT8EtwKpilJlQf5iunkXCZOjDkrT4GKJ5EzAAaa9SOwFwheMwAAFXSvnRhQjQycAHTu9XT6
ETu50nkvMupg40PIu77CLfuvx1cwfiaInOKyjDS4UX1q8riLfcLSWT65LPjpw6VkZSKef/eJFJJH
fzpdxVp75KIq0WBhbsPBXWoeGHcQ65xzUm8g5rfcwzzVyp6/nfIeZ/VKDhrdIgTacNMmTTnXpdV9
aaRZk6F4xbq0JMvLlAgx4UzBGOhVvp3+oev4rC9r34OHNrckD8pJf0T9l/UZvyrBrV9wUyiEEFg6
WpoA3uUo5rIpFb3Snxlg+QOUDKWXGquB2bmszacsj7FzkSwrqpgUDENgnXwaEsYJE+NIufvMkxyv
wCSOyf1esepUXQPbJYOQ3sZg8dnyqVbr5/9aJ3p7UD1U6B7iEm6oJw1C7R7kd1krM+39jILOw0C6
hGqPUn8HxldfeXazOtDbjeZG5hWQeyUE6WoMJr1RfddEP7HGKP7qaUfRWzJTMSAQfAln+DlFXZgE
3PPBfBKWPP547O1QKkdDRZlAuJN9kCnIWZW4edu/smEwt0UoItWZrmK2zQ0Kba+mYdD7VCrnCOMY
zGD8ePl/6K0YQXQFhxpHYxWqZCM71USr30qI89EYpxLiCIIVoIvaaAwKvD+FZmLDhqydRfD9bEwT
zE8bmbYBCs/14b7FJNQ2SWBO8ds3NVodjniPMZVpvAQsZyU9fx7ckNaoeKQPEZQxs/U4sWYE2/zb
dVJu028zs0qf6fcFVK9U6vMvutFd25nRS7hIwbBXRY4DSjoM5xWxEPdkTO7w2/eQCQv+baSl+PEo
UOmzdgmuXcZaOftObz7OmJQ40AOKG0VDonl50iaPzmn5W204UQTmMHjN5Hnw87SVKfCBtWcoR3dx
Zv86okc1+zrZclRYDsrS/1ltM8Hphh4heJbjc8bn8/0kzsLKlufGPLnPLF6t0hIBp0qEQDJraVKL
PkmphJmaynDWDaZ10rGc5hNq+pF4pl5zVILp8/f3ZFNErHSRFInyZ8vwq6hz/Kk42BjbKarA5nMV
WdLVwSYJOIdGphtkiuaYQv/gcKk7xULFJf6ybMA2tZuMNpHyWGwQQnDGeRyAS3RBHvjEVHro/Bi7
sMcaeUdTjRqamzBqMnWeNb83dQPWf5IaxHXWP5AzilewtAgGf1KdKvrR4NU4ETqR/WjB0abwTYle
GewZFIK/JV2/7l+instRzcINZS/6imFQvzdgR0KTR8XHGKuL3hNYrRTZuTZad4NkT+wrkjMr+zRs
y/UmLngCIZxcrze+5NcQIGU+KjgsX1aorE1iAoqz4xlSbP4IBH9zFQq7J/OzS6N24p2zsNcafPjS
OMoGWEIR6AAc/UKZwOIdZfBWoEXnzDIE2UcnvfPceD4CKe4OQT9QTvycS428yzYfr770wzlIt8Y3
hr1Qz/ahzmhKUsjYreDlRJXKPHMu3bHWocIIG7oJvFxwSsm/g9Sz+XW4/ZFrbQ2NptgJF842QU3I
y9YZuigsHq7PauY0PuFkiZPUiFtUM6RNIj+PLjLbWfkYg+hGfiN0iPFmYybJuUR3JODWsqflv9xT
SIpmQoVz2Oz5eEUDvKxuQMqb1gDVcdYdRCwWT8u1yUd6ZFdJ0NQuxL7ydgN9N5gRUO3k8Yb1R9bT
nd+Ad1/8swwbzQ3QNE+CfxiFL0s+aDvnoweyFft5WnSVkk7/mubT3gk4YMmo/DJGGPrZIOtUdPcA
WsUfCT8ksPV2uhiYBv8KoE2CNORzX5DSroNlXe0LCf9bVobgmd8nxMXHkiYxgY/aUUx8XrakdfJT
Z276pm3TNUWp8c4IZmlwKLCu8VEFNpU2zroshLVW0jNdo4C6tWeEaiv0h+79vfphs7a6GdW4aHDz
9D2+5E0OqAT6lzUyR0gRWDAYFloyLWRTW2hH/h/lXniGG9EkiThSGb3d42E5bqv/rXsePdJnIyRi
2ZefMrwdc2642dMocQ/ywUmkDxaZ8ahmEsIxpiFhYWifn9ZixRGCDU5fI2mWJiJmRRnUbUHMqhB6
JgxxhQagNgTG1ptR57agu4ORssDGOao9Q06NUxFJawif+ItTKnQPDatxA8sBMv7PkUuffRqeNfC1
QvIZ8QifqutCt8GGItTLx0ePvOrD//vicvA305SMGffksaQk4OwoZm0byy8EfI23fLctTB3wVqwj
IGdbHb7D3RSnRWzwuZ6iSX62UFFp34yCDQRM8Dz6i9s7xXIN0KtyTImy/YdqHFVIcBuc/Tkro974
Ftx25YSQFsZt3yMA4MCeRLvvws/ZphROA1BU2e56CxKMyxCAuw1e14MVO8E4R2RJ5hskzidFqpll
lNGqgtnW83QPzko7WHnlJztwTApbpqeedZSOtjBazyV2z2igmSB96GbKOKXY2hnyBJMKiPl2jNZv
qdDeHmnC1FcxyTILTsYyK4j621nZY9xdW21HrHaLnm6Sfbk8WHQf3DlWpUMe1yWJNyWrn/gDiaa7
GwzPuJrqrdKIB6dazEVIGzYKcX+98aq1cQ5Xa0FyYDUc26Bi8k3jrSr2ZUYn1WzrgNfmjZ7kMCj+
OGGkqje7PkMw7R/mgGQIbbwjRo91tQNFNMAtnsS1Plmca0RWyUU1kbrjwhsIAps5Jtn0gvAd5Rv2
NqVVTv1GYllVpq7ZyskyFF1nO9tOhGKdNNJtnVw9F2i/I9QpwW+CTrFbnve1ZdDCsVesXWSVbJ5r
xhKmZr8MrLvDF26JMmPVjvfA+zJQogA//jWAsT7GSwcS71vlvmEZJtIhM4VT2vIRInOjnNIMDEd3
mPBptl7bjsVL7K3ipWPok+B7A8fhPOdDrwd04ZYLMS8+Q59k3XSsPj0IA8nJ86QZ9XaYOwVzL/Nm
ZEMlpg4apyJ7gJeeP1RzrXGovpem1ywnckv0Y0ljc94d7XzHIKEw83zAWEMpAXnG8+KyfUqKHKat
74hbtTZjhOPazn6I0FFG19ORtQpPgT6JrYI+mUR7tLn6vPod5+wLTsqsR5KdXnXmENU+jfqMh1uj
gfVpENZILs6xMG8nzbbaOAGatApE72oJ3riakMBXrOmaGV4vlX9srqSAdDT0eV4Dv6OHvd6tigEa
J3r1AHnLkIJVSzmFgaDj31gtVGCZtt6QpjtqDJ9noJWyPvBoQ9v3yfEQKu01yzuu6bnNtcyw8o9p
IERrB3yVBIwMJbdcv02optEdhNxrVBCWzOrerx1ZEdmVVyOVNhy7s1ysLdiBSUwHjdw8pZaXWOSQ
VerGwqLEo4YW41wrLs9T7kPdBXfyHmKQxhwv9k9gR3dk2UYb7UtUsk1S+cOIsk5QXYnAlq+l0Osm
rWEs1orHzqoMxBGg/C2ORC8HO4UvR2Pd9VvVuyTk0LTZ7IvU/5khmOOEwn66uIP5SmHNu1EVLFlG
Eeapaukv/DMghSEXU/irfN8vaG0192X3M1RncxfWNNaFcJYaLIV8t3W3McOap9bz8mSCLbFWkhAx
1Wjs584EHsJkS6BLvz9R4cfDHGyThklbOy2cbC8HT/xsh447GIPbFXlEJnMMMmyojh5j+ZAd38Hn
ceX9J/y7tNCURBPFvk9fM6oZbMSNH5IRTeXL0fED02UOMyr+RXhi8MB2wS6b1pBxvX1tPoJ4afU0
qXctBlvxcX7lF50FxHRmSaKBc3qwKxDBUxwOi80LnADvJ/Eg5AoBnTDJInagKeIKFq+EtLeguYrw
S3rxcx6N4e2PJi1bKa2yYhLxjxm8nd6eGd3PNmoXSJaZQL3rpfdtYsdX1Uam//bC8mx7MgYS8fjl
w2Ju+QYLczfbwO6mOE4KrJyU/I1wgFRb3r7Th3HN4bEzZrMg7KFyam0hMyU1ac0XDF6RZnq4q3Eg
mH6ljiI/6sbnbnCxJ3JHQAtcxhUV5KR2e/I8q/BswSFjphvuvfyPlCF+3eWOi3SVriIGxX1tw7p8
oZn1DCy8AaPGJWv7+OS0XFQ2GV7IScM+Rjtn6tBNZUudTM70zne76sfJlI3MR+FSBNhUXD5s/7ZB
rFrL+foFs5ITms3rdFAyC43CqDiLL4jDbZA82jXh58xDsvRHEyYGpianlsS0jXzrIQ6RnCc1m5zw
DD8QJH3eWfWPEtQSIebxe/H7PET5fyEUlYkd6qPGC+xxwdqalJMqrQIQpGJnr08n+bLyD0AVf6gE
Rxb3Sxi2+y+FJgGUbEhr9gU/n52VyG5J6EHQg2VOQE7hO3qG2docs1Qu6zhrzruHaUHBWxitxd6Q
XETiPp12gi6mccaL44WqHjDLs71vABpiO9oZPyGy4dkdUkMMBrPG+h3LodG6EexVf5oYwuveafri
6CGRDqSxcz/H6Rn5ozHHPj2SuKQZHEfQeHuEz5CsFRA7uGCWd7dFWCWdXbytckreEP5FM9hbFfTA
k7f53Jyrzl6XTMRb+MXQQce+j37GNvk0VLTCSUDQr5tl928LDWSNkXRtBykRJpGgbFD50dlJLUdK
XNbrRsKBpbAXtftY92vzvB8toVLMWI2jqHeyE6vdJp2jgSpnaiiDCH+i6Rx2oRRGc8HEHo9TSo7n
XJGk5oO8xP8k9QN0kzhUDGhZm9CKewwy7o9a7qgJe/6f+WfxrNflDsv5QBtiLtwfAcX+h2int27G
Pu5OO4eJyfAa3eeSelD34AEsFkw6KxiMvVJZV1etXOI4E4ltbquZTKV84YEFvnIHzSAAygMXZLby
FiGS5ttcN3OoXIRSKwKthx8yq5U7ZtzQshrffn7t5gU5yMgsmGDamRznrAZNommBEcP2UupJT/ZJ
FlqT2El7Cy5mgIgkLuBR0dqwR0Ls7qpPTwdFfWESD4RB9Wv8XxeX3+C21sQdeoqWrpKSWGXOfeTw
5HFozR/qYJzOd//Lu1d1pBoMRAeu90ewadv7KMGjbCxTUdeybtaxQ0mhRjsPUj7jFolDF64yCLLx
a2Uc5uo5kLtO0J8O1Cm25rWFKiTDjEK+NdrtKryDqh8oUivN0hntetowJzXjcomgdF7x4dlY8Wna
taY3p6/RXQIxxJ52s9qxGxreWJ6MVqNySJSE1Vj0QYT9KjXEY1uOKVEShpq42KhFlymYMXT2jzzN
6o8ePcLCT+uEBkqKF0XhfX7HUdqdBtuL+xvE90wroQYxhkGHI4K5EOxCPN+kU3fO5M+oilzFq5Fz
isrYv4UaigyV4jQ+JWt+QUMSlXg0oS2K7xwzTRIvyGZuIklr/N+cx7HZjV27fK+zV2xUzenrOU1a
qf6Vao8LfX/mBm7lzJQsrHwKnMa8DsrqK3jMOQlqfy0JGZbw0HAdj8QSrQep4vl3wbDYgzQceDii
IO6FjHCdRyXVfCRnj5WmdFtC74rx2oYqFkWIYpTiG0v+MkpBxbQZZ3iFtvGhFBeb/3jQyqWM0Frs
vghkml6Jl1JUu4V9BAWmv618I36RTeHyylO88Vg3ALSO2rUeR0QhJhmpo8tr9oQpj6pfX0gkILke
bKczXDZuBzcg2JVIBNTPai7s1cnGfDwiG/BhqwfS4mxzl5zyfXGYdURmECdOsvi8x5HhXTHqL7eF
arrgfqRjLq4m54gq+yiQq9U6tYkPu8ks61e+6uov5YDqJihtSgUCWxRC92RqyJWqYwk9IBH78nRN
gvrYmxRRsjvrK1jrkyNDkdcJ0KXuXB6q369uyLa9KBAC26vOhjJoAimnNo3k3jviRvHi84YCzBxa
pM9Atpx7gYUfrs79uS4kgEq0o5dWtmIfxuM2Lzv0Ef/BJIvXT8kCN8QOuZxJFpld2RI0xN22DzqM
o/2Il+Rw+9dOvurcQDPWD/XYx4FlVWe5vZVn+lmo80YUpPHN79c5jRnojcMWobMd0mpxRMn5nCs8
b5221F6DBYTc2b8Ussk4e+inbh4vse9DBJrs4f9MfljLbwqudLWK6Ou8cMQlFS1fKLomcFnzEJAb
hYaTtyiX8SlQxef+pdBAYuPk/Kk6EnzMXjocamPYMrbkzLnihvudTE0TlsU+HuVfuoudEMa9u8DW
NvgbBqkmAiqgh0OZDpZqTXE+bbbiuqCks/2oX7Gsf0n24iBk4GalNeqRjOWuFO1d5VtAtStcCqZf
CX2OQK3dWh4v9H02MmIWcPwYlqKwU1SNKyAgqrcAgE0sm69YD/Q53NxYis4sP+71nCXPeHNehyPD
SbJJ5EIKMibM7kF8pac5JD7H7JNa6g1bmd3dDnhIWUt5tBXwxl5IcuYss1sfyN7tI4b8azcF8O1j
L5U3Pg2hSLBpeeE4D9LJ2c9CR20O7mbW7AFmhdh/ghT/635OxKmalL5w5nFbgTNP2WdwaG0+s9vY
XPOp53F86VnX8HppKt/I2aeDC8IkrtTew/BeWN0jZcfDT6F0dYR/MCdczwAP/U1fyaXiCRKlNYCz
oovNl6UsS7ynSjUT5LFwjdQuwTtiJKGrd3jeUmIHqFTztyux21PVNFh+8sYoeTz7W1wpnnMnkoN5
XYXpQlMQo0o6c2cOALUPb916kB6AeIMqHk9oY6aS3A0iIa5HEH70VJdMbteTgggnxpWpN47+Dhi+
DXU9clQhNSf+UkElqvgDQJTWM/Myqe5cMqmiSLUQpK5e24FzEB9QB1fYf9XOMJZYJLK9NQax5Qc2
QXARUoNP/rkZUpopPO3QHbZ2WVGzcizixrlKZtW8uBTiBhFkJhWTFheqseLsvtvOMKuN6UYmb+et
eRL4mMb+IMnyRKcxqye53zHAgXKdrjIjdOL5hsNP5oY+pPhJk0Xvfb40ePlB3NlyoAabzxAfqLjW
yatrbQ7pGfoaGLAnVHoJ0v8jKofzmt09nAQ6nzh9lrnVer6T3dGB2dKtyS6cAn1H8I1FVDAaQwAy
p2U9CikdyypdGbJRLPnr6x6pC/hJoconvc4F6qXfoCO5m3j+oko6jPIEpsdtCE1njLCPHc+AYZqd
vLQ3GERopauwjEwwqKsc5g/v+ypAqdI40NP9558wcRgDGAQ3ap5mijv5RV6QPiCCsedktY60WcUe
NzBGbaB7IYvLxbVAjKs9h/2jAtWjXkoW42mofz8TJFEk0+IIGvc+mYVhzUgNhVj8uG4tgAWm04lo
uv+zUZJ++YXuNRdZD0zUFXRfZMZur48wY7mZ2EnQIl/OUxYqxY1WscA1gHQcIH/RiEBNX8tnrdz1
5Gg1FK7a2QRm5D6HeAr76aVZLKyt4wNrXXRXOB312M8XlCvBQLU10VmkYn1i5m5/kofF2Qy8O8Jf
SMmRjRaW0Sywg/mxdFqMb/rVWL2dUqWWo0HnSWquICBTv14HyYz9JP4yLVLqZyvR0UEnQck4+uFw
gdaaW8L9M9E3zeCTadUlNGOxiaW07oMIvhRGBTFdB/kzwICLvD3HMZ6n70ygqdfM7WysImDdkkYs
z5G27PNMhk1C0vIQFfHFrfR62enTVPMMy2ml4Oxfwm9Fffs+wN1a1DyQa6HYaADzvPTWfnH9ScVo
KyIphASxKehL+DqhBxbWDR5bbmNMo601+NscSJSd0LhD5xD0L78sIfsHcYBK4PQfjwjE1N2e9iM2
Xt8A1ZdKpGlGNsJ/hm04VzdSPcsdfIEZWWWzhaiCNwbXA9CmyvFUAcVGZqmS/dLazA8u4fUZugmn
+urZhL8lYuVPGhEdGu20LS/Ok5+9be1YoMKtd/m4sIHpky12HNtssDE1/iNI3KQ3tIi6Sy6ue7wl
bPGA7yrJvIL5J56o2b6r1CSwrhxxUEi7zPdpkTC6yqXCR7s1hs2VIAfTOoe3HiNjrsQCtl/zTjls
pNhERyCo5HiD8KjnuDia4yW5WjMfL2NmJoHHM3zmjTvxh66jAdf/20gn7JMqMvDg4C0C1v/WE7Pv
I8JrEtOUM9fXHK3vkdCFjTrld2K2iQ2QhlyRdJGj20VfYg+pCM3RXOLOhbR7vggRJQ2bc7ht/un6
SSNKIuUr5iETn7lnjJ1bh9+wkhcp5gq2BLy3GoY8TwIdRO8Hm2SAm64p4z6btWpZyViNrv7hzHjN
vsENhAvBx+p6aaZ5OMI5irusxDwiAjBsbROugjDFkmK5SJnmLYr5+QFu1pMKRIk/uKzXZqOxyDDK
9BqMHel2OScZFZ+jlWDyiAFO4ClKw+yWZ+55SpyA5R9AVhzYpUEt2ZjmHMidgduGQz+Uq9qy++hb
ZHer56mc7DlbzmuiNBKIlIOzo+42RLKNIBfJP/aeAR6fgXZbDrthM2V8JcZ1TnrB01aob9k4BUU0
mYLxi8L9D9LU+9wKD/2izbl6+h5RlCwPyn+aB+ZmePXLaym88SnKNKB+gne+fWiIP/rVePIKlOZd
h1ERYondQpN7uqRxICNxwW07FF+g5GnsBG2rPF/y9VjWqy3Bj2wUFfpowcrBCXfm9j91CLXkMWyy
z4Gvubo40zl4qTM/TAS2Rb5RZ9JcfkZA6xmvrrMNVPH34cD8YkUzaOnl/KYLWNKlN6NTQRasGkV7
jCpk0pnLCt7+Gje/nSmPT09vdig2wQkiHMqK/LUv0dO+sJO2WCM+pBl8HrJDPh2fHjAATxiO3syN
yx+onaCAzsDl00BRSChqwyWNCgm2neNXwAIqOBbcHTCJUL56cqz8BP+bim7Nnz18mpB6oMUR8qOY
F14/tPf/FlGBQvhCmAZ0+qK4atXoT5M/xDC0pkyR05nfS0W9SU675yPaK8QvDxr9JjYrojZVEWko
Fe09W/2iKnAFU2WfmGwAYOXVOADwJb4cq06F6yUsIEQb4EQvesGbNaSedfqxWaQqkjCkfjb73OIV
QQ/G7xWCgJh0fRUl8NhvVtn0ZoENBf16WtiOzoAnrjUWgtX8/nUpxAT2SsUMZb8/wMTD/C5cEMvU
/iTvu68+fgtZ91u0GMVKEMe4eBYLrfidG0dUZnNU2QcmuBDGk1MRS7JDsxShDXadFQ3/CZbvxBw2
FMsrLdTfztQM/7g6udv+0iOIEQBI2fBYer+b83R/zVSK47tMHpFvCnSStyGuGGiJreIA7/mz8Uee
yEPWDCvrC7DlZLxlKgG6Zm5WbelSFkmnxFeGLZZq2+za4ndhB/C7H9g/hzYCI47+jvDpMtKzDgKL
2E0mFY43RSzEDptbheHjPaOIqqUCsHkPzBt2iwPTaBIqaiT4iQmgw+uP3NvIJGM6pM7Lj17LXzvw
1qlze+fk7f84+hF+tpuScNFAXkUXJX85eu1CIsN8hXLV/JM7cX1hEw4WdTybBCuca2MMHCaiybEn
+PiXHpRuCUstucnxxXwdgJOBdPbKT4iQWhOvBHTwn73TPUXq/w6osBPIWwQhiAPty8SGqPah8gLa
gS7Ik8oh4F2//Vz0UvaoKO/D2znE5QEFSOxTvTfifP4swpwZodmYzy0//fVJWhTlXVFn+BXAaWVO
o3AwxFiGK7spBZKn8Q1Q8JUGj0lPMTB0tHXhwsQXYO0tHslrdMuEoljg41Klrnbe7FVHDfjAePld
DXWuGeZquU0r4Mxfc5c8EykLnzbxpIXS7kt3+9XcToUT2Mjc0R8FBes9RO7GShB1h+NgKphdTvvi
GJHGfFNl5hhuK2/RY4B3+YvSf87ZZdXqBWmxetIAIxGsYjfH/AqqHrOZ7j6mvTm72A6P8Vi+dYHH
x6z7Loh37P5G+vxmHiJ8jeFr/tb1NtKNgZrN9EXP12J4keeAg2zcxvs7ZH1ulBlD7LjpJO9VmqJ8
njnEdx6nTGmX9zPL/97QNPmGWuXIqFsi//vvpmn38b+S16bbb7poNhj7EcT6pb+TXvzYxmDy6Ckz
xfZbk1zyTcPdqzJyU1A+V3t1AWnSOtVYJDTB17SfkhhbBr6t4UZrTD7gEOD0jlmTTZf640bAi/xP
H/jua6VaDLfZa88Pjqr5rvd4Df78s7Mt5dmEImmv0uM6pGrjFIMqOJIma2t+WVzXbUs2MLCFg03E
O3dU4uezcx6aKfz6V80OBfDNxvK+/7CJ3oEF4Kjuyw5dQz/YRfHN0lYVa8owYhdskWS36JK6qrhe
1KQnJ3RF8l8yXSBJZQnQcha3Wu2rOzE/zeTOgLSUp/qwbJwnmHU/uzIup5oH7UiZPwxw4oYTx4pA
dQIswR8O0IoimEcHQsE2qy/r2D9Av9FI0SyAb6k/Wl8LWvwr7/7RT5uNyagl6Y/B1Zm37xK8KfYP
17quFTt2MvncUPZltS1wip5yyDxqtl6ZBOp0tRifz6soA7mQy+me5wVZNeH7uGkhBGqBzNRJ12pc
lONuca6sI7TuU2rwxIvu6kGKCB5PGFwJho4WVOmGKvxiv6iLwA9EL8wimxg5kDWoOI/IGdhDe5nt
mdKf1Y+L/tpNEE6rTKbM8Nus0oaMIyjVfVk1Jj2Xrly+5TRXwJUm+4PjtoCSnC7A/N1i3HuAi08i
OP7/XrZfYDH5MjDesZ6Nyid121r/LCwzvhi7nl5qdOWRDnhpEyPwGqUmPh8iHJ+Hvr//ruISX1HK
6QTL+OXkFc2t7i1S++4tzG91RLN7NcBgGBRriWbhHJ5nSXNDTiVC0rFdUQxOyLWA0ede/VR7NTce
5tGso35gsUYKxdSNPYYqbApT1L//LnQ7yUTyD/EFZu7tV27vu+g86LmGo9wCrDYmC4pb7v2zJHPr
A5Rps1bnSjuFKLZwqU0Vpvf93D8QXWn5JTljdGihfBZ/QRyY48aW+aIjr4Bb9/loIT6yj0PwRKB1
zSHydtGGeJpz0vXtChtf+Sh8dQ8TKobCz3hmJA/3u3ucRxzxNu3pNhkBLueu1CjyUMe2xKved6wz
pLKhRgNquiSoyzQVINZmK2R+iKqhkxQEE5L7C7PMIelGb90kmJSleVg+GHUmCp7kBaJzlfPnN0FQ
V3KsrvWIrDWvmGPrNjCw4Dq//BuICPJKrQfdTSKjXAWJAjDgreCIlOiFTIl1xr2Ia1MxK1geXNlS
TR0Q4XDB+gfi1ywwh1xyi0FbaK+NZQngQazpCGZwXiPlr/GRJ2QVBFKwogTSLr34/e4i8QSSQZrW
fG3vTWWaxAWHQmY0JBmzMQCa1pfhXVQo5WLDgB3yXWiWNkDJVMWktFYc9fcGLZXcF3VBvRODUygA
7sJzule7JQaOSFH4FIQKBAg6Q3FgzJ3qd2QPw7DWIpqH7GknXNXe2RbnQPDAIvR8uFnd6lb+e+Fu
DovQUEE6EBHqLdAq+XZ76hcxZa8BN6F6Olu2fTWCpAC95diTnLuvI8Rov35Fu+rNds90XaNoLG4O
4T/EMzLYjw0HvE9JN9e3gZ8ai5hZbiVcN+lnCDylZqP1LmH+nuDTLo7L7gsS9FWbAgpn4MyC8ZB+
ZOi5JxJrYUrewB2N25lYtNEtaPkhvxZzwXDGX1Eh8weHY8HFuNwI8wRdrtdsg+RNcCygVK1AEr2W
1zmDfyiPvlzYGiToUmp2M29QmWbHzi5+GIYjuYOdDGkTdApjSBB20tFiA2DNYOZ6w8NCIIllDPyu
6MNpFydOn8Jmwa7sN0DAwM0P7CO2mqOR4DkH+jAe1U2hj54669FbWlTdMz5Pf4ubkFidas0E085K
6rEzCFM4O7ckFGz/20kTPMOlLs4QHvW1AvAO5vkjIBHF+OplJegfCKz8fdJPu+fYS0j/rEuJ+JYr
mWNeM08R8vcfmVFLOx5aWjnAxVIKd1GqoeJAcUES7yoOwBxBGr1Dv3EOvUPAHicYxXWqbVL37sWk
CImLg7qVRciPIDHpLaXaEQmmNGjAs4jD2KBNPPjtybb1xMoNKTLhl7oTvXvtQtQRnl1FL++N8g/1
F/ItMknEJK8vx3YR8XJaxQO3FgOCxf1r9H4KgYGWlF7rY8cgplTe/waVSaSNdCA/JUT8NpW6vPRA
T7f8LBVvAtZ5Oo3rb8VbpYcjlIhNi+5Hj+MRYSWvnQdYKMOV0LM+moCMsiR+rbEA1xKYKe3FaZ8v
naaND7A16rVg94xFGCIakCp1+PWwOtBOd5r8vED9dCB5XK/z1ujywp14AvvoX3M+D8tKvISvLoq2
dEVp6d0vZ437nA4dAfuIsqc5Z96HubBobmLCh5JQR9lS89lDukdJKhKJGfXg4ilWjKK3GJ9IQpMN
aymowUDmhZDiVkSRekgiQWApbx0EZo6izeYTSZyx5Ck4cv1YPsKJiDFNIVGmEoNnJzb2qdXge1FX
iPkyqnkv5MbaMemfZJWlLYek40XSp69EPGlfu+ZQmEyqJK069HGKUggbpfAtzcnbEchppvaRveM7
FFpKK9loxtA02f9IiXOieJo97TcLVTbW+fl2yaQXywz7B2+BHfskJ2QS00rNNtytlzcaN2X0UOi7
UGCLXfy/86DKOxZuN+OceIqEws3CMXfl1zmdlY6ymwoPvEoSfsmz4Lc631xOL8pHoD2Ay6KOMtep
uE8iPdSOUHrpKmV+D6gnF9jsiC3SByYCPbRMHitkeO5raoiVlstJXOCKGgRfjWpDhQ3jYz+DIam1
pDXvS+t7tGIHljifVoYGwxT5PrJFaYR30wueVN2ED7L8CLdS0e1Abqn/JeMaesyswE440CUHUP26
4YavK39C42gHqmoftwNyCuq/JFHiLByBxptDYasZrn/filUHmNDJaAw62ld3W0y3+Ua00PypJJkx
TKfDi3doeefFpnTgmbnbEYyrQ1hKTUwOy5ylCetA43sutS9P/czdHfrWnbaNF0vPvGs3iYnHlrYj
q3B0x6iS0XANmS6/m+JMCTdMJKQZ5LohpZOTdT7u5EoPXIMzrUqR70pNWMvN5I7l3H4F5foAmHNw
hAd4EH0cCNWDT9gd5v8PtppnGh/7hqU4R0AwHo+DCGZd6+K2ZXuZIPoy2UqXq/3Z0UDmuOu7psF8
1LtJj6qTUTgPal9NEUSxV5qZiXTO/Abw0vsZ+BDekhJ4HwN9vk7KVZhaF+YKcOvdwahdvToepzAn
jkFoBvBVmf9W/1knr2bDBW5tfbCGuxLlNZ9FAJXHkAqAEs+Az6g7CLEnvxH3hojc6NYqFbJNqTEC
Qd9Fs+oenM7muDeZ8LzTnrrHYp7rr2Sb/pV7AV4T3m9S6OY1S/jLfW6tNJ2iP6hPMGNeiqzF6lvF
o5LS9z7cRYOQX1cszO2087u5t/+1gVSXD1eEoT7LIS8JD1otvMkMS2v/DIXXeAautLYrO5+8gSZ+
IZRCHMFyf2HBO4Hu+M2fMJIYqjQyc4V8X3GQEHG+hXFwXY2lAunPkc+1cohP3JaeVKBvJwF/EcrW
jFORMsRpokBbytNkS8TB9bIPan2ZjPhMpx8OHgWal4z8fdFnzJA+DnFQ7sk5tVTkVjEYldPGrFh/
cbLawa3UxJ2dffwzcvLt3qPjSbUlOIMJ2f++ow0ftCftjtpmnijPGgjj2GybYt0P62yWfG+KjBsb
sM1yq0TYoMyVhJAYhxs8gmzDWdus0F8GnsQJvMf6f5pHA/em8zfs3XsYGd60WAxf6sON/RAr6jxb
eJr27Kqrc191wMmdgLFrVtAgOGONWqz3V7O7r5SZIupqtppnTsw4YlQSz1hK3JJJ0I+szcA9InaU
nnvjCGHbP1nCLmNeBOt1hCZCbhs0/CsQkB19pZgddQ3SFOMOq2DZJ1bzRFzDK38M9A8eRd0kDkfM
pOSl2XiNnTr4sZf4DNU4Zzmk/emLK4X620mwbAkWCaUAdYCkK169ChAIdjeD//QZAqQ8D3HdGd3h
KJk7CJSY3XpysAxuwEMPjFFvjrAkShMASgGkhQxkWnGJUhZfsbM/F6XlThAnbeQfZsyH3bc2hObv
lbeCR6QFqpdsDreWNtWg327yMevezMnjzZw4CAU1DhmA7zNVWK+hJxrROJkOZQFlEvvs/DppW8P4
RngXS1HHdFVtAPjc4k+5CrRmlu7L8kgotDNAcUPpzdmxV1OKHlSnII6cSxhyQEXgUWoEGqYq6lp8
v1aCxOoFniDR0JDumbRTlBNSlnO0eBKkW2lYtV3KRyBb0eW1V4tmdhYJPGOQ7vVgcgsHxXqq4H9r
PoqHxi1paRkyH8atzTMzJkv1gM5DnLRIgEdrepUZyfT5LYMM51Yy8A9rEbwvElNwpZdecipYtI71
xCJVvsQu1pSJYp1+oedZqSvsnNCIv0UHkbWoGEf3tzsnoUjluDNmiCGaDwbikl9edrdze5CrQY/9
HUsgKOh6wmeJQQa3h1/+v1b5CayooxJ7HWrw3ipdU0O5OyLgmkrBQil73UamQgmvmSXJ67fvAmJ4
NNaf1eGsuD4JiL1gYD7HFAeNawRA1/XqSx8mml7mzsRndbj0Kppa/7j2dSYj9zkLob5pzxKe+PRF
YlZ8ytrhnH0wVRCni6S0OX9uGL8wIdsTp+huenEc5h0h98Cu0tt4Qe9EnAyML6f+2Hj1G/avA0+5
rz6zCxmCWHY1kWnEp/Ab7qNSuyaeYbBcGWWbntRNGw8HSOev8huv8QkjEDJQ+DVg8kWBlQrPUy5q
qrq/wq5EP/h/RLSMSlpGV7PE4kSsdmLNbvsL/oDbh+borotx+7n5csVijFpJStNq7MozylBBd9iV
qFU6zInPNjevJKT+rwXUwkxBQPN+TEtoagkpVv0+yjjj9J2D0jZB6ieBkJo/oOp2AE2NzvtmYwO1
tG2C5n0gWlmJNpIrwtzuOc2+bSnpoWeeS6Idft0QHx82VGPlEhEPfnFS/5+c4z0dzmZEARgwPAys
AVy/TkWP7ryjW9GRhK7jL8L9dtryzsui6TX8BIMRKS0MwmPEuy+0M+uA6w8vxKs//jENVp+/1/aj
OrPQAqs/qUeFKDrLuRsQJn8yzsrS4vrPPM3KbEhcRD7vLkMfHbdoZlafyp5VWbYQ0WnnFuYUT0K4
cflvC9s8cDipYI9BzT8CmXZ9QTEDxKSy3/w0XJbxZuwgQ/m6Zaqids4N83QqAiP3GTQjWALnbVux
4tJf0YG1x2l9j35Du6Cx3A/KMKbTvD4sBC3hg7KvPYKCNeM91bq5p8AULY/OzRsdHzxOxl7Vbp7N
tPUGqrOt0QCM/V35SpoReGJ6bHHOGx0hE9c4EQ7AcjuAenU2nGrsHWd7BrwekvA32+yCA7i17sW5
Bvrhuq9GSzpDEeapivCvJn9F2HEaLI3mvk1zbeopROw7RMUdUYnF+kc68/wPN3SDtNl1OM8ATFUQ
VazJlhzSANPLeg90dM73amwZ/8q7YxzhghBio5pOpFUZ+m47QIIxXKHfwuOPKMaNaBRIzihvlT2q
KEVG1SBQhqBvrFyQ/7mIlr2Mhdt/BRV6gEPXf9FevhfIi7dCkJS+Dfct2fNczWDtGe7E5NB9uF3O
CQ+XfJAZg5QLbv+aBdc0j0QjkADL6lWlczGchj/WmrngGOofSx0KkddV/0SW2JvQdq6OtKYsByzP
WbUJhpIdVDNFgaNyg9jRPtUEYJBggKX5/MM2azGz+fNTAUo++3vUNhrL5aCllrtw0x97CDgTsCuL
hT4iKoeCcINqACfLFS0e11NgDSetfL2qEf/Q0HwOn9KbIDa0zD88lBTDIXavy0XucCApncJg06J3
4XbJt2vArq3/6Hez0EHt0BakJrK1bPpiTtjpIJe6JsVhkVm1NeJqvNAGcUo6GM/8ZyhFmDxGPWVH
U2/gl1yLsRk2JrHA6WR0JOWMa6Sm1PUXOCZceCQMeHZZCFUm62M7QsAvK9EU3rZ0wR280nMwB3IV
rAaSNyhQCnQca4DFcR0FvfBJobn+Twq9+PH4u6O1Lncm/TNp5qpKxSEAWh7yO1oVabPatOsloWCG
hlNfPeZ8JUIhkIjgL3hk23eapkhEIDlHds0/h9/9JAvWBTTfSAwGCLhUuxaryPL45LCNR3EHgty/
suRgtIR/VT6M6GyOwpJjO6ylJfDqLptUan7j9gQqGvJexO4NjGAey1o7MF0oVW7EiTkJMkltYJfd
D9S1Vs0UOqmhkB+q0f+VYo7vky5FU8XxJgZ8C1Tpd+WoY9LM37J/4Xzt7dwEJezJEcba2GTMCEBb
rqhKI/iXNT1LnfnvLDG9jg6yHfmQNJKov+zI0MWelfFLYJddtfe3zzfFOxpKHaGzpp+TZl92PJXr
wfrKkos6BbMKKPZaDREynpAa1jORFl3tiJd+syIRqHujNGJHP1Nub7kKHEmkkt+W322dSwK4cxJG
ZBzBj5zvjDz7fKHhpXCC4tZ3+lPXcT7dTmWMowy62sZUe3JJ2Y92b3U0kAdQCEuxBRtLsP20O78K
RbBaEOvo/8XwG4CLWy3aRmjvvt3/aRAYPZoN5Ia7RKUJxhiGVLRd5/nee2D6+9s+yYTpCrIeOgDH
OhzRDL2zcxfGoPeNo6/Hezmh/jr8rGrdVMBJ4oYdIZDLRuWNhA3jC54dUOVgOrlsJ14RhgeSYMSY
9EjfJmSgUhppr/YwJmw55RJSEWSSLLd3tPRz6MbYvB8LhVs0p8RU5JQhqIF08h+9dnDESo7rDBhk
Jl3nrR43DM5JFfViMYBw4kkqUoDQNl+PsacJCJvI6utxbZjjP3ZkpzGIjd24tE/6KK5mJCH6JO4O
oz/LUG56cYGNkLi6O/JYxQ+4QTedwbqAn5O7cpkUagKl7cxI5nVGA1SsFWXfJSd9rYK9aFfvO7u6
bvdhMtaTqvHSl/kKN6mi/MGLKYU+3gCqf11Sg5MPwDn0lYi8UGJozxuqR+9xgNEcknB84hJGqTvH
jQrlNW+d4MDVeCvbAfSE9ozysU5w9Jd0C3XLZ294dMydelMZ6868u8gvXLStM0mwPN9oHMjmc5gd
7HMND+Km2nxYk0PHHkSQIAxq33pze7jzpoTwIpYdDanU0OXJ02dcnUebYZnoMN1tpiO+Qn3qntsE
OeYepQM9a7DDRvuLXwdQ8ofohZ7AlSQuHE+Nr95p3w9hdheOPD4cI1S/kVE9QhUK/TwmvEEuWycy
VwxAMAX+dZgtubDJUMAN4V733zmHK8Zs8aMYQ5ZOgVydhKcnZAZ2mNGud+Igpkm2B0VmUqjHb04x
LA1Yz/cgEijlRAoHyTUrov45xNvbEoul4XMVicITSNvJexZTFs408LIzO+oqC+QHnEvpgHVqREch
omCtl4UbZNA/rokM3eRrMT+Y9B4Whnamwqn9UqXCSkibJ5c8OYbdJeEQwnuV6d97VdYjzVitl+mi
JNyrfFrg+TPDZT9ze1UE1KlAvadgcLQfJz1mUUnRoLqP4OhpqJPBSQk35+pC9BnVm1wZK42NitGq
XsCzPUWjKDS9FWV3swrZctU6MgZdlQ1w7CkmTYQFvvKl5gAKezeUA1ir0azaq4np6W9EwG4CIWUl
luI6zdyRptL0MDjqpjSVwRLdr0V7DZ1OInhlpBxQmZrQknLwNSrrh7znfmLced/JWWHG/+3+5aAe
T7OrQXJUG+B20+GjBm/Ed1GNGhxhkJ8Wq9stdAGJbeh/pkGjMS/CXuwYrO93eIO4ros2FzHcCvkf
4TuCCOekus4PmBQ1EY3B7DxhAq4OqjhL1QJ4TBt9FHIyHC5N5neeX03z5YfHDK+YfYX1vy6QYon0
VNVb8PTOCh2Y9GkVP062YCPDOAVoc99fpTHwThxvO5QSETw8JOMK3iVXrIJpq7TPi0A1O5SogRfS
7sLjFyZfpcnOTQ0738ASHraiTnpfrtS5nhXxIcjccnIe5puBjAPzFp2+oL7BuHEk4uCxBjyW6NeP
hENd1y/xaf76W8iwVQZ4thTS/6/Zerl7MZxkw7TzVBKK8Y1MCC4sMKOS2jzE2F94US5kcHDtv+Z8
EwBp0RqR8pnMMHtyazo4O9MlPxOeSzGq1Z6mU1wme8y6mrRo3K6fvuREEhrc08OwJqn5Nr9Y7Qc9
OEI4Q9r+7P+Zr5aZ9sZfm9bVNH0dDsxtgZcLBn1STOrbm5pOtMjx3+88dFE/ly0NJjv1TVrqKPsX
nGvO4vX7R2tkXlrYGD5KfVq2/U+3yd0POG4vEwV7VD36PhLyrgfjUE9rptb2j/1HyHaaGXvyeOcP
beIqsdkasdudXDc/7SrZyyFTkdvreAbIIXjg2IPc0JL6PBmH40MhgA7munQ1SvuIJxZ89J7NksCi
NbtIYhngMQIZPybxbbVR28hE5YcYzOWcmn5r42abD9gNpR8fS8DjZPmJKuFRBhgPnGjxbEljo9Ml
bWRinu6mugr92xzh+hHdwx7qHAsadjEE79H5Y/nzmyR7NRfuPyzCc42LBl1+oQWiTNSRd5sQ99nM
i6aLCscTPEF+Ya7PuN5edvbCzOmPX4FayHj4/dOJ5EN3hDlg9p4MD7IOFC5jlC/N6sYuFyKxpY1c
0lErwSLBOb/6raI4+Eaezu+AQCEClQJNFUcHfLpvsUWB+QDNDaTHvjLW/1/JmCGkIefTDSOLuh+I
3d07RhEFxzkMUL6QyKuVspDeDmpk8qK8faTNqNXRMIB9n0hchhgw1g+7SljlqEibOKHDm3hej244
38HjKxIjVRJhg4ZBb4FjPWLXBFJQBtUWeG6RUxSI3iK4APaaYKIhXY375El/ZGHjFZxYp1yqB4Rz
S1+c8OvE1Qb5MDCycrxVPKnlYrCnFXNU+5yU/datr54/JgHEb6wDN39FDaBA09ngVQtU9WUgmxAv
IaqO6D0agO3LfuMUwPLx1zzR/mqTPR2ItP7jiQJGPfx9kWXRlS9j6TNtvgrz1shHRnV06cc2cres
PA/WXQOU6B+Ub0nvY3WCUk3KjGyghiFDQAjwNQX+HMb3qvdc+yyK9CErWgg1W5JRLj77rqScqNgj
3DPrGomh8br7ZFSlXlbXuBWcgu10iem53dIBspMvM04demlvH2pz9dF0jmSRZpzN6qtoMoQ5ZE9f
UQRiBvq1XSOssCjzb3NQT3ezlXYafGACPYCRRzkgBjTVikLKi2ssOz2p2ky0dkyD32NR6ENgCO1D
19VTOh4FGwrRyzgPBX/eLTNbM50mG2LVX30QSVtD1HkIIpXb7+0cm4vKORAjGYbSLYN6GIWbCF/V
Vv0LWtLcle1H1Dcf0xQ6Mgtwn3Wc75Pzxo3V8fINFyO1M3MbXIomFmRqzxJg3tTYcfIuxkxfie9t
GywGssGXyx6snBQHw5w6mxniGhi6b+ar6Hr+zSsmF3rPyrF6a/qbjU+76TqC8a/4Ej9HWnnfp0iE
PjC2W7ImeneOHoBHsl80juEpRBS4BUQCQIIp9cxKGjHufPI5D60jNFoyfywsziSS9WA+/9oXnh3y
PDge4LtfOKHAF4EStPW8OIl5GsEgdF038q92KJ0eHFcsw8chl7HT9EkzJCvJ4rT7HA/9V1CiPgvU
YoiaJsM+13epuUrf4x48lvLEshu7s+wmIcWM2+ns8JdatFhcZ5abxEnPEvE3SuMyBlCDjpzMLir5
hzl0EgwSnMQMs+/qNJ7K3DW4gfzAwR04ZoBJkmPlPQtEa7edjnYRzolqbWucqSn6xYtnc1wOI3P7
CLBLyL0utNRJryWWxmqcylzBPg0B0XChp9kV7kIOcQdwqVm43jKzvet+u0gOQzL/fX3ssL2LS39w
ZKNZXCf6P3tDLdO3+aX5En0XSNrLqrQKtVLd7UC8/jZwwATitbCxhDR3i9fR+5zap8D4n/RxeNAa
t3FHBTYMXyYm4CZJBaYqQjHC9gyp//KpsypAdbPD2Daf3llYSHa33OwPkIgvJs1se3azxikEMWw6
4xC7onNnQnqjF4Eu/w2EsJm43a6yeRT9hiribxuCyk/NxljJ5pR9FAc7HdNDeWlEiYgX5/2cYK2d
SltijugbhTbSOXadvFFRhcFTGzKjqh0Jt4TLPfEkHjB6pGThsyCzLMdlUBsWF2fSrmo6FqMCkt64
29B+sYqzZViQGl2IrahBraP1PmqjlqTF+yHeC9jzN4uoG4lgI/oQFutEg0okr7tLoMIbDUx2s1q+
KtmcW8lExJ5OjnhbrMIq3TFLMDPtppiB0czxijYhoQYPoFoVUY78BN99sjTgbzAVrs3uFpo8qFbn
EpvJA9nC1iHAESVw8wxLMJ7Y4dTdSuAcR2Qqc2hjVXjb4vXVWb6RG6SDczG8gRu6GYC5Fp/ctTtv
Hrf81o/fpWIGqcMptTadRfZO087ljX0u6rzDJqoFWRVjetEWRoBkHoa2RWwwu1HoTT0vFNdKZQgw
rmsVraq4GOYyqCSdm1IR9tRJJoLpcYNQ9BBt6O8i0D5Ijb7R93V/d/F1T1A8dpBm9saW36KA7Mko
P6qQM25Ppov/X5miMC85jfWkcnd/3reK+wJsANzYGCrWGFPwODr3rno3Zgm11izIJc/y1UzRiPqj
VyOT4QoP/UsmrL/K3TD7o/dhAc81qv/60F5PUSLyXqrvdVqgpG+lpNAVMPzJbg4LgIycfwnuVlLt
YCfN0Wbcyz3itiqewl567ghNjpW8qCwMcr2k1yxniZ2HvRrp5NdIZX4r2HH/eVqM59ru+rteYGKs
nnxVFoaMt9eVEFaalRH9cx2i8FgEWKbKdwyo/6IlAm2s6QS1oM/pY4ZJCdn3gJ4iAmQj40vyp7Gp
vBK/XaaSC8iZAWMKaT5OkXT8wj11GYO3ZRCNhmHVl1Uj/BnkjiJjpClCfB5putS7FVncBbad6hkz
yh/S07V3AiawgRgROTjXLhp9jjDbztgzFuwpkxpbsXPxudATuAEi+fQZ47x/ubQ4OHZ4oNgT//yV
S0+GB5iISR9KrWvrb5YRxuDvMmNM5uC0MAuwahcKfxXOK+cNTDHKCALLMlHzdKqYbEVknvruCiyv
r73CLLW2NhaMGiCFb23hU9+xQobwC8h8kEzaYmphLtwDVOe0LV6sckdPaKX7E5FF3CcLbItnIT7g
EwzlS47Z2qWdJ3I5GK7fgh8PLfT/WWx0xcWMK4zQMfA6KVdoXU3yVoLuRi4sU5SvACmmXvK+7j7k
I36kCP4674yz7UrRUU8kv+aEkUyo9BPoPfwagFqfpvtZETHrRxOM+ZMpQqfHyFdnNvz1eC/Tw0Hz
TtCEd45kP5153LUNCXQ651aEoUI5UkE82V5q5BjfAFeBua8AGZLBPQdikGEp9OBWmWBLYapkcvGL
CL+1foMroQt/LL5zHOufJNzlPhwZJDEn22p51urzKPLg6K2tmPakgzfeg5zmNZXksf0V3VmpGMFn
r++JOWdyWu17Sbs/wUzn27m4U1QlMWeGLFFTnLHIxzbttav7pBLZPMy9ljZ18611NvuvOcfTQQyV
n1zqJEBdtuZq3SNY7aGLuv4ChBeG129RiVn8Wui5zmRoJ1F9AgiGhIgPLW0KdlD6jzb1Cz8RIVLL
8irP56BedscJIsmWVeftJ71oct4M1IJOf8iSz8zb8k/K4bFDHohnFHpO7Gn/Ux/zmLRfKTqV3Lsh
wBeQ6v0iSrs99+kvx43D7XBMsxEeb/UjgrhergRU+22pKm1r0n8mlvHapIQmuoHAb9c3ipKThHS4
4IYoQILmzj3l4pCOpmjDO2SOGM6GjPWna0ywJ8fBoCDeUwWqZhjRegvfRaHu5i2oTO5hoFvcYQ8F
/ellKUgOyo72jgcz6ebjdAbGrodw02vrQnqUxFlcz1zZGTRf2hHKBTtbU+fgIgHtCLcpk8Fa2BEQ
yiF1qsKSZ1QRBQhvmbAG7dcRep/lojcjEzb8CfnX5nsgHN1UF6hMU1htSaAoMppSM3nPc84ukmu8
EQBilN/3u3xDyvJH+nzfJ2yfDBwaErIADeDtZw5FFpQpwhv9gaIn23Cod11B9ZoTgN3ZiZqhMT3X
JO4QAGm30eJVMZBAw+vEERHZ/sbjZ+cjDtdgYytvLD5oziBQXvVjvvLz/mDEtm1/MXX0y1vimwEA
AocHSRiE8+hs8DXdm4rPUDM7T9XoeHiOHs7KC0NixHTuG1e5p7HMPBBq3SNVGRlp3PIzp4z7xrWK
MTrdRMRhpEwdw9wSneQKi4ZMvG/PImBTbEy0kyDcXbsHUQIy8pUaoedF01akSuMhLoZOs9en1WFo
Bc/mmpBgxbvzfWVRva0ZQpoCMsG7i1iX5HzDdvtbinVcbRk1vaG/KuRTB4nI2HV0dFkFlULu9CF0
Rd6QIGOown+pCNjK4hm8Jw26wnITA8PgwuE/wjL6UsS2ceMObjCF3FrY93pcC9muXCNYS4eR6z46
ri0DKyhY/4DLeQkkYF5CnYMjs4fkLXW3NKZR1zD4pPodZZbnO4Cot6dByCvlvqORnSrHF61SR3X9
lFuMix1J4Ma/IXAopLUJWd3SkNg6xFiJ0Rv3bz79WWroF7HV1wVdQL5kau+oZyRJwidvjZWySigs
QPE9N6sGmUIdsbAzKC6SjwjnypIjL2ih6IH8C477jTKbu0zw3iVyp+R3JbwDgPlgDCCd9ESqYY0N
7i3m1sMSZh/ZUKpfUopnpNrLC20aXWqTgFcDYl7dsBE/JcG+lYsfBUyg6oHkGj9nmyLUaj+87Rdk
PL4hvtBH59e/CJKiv+16n6l2KnYWgwxi8xYycQuqa2m4h/hOEQBT0LKNbBgq3SG3Wbkqx0jNph2j
50qii6CeQLQIM+7zUqU3vqqJ98ayaC+taJX16/r9F8d4ujDMOE/YYVWpsL811v1955MCfxcvochL
7jwLg3Ri7pseyLABZUYzmJZxo6OthQcbP2FJSvihezATi0UUjAVFBn36CwlKp1JX6r96zFqEHw2q
sgP7jp4ZOXw1cZBo4fC++aZMf0UWTlTPCOkooO71s57fAJjEMSiUE72We8muQFWWiW39znt8G4ZN
1iBVoRTz5p4jwSurYBAjbc8jgym9Ar6GrR+U8cPHKafJpqPKnjrsd4C8/WXkGGEsLLzPB2+ogtWy
oKS5cEbg1ufeDXSrglwh0K5jlB6RtS0qZp6NqjIhmFydD1VH9rbnF+MYCyJAqUm/CdJXyP6zOd4A
nfxXEfcBM1t913ruIvx9xS/9D0BkY7f6f6c0EcRrvbBpWdO+VGyulhBsZvvro/uTNfSaBr4QWDeV
btg/EDAC+yHvouAwYoUCowPSiJVmyet2gz8wMaXWkITPet3IXKocZ4gJnmTRCTAFTYuI/0YvDP22
tA1qSSO1r5aBJSGXLiOPKmoZ/JflHeXqLsuoE+G16WdMQs7dBuQ1kgKjvY+5Dm0XJOFUVO56gfDd
ktiVCTXIdmCuH8453pknBpLIxOqR/y8QOmkjuwDhhliPjYz/+FgugnxTYwU6CW7QV3AQEuaF2Oi3
rUHGANTiOur1WccgWcPNF4wQ2/lmMFChTcTzJjubVSya7Yo0aHjneVkF2lSiFG1UTLXSPi4r4EVa
9Aox4s6LkpMwtm/zsyZ84WgGztRs+WRsELiRZKBVz3U79HjHpcaFdrYiQDVhUMer08dpUjNLvkpK
Q4VpDFuoz25jWAktRut3yQXsvV0qrPVBPZIGiGroJVXitYcR7RlM2a9Atzvi9xgK7Mma/G+V5fdH
JT+0OVzxjUU06XFdSoD9V5Wxs39jhTEJ/lRwfm3uZ4UG0QjQlnblpL+U4hoYmDv7fEBCRr0SYuPv
8KNDzqVP0b8O/FP6JWianNcuTqNOG8IYMuOIjipIcjhlO/gZUwtB58RDCAy20dDVx3INR3Sb1TRN
TZ3D8ZuIyrkt2iZ452Qxbu5bidZuNohKxf0IIGNHpLRPe5k4wI/luMIfQUhEW6D3HmyLF2pN8Cgt
oyr9usUufedO70taCNzCDjIGpU4MCFgurClkWd+q5dKHFvIbhtQTxZ+EnSt7T6ZTREYv0Yai9g5Z
aYi/GCSQeYSfmSBTt1iz44pJDJ3UvVa6bcBb8KIte5Q+XILZ+kMH2SEdDTmVFoZfYNRBd1HqScUc
lCRAPtKp9r6ytgEy6gl9r1AXr4Kax9wlIdfQcoHdBl7s/XtcVVoNXN9dFjy0tkgNqCjnkCUHjdXZ
8Jliw5VB/I5kBaxKbyKrcr+2H7Ovah8xlB3zIgFLf8XpGs3AMs3gDndinH0XjznFYAIxpH/a8+gR
zeZHnCQpYguQVggUNTwXiTiwLlH25jPIaFT5tgqSMgS8p4ZSCvuF/BJ+6ilXO7Bs/vNd7pE/sPdt
QEj7OLMOR3bNzMaRBL3PRekcZiuW83rUF+AfD/kwa2YKO+R578x2+5yc4J8PjRku5gdNzyLVAJgG
CYPWRky/zCvCjjPNA3dWCccAw+AVk3OjqIHbjEnVCy4WUAD8XvvHDYHtjZg/1+c7lQfmyfZvoOUW
sGE7QFOJ8PfiE8UMZq/su+HYwrAZ3L8Pz1FTMDq/nz10PyNshhp1uCbUCOcyGdlAPyM4hCmBF1EJ
LrTZP7tRNyZz4JfMiaW3L+mG8GZ16blGGJFVXp5UM/aPfLSTD6gFwAFhnRFj4pk7A4dnRO7U9cBR
VLh2g1WD2nCf0JSgrGL4T287nRYCYv0gijLqJMogAB+5laXN0pZnplqNZQ1PP7n90RbRUw3nNVsy
fi4ESssU55Hk0wX3kfHZsQ1BL6jWqweT55C1eQJa6pHj2A2oACwh4pYuqAMeJp/1sRNpWty+YyVb
yEkmF9w4dH43aO1fT5Eewb4TbQ57B4puerT5TimSiP/ctoEw4V9gZV7wn02BGBXdh2Bk7gF6mBXk
0Ox+2bx5fL7RPQ2zSU9SSJxeWGsLCNQ4vbdnNTy9+xbLcrvXlPmk5b9w6uZV07yzPAnRhKfwPLUG
NR/tejy7PLxHF3YRlxbunWnCQcfVv94+6hWwEqLNRzPu2fBUdJukbYrdoJKWTaVqiJuErxBSSwvs
DwqHCHG5ykLwi4nt7co30tpDvO4eqm+99/FhqUk+ZRoTjCmB7DVltDr8NNlTpNaAZVg9bAhY7YzZ
UDkPp23sj+0GytCGt+5HUMw1gWehhAXSJxkxHAxrfOiUXy2YXMbAOzR1xOwpczos5n3X6CftOcm7
kF+w8l64/mWNp28ndkmsyIlRgjiulJ8HeDSfFSo0wY+VkJJZsTtww6gN88kkJC0E4TJkfY6At4fv
aoe9dTuRit5RcgJLAFN9cHk0yhVU+DhDpsyzFS/r2FtEPxVUUoTcASfnWuvSuq0EZynOlTVNTzEA
kC8StjnsZd2nRugm2wYz1F3rYyCu+nuKJxM1UqdEw5deJj/TPpM2QMt7A7XY9Q8a/OrRZFHLqXCE
6nx1sMOF50qHKFQPdtCZhljQf28u/rYaQgKmbFveGf12YwbziZlMe2XOyvqaALd8Mg9TSRUbMjEj
sfNeV1WqdvDys56FYxyXSZ0+/J4MTMPKkkQYfbrR/FqOWgQLI9VwWKZIcBYPtBBlA90tG7aHpN+7
3TQiRL/zNeoVJ+72yfL+nhqIqLpmLEDMAHCrIlguQ4vfowOLbSSs8AIrA749uF8Qjkcrhx5kUTE9
k7CypibaPRihPEQbRh29ANnlU60ZAszBbEFi/Msf/IjhYyXHcCc5+PaDbZ2K7Kz6OnabsFsiHoM/
ZjM0CP3yB+3LI/s6y4+fbOeocZVqsb+4ToukknTIKtZUAGa2sB6d2PWx4YaUBTMOd2Rrk2i2E9ul
NU3loC6Wdz3steJYA7XtAXRpuKkeZ/snkYXyXYtKKH0Csx0nLpMxBp9urKgbcHy9SbN7l28/HlZp
GyAqHE1iK4DgooVy67R8+/Ar96jhDlcPxniEVv6eXniI6FqTPkB1AyYWkditsDNjun1ah8nYOOSV
LzCGJr8ZPGPwUtwnKSp38B2lG8eL8YIuzYsCmQPmSCX+9Ti2Gt7JN1NBTPtoyEE0fkFHEb5+uyiA
hGCBya9yLYVhDgla/HQu7HlroIepgk0YeDsUUl9Dyw/Bix/TlRzZkaF4yevAGhnGnucd/clpP5R1
YktPXw1Xn9tUxpTS/n5BgaA1M7eoTZ9RAw5bWClT5stWZb2JuXBf17UuXMtjGy9K8ekWzwEKTB7I
piPyD4N5WFQSLQm/RPlumfC/hPkMYdiSqvPF+MV2a/dVmaysOmVH+7mEj/t9j9YFj31v0qLHzMGe
8ln+W0IsgO0ZrkN4eYJaD3/GtahoVDF6kbLu8rZPbyg51dh/qArD0pM+o0ANTy1mCA/vHkITjiUM
3xW6YH6brGPLS/vU5wCRDe4/kjVByZHwVd0Il1nCv/MpI8s1vdVHfw7W8h8MzPKuzv7tbOsJ1e85
Z0iO2C5GIO59Zvj2bzbXmYDziCFGCD7VEvWJlXdk2PXDAdodQAW+e0Rc46NIZ7pHLYomZCBmvVN9
Xhr6ywh55KT2iIFsQECqzBMiz5uO3GIAQMIw871HTf/5ZiqhlHWHhrFIOv/luu5+8v3yk0QTa9EC
z8Q9ONraybbPFeKBGqaaDVYJDK825nGhjt0TYBUOZFqm1lZ+20u1EUQ7F54RzG1WF+PUzzpWmiqW
HPNpn2hEsjzFKigY6/GQan6rhFph1f6reodVOflWybSdegRHbzSR7d4FNxRFe6iAWrVo3KT2rQEp
lL1puJO8y3hrnlqW5x4virne081Qk6aaRLp+aosiyO2wsjFJy9uEEgYzF0SjR+VHKq0sEMcoytEq
d8OuU5SGywRh+lzBru8cQ7Q5HFf0iDXfYcYvFNMI9Cv+AUl5w6qgDUjA1wjjz2Hkjinkzf7GIrE/
lv4+skXAknm0thfcwsjLsE+e50t8v7VzrZpKZppvMLEvaDxF/mIHfKX+QZgOoOiPQj4rzrPO0Yw/
78KiwxxQRHub+0T05q1yUmF1QI/Lv/5pnPMRJwMiJvPu5cm3Y+UAHCxBVgnO8DIY2QvZ1LYAgg09
MJutxByHScn7oB9QvMq28HVV7X5EgTd7bbjrHLqqAg5X4U57xQ6Ry/L7SLiNkW10peyyICYq0S/1
yoDI8vUkyhV58K8wKY+ULEmKmdoiSxEO0hb8/RQopNVmLEpJoqVQ+JCfHyPCTk20sNVD7gLkJCyz
ix/rZQa/8Ddjr0+xSHZJpRbebaCh+5YSCdoUqMh6Fv9AT1aSk8e5rIPdbN8DpNPVL2H9kSbKabnO
i676/S82lwSio0b10qx3DCoQnK8kNgCY/Fn8/lbVguEXdgwSUa9Ej7pmp9hshGkZkEq6TRQ2wqyN
qDO8FQPWpHVITnJRWezRpdfK1UYVIRyAtCoCOV8xbrLsMJYOP7hIHJPS0PTwUdo0bS6VmojTLrQ+
7vG+2uQe7DdHb51wD3B3E8IcWSVY+7OE7H8nSVgYUH1Z6Nb195ryBLsx7eDdMUvKUNwocmMMU8DN
x2ExfB58SqwdcEDCSChy5h2w7IUWRmp26Jo3Jq0ZlFJMkjgJRz9IVVw2scokSudG+AWKbXQtlx1j
Pwt6s7pfcGUqEbG8FIB+m4RqhqqRmw1XP0ojtiJRmEv6uLQntX2lprHT6Y41IqhZwjUbyUC/mYnI
PC/gyFqpWWkyzp93kI2khq78DVByJTQnzVmF6a0Gh3GzIq58kkBhcaRhlewx9JB2QegCaE8aWsZ3
OE8bPdHfUequs32EY30vz0bCho5YGWbcPYqG+fZ/GwkX4+kIzgOB3H7Dhm0FN4cLpAGfr/ZMs6gB
TAhK/xg98YyFVV5U+w4UeuPFTeLjC3V4ar3IqsrReN1hz/2guf64uf8cwackRCCCkRdITSEkUb4m
hsSev9ya+g3nG/5hbKAXc8ac+YPIq4ldAy6As7yGH9doPUKiQIl2O97WkSNZaJ5P5CtcyPPVeOE0
VVpu9AKQrlb2npLG6ICc9GtRfcOzhCNdnY91FEjlW5ivovxPjtaBxE0tUF/RHyJ3a172eMiloEEa
2HOg7+lKStFl2wkfnmi/vokn0pcsjkQ8M4f5591ulFf0g+LnUz2iHnSu22FeQZ9MMkkLDURH7uIq
eIYlk22WfNP/JudYN3QRJipl27UV9JjvJfLw7CM+vYH0Lv/qxNQtB46vPMxapLX/5Ika9avVu/fL
t/FM7E5ZGpvNAg6fX3S8YWOuN8bHAFWwSGEza0IXqxJd5wY6mi0ss0TfxBotjPzfKAJ2YATgZIra
Oo1xO358ajGYXeaRlK6FKOloOjsNiTr5Te/lBosbYoZuj681GCOJ4HJgEsu3mWctWQG4mooXo6M9
3me+q3LAjjgyQRcTN0L7igetJEH9eGBqz+lWAFilq08ttc9emXfRbOyOWGRRx5Ygi0HkhRRdIgTd
JUbRhXjodNoUuBN6yTedEMPM4bt7YAoQPvcbfaA7JvaWIhvgZTVpHfcrX20bzvyD+HCabuyN2RB6
aPuaUTGKvPwxicMfZ53a24FUJ6kNOO+YljT0c8uG7mcDRb8yJ9qaDy6nuh69lRu9rDb6EXjP62uA
1BGlDY1nZb3cbGJ0z2lPadbscw0ExukP1Ga4VI9/pNCFEM7DdaxDRFjTYC/zIMguth4vwAqXRcLR
+1e5t4OJrDYAOSoE48Basf33mIkLKh0GCopg9uEmB0SjhoQ91RIhQj+QjWuAKtoBmx1h7TVvYXFo
NeAEYkFdwxVhz4ILpYZKGLNPjSTLFQUsgEhcUEmI5rm03ZqHUwFuABHY7ZzbnugUhNUbB/xkGWid
xa6C7DCocg8JbVK+EXFVZm75LLlEogqcaq88ZWMGRKsfmprVIJKWwm8dJTaQXlRBGpGfByQJMA7g
vCxN8n7AHEVnd3Ahq2rtFUJQKCup4ZXZvK9wknNSY8HuJFCbp4MbRlkN17m7Giurs/YBFVUda2LS
QxfTdxBn6FLfOuHZND+N0HdSVfPVeFELSd67Hknr+2OJbGEf/88xGX6SUZG8pYDX+d2YTSqmu7Ts
8HyAJ8VWPNYFftEvhsYvdQNyVcdEJfik8yvnHmFqjFbs8J+8zuT5n/GEL9oC+WSOULhcW4v/Wfit
ZoHIAfr3HbZAJK51QjHWK6xJUhI5nLfQBuJfMnpRwZVzuV0knMTxxwKnQToRNXQa3M0XjvjMWjaH
yAvYH5VCw6dgzrzv43eN/hPNZk6CT7tR1gpps6Wn6Q7fFu3PzGLH/xStMqKFBrV510Ei1hZ4EHFf
+DrQOvX528OMzaDaHy4OMpk8PP8HjW8YB+5PBB8+ltrdh20fSZE5Oj2+neiyPDIVob7IYmxqTW0P
r1Pt6tOMjb8YPBmRpxmPrSb31Rhi+xUyaMZe0zuP0dqNAh9gKhukGCg5OALLB2owrXj0q9XFO5U8
hrbz2XpzqRfOwZYMwU8AGPaK6CWexX5Bx/KwLD3rtEis3Ocr8kzPaYyAd3KHtRcza3/tT+eM4/u8
xtcc2TQuC1wj6t8DGFIlkHoFuQ6KIIkIxu/LGJ39F1R4eDIm/nm5pmU+guHq7w/tmSOnkVkj3gmI
O4RjgZfcbs/O4kE0XHU2UfSNH2i/dNAb3ujNKZiI0z9VJF/GyOdvrdPwJLTjBTvf4eHF6s2ErwxE
mQqVVhI73r2xt+DQsGCd9Ql7SNyXB+TJmIqEVjq7Mh2tQx63FuCfXNWQCEIlxISKolN3gj5Lptgn
hQx/37VfAF+yx7UdU3WCpLrkXv/2gkkuwFWk4mi5iHhr2nwQIhbOlp7cSHltwnKcmL0TICT0bu4+
hnPLQcFfaYXGdXDD0gAOzWERs1jrV1MDNAVXMSrq52bx2B9+6Kh02wfuEwQgzbykEqW+jEiXqOro
SrueflUKRJrmksEozkY0zfTyyTjhatN0EGJRb5ZOdsIO+VMzIuEyxLwADP2zf+BtXtY8wivVlJ74
St6jUlR4WMbD086m60gRfHILz+I1zIuVZ18vt/EOzTk0BoTKRHkq7FYJRe9NL8qQ9vUROF4ZHWtq
/8tKYfM0EN3h5nAujz43m4Y3KiAEpV6Ps+saVzDrIQI4lmgqv5HINSvXqsZC7HcvXJXbtGmMvZ4A
0S2ZXMOLnSLAAi4GfK5vWjb0Io7fjD4Sk2MpUv7SiTsWa0uG+IWAklafChJHctYtvtnwanKMwJOx
smIb/jgvPXZ+2eERsX9yqU1YbSvynwCwx0ZcYweuYe+jj9RDYmnWz9yBR+N50/kmDApok/GC8fdf
GXjHaZ8ckSVCysNbNuf1RJsgbCv8TBVLBI+xsQWYbRp4b+P/6jzuZZLljEBoZHPraere/QjC9+Z1
QsIqKQLsRmEfMRVJXBH33oQIz+vfuDMrnBsoMCtSVc8Qxlut37JTfrMZ4SDNlACB1yx5XZWEPbtq
0pq9ko68nb76A7Zib7x3BKSI/sEFgQc7uomgJw/+BJnuFxZGt0pQyhlcHXsilhlOWs1df1xqDVMc
jrpTbB55lHM1EBShos2aMVBJ3d8sZ+q8xS+ps3sjCwtgEGE/x9nRibqX6Fcqsfaku8GYmUYqQ5QP
Dw4MQfilWcBgq3bX/9+hQb1D9Hf6lj06XQ9yXCrUir0tZDSrE4nfuxmvBYaAN4izQhoJVJuer7U6
dl9RrN1ssNGSW5f2lMcszzLYYqWVFTPAQ07+1RmSUY994PW+o+wzFPCDZkP+YUMYeMGDkDb2Y4mN
VtyGDtJ1WdKzpg27Ny10SFzsAjCM9nReEpnFBUsyrUE8xY/Ky7LCL/aD7rf2IosiG/JyawmQKK7t
dpXJTd6sVdfswyjti2CdMUgQV5sYu+dPcTW3gWx1z7qoiHBNOEXsvtNwF1ar43i4E6S/EeCMphwA
+DdiE/C/5qkt5UTCBiZRf9T6HC+EH6XEGPguF/RjMaWIaDDzr1H76i+8cJ+LK68ZbQ7WaNs397fy
tVB42xyEAKliQJcIoH2e4TyDhYJ2fwM28YoUc/PypyLAHXsE7ezZAagNLKk8dmqgroiOA/YfQTHW
v1KwARbVC6G8sIuVBTSGos4LscBfbS40ZGvocXGaLdrYQLSSPQiHNu7e8JOaVzoNdEkvCurVYJwd
Hg47l5WTcJOpO2BoPLvMhQ/K0/IHtITgCOYKVBOQrhpBTg5EaT1wpdFvX6iDJINjLB5OZixYGxfe
zRYy1LPSgW2OzTMe1Yiku516jj1XnOJ041NrmU2zsE3bzNkuwxLaEqPm1lkoIsVpvqjjdL5hBUdP
9S9pbqqCEd+Q0G54XoSRpbOTh/4GBAG0d33WB7BOuegxYv0K/t19EEjC+34i5lvik6G2B+nTCma1
9uJ/Y074dDCk17KjoTERBaNvgdcGPFeuDe2g5sJtuYeVlsX5Vs5T0vqSw/pROk5ghLNb2IEcye9F
uw7y/omZAQCtxNAI39mvQNnUaUWwZ1EcDpvmUoFbHxU8Mu8/74vaQCKC6PN2UCKSWfPn8IqYSeZx
sa5q1lPfg3JybfQQ0ajY1fH3KydZYcAOCYzAUZoemPVFUkd8CqbqQPfkxA4+vUU0jeWMlkdV5nT3
n/DkVRmEpf1El/+NARFX5nnefjuWrID3HRQZx7nIuNFr3XCW2ZE1xA/XXp6IxGG0eQL8aBUCCWqc
KDUm5j2RsotZxg/T00Hds9dIKpzF0XtBZJSjPueIxnzsGGCoY3z4HDo4A3kv8J74FfbPE9sbFDYD
mFsfLGZ0ixUrvdLdn1614f3lHBZXEpekg8JBfq92D0ss3EpGSBfxO4hdXv0G3tScKGOAiprGgzUx
vN7u/fsinHgrhNv5n/cbhf9wyLYqkOcaWIKotcXx8NTw1vlDKdDWUcrHwPg3jB71kV47CRnha84R
6iNs3L9zL1rztp6YyO7meQEpDe5MPO8pJ+84yx8z669axNOLVtAYN0dAfYX7zjCvEdYVS2UcZton
xlKKzOkoDeTDtHCMG6HSw+cmd+BcZTDmL+tRCImKxtrvJjYlLRdYJY/t0IB/EtE+lO3lD+YcEs+t
td7qToG8M3rVsGdX1VvAvOupVjcogwwbruomEdLgnYd9r9FoTTVkIPZOJmSO/trwvX1ZGHFDbR+h
MxgUYL8T97VgF+ARht7u2ToEXW8yoAhwvdmtmdMTU5w6g4/BNwkqds+FyXzktFWYEmIBfFYkuLuq
gdQSWfAaCQtNujldn2PFpz0exeOp4ECX8W89m4EbICUUeLMQMuHUR4GVJFsqKKOCZNHwJPTA6Th8
9GsLdD2ilAu3jKf+5xwNXmGH99RHqtVABk62uyFiCX4EdIgeFuaKsIe0QV2Np69tnOG5xKsmfilw
hjESRuTzNbElJ/+B42HWeTDDRlEYOfCygjsOyvTBhYemc17cK5bRTmWKa4jAjLa+Q+Z4ODudMlQG
gjpgAGSGeP8E8d0BwTkYT6VJCrAvVbdkp8+puddEmMuJKkTsMNsYWYKt/nkLMi4NVpze1LQeCnqK
AEGrG4LNYD0cN9CsdfIAws0CyeY4MH0sPaVmFYVYBkiIZ5QcdcnVykFUoTjz98QCJrii7zxeAMNb
KKOCRNFevwe/ZkLYrzEwQB/udh38A8nhbtdcgYLRDyrzlMCkUL88nTFl9Ikj2qjlmFpV71HOY30K
sSDQ+tOEJh/K6YFAZSedCL/j3XO8sKZkqPAHObisNOwH5tQ+4GYHVxWsLHCO76YztpXZSEr9MISD
KFGaoSavbYoz/ZTRi5CekZd/b1i/6Cg0/EUHw3cwJMJkgrbuBnAUk/Cs65C/u2iLD6rvD3nSm8RP
Ek9hfpb7x1tv0a/PQBPGW/SZchGZJJWXdx2bLHcnB+7sdkFvYx52h5YBWHWI5tqjn8zmK4VkIV5X
XvqG2l6G5xqqMyz60LrMhywVs8UDAGCKQ8tfcWKqzMC23ZAq04GXO9K2xa23Ect9gQWqlLGbFT3d
33R95nFhIp5u7Fwgu3kSIweB5pyEtYjrkFznZLN9vSojwbP7TwXAJwIKyVquCYh0y/C+3i3tWnqM
vzWc25D/LdcVfA7wC3wYn9MpvH6NmapbZYq0oqCmoE7LCPjffrpKaru5daQNOXQRFWCNgfHklQSd
VlYm3sFBoOm3Hq84sp5DyDYlO0QBHVcHmAZF6bx9cuJ0eL2qwn2jQWqZLiL9s+bvjmUMPpsVZo+U
hHifPA0KT4ktwAAJ7OkdlwIzysmTfeBMirDD3tZkA5WDX8eh9NWcju4lVG4awXqhuv9AxQ2ljHZd
0mJxK4YySvINThMxUfENIH+CkIaumuADC3yYoMnyI7L26MA08eKsU8BL1BHZsULsJEVuEAcPyj5Z
hNbwbqrr2HIJTpCBD76Csu4e1OHrScm+FzRBU+PEBkEsj9xUuSAOYgGDSeZJ47KBBNxhPB8gqd0a
LsOA8zqxzfV773PZk2z4F26Wj2GuH163CMF1gAUHWMoVUi2hSWBtSlIJgswqQM286UAcyFCWDAe+
BRqxcVfTeiqCRvf4k+2Fz93sW2EM9YQbeZAONdycN2fxlOcJbdVFiaxJu17XdZptbSrmhsTkR4Im
Zn8+CLzHaqJTqqsgd/0b+yd6yWayI7EKuukyl+p9/VJVq2IrIzKXDitV5FSdkMjySJEkGIq/utgz
FGP7WyWwmkWnzipSqzWAJnD5gX9hnOpjJXVBeWXjARvmVktI+7Mc6IOJ/UWz9eGBcZBcMLFyqa5R
2RCtL7bjPjMSrni4peV0qYGMncfNRvHqebT8Ibb0KCo+DHaq5xkyXqfRkSjLyXfeBWxa5XtJCOIU
9H/jEO6OWFfmFkocxNCm7KnXYe1LrVULpGmEWuE21wWBBA8X8wdohrTiUj2ToA2Z5hE4hEgz9EEL
NJAexpMVnUHRbsY1unQLckpa8QieYKYTpPcw4O2DhHeUFplVDFepVGn3vmlH+A9mJhGgpxVd3rUn
Vm9OhVUY3zS6kgmbZFgoLf2iRbBEu1bwB0Oh0t/nttUgGfFU2YWGvM/OK+lzyfNeboEdAEJdvd+8
CbI/Mc5qa1OqR7fAZIwXdrxyXyHsiAe19khDDht+EhFQnkVoKWDQBY4cealPSHcF3iHAEj64zdqf
RJouHMHFfNuBn5VILcHBOCK4ahPTfHxVd6UhdvLi4IcfX55qJqav0R4ZZtvCH0zqifbvhImEy28E
TKOonMW9yeUjsBxUAOUz9VnLynLIJJ0gsZjVxGxaX+/IVU4Q4+7TWvt8EvQC63vpFqS2Apgo54so
4Ga5OJq0we4H+9WdnRNyFihxwU8hyWjqqthPxbEOlIajvuFpCEoBnV//MQmC5Bh2KjCfBrqjllgt
N+TaPgHml1qxbsaVV3+512+DpogcEJP9mAzFRdgkfhgVBebwOjVdnQJ6oaJ/G5Qbra6x+ViD1Zx7
k6Ln7DplaTAEbWibq+BaK+bxgp/lOsor8X2/5ycGbUu82x3ZPeAfPM5m7WpctYKphKQtZB9CLnlA
F8R2ecUsymPoPP/3JOxbUPLuqwQg22yM+FDiXx89vgBR7K1fnKcFo/geEK5682h5V3jndBOlGahF
dZEU7VIS8Ul1I4rwVNiXEQdianTIrdC6WX6+LHmrhJktjEcjlFb2srHU262pI8skfcLg86Jhgla7
oE/cyWrzTsoh1c0q5ukIOSSLRtu2S1gsOtk1So75x5813FzUwVMi/FQ6sHHJHmc9xzPrDFrrZ/CR
Q2lAFdFnj2zCxC2ualsZ1Yt4Qu2R9HcAwv2iYFc5WUQDeqmN1LMG9SnMCVBBuSxMPkO6mrf/O6ls
ygGErTsVQrb4Vt6jNUQkUbMkmUh0Rdo4WRpwqO3EOUkTYbmchoPBtro1S+3ovkuFJgUddCGG9p86
1jccVM+nQyqG52E57bF6b8/Nu/A5zTaUREk5CD/Untxbawk6aPuqi3njVncjmHzi6oU8vHWDAaZn
LYzRJ/NET9KvM7qYfYdQmdChaA7WPXM5yh5bHvRIMMwOoVAs5yb5qyDtF9W29uoo3CmyBcA/PHVz
rJ0ylV4UxwjPwEKKdTbzzENgjgjTlqUpqnsxBb1/o5uCQVBrATwoOT4v9uCzmeJCHk2mByVG1gcd
FVgI9XXG/2rObzSPETlWDnWWb9N09tLi8SKfYqDZdTjwCAlTU6/dMuEOXnl213/2AmTZv3ryuMyw
h0u53BJpa5f+3G8rhKRaKnduuq0CQnnUA+/3793F72/7HTMyvmhdIWYJKwhAjyjZlcnHzxOINE9h
wjND61+daJf7oQCbCn+UtPFBMVY2AjzWB/wZ4s8WFt/R3Nj+oiN9SnPZhVP/CcTHgioniFJ2GI0h
/wWV920oDs+2eIuKaPmcZH3GiZynZT/3gYRDoe2cO9Bp4HQ1kp3Z0afF+yoBs4SggkqRvQSC5LLD
RnNAldXY4tn19UiXjUBnGPLcvgUgQFQyW5FIWdloNscrG+tFjJoYNNWuh0H7tFE/fZ0A1jgzwNke
OoYIYuoQV3W+AfhHFaAqE3t+IuW3GCh+fxavWRMqtBtluG5mcJO0kDzoJVZee2D94afk/K+1eTU+
QtMUjwAmwly3XZPvJ3VSXGSEHq4EVRudW0HYh6hWtNrpjA72ZJ/FQiAsOLfItZEnLD8Gp22iwXs6
eapoRezq4cvqwktz+10mj7sRyS98zg0Ee+t/ADQrabb1Czq3Jd5dUyuogQSlkrrqgzzmcHdf4C5H
QQ2zs4vOD/ZHkuiGMiUW2/LRbYgfIot+CW1G7gckLsmWWN3/4fbwyhvEXBFy6eb/4NL50bYtJORf
gV3WFhfDzhOI523ezAP2lWglSSZSzUV/9Mdin6CzmlWty7UUqrlRlBX0IDYtCcmCS0DvbWD15EaP
9JaokeQJWRblaP7mzrBWAbwQSOjc3vm+NOYIWvaeAnPkAqFChL7vWaVZjtFgTNqm7EV+Mh5zJtrZ
jES+xEl6BAcW7HNxjzRZ2ivLiqN1uEvU4iUSoqAzgBxbiVJYjWOOnk4SibU45J1+EvflgIaVk7Vb
Iy6JTgm2vyoEJMQDV8v474kUCfztl5Rb+RFbhhDxlSXIepvxe8nelN2mj/6VY69DhPOnGQI826hO
0I5nkguOM3jkeuuEmMvOCFPg+6v+5/UJYTsrrfhOrZdPgHbLUwZhcGTGNZMkG/DrlFIdm+vPV/gL
QDG5db8q1jjitS58LIqdV4KG8ZoLrO0k5EKHEYu7hfwU6dLPh3LAnDj6LnGnskZQvJIJoS3tH5p5
zr/LrAsl2rvznSXSCPw22Qvej9Q6JScj50TnpBEPvHreBI0Vog7KRsTYkpHLnR6bX5FF7wA5g0gB
mMum0Mc+0x/Jln9kDsm2bSXz6AZeS7RhEpJG6nBY+Q76abMC6s9tlw1oqHIYYRU/GSbTB449+1/K
sYgc31dgz4nHxY2+/vgfpBncbZ8YjtRmaCjPVlXdekqRpM5tMlHL96DSV5vjHWGHlF51qluQuIG3
05L8bdX8O31O+j6qwvkDqkPnROdbUdAcY3ltFCjdieyZO6v8jW/M+hVvA9i9OenTH0jUKiS0Ic36
fuXSTNM21hec5gALsCtJzUALsYZVGos8SCZ1ANda4PZGgf4Q35zBIaG7VVyUk4YNAqqv05+aqeG5
bTy/JV0cGRJVl68fWSDuhSZKTAb8bST4Uj0ybG++bUrT86pxYi21SQkQ5P5HQyy8K1S8453pWPc5
QaKVgpx6xnmYA7vI5KyhwRtysOJdQcomGs9hZebhpd0g+4DmRAJW4QUBdy8lMIbd/UNt8Yoni2rS
EgL6uvjaYydC7YJCwzbN1DqjeNDnFlJdsLqRSE4CtQcCyDm9GR2hYjTiqN4G6uvMY7RPiBI74XAq
3f1H3a2yH8s+XPqtu3POvLKnJqJ/DanTUZTGMdWF/F7FPwd7EXqfk1OVzqxn2Ms0VA47+prv6wiF
wRBx5rA2Sf4G9n4K/MBl89c5193Lyia7LE8OgNDHOvZqFoUgQS95D9dsn0kZl+lDozsSbqO8OW6n
N11AthXb7/o4qcYX+QWj7ATjfgUWehCAjI4Lb2kShrZ3TgWJ2UIiWKYxxAfhr7p5nPCN3alei/T9
0DS5DVAfX2YcekXLxEeq9qIb6u2CZUeQIrHLVzO+syHHW7rFD36UavzFLRN9a7T+ttUK+ll3p2Ng
Of+T5APvcEfGrTqxZiEdGi73Ex+OZ5d3L7HX9XM6jCg5yLZcPOz2Uoq5iBy4a6R4E3V6Vwyv721G
3Spt/mnxcuhKrGhHOZQ9vWbDQSApIBZMZzzLxHk21TUdO5o+FRkqfkYX0qVHdIVkowX3XG9VrgsK
FEpce948SptF7dhA+InIbWBOOxROQREYdCyiq0X9U6fHSYIFvLP1CS+02NCOASjfgCM2YrW8CsVJ
Nep23e/iQG2mb5sSImS4CIMlgqeY7nHjyczeuoOVdoh4GtXDo34o/hUa71zG/0DHlr/7/RTyhEpR
via/MxwvBdV67aDcX1Xdd1Nzih2qdF/GwuFcVhev1dlgHBPwkq2nglxB7DTNPwsULpgmzKNGNFlN
ZgLmaFw+ct5cYTzF7IpghWI3VPbtsFQyck+/INXXb2iCvY4EvRm78m63EUY9eo6Kk7HLa4CPMU/H
hwzUa4+CLa+WhGHhjw/a2Ja/IeaqTND0ielWrCo0tnfuCMCrQKqr7rfAmz0EQIjJ26z/Mr3lwu4e
iGVJEMW415jSLRZsp1q+Ca9iYrXJzl600jrvA1vrnWt5vef51ZXgD8BMaTCXkRIstOUo/LPXb1U3
or6uRhQZgQWf9rpmGFwlHEute8jmpG4gjl6uY3mNzjfodbKXhd6capj0UZiEeKzuRjiEsWH7H+n1
yoGMaa6bdaBoXwEejMzzCa96ya5V9pyQbvOH6Ntl3VVreek0HeDVEUaHNJ8yx9tSwzxLFyC+iAJC
OayjXuejcdva5u6Ql8iVEbcL+WCU592JvQYPq1KGmq/CLxAqKCSoMFqo8pe+C7oXuy1GX6guQGg7
XwzuZ5YWdKf3zNiD8OPMnDxwY2aIi0RRoigd/ZqK2oR3RzTxS4hBgYsOMvNtublfUU/CQbYr107/
50+Lp8UkviZgH7+CwhUxGSgndg9PbEtxtJ5tPY3u9TRQT3iLdkIcp/8wAKxC5pAC1tdqJSTjBXa7
/dvo3bKwCgYy+ZgtbeYsVH3BvzyDVnb3JMO6m+4j4DL9TOq7nRwAfAu6U+SZX1aLjIJ/OK7vlPa7
HcLACQByMdsjaH5W1WC0FYeOKWlYR4vg7V014BMIhwKL4fTrhE0vVpB/wPDSgHWUBAQJmfKgQq1C
RfHUUCPiFS++JLsk7p89fST3JMHl80AtavHKzTEWmGHLSn0haC9xOTRTBUMKbFhq+kqxTL6Hsye6
9CND/7BeetzMW0ZlH0I5MkTosXlvL25R7huxvHSSfWWy5OnTgrCD7wy1cNe5Ny6cBctSj0S9bMdx
v6BbeInojRFu2XCfX2LVr17oehwO8VqmXf/TjZe9mXou7fTIQu1qMToQAQJxHffAs9HrCd4Zf0hk
VnskY5pl8hFlQwG07o1xB72E+LM5F+7bj77IOPxla8fvY5r9x+Gr0/md+S4gnIALkKFCKH5GRtq3
0ims3/HbDxGu1A+APtdzNGZ0pk3vRvybhIIuq/bkvg7PnBvRapKZMan+rPHtx6PdvTqNN9oRLRJd
3JKxh3n2q4+LovKh01loBUZV3vDrFlJwdvvv6ytDSS1v0C4hVi+GCJguaEEbYg467k3jrYJYyLt+
StZ011ulVGgRXi/Owr3q+a8GxVNAsI4OdjBJls4xpkrVfRZjCnJaaatOmAjoeigFtM/VZUQHuDqN
FLyNXo5wpzcQn/02RZtcXybVXebp8naCVUXzSsOROXfVrIIUBx3NIBxl9o/DNVoeTM/lXWQN/pn0
b736dtrm37weB8JkHA7dFBs5tSJK7M4Hl4aEVWEAyyfNobHZfBW5n5UtqnIdbprbB8mThxxPZhtZ
yr8uZYlqf9p9tWzxxELCemAok5UFkQ33LY7/d6Gm2p1inHuwy2ZFq2bQKTsHqaCORv0jQr1KX572
vl9yk2Kh5g9V7qCCsEU6Il8i7rfDHRVjcRTUhVeVeWKYPoyaMHHLWwOg1EXAVDdcHd4ri5eR+qL7
p9nrMgwffP40mQ9sLq7GybnDkpshQyv5pgNolGxIE3eNqqmSJBVbX21nJ1umPw7wcFwEJ+6tH3wu
IFoqiO8/2myX7VsY5xVfM+Zad0LiDpV5ajk/Ol22VqutGEqPYVJSah9lUTq9ZvxbgV3I8lRtFa7l
+mMcYUipjLjzocrvA5SE8XiO9NVUKBzWnNNsr9p2ObrNL6MJ7MjopmOoIclkxOSkw0f1/VK1yhFT
3bOhTJXP9+D/lO/AREiwEqqSyKKSDx0uJYSM0YfoRS2FdkeRLMSUVWWVHbIKZPIEGjWMeaR7Wc29
uaJSYqGD3+pGgKv8jUyQ+IIOei9qhKo0KfyL8GQPEwyYb4yk2DAD8A1aBdU1DYyCwBrR4wGVpKVt
opmMlDHAmBXrlhSIyD7maR8zWoGWRDdgbllNWAxamtF+fa3PotqLK7HiE2xnRLHr4NJon3OtINnp
EVjkOqzxxwLpDZoO2bdoo+lXaPozbjVFgW3DgEzYWX/n/vGON4tkFm6E2EZsmIzmfZrG4Ap9kPHG
UZYwy0eSuNIb8+Wrq+q8sVxjsTZq/zR8i/IpuiSGDhtzPxNJRPFj4WyGddFfqS/iybHBqvaxVFe4
9xoVTDFZkL/wIbdXxCtK16i50JFVzocvikOA4Ixlu4599934fDettpj+0hjEuMCRrfnZaoBJjpzY
xNw3rN0KDsFDuGkvFFYeuq5ByTnYwjj1Izr0wVRflm08SJcpq4DEfodfBRSNVGjkm/ckIOA+jJ+u
OqKjqZQgH7nph6y+JPCHneta2EcTJv5vFBMEiru7kZVdZYIlyhWwGyy9rZntJkgSN4RKwP+CiOES
Gv4UhRGk/JY+bkLzVB+lbcF/v712x1xhICCcjZsEpvnMHzDLTstBL5DWGg6Mj5ijLm7ySu51o1gd
VkUpNqRR03gGS2ZPHYOUH5dRG6Mj599H0KYAxE2/RpFiFxDfKPDlmFTS0g9XESaMf51Sep7lmxmB
uZPUIsfbqJrD/psEiNoLGovB/SIBywq0GZf5w7a4FdfJ+DbpIwdEsDDi8tL6Kr82xCO6x+SA0WGq
uOQ3AnEAkADJEbbV9JZAWeg4m+OJJ7CxL0K8uzh5nHHE/LNhsKtDVR+KylE8Q5Pf/neDgK+uSwP7
DdIMswOy/ADTDwfQPdisPSaSgGzf7yVFTnNXge7ChcEcKk5YKcSpUWNztIlZiVXKKRF3UvTUViFg
5mYfjiwUxpeKoMLJLtk59i/1mwNsnurBRmQ9TQ2rgLxiiDndSX1eYLvbI5QkwJwpHmeZ9g3XQP5D
mAFopqrIMc84QjTaNt1N5J9y2DhyAduJfumv2KluCDHemSOn5nbO7GBFv+bQvVfQd7805I3gK33m
PvYvaeGnYvxzIyxEoBqQcA1fq3qwb0qCYiumRVG7ZUtVyQpTGytL8TFziv/JRu4Bf7niNJyh5erx
KT09BEzQEiRvztN3/gRaQ57iHJNqA995bYHMtXJYiBT/4jBASBpeR3EKns/nKfo2JKEQtHaC2KRx
8zhpeFExDRSZWOEVRacykZoWrRz9unGD52MIcBp0vkpY4h2ncUQMBYRuB4UVRFIycNHmCytrhwjq
AxD8mBiES7mvn/+q64SOwXCj9olubm4EkQ4+NHSg8Y3pbiK/9lTHCiI/3imlTV8zzrPPdbDCtb1l
jp2ZroQiJu+6v48+na8hLNPNSpqJIVOzuf2zMjwegJGKfuyePHHJ+g5sD4MSl3VxQZE4xU7zSh4A
+sYn7QcO2oojFnqbbOnfhwk2S0Xzl32r9YxSpDbRHa4IJBt1FYYMSRMyg3XKxPtKZ1F0oyWasXLx
/sei67xLZuoIOawZLyAGC+x3BQOtLdb6UbrMcdV7W+EtSt85pU+Nl9wq5mjQaLRGbzq6IV8VHKgH
HTbrJBEivxGUhnQbH9O/aBNYWkvMlt3KPGAId3u6VEw8nVV8w8+YqfJ50BAQ+nJ7BXGUiVtlfX5p
8+d++cvBZ1O973buhUF4pYX4d5dFALxaBhmEe7aETLAZ1Zf1Pf6L6rm/GeaxvHflTvvjgQyWFEeY
cfgkFJkW8DTyGL9x5pYCwdShDKFcQcIuR+QMyzkt/3051AM/vCOsXsnZvwC9eqj7IHGmCJxgGfxx
OwLxWgERXAXcMpFVvSlC95Uytr+NWdCa4CFQTwFj/Kd/antxyZbcbfvWY+hYM3Fxypt7HXO2x2EE
9gGCM5hdT4x1GboIFqOXM/DSldlKelsE0m8aF0e+DqZZQT782lyID+RZxDs9TKwaCa1mO0Z7B5Sy
W7quCP/Lt+vf7+eL4h2zh4khcNz5usVkOUThElwOaVYMUUiM8op9qPjW1+rApuwu6NKm/M6KoNt0
8kddWsL7ZKrC+ApNrO2v5NfrFq/3Lb9g82c/rxI1E0L5bL5Fn0AbyJErGqO8I8G37ix1XI+/Eklh
v4ZLXA7BdSZf8Xra2g6X7T6OOCqi64WwAmuTPTrq7fsA0smn+qMBdE++6Rry5WIMIiwbdyhV0QlH
iwf+9Ezvg9O4j2gW9lOn3eNBW+JZuFZDLgulIDa633Q0SQM2CI39weN+tmJ9o+hq+D68QNXSSjcG
x6miQMHfTWc3ig9VUy8wIIa6nuVDRP6OD2XEz+pmkN5YuwP+Ye9qQ0TfucE3plHZ872L1gGsYk8H
fKDXd41iR1+/WPj1P9YUsexIpSk0T3aAkd8jph0eY40wGCdsgiAfjPCxOvkZi+yUBfMKRSmrI4C9
k3PRYmDGreCdCQ37V9RMmsHj+DMKk2i1iCr4Dp5BECdWpfnizwqON4E9UTizqZF9lqfKeoLueXDd
GbyNp93kaB5si9lBWbKynEOdn0YTTXsGtxEoQJ4Egkl6KHptNC3Cj8XNJuUdz/8vnr8KiAjnq2lT
loJVtbhhWJM8PR6kXiRpqW7HHcfz81GVLavnqsqfGW0cHN+uRf3iW6yyx+L7SV8ysGKC8OxQbl/Z
ilPukhdpmLsEp5GieNn+oClrtio8NTLBurDb4wie8o8pBwpUWHwz/0x7O9h4z+mPN2c5xL4CJS28
gL8phdDfwAktLjzj9vY4RwfmvBTGjOBTWwW+6qAESuAUNzTfkx+uWfNZCi3TD5lzLM/WNUKJzxie
o9DD57qJbRLqEglw9b5or/RNxoR9mAVyPk9X2+7bkvNqkXXOEcxxEgUxW+pMqWVcp4BVSebQngq4
xJ7Bhj1pwTJyig5JscVXV9NxS4RrwsnUf+U61n0xpWoSX3ux9e0lVTlQ4k7RS+5N1HWgkjKemICl
ePf5XXhCu9mHuEqv9ojWXn7VHOySRpQpI02Rd5fhYOmAyIaemwa2V1fpD3DEkptaA6YacxEEDFMp
4PqHWcj3dY6zHFxLZo9COyQT8HluT9F5csr1t5Ni0Z6Q+C5xhU9iFzhd6x1pr5p7s/oSVVEDRQ2Z
V2eaF7HRDGJdVYJ9fIv9E5UPd59WGTVP/Esn1LhFxqu/m59uc5LevxQjIQQBw0SGT8Mg1+KOJECr
rkvO/OCEkou4endUcQhI8K+ryzYcYtRsLMNb7Z97wZclyxKcZIOnM2rXkeqaapbM1C4LrsqnVrkQ
+M1hQFJ4DpxMTPT0C2xRIvzfUgnyjEXP47cXtfIDZOAK33dm9dJcDh8PQE/iiRfduQNBeK/p+hkF
U1Xb7zgKu3SNT82m6ufgljLTYuQSnDQGVeMZGxv62IRkxyu+s723+tgIpcaoUQdpgb2D3twk1XH8
woOIRmjHTEzQ4Sn/trftmNx105zdDTxd+nvtuPAgGG9v1Hs9lF67iCBuSzXmY+h5KJsMOUqIG2oU
+YFXXYdBEEF+HCP8o5+bsSUpA8Lt0bBFd6EA+J8lP12SbctPRRLup5WFMwL64BiAoHfkI46c5AQ3
Cz/hktbiiKJ42nRlI9VnPzrkEe0KYLdgNihsSAxqGOfxFJqSv1GiDvSaeP6b3gKxiOLX4CVX0BLs
HBiWQ1S07W9k2u6GFcT2CDIP3ACZ0e6NfztS5TufNDT2i25lnZnirEDBwdSBefNpEFwA1hi/9oMp
In/JKYrAOtuo/YjjY1THYS8nDk6C20bLXH5S+rQevmAY+YIJgkd1rRlwDRVf095UULg3EDbuvnh7
8XAtNm2F6bG5AMCioQ71S9+GUklFIcWrW3jL6W87Ur0CLDiJJV1o4KCN4xpBW4cWQwH7HkiFtVfy
qCYSAsu5c8lpWQ8cdldJRi9ymyKE+/U+s8KvhMDlB6hLqn2te1XbkNEVw3a0WqBFBgQkSQuFDFy8
zZ8qYUnZNp4XnaArGhcC7QZkHVRyAxlV1ZymWzym2urpwZqjUL1qq+4fF8xA1DUY0FkBefYrjPd/
MP6kGI4CLqqxZ+4jGiMVZwP4va1Z5M+E+nJx5n9Ex8MUERqr+YELlFoP+zHrTer5ps6Ei0/lTBXg
pxmZsayjG7IeWLEENnTN7o3FaWNZOR3dfuFcgbIOI41eHC3i4oKMeOgrW2bQvi4/YnFW+3kIiH+n
ctTbUTo2UU746YWVRPmsiUJGytl93cZ0GoR+0ZGzylWBI80rO6yNrE1s278rCDfKrK874koSqfYu
meCEG9vgZ7AUX0PLRyxqFO0MGIBLcsDrpS1HEnOsYbUma08Kjn5EeIE1AekW0TV/U7bbuceoOzV+
DBCn3/sAHNz/lmpePglsxpwrxB0VT+uDrIUgf+EGLu6dL/jhPeofx8VIHAHM9he8f1Omdfjcx5ll
i90AQtwHzqq1xFipP2EtF/udKurNgR4tw8qBqVVPnPdHsC3O2wsN7d/uOMogFbm4fAMx9Am/w0pD
vypQGJsmldGfWYmMkknJbAWYvf2ce4QOiJsdq4cC0zp3VFBjF3EDkfcmhjIWVyfs+KdUj4Ea0VvX
xoHB96PpdNUzv/8pnynHjT6vjKggl+b3TpdVV46Vqv7isSVgqnSn4bjmKktfACLPAwQD3hQeENnn
73Pbjz74+2DSt499KUFBHCCt5Yt/lf0TsaZXojaz9fhZ0ebZ4qiaXkJAaHFNhV7+1PsoMiaqQ2G2
T2Gc5/5K5aEygsgGCWMcEj3F6VjK/Zbmusj3CI2eg5hgBslcJys9OGmKV0iiOrnegbt/ZEBPiZeE
IeYy2ecAkFIMIOBqkq5jbY/VQOBqTPUEkAuq2WlGljrMuLl6M020T7iqEd8EQupoDGQsg2Ii8a9T
5pNVvdvlENUisJok0OrAwAZLcXts/jAQP6Zu12gLjLDkfAtYbnHr+5JBhOlkpPMuFdPCJ56OjTVO
DAmx7ZGvjxFo4rVs/gQy8vc/XhRKvo0IIE94yn1cqovEb0udUSUMAY953K9b7IUxlQ7BJdMog9hS
p4GKoY5VlgH4hcRc59tXmGg3NaFvom0er9kycOye/0eLUAYmtAtPHnqiEE7NPFR6CsO50b/jH8pZ
7m/q07rvEdrf+mg/JEP3k1RQ4hkTry3Kr0ay53OSY/Hsx4wrhLoXwVLlrT2BxztT0eHbNVVpdYkU
26dhii5320axoRaWQzM2Rn9HuXeno6m3lOjQ8lSCS9WMuOCRgIyi3VablRES8ZMG1jkK9TO9EJYR
nA5rT8wbY/Plqm2hDZMP/5LbczIxvufIfzRbA/lOVNTfyWoYCirL/vAzl1zFK8AvnhY0k+dLdrk6
k2HjbJHBGD/PD6/7bcv9hgWWAc/rRY8ZtyU8A2dvkbvHsU21aGb0IXTzKMoZS1nmYTtW5B1jE7Rv
T3M3NF11RMCF7jrOkqtV+w5g5FCvuHQlYgqgRvmyAUm4HckhWhfw9Y3pryjAtQewfVVsyLTN6Nj/
pq1tZyPFVhqZ5iEjDtw9V+zQCaLShSh8WnP+7ka3BSDtALSVCJg6DKHZyA1elLfLSqwJznAhI90w
3QDtyxGZik8Rac3OYvfEBhFYJwizXx5kVeLrH9kfo2eY75ntoH3hoD41bsauSVmxz29nD01/khu0
NVP52KHRFbYuIido2U92upDKnnJZTzzDjRUIwho1Fj4jj0AXWn5WVR79dj6KjAOoKDDdzUIqnsCL
D9UZncNk5g6dFcQTGHUSVcJFjexIPhDGioPw5YG3ASNllfvzhPzRNqC94vVhwqu8u+ElL6yiDrFQ
fl+9y7EWnLyzs41YgwwQPTqoYfV8jQqHCclm3M/BASxnLXDBw/zGm5VrI4SKxtvAiEvFfgpn234w
TxjZdyce135pJcoSkWxdKU7xe0bPXOxUzV5mcEwzXxOWG9iF8toCezKXr8v4kQGy1FIKVwoNzwj7
HzyAvq8Nt9p7MVz8u61CK9BMoLZzjkqIYG0NdDT/Qj6Wck/mruwcOZC5AKmX2PxAUQzsdZKRHhsE
XAusYdGqWD2Beyl3EoaS72bsiYgKBbJH+YxhGhCaP9OQ1cE1p7ishPuSkLWJjZagupUwg6miSoMQ
0tVrRR3IabG9tJWEXGLWqi052/Hbu9MnuwjifJrPBPe6s00tbs1BpYjA94tK9Zm1Un/FRQiPr3L3
mJq6MH7IQ37Pv2Y8Q55Eehmpddb9/PqmWzLLkljOxNYL7mtsknJO0cD+repJXjCn8xeYFa/ANdxg
o+A2ZrkSuyYrwaD1gTsEr4NErupPMo9pdZlW0v4S1ehCSpKYUYcqO6q24VDk7WB79uyMLI/atWEu
XqflSHsBaRyZrob3IUWPtV0K79qmnlX1bUJ5tShh0IhjgyAXqmeyUDE/53ErEZ7qX01ZkLWBDchQ
q5F8YA6eMM9Aj9Fg6GjgW6ZMEL3Q/1HuZDMQEeWAPvNDPk4XxyAo8qYm8Wg06/9oDuWF0McvHRfG
eM54s7mI0jzps0lVAnoiO0FG09F72nP77enZb0eOpiZltV/c7y/s/fq7uX22ujwXMZ1RX9aLfboP
D6cVnm7OzMg3XCWICzwHtbIHgDN4Nn50PjIBAxJrGDKfWIeAojucCkSnmYIAlMhXImzH/Ibqueam
3k7+lZI+TJoyEqzEADT2YCLJGFbVkeW7vRnRjV/Hnq/2sQi409z4A/LIOr2nzVmQuWIRnRNYMsbS
pMAKRRK8Q7GCxAe6EOAAOt8LHcNpVxCyfn/meSSR2F1UXBVtN8RVpVznaTPWKJ6FFIHa3wwzTYUq
I78jhppgobIq0/21+Lvtk5aZ8Njrh9iuD9OeI7Td6LZq6fpItyBwVkld+TyBd1GfuzcZse+8GMNS
UB2v3ZQ0jfIearqrxDuHB1I0Pc0w4yHFzUOKKg9HxKUmpN/qN3QXjkcLnr8tKLSqKeq2OxOe2U/l
3fRixWdccyV3McDCb9zkrcPTkjGbrSsykfpazV6id3sQ+mn2iS1bHnEVhieug4mplBK/zuPfc+5f
yd9+bJeqo23kusOvDhz3ZeDFzTnM8fcrVQSPqf0W3Jh9jNB86Sqy+vjXqf5XK23oOdRR35NtT/9j
+q4kV8LH3SIfJwZ9n0GocDhnzMnlCYSMtairxWoVBWBc6MFRQ86Hfr/UXqbxi+Ip86HFmLtXdopD
9vCwMi+EWZUt3MSZllYVTt1jHRwq8WQx3WVrn7e929fFX/vP7++4BghgfdA0i9ac9RGqgM3mgnmx
FO38RaJ6S8yWCNVwWoaqHQq/50uMQ1g2TNwFTm2Tm+o6H7m4kzqiH7I6kURXMFAmJT/TBj26Q7l/
Uk5MI6ILEYnwg6rex3uNAzvvVzhJAYmvzF8pN+rDFw9koXNCB1QWDuKWCyCsu4ITJrUUP3QuALWr
2neFz7CeqlHSjJV1M1CL5CC0Tj568bgXvmay7LH06k59G2RaycIuLe03Mnkif30mKL8g2qm2JNAT
Iqj01IDHBi62W+bS3tGyX4Dd0psA3d1lsx6O8wh4z1C5W4l6F0G+6a9bo04kcAAiNkviDOjAcKZq
H1uugo3cFE543UUocIy2BAQw47M1xT1/IdEJpdatCnRVeGnduxg2+GOVK17ezfmhkFqYHqyivZG0
fMOuCrteQvlDM8hyNmr6KqVX9wSNQJUNPNrR2pWOTN38fmte4Vvop2QUBBOzcTohAT3sNYVUyCyv
SeZnbAvLz/w4Gw6PSSIeG4uZt8SvKCBp/tj6H9+zzX0hRlZ6mbOx2HS7MVCP0Cv/zBX18ikQuU7o
3Uejd35CggC4QUU5EZPYCiq+YIZJ8weIzNJl690o8AHAT9gOL/Z6MxX9ZYUZh8pFyhEqT6103VSs
QLnO5hRlJf9DKygeJ3aQFaOEB/dlRDQfWpvZ8HV2w1zNr0T5o6rBzVW9TBSnJXgSaNWlrlgCKpJY
CYoE+kXcGVgSDC/kTLVPobGkJzoxl030ExGsZ8RNRuKVaeqE6vfQdsffPYD1t0m2kNxONDO+FEik
utgrfdtPLIBdaA3zhw6ar9umtII2+fG2pUOYGPeB77tZCdpnpav34KbScEPodB9zOJ5a16QBUwWS
xN+7/hRJpS1vU2wea9S0KtRUiCcMvsJU0Pv6S1IMeSFKaJv6S5etClPE9SbdV8VGSucVHXJyNUG5
YvVHv5ozljDKqqIDAVM2NhUpj8gsL20WbyIeQSYvobKjCdiDm8mPNLmgGdCjBTA2KlAM6hlGKd2g
YxmYpBb4441AznHiVUkXKAlrBZi1TlTQbVGHMjaezNzIG0AXPB8XagK97XTf7KV1skqIdGSBibXS
TIEojcIMkrnKYEoomTTLZbyR2TwEN3K39vbbVmxqEBm+RzbeZS5PT8jybWSKE7kPAiwYYdDP8Kiv
3PtL9iiGUZBQrhJS0XDgf4hOFwoSW9sOE5R5Un0tWSelK/XYS5pt+e9CfXkLrOrxrolZgZHNPJ2Z
jG/u80qtVEvSNdhMuStCh32t9s2qzLXjoVno637vbMKJmb+nRA4ZxJI1FsIkJHV9wd3IO0sTS0aT
S/H3hTwfNleuE94r1nVyUo/WSrbWegw5bwQDtv8Ahvnzyq09Wyy4NvLdaErFiwJoBqiWK0hledqc
y0wlflsA95uDMi6jjPxmK/rFULLLA/iZFlztqj8By0NgCZIKu+r0OjDpl0W5kUAxv/wvjIE6Hcsy
C7IFt3u/OzrFizj8UcbY18igffc1HTja2NSOuDlO7kGbaWbPS/mpjgVBev23XW4HnQFdKgiaIxwf
3yqbQR5HJSJPd1kInYUxW5hyJtNQf22jHt9P9sYCqW3ciAKMIAcZN9TCdn8hYMuHk/CWhCaK+Y2D
uIuTE6/UsAkeIxoRQ+AR/e8eIBc9uVK5u4MrO4qLFvuvWqr9xfvbW+wBN7DpUE1xGFYwNB/O8fnq
/z/OisODtpPx8lpc+E6k5QiQtSetrJFHtXsPEiGORbcHtM3PlIHXvmLIbxNR3viNuR+A6mlOneSA
qlmtvUyNx95hGYsAt1WtG7tJUp7vvAytbDZOQ60mdzl+46FtD1F8YeLjtt3pDKbj8SjSl31vOG0l
6j5vK/4ya5pCLfgSWbt1AQ1X4R4fHCuPr/OKDUCkh3xCl17M+tiDP6NsRMVljrOxKj+vVAQzxdwa
uFjUYyCfKmnX803f+hyMD+c03uZD7XrlNb4e/jAg7GGQu8gfdJxuCg4Xy2gBN/qm4JxXBdyGFNE2
4TzpHj6HHLZg3pGChBFepadniImNO3EetYdh0NHfuhYqU6gpSlWQX/pfyz7JaP/5iOlpkectJDpS
9yUXduzGNtl1Fpcr5kwB12Jgz3uwhIcJ6gyFfzM/LLFUHgaP90/s/GYLk3Ung4yma4gdvr8KJONU
g131efzVeQalBhnXKRB22zs1k5MJYuDhbmTfq65yDrI6HMC6Aiw2ov1YtshOf/IF0LeeRTovNLii
givaQ7BfkGwjjDkdzFiArDyMb14nE2TZUSfheM6beOGMgyde6AQ3i+Cf4deYteqdYa/pzPYiNji4
6DBL6pJuPu/sNtO6ge+bDUVboak+/4xLOwiimuWy+k1v5IR1AzZSQ+FIi7NWV62nPS8BozqjmzfT
WGiUEJWNsFDlqJh4lNB8j95ayxy3EFsBKyf0J4JkDXBi0W8oZkvcZdKiEn+aQ7oji719t0m8ywlY
yvzQbP2ZcDx48icvki1ir0O/6eOzSBhkKxJdWEsw68tvIYCyTWKnqZAi3CyxSbUT2hburvvvLjRY
jvV2Ux3Xy31g/YpAFzay440f3q1cXOZ7jU+/CuEETgSOyE8ZndmVkQpGe5gQl3zRiALF4WV7OUi4
fyIwNH+/zt5I/sW0bgJZzqT2zdUJBi0DVG24+lHQ383buS91Vq96XMTTSFVt2PXSfNESCazajQ31
1K46amhKJOeUDP7Utayp8+x61XGgtyI5ZLskcR36sMSzBu7W2rqAoB8RktYuVxlImhwDkqAtdITM
l+D27q4n23uzz8yIHdPI7vvwFgzB15y0Zn9Klhearm7pV7ngZufTtQ/fSuptRmQ+r+nqnJTubdkD
yoJ5azZqkXu/5nLactwOHRWhDhjkkqcqdN6rrwxLxt0ukguysopkj7o6i/8Jk7jzjSSvRN8o6oN8
2B/Tk14vqdeacT9eBZUXfG2msEYchli54sxR0l24/zI0IiSf3PlnHR838cGCNh2rckfXbxjozX01
JvW1V8pKa/CwDuLA/zeNywIX500N95QH+WA8QTf3dVmPAgTRINwdNFH1h9FjpMW3pYEXZ48yKdH/
AmalxBAT6xXUZWsq6OVlBjqU7vJACaWsaL/gpzlCIK9cN4f2HpkrD6/kq6feO62OX5iZ+zOnCXrR
/Wem9L2B888aBv2PCVBM72iGMCXe3L2cYYXFPvAbnScyADWoyJ+y7IJ4AdwzqzH8VdXOXWjQxlJn
z28wj8Q3oHca2j7ZI4clhkUdLwrbEOb1sjhKIyP/ym6dz5XSZWW7ySIlScbHHGhtKHhLnko7JjfE
80quy5IP65lYbw7LICc22vSWhGgKYKqZMIa3ml+vyKr/oUCZEQKX9gDcrz+TQq5mZ7C6b53dGqmu
YRO9XkCv1SbTGkBBfFyKu+l3fy0uepslfPUMHdnTUK3KBqZWm/yqdeqwg517sNFvQR+/cL8ATJCP
Muq6rr4sabMB6Me5XltVo2oYBCckTWt1S8V/2C/x9eZH0NEufwSVhJDvyCf0mWwL5CFpqFx7TvMV
5MzkJ1fb5bAev491n4KVcxRv+EM9qUcsvvL8g6xlfXBzRmx5DYKc0oL+WEuQKgeD06No1jgnSEUm
yBNhVruTT209033WlP+zQrrjWmD9KYSQthp3UOSheBvxdEwY2Lwfaf3guAMtITCUUpzeQbo2vAmz
H9REUCse8BTHchQKK+TeJC115Ajpk52I5dujrrgKhEDSf60hHaBehzr2gmcfqZwDzQFNLpcF/XyP
XB0YhoFJROSDVDOk/whJ6zzCcj1FXU3xGDZjknDTLY6DQSDOVzhRhCV5UZ7lq5u9K7f0HDDz7lUS
1VaZHjDw8541e0eO7QYoZfmhdtFuc/whwtukE+m9AwphGi7oTbrtO5lMu7I3yCQmPerhQr8h+xVQ
ZAK14Eq2nCTTpdfYPvJVbwDEibEG2IuapcJXbcTYcde6JOZec49cRFsZt5wHsTPPh6bxKvIqMtyu
WVPqZ0cq+kl1ZL+/T17O94MZNj/6D6jx32dAoznF/3PmZ9RXP+yinQtg9GVzwEg9jhYmjRqHi4VN
iZveu1CnZkGxnjYVKwGmFgOeC/vNg+45csKZSU+e9uO/E25asyW7GDgQOpTRXeasgyAerkZaBW6B
EquRnBToDbLULI+ucHUj7LIwUuoiS9ieBsdVInGliHnMjGmxTkVGbYaQH0eYnxnrg0TubwLCMfbl
WvPKuS9FfKznqmbmmtIGXEkDOmzNPthuCokli+FMEgt6ZeQoRWF1wgrUqSu/yluOPr83oYaI0659
cTfWFwyRqvRRl8kGmo2V4CHLPpVJtVH6BREUyH1T8jEDDZAPsJV/u8NAc7s3HyXKQKPTxSbX2gwi
mbQ3+mYqj1C6Fqmg3/3qrEUwovHndo7S7z4Ei/OTJVoh0wjE6Ovf3PtNryQYRVNiOaXEDiUwWiyf
HLLEXVzRt7MaGGl8Uul06rzirkkkgJXiE8fAMDAJHi4NcR33tWGID5YzwoCykU9vymZ3ra0+qMG8
NMQ0tTEsoJAWJGktbAbT/Jk4kdNYM3Xw/ntAl3i9gKaoxKKBFhlc5+fZAY3JgfJeFxl7E+KRV5ea
idk87Ed1yEyRXWnSBguxBmZOwp8n5YRqvNRwgoGL2Svi07uJsR+oaS7C7bAbcQd70T6Vtp+raH59
Suu7pw4wHTc0VEP0hmUTWG9MRy5mi4/KPFeXKB0WkBOXowXJnBxf8IZBZzeO5WM4K+fbniNBiyHh
dJP875E8TAeNkOVMzKZ+xpgUsTmwqRwu3UveH9cN5TY9UQa28aA8Pwt4unP04cpcObxnrUc6VVYM
6UaXAIugiLXihdIXxh6peTturvEam+E/B8sQQRWfOra2qiHzPWycuGOhSboImoTEiU+EMEtdnNnK
nKCN+Kk2qrcGaaTTHNk41qnl1y/t/doMuz92TbpTu3VcKrgwto0ir8Phf6aHuzPagTZsz8g2QlV5
/0GshNiP0uG83/WyrMvL2PbJIVeu9t97ePsrcvuKLaBwpcNZCGes94rmvNQ9fWyz6ZCNmTwQAlgQ
qagHxWgg3ggNeJFHleAnWfXjOJHpjgClxtrJkxwm/wA3ehIkI2nwtikbSQwcJyUUrUk6r06FRaht
EGM6hOmq5SjOaAaH23frtF7o9kry7rY0I+C41LqIOvFV0ZZLIJHcLp2qoRCuW4YSD7KRHwSZbNp2
Y29cICNURs/9lGvez8Adk5t27klwr5Ti2OtEwQEUmNgCbTMTo9zCXtN9xPSzNI5CNbNifsdB77a6
W6YxP9IxrW08av0g/TXY0F9HiqxeooMIpkUzXnGbu+/FkuGM4GwpSN2UtsuQTy/PqYMop/7kfVFt
CDL9VA5CwGp73Va3j/sEnKpeTZm2vOov2oBGk5dS3NiSN4f3YZ86f1DKO9l+vQ7vQiCW6RtKUE2e
8eIs3PHjrwGj4zUL9+h8gU28y0fTrCfHUmREJHbsqhx9dNhnGVbuOxz9hq40FdHwNSk/hpQHnudd
Vvn46XIE2rXqBa58+jts8xDGdonBK+08WuoBEjfr7bcdNgzd2McZEh9VLLypELuiejZzJsNW/cRM
FH9/jK8EEKfrsql+zl9Ypn8PR5xQLf1dPqO16Cx+9QdRIilStIv9OxTooz/4rAyq7ytcmVjsz8dF
2Irt95UNcZr1EQ+V2WyrW8zcPJYa/1bemBNm+132J/WwUjUwbnS9tJnIkLoi0cNzzQciEmUMK7AS
ceGp0oUYSGGneTwSN4EOO8yVKXQGyzP+C5zpgcgF838TTiBpN2qXCCCc/dPidqtfjJxGYUlC24UF
vlO4Ypms9NBoRuVQnbuKk08iYSq1N/lwK95joSiJrSv90IKUfzxP7UzssOdP8vAmEqAhlaicV1uh
CDTJi58DTC3hwVY3zprgTL9IKqz4SvkQ6jCJ6M4MV8my2p2W+PLq7nzSUCHb8MhoyvBWgvf8AHrM
v2PslaAnzLN5Wt/CwD3wHt8HNBZ8Th7IhG1toynM2m15fQJ9wOEB6bN9K/pNZFYAfo1CLklfEpCl
mRunjy/IXlxMOEm1HKFMUwUiMQ+PGrJEko7FyiVT2ePoQgMZo+OgcQPLDE3MoQLYSHyhR3ZK79bG
yXl5tCN5wLP54WHEoGZyWJx+Etf+SUzXWdA2em2EZ0TFKqD4z29maFSZPVAsCYdqGJ2xFnVGsYk3
LA0/Bt5cIvvOct1UMakoZ+H24fcMMUUIAgAbveG2IXFERIunb5/lPUzQ4EQmX3lOZQ3hHAjfgziJ
b4+UuHeGUuFjlvzMN9oG+t1+hKL90/kTiKCn9Ina0NCIGP77DVcJOMJV1cy8OsxQX4iUgk1pX5Ec
ZvD4MGii7s+dybEtiBNGAatApENCV5DRp5a/bLaFYUIXOA1vzMjpcL9vuQbpEm/6q7QzUJEMSW8b
xHiPDdiREkaIqeSYoGgzqBVTiFiagl3+nvLX/A/o2ij2odvLvvrqr7ORGJYuKfSAYjpzJbECnz1D
S2J2WpVUL35s0N0/COo3ecCaOsBHAXGeT4L82pJLpJVhgxAomeAjhwhKJA1ML+WqTsLgIL5IXj1q
LgBMT1TcD4UZMDfNhfhNY/xdhw9yNnnuvrO5MSxdcHplhCXGrZNNOFjrHVpFwrEXJy0+Z1gVTtU3
8wL9f96XBawhjpmMU2PpJnngeoIjm9zrnwYGtxV0l3QpedP8K9hjRBaqvo1UuWoFPIzizOeJPYqi
wI528s1kjqIsaCH6HKzIg0mTOfP8woEFAMhmWvoLxM0zVXSXKzC8El8AtipbMqdTaxAqQusHnp8G
oO27aH0J2g34MYY7UXAcTMkQ+dylnPczuy/2mvwG3Qq9GEUhdArfoFHUcQMjX1T3dLm7bDg1lAil
ahPiccU1eXdqON+A6thjgMA31KFTImeRso44xApGXgsLXfeqdsqs0IJQgiWlO7CozJFPWuSnnRE2
RV9wseugPY9VDKuBecWeF62u66QlB7LbyOiqBFXYDdy3va5FRDD5s2eYS3Z3iCrMr5XxHKGJ8onW
uo9pqyhbAIIJAnXpsLovumY4chGxdir9IJZcJWikrl6ATKeMjH31U2lK1ZUSS/xlTuBB6xfJ5z8V
6a4cB06AGqQGde+3Gbhz9g4jx08fb5ZJjnBd6qQ/L5U/gCEc8AfS2eYBvqQ50egOGxCMPHmTS8h6
CBlYChiLNSL6n1pr55IP62mMGfZHIfiThWfyq1Gxg3fa1aec9DUcmhlO8F3QR3SS0uYwP7OQxHjQ
RfshDTzFSLp3wzs+C8TBE+638Fw0FyxwTKMlcgAL190srsFjWDBnXzYZOSDur9L4KaUNzc73Arne
sZy02qXkHa3aHq/Mwdr50kHJzvLEAQMKfqHtt8S+yrSY4hEAvkoZ1iLI+X+D+fSLBUVR5nTXNls7
5xa8GsW7MQTkjqh6CxpUZLvXyLJFo2EcThzcLC2sosUuhfE6/6B6bDkQdwh+sOyFIywDqI2M9OUB
IIkteZ1y8lJt21whua3UOH1AUWojNdxeomThNuz5q+z//Eg8bNIIqbWtDXMN5C2OaHsPEe14Rsy8
DBTQDoyIu5yQVLTl3xDjv9GfEGyw7jCmfr7PoxS4XkQm8zMKFf96ghhaHrZSI9kjwVKdxlXeZJWV
fEHYwEeYnbSF2Tf1AGULOfnd27Wm49t5HL9ueTwdJ+hhIr9Dqf1TreBrBsEZXy8pzgu4qMbmPz3e
Ro68xBBCTwh0f1gjnyZC+D3fonwqz6k15OgCc/MIfgj8vVkcvqKelGO4Okn6dzmXAocPZmKfx8Ep
f2wrNyviMYSwPbYYdYkCJTGdSN4CWb064g4OxiJL/Np4Au+PdIlZJvag2nzHVKLkgTCi6PEaBTIL
oGgzZ41OxUWXqdJymBWmd5ECtyfIuYuBoUD3bAiJ2ASg1aq4/DligJIlsORicAbKwwK/Um/loTyz
mybJDmo00CgA8Tw6BbU/sEucjABWheVt4C3437vrN9W3as+adLkSdyfoN2X3iElQ2zCE2hBfVh4L
kbBknJs09i3aGmDiI+GShqXKT01jvmFRabeeHGX0UKFyjMAc5wHjxuRuxOp3+yeQWepsHP4TCqHn
DKoU7uAa4Ct4EZymihcm4JypHVFQoX7vha67urOaNiixoTNB3KAGRnGIWDTrGDUQkJ/1EAf2+Tb8
zTaii9yxVsxK/VX3UyvrnKYAdVgmPQcRNPLR0XQYxls4R4g05wBfvUQcI9QmvIGaxYvtAU1hYDF4
sQpJxJiMPnLwlHRbOyoknSyoChQFxrZdAEvdoLs8Rmgg/7wEH0qV5K03MZRj6+GKQ+AZIK8fAogf
0GSerFqh0ief4Vp8YKY4+g/VmwC5L/1O9tTDWbEZ+3e0QMAinKKa330zvtz2a0CWasGn98KYGx4R
9bZSKmweM+EBeAEkojWliIDUtYYQJISPMRtAchQC9kho67nZFSPXP8jUlHQJ076NFTDKzpM/3rT/
B1wXN5Iyrn1bYw2MzTrj+zE/v1MAR7VFMIDlsn8lIp6inNDyuvXgcs9EkEQf30L0jcH+IWjp9A2+
HiBpc9wk/3oRIHTWSN+iuBA7akT7yEPipBbgIOB1A+xpo5vBiEyT2p30eETCZaHrUV+FqHAW7Dba
99ArTfrWoBcXdnWdZtHJJN1JtMKRGtvM+A/7UUDZdzEQD8SjsONszqSCLujUA7b1CYnT9fHXkRim
U3nbYqVIb5pSNGeqIyMynujJLAPTAJ/cxPsc+AWQUTe4nRNly+eVb4BZWrDE4m1fITJUZgx48eK8
tU0Vgd1HZX096W2Gt5DchWUxEX+a8ZABV2fndC0knHRYv7sDD5X1ca5H5xyJj1ZQ3V5N3og2y96+
Ddy7OC+6lb83Cdog4b8YziZtgniJRx759BiuEnQ0IbSA2Kyl+NmTbciCiFxQjpY201c8CsKw7uW+
rem3+G11kG4ZS0GGzdqQRlMah8ErLgEuUq9qVkRzwlJuQJBkX3NwYQERW1C4XGneQoV1gea4pgBo
9DeAa/RyFgQp2ejqdWmW+wTUQ3Wg/43g889tWFFoTSIhPyUwc3xYlsfP5wFlHs9eOjZlWsXc1UaM
DaMIJlR+hhaAxWoVyJXjddQPjlUXbSfm62Qhe+/fztwxt9I1kgkJEmIp8P3XsOAPW2atugWLU9t4
C5B8SlPpV1iY8ydw0K/7WIDijPCGcVMTb6nSQFRkrIlo6nze+1cHsMG+BSz9+bxOvpvSGSQFnvZs
EnCT7VzHB3YXztmxeWD77GLRJ3WVkWt4LGMFNaEsrjiGSkb1sI407nvyR+ti1yIrK/7X/cCnenGa
bD8yxMRNNCdXl4RWMhqrb9S5Fag6D9xjKgVXOOgO4QI/roZ59c+z0MgklGnpXiwCcFB+fNK/h4gY
h3tOKtD3BKSkIj90P0uUqhQg0jKS2ckjzTug+KprOey6ER7yXDC8vWrKqY7pOcvIlMtEZAGwaSqf
MdnsvmVSVeuDRs0l5tVaNAtVPfG/oQrbqnkiTkoSK1oUTep5KvlaL/CpXknifHu3QRVzbsiVGphk
W+IOMx6gENXt1B5a6oApGK7xfzIb+qTs8K4TGPWjqqGsddJz1pOgUk29B6km+jp+nJXyaUyX0yGG
jjI/5P+0yw2rc5oseEVzjB98sKUBGT/qQW+Rq8sZpDEJyWvWouKvaEb7jZO4aWQjjjo3wc9XU+Vv
4BhDKzRYO7/x3BBez95a+nkSfQViRD7NB6wP/C62ylubgcPXFtuHqW4535caTcAlUojKnW6JeL8D
DTD6VoKXOy0HBSbJD6sW4w2zP+JqC672hvEFOfPtW0LHanbvxWbi3V/PB9ES23oWaS1rDQI0wmWw
GhzqLUvkgFhm9pskkmOnimR0Jk6eSuywbpc1d8wkG4t956IeWwB4UF22ASnnnuGyR8yMT5n8/VUy
T7gJSaTZoVl4cTPPJyWhyZpyaFL554uFp+nZwxnSuZ8xf1ardAAc+SMW8k6WGltZNN3dq6SNPEEw
teSqlgUQmW5mYPG3aM34zrtoTFWOcTxaY6w5oTvnBSSyM5Rh0mhppWpohExVpn0fpX4k3kVnyz8D
mkXx+HVgDkfRFL29Jyfx1kxRJePanWlNMPZGUhPu+ECH8TuDmy4QDCSG66IQ8o4dAWfH4rm1q5Z1
xuBi5UODUlLxYA0UNliLDnh24c0eXTCOtgCZAJ4r/JYsuzTbVqv7je7dWA88NcnOsB/nJJCsmbAA
Rujf910y61A6ZlPOt3qXug633VBCINJHwpOHyjNc8cjMoaRREV+I1E9zmqo/sfRrB6SM9UxWsVjo
+idy401kC5mE+Asyid/oPJgZyBaSEN7vPJXbUoTvmaHOtHel4W8YY/KOFJfzQQbNWBoihLwjtDcP
9Nc+DNEJJPcpsyGuj3UbTWbMHgvs+f8g1jnXlIr48iLP4h+S2ziYlJ/ZHD80A3u177KdyaTOpFLr
XaTajagYR3WvlXqrLUT16cBFDebAiG8uxYZVHrgaa7BkGqvcpSohKWnYlLYY6ukUxfr1e+4xZWyt
0xiU1xSPMZsl4W7dpFtB2/uLF4lvVqADaSujqTIRBwezqpdUZoIiiZS6w4fmjss6q4ggv9wjJqRK
n9p04rr5/5m6OBIapsU73hAiiDMGueg1fP2c92f1ZB2kUeYt4pUU3o599PIAnIxBokePl+KzTW/z
bli6Do73W0IKVY+BtRshFiAdsw9PuL0LWkCnRmhH+iz4OKBB4I14aK/mAzQZjbnjM1Brt72cyEmn
mN+ai4uoIjEs/RXX+0MeKCTgm9HQGlyYQkh+JOzz313C3j/YxmVP76tWa81tKI2gbj8xRYH5TVME
/t2fXfoA+mLjbNfrmbrK2R/089gLJ+lPNF0E0UUF3jVennARZB8xvHhUqWsZ8WkD3jSMMAs3XBmS
sgyT9CagB5sZjEQip15GYTZ5QsqFGRPLE/99lmVa3ja0D5Uk1PfRlxi1hoL1inqQdyrbKKFAZTXT
Gxx9a1sS+lsTaJdY9w+F9lq57NQrzzAdPOao5YKJUbtDOpTDKC16KKn13Q4UUL1co59tkDoGTRHY
wK8nNm9cMwh4lHhC75Toqm4WT1GvYaq+00w3/IovACqKo74AkSJ9IcARWc9HuxzyZQNAHvnfRbfA
nn6vg7DHp8epzQtLnq6zMbPVi3HtA6VLDIJ9uVTnXpO6cCnYFmuIeA3vePI5O5Ss1WnQSg8VYYsa
/GA2vfUrrHV1XTjUPStW7YYGBt3Z5n+Jy+dVxwma6LbDbZ4zX9G9zQuNbT/z54LvJM4gJ2Ggtl8M
2Fn1ZsOxG6fUVFJMYnTQTvy49BrtQW2sHQGO/FXy0D96DEDl8KwUC8RqraeCFjqXbBkQ8heezSbY
Mzr12GPYAHA2G0I1lR8hJIRUnw6ELoAG1yl161zXNOHAcIvpl833GWgYB5qdueM1kGhcKfBEtSfZ
JsBrengU0Qq0SBTOcJwFz3EoL9pnvrBnvw0X5+dfwYNEkK2dKUDNnj9JZtyEpNk+BSuI3zF0YuyQ
SKFyEE/q30QQwKC2RDVecgjcD4kF0JJ9g99gtV2k+arx6oKDA34Dfmzp503xoyxP7snTXQx2DVyu
eRBWfAI04MGlnBy8nCW9WXl9SpfoNh82MkLqPUX8WBMUYPZ6agB7ZfjwBryEKRE0jiAxSytE0Eg4
2HiEM8xon6PnamkFtBdlf++oHTPJFMMjj8V3xSYyk/wlAQrzEClY4fI9hcKi6TJn/BmgxKhxmW+2
ZVbgQ7JJWw6mqJmhZ/XFSE3Kgm/gYL6TX8GKfMTpKkTrcKz2C4gPkzy06gRZqWBbSTgM1bJ9E/lk
CHs38Z8P77NWuNExrjcQUpeJ4Gc8gXPioL6W22v77wkii+N41XbKfnTcNUEYJl4mulWSdbRbuEB6
j3xk3FExBvyqQzypH1SvHdN5xCprD8msHfqP4JeyDWsOKiVxbXiZ81Q+Wh1nmKtCpryFpqkqeqFq
S2kQnrrl2TdEd9EnC6Bda9ms06UnH6cuuJh+IBLqzIoI3ue9GWAB0ghfKAN9CtOqyPtQnycLUVo4
RqbEEHaKxk9kdCSKfFJiT2dvfbxW7S8fMgnsSewQ4jI5S1vxv16Xf2c3zidQ4rO/LXfWATTak1Tu
F8PAdDXYHpEpwxXGxB0SnLjU4eg25cRCLX0fFUv3nYGa45+Io3qSYrOJlDfS5pMIKw4xLpeossWv
3odcAYfGySGnzUt1SKkT2sEFe+lCjpHlnUtcrj32HOtdnFDskVsGVpZHaRHajWhDY6QstkHZLeme
H959SriSYas+gsnzFMLwcLulKl80ueUwPB1cQrq2GlqDalac/ZPWzOw2Hz18Wn45OK/hD/HFoCtl
OY+HL4Tol6rR2VwsHdA/xKtLD6PFj6LtW2ZnOmWH+joXbFegiN6xluXlqxlHkAy/6P9qbO3AFNw6
aBkXtzVYT+CfZJ+IEImaAeb0HUqPfUVA6ZoPHueY+Crw7rR4VTpHRsKxHZPsHRr+iYNu5oDXwR8l
9Qe1po04b7IROMBe9glOmX73Wdt45fkVufMVI3eHnvUjjvmmMv0uaJ6wo3yIjqfj/dCCOancUlys
6BWq/+kG0TWJUD6lexbz/ABSOQqgO/HmVY5hh4lzSs5TosLLw9DpBXwqexJaNH5Tr7Pcor17G0Z7
QU9Jia1YIlb8Kra+FEEzcsXqIdxsQix0PbXzu9sf99ybo0MA9m5NLKPHfoEkWFPhTCJLpLkDmdge
mkdMxKQYu7+ALFK8SzKqNwD32MnY93gISHPngjCAUnF9LOj7D0gXDBTZ2WXE59SoHBFMLNQF6PT5
k+aE+IB+Y4iMKS7Z1PuaxahD7BzC3anbz8k7vM2f/4ex1ElBLf20uk0L5Mi+kT5J4tdpAt84yjF3
vieGBj+5Pg+dDYH/b8BsGY+QUM3Z9exowWpX2ApU5mL4NkqNskuFljUPqzsAFkR36rUhflSxX5p9
1wEXXTAymQ3lqf/ARb2L5CXZZYNgM1YcK9nQR0nUBU2lKMydYttvytx2fW/6Ro6KD1Z2WhbObpc2
/C50ziNSwuMervzHRMz/VatfzB/9m6L65iC7WyLGslY8YwNzMuaPwVkImV7Mx9F2q4LARwZAtU8B
kESU1NTfBtWVi/5gfdDxzZWQvVznNLXkb9ei296vb3D9djC3BXe3BFn5aGXd8TQtOiHay84vrKyr
v4am+8BnZial5Xbh+3fuvJ90f0bkYb3dpWjYL8yPZDSxFqcBO6JnMl/ao3asUJkSjbmuV6JAGHq/
AFgI/NjcDwHnuk7Bt5AfybBPiwFPhxyvws3o+cGJT7g1y7FI781uiNmKjBb4SkQXHzobIxIVl7WK
G2v9h2O0Vco1gXVo6xvKVuXT6vaXZk74fRUdmP0VPY18kZMXpY9IIc/eMvStLkzyjf+/9lgw2Kx4
PXjCqlzGdQAivw972Qa4/gbTLcgvSNk6rKt4hhlqKPBJMGglknJdwVECj5JNh3hBwhGbihzZ5DmR
J7LIKMro5ccD7XUoQT80CY/xX+vtf96DqZUmdBlCmhaXrJe8s+wPONa2GC+JYfH/d6CBzhRXddjK
MVrGgKQ9HFYPwfO+uGYA5rXODuwhOv1QvRbm6TiVeCerOiT+pfiI2g9+IQGjhUswUVZsszmCim9D
JjBA1Fs1n/0LJmJpP/YUw8fjNEzUkXuSUNyC18QHF3DScpRX1LVGNvC3SSYSZlokVhwGHc9wB7qz
XEoiMpiWSA9MQLsX2SleQ+CfvPpRWNEb+YsSBYo9UtDhEYnjSrnYsCfAc9C0nxoEiOZ54PJUB+w1
Iyybpm1VBB2MM7uDA9qL2g0X3FlrFkToYKOFuUXU8B5HCb8h+XLcfs6GAealqR4iwtBkm4zb62tr
N57h0gPPDvRwwz2yxPRUqDcBEGi2xk8wInHsj7oT6wyPuZCGu466F7Ui2lJ7/RgynJnygquQRLTn
7uuz36+z8irVDLj0ytZwMaBBOFADUida7uWrhty32zXu8A7If/ktJ0BWE7etAN8leM+C2IhiaOqf
jXMcKPrqZ4FXVaKnTLa14MsQki12blMaI2o+0FqWjN10GMe3qWxLidmvuZ0hPgXpT1L0tmLM30Xl
auYGSKjqBAvY7qouFMc4kVzYrf5oZsPbYlXA4L2b6K2fEdSX0TAcdqjoZvhUaSa4z6B2nqxUQJWv
zgfT0/fO6tzimIr28KhBceieo+P/tf91EfEzCiv4xXZncYgctwQO5Geb1M7oDYvVOL6cJHVQ5kNl
bk0BS5qO0WcJrbq8Al0mbD4FxbSwfCE89kVS5gsSOyEQZGWr+VezATy6Uj+axcXdRbH7n+obZIHo
Vyluxjt1H4KrhHTSiQR5pOtmIOylDeubWbzeEXUJg2JhFqhsW4KPf/88sC8Agno02AYthotxXj4h
WwHEw3GeehsNUJ/hCD6Isr3QKilEifQPTVuDGILhdJy05vzCSv0AEh5+cNWzOUHwT+nEB3AEnkVh
4Uxt/65KBqZQNDkDqshGSN94u1pOgUjqQhi1VhqnCfiAgW9qodcWSl1C0LxBJxPXclb5VagEyjnD
qJxikBz4R8ITP9yS30irjZq4QLGMSRw63VmkMgPJ3YurqRZotdk6XSl8/9jWSyrGMmpoxtZHE0Z2
zEWZnjphI8NvAHgdtfTh8ADJAMKLeQtSflhTqVwnz9LjVTTDhSGIC7PtsLpsX9YxQfksewJ448bW
wRu8WQOv0fDKtldtKWawp0RSnM6LDmIjK8Zu2KeoR9iIIFhnwy6yc6nhm6YX4XC7HPhGlxKTz2Nu
n65DqzJE2dF22nMer/MvMkRe815dYS7LMDiukPp8pJ3PoWeeAU0d7PXvijXggl+EqRyHvcyCAzc5
muSchn8yZzDJ3HKMJ2K0Tq/Htvu3kxLVAWEPcT63nuGM8/pwJ/W0H20q0lzKWw/nV2dMUq+cc00v
qV/yVlzYmci2dgMptnbVr2aX/GjfLParEEdaMnsqXSnihxxdvKPXKiv7nufO6c0plKJcFMivrK3p
VtxE7ATa2c9FY8rKnaG5iDvmUy5a5BYA5y+XAPUPsOydkk+8L7beW61wIwTigeq9nI9wOvW2c0jJ
gI24+ebMBpsnYrNiREERe+NHv11Ibj6FKqp9Yl1yV0x/o0yjVc5OUKMNaOcC6UTRNMTPZVkCpZfN
n+tyXT65LzpqMHEX2jfnhp1Q3AG+/WmNdxp3U9sdahiLNNsqDTgSVCRM2DRDtdB2Y3eqdXcOnr+/
dVrU93+UFHgJt6Ovlr6jnOZuMH8l5PiniF36bEF2YcDYQjyHGMSC13fjbtTDZtWame/57hq6ZWqC
TQAzSwyFncCkSYNOVQc357aYvojwTEa7lLtBmDOaMMUNTBCftt+nqrfaCzKfI0ZmW7uas2Qn6MBY
KSlIfoV8s0na6zhSjvjfeDY1RgBs3fJBf4fELFfCnBSBkKwhE38D55Mndgpzp1NkbXwqIWAWpEE0
cgrd5n2ycCJUJ5hjhULmmfPimkaUkEzSA7RbYu4jpqnc0RALji/4tRkI6p1/2/tfz4pTrwFkbQI7
kTVhjTzi5q0MtQzOEGXXGa6x6msn0XEYAI0O0fSi8d6SvX2y5E+rrA9AhtF6vKfZosG+mFDzpkdK
AfPpQUVYTrnxy3uTMdOX6J4WPfN0UqwdxHvCgHJ4vEG/7JQemG0LvnDPpkUhbLihsiB2ivclQGr9
v2g67fC5OBI7huQqtsu41fs0AAzvcOCTHIeGzKvDmgEfllsvsOFBgIEgmsg72Xn9YagzhFoFz5wo
p1M9DPxdm4uXwtUOQKjQN0OeZgvgdmBEI8JRf+Gwqphx4qMyGurxtAhf2o8p/6kHq2n0DIhPVRib
lEqdij+uwafEV2Uk5Ey1oSwPWialy9pyJIagXcgqfosueWJA8sCtiU+6IAij2mIiPHHveIFbAsvy
IgdnPbsqKc0H8tyg1670wPVhpzSKReYruRFn7IHIW9VnVyFBRQxQf5eBv70xF1y8psH6QeaX9o/a
hSTl6O9BfK1SVnYbrx5yf3UsqBvEjBsOHAyeOWBX0MQksPf32nK4jC2Z3YZ7mMZS4dkyAQ9eMn8q
cq0cIjXMk7DYi/8C9mIKJu33ALV95TXDzytGR40pzWiBWXuaKuclDbuaiBGPZ4WzMcFLCt6gxn1m
n17YioJzh+UXHGtuJViWqyD7bHHsuJYGxWGj2upmFXVSWbIXdXYeT7iifJBEcZ2Opje1vwpBcRl3
FvmyKwt8UHJUCI3xneNPFv9GXe73OEC3P1VFF6xtg21TC8Q3/WJBIWPkXJ4VUTHJLAdQE0erb/13
lSQUkO6BrF6rCfRel/pQTUd3zBPrlncv5jf7TTpUXBQtpnwL+mvdtIUeGZzRA0rXvTctihu1qxlg
r69UIK6mAF9vvGTQ+cGUFHw/xrC8ongz9oTIqgEw/Nkrl/6y2O1Dq1rlTRi7c1FeLiONdNG4Lpo/
rO+umcGLRoYgJp/QKNDPZpfkusXphdedNzWTJZMtaO/djfmQwk4GSX0gyRoSMyieLi+j8q4wDeOE
cIF+CHwkqAfi/s2PDdcfzOpUb0OwmLmlMyh/a+rFWTmr93rbb5lodphTodJN0EtdA2XJRCXsZyWj
P68hb8UECB7J/sdx/4wZchmXmPuZTCM1MJNQWM6j3L3EFO4mES8zYLFRKEQI5GYhADc1eJTlrCUi
Um43fosIX4H0y+oNSrIs43JZ1ty9U272vSnQdRvnYedQnJrRlmJMMXee9DKaY7MGIKyKBieeEYUt
uB8qtvRfdrYkv16DH11bofGVWlQO1emiJeitW7HvDzIyQFVxbhwj/CCFVwutNNSpQMiYdy9PahlS
qk43EiafE6esXd8J0PEMwD5mEC+0kUKoxhn3F0ckTV9YLHXtBZZ/NXZa8f3GNIWNYGyftdiGOYrm
DA3UU7LLRp6wUWVZmYQluJSBYMCj6fYPpwwbAd4aH9yBG/iZerakiZXEnRchayJhWYpeMHvl2srs
x6uT4VKsnomY+PUofH6vAfz1aMfEwHaVaRW7wVWaBulPRxLKEsGK9ghivUSl33DPsRsNZAVycsTw
wu43lUedW1vV8vGhADmsXp9RujDiqsPUA2u8IshejlsmgM2J631sgB1FtyHEe918D4E8IA6ifRdv
kd3H9ihetJv2PjuY7IxdO8qfqZ/Po4DOXEzP+qLqen2kJVepHqx9pwjzdSsMxcPRgotmNNNVTqb8
GBoE9z1LvlyeAYMYpsYSxA7df92OKpkbMS3rYfY0wSF0Nw04JnDqZ9V0k5H/hNy5feNTiCkGj531
G6G9G39Ui9MpHMEJXmA9FkZ2MVb8ndm6f1u0mJCHoxk+VH1cZgCs0AXlksEYClaLS7mZ2W5peJ9X
wGdI1y94T2/89IQ2+Ft3djEW1UrFG0xyFZpx1m8eJJtpJP92riANqLFmWJZmXCaVxORKGL4jgsMW
//D5RinwghBJIuTD7QUrBK/+I0LDnpxLa+238WcIHk67yMwRUDSVYELCnlhml/yojU638pGVSvEL
F1KRnK3ArQsOo11Mqr/3/kubVDuP8sDhfJugcSZnaC4NPmzM40nH9x0fwKrR4HLuvXrWKf/hnnVv
vDCyjSdH0Li5F/wBJdrzFdWOMkVbOT52KNcfMPoT5+N8QWICdN3NynZJWQ1aGnSwsPz+4UMvQ+hm
c9cEoMmS3wH4+IlCdqvS2FFTYedJlnPZB9+aN9BK/Av8/M25tSp62s500jx1B4rmjjDnDEV6t52v
0Pu/9yHU7j3AFbBDlYuCa2Z8MF9zhL0X/7IXlNcw/ZaqiLNxDwqdyVSs2/zyK+y/khx0ZN8afqJH
SQGN+WHOSz+Hm33g3xe3mLKYp5Bdmx57dSWY8maLet6lR5mYe3lYR6tk2Ay+fHR4XFasBhFubPnA
z0dwfHcNQNwlVaDshvxOvykT1izjUKngCAzVz0F0DYut49pilQx6Ncni4JOQKvKg2gOftYWEOUeY
kvJ3oDhVTkDlUjozweSmPukSuhbetsct4IneemTweVXbT12qRYB9tcCcKLsQzevXBeHesJdzhE0D
d45d8b9ZEEhpBBLabF7b0T6kpG5GbMAxJdEKwEnx1NT9CEAigOsAu6wXcuMbFXPj0yNPxzSUMNuJ
IYfdfxOYnRg+NeTXP1u4q6yajPHXebolbuFBlT9TICKSTDoacfrzd+Fes8XaRT9z6YspmKlCaoTH
248WcsPXZUX2hZd0EZbBt4GMmkARU8rpuOgthK/VKJW5052YBEMustIqx1XnwkR8jRWsfapScDkj
EQo71WXbUA/wDO9fC/43vwWVk2Y8dUI/3PqEba70WK6BL0/r17oNfqyqXvps+6yoWG2LrE/2Er3Q
jerb4pP4Ak9rM8oXjbY31wIuxNtwRWGb4hyusCkMakWbfabddlyjRzVnL2tdIsmcWQoenrax6nJt
mywDAK8MJa5/3Hx+m7KkgFlzBfFu4yIAWhZJGYNXKhjMKqTDXPu+Dk/3+XsaQOrRVVKa3SsNGiME
DMcKY29NEblvU9fKXK/gbpkkn9xTE6uKrd97DAceK9uo/TKQYfyAYdQFHkUGZwHzjIZOwp4VuGhw
3Srs5k3CYc/JNbEgi6MtXv8MXD5uIN0BubIihUQnBe399F+SULDTT9UKiOa2y1CpCwAoPUEaUgSn
bQScd03WlUaVrO7VPhQMvI8FxgR5oqZNgpTEwmXDm+AGV2gLtK2wYqObGwTBigfbkDEDmwl9Bnzn
AZwvRzGsS4KPsDlVUv3UaaErtbknpYfT7yb/zlYgkZlrbW41jBnF5JJUu7vq+jFVeInvr4CEqHCV
JCfjDLsiaCA2HheJomXq9cIQe/zk8xOK1x1yr+eC/h7qjSn8YkiDs23ikA99eGauLGL7KtHV8+/c
ypJTnkw7MPN01MmZcX7o/xDYvxOwHjjivLt0wAYWnI1/PE6b0CNmT91jPKYSGwkU2BbO+c7fzzzV
rdx2ZkbBRXViTS+LY3j5zxfcuI0c0Oi+Ymbjs8VbTqcY1S9aZTZM6Gazk4oH8eY6OoLuTByr4WEq
04GL/o687tP3eS1Fur5ZFPDuV7ryxiJ9f6xeyeusoSPzeALuZBk9TPvIv7LzDzgqN2/jVSnCZ1iB
wL69fwzvgDvqhVqebJOiEMc06VgZsg1+8xGtr1enstktlzaeaTbsSxvcRvDkEKn7MdA+wmfKM7Ud
cmqmVtt3FKeONQVtgsZmJiE5QwLamqyilDhqCdBuMnXQnHOgP66pRpRx3p85AWOsbMd9fzXnAcXs
IgHVK9F1qCHrihQPZifaW0pLgqY/U9MeY374+CRgYZTjyPFI1G6z0abniOiIUPOhV1g4OMSlwUFG
aedmvtKeUdyU39AKo1z7tONt/6XkWLKFHb63TQAZo0qFId8cqHGy5ClUTKIOYj6UPFB0Pv3cDHCF
s/y3hIWdgIHbl/10BorXoHcyj8IHzYS6KflQxRJZIRVTR3/yLlK1fxKYUEWrM5BDtW4pCzBQCEDX
L0B/AAC8WCcjA2J7k2GuPemWxoLUOXhJgSxLDopdHP5Si+FKjj6jFdNEX93lMzOdL3WBvQMlT1Zx
b+qM7FNzy9LtNAwTqW5rg4aOMJjkYbrTtRypS7pWtTd4dcwdiJVrtn2Re2QvA3SRZi3uIBuyF3tq
gp3PXEKDfikPLUK1wPmOfuP9BOZ7fQ39BiiQJiZdfNcvgXAVtYOtYURG324Reb8mHs0avnvZXJ+2
xyyYkxlCPAs+iblQsmRbd3pYpb6B4J/oND23N0F0ZnO0BIW/JDQRnJvEMJ6W8g8N7EeNhwwpiyo3
YJ3GHdI+CZFIou+555R6xb9JBizrFBJaZ7jt93UdgUJjiQD+FHz9JSjM6wLUgnGDdBeg8DTxeg90
3wtwrWVyR3qaJgvPDFaSXKDmSQMtaCWvqyhuWXW3FXtU/Cf9vy7Uv9Rc3Fgz9Ep2zVSU0pQmkINm
iYktjKbiDoHEDr5f99PQgWw/Ap0pmv2la7/422VsDU5jvnEZDqVw/XxChI9bUQ4Mh3DU2Mp3tzBr
eatGHJV2ilK7K772CDHpe7V87+1ISG5mClRAgsPqJVDBt8UMk8qSxB+KO+mBQ1eprK3wviQCXEm0
PPCWKpNBuJ1LMnSiSXPepohG+J9Cfaah2KkCc+xEbBHhzSM9aE+wIyJxKwN0usJqYV/rAXsahchi
b6l7PKzjhUFyhFpodxg4zHqaB7BpQZsP/DVRc/Qys/MJPOY9SEzLSX/WqpDwNIsmPjbuq5Rczzl8
/KnmKXhdEorVt06pUDE/Zb4zgBJ3XhXPnQUyxvcTeHZnjB3bEcJzmL/aqS+jWK0sQSXU59ZqvmwQ
VarWOUdG48N+XQYeaQSp4CuwFE9+zZ1BATYL/2fBHOMht3opDQQ/C6whjuX+mw17jXhr6yXcyaBJ
eODjyCoQW0LtMlDvh0QWMzYMuGepDMZzqAYoRWpihkDnzK9YBeM/UsZzoyWaeIy1H4n7kLXBL5al
j+iMacTTOlBXgVL3QFRfXIDthCQvjGWG+2iG+0oOe9zBIRODvqnWZwsA+jEC9PSUUX0bXqqlO0zW
rkCsC4u0/zbdJ9+AaaY5VfGoSecS63lrw7qPCe5Z5ETQQ2S3Z/0IRtKxjJLBDViKniEW9EMZcF6B
GwFEdHBqYZYE9ycZ9eWYJCL4RSfhe8YKjay5XYKNxLJynWNbU+dGpy5PNzdgiXWoHBRTwwmhHHdX
krXFxTHXC6ieh7V5p8m0Ad/O1qyzaao6lD2be8RmbwnMRwfQoLbiSFYdKHDBqR2NMeBmQe1Mzp9h
z5HT1qB3YxGo8SIqePwnKg/ctWzORbcw706H28yvpDAs52/MPW6VN31F/woD2KMHye8OLHSpgfSM
HQLiK4KYs4Hgdiw2dy398+8EjUMH33n+gQS4OnpHVuTx/uYVdJwHqS1JeBtTQmOG6ec/zt+We/tL
m/ckrRwD1PBad0qedl7OUCnxM+GJsID912oKczXCz6xb9AjCCCDqfQidzIO5wFFwKS63tpTUVQnh
+Bgkv5KRErCssnfmWZGXZA2UMQRImJTRtuKA1grApQ4Y9LpTPU2+NgaQ/LIDv9Ii+DPM5AJ3SGCc
McBAwCCaSEu3kLw7y4Wwl5ixL5q9TGjPxy68eIBw3VcwtEXrMLrGXERcGigRUwpN1PERSTdaKGI3
crpKO4+FvzBy60iO+h/Mift0joeqCgkvlHuQRFjNoD8Tf/Y2c+2taJ8gXXyXnwND1VU+5f/iOZty
KrNv1I5aLfp5cTLwhjfgDyhZU4RnXGzpMgLzeI7bf7aZIx7qZix1We02J/1VIunwxjxu+P8DLgMt
LeyWlNEM8OSzynfrd+U8n6tRB9M4AyMvwumDDpjKJYK1GH5tIQP0CElcYg5txfqm+GU0FvQP80vv
wYt7yCJARB+D2rgKDBaeVbjWQ3+tzrQb5K+uBsH4v0w2Kr85gYiLTosf1gURZuhHf8a7z/wgOiqs
i1SdNGIyFaut68D0lp61VLnSM22u5BgW5yXnumRpvitR7x045WR/GIH0l4peBtPOHjAJP9h2165Z
IIoygf6yaNOhUEAY+EPodSElb92UpKsKZSg1yN78sdzN1USO5IsAe/1LEtqwpCny5iI2reIxgrZ0
pcRqch+yH1MTpO32sEjRTnDIkayN6l++cT7jiOaqoT9m35kgJlt/dkZzBl5xfMCGAqB/32LQLAEF
og57uYy6ybkZ2/JVKrvxu8jUntSyazIlpIlo5D4n6XuhDd6C8wnWgKcWI4Z26VHtNJllTECOyqN+
fNpmHfZpFD7UyVWmOucdkMSbuLLd/GLTOIzbEmfX4VgkAuYfpFwLKjos9N6ukaCrmJocUmm7SyJT
dk/ufqYlEGkxrfFw7khEDTcrD2PHK1yqw6qKw0IKLnRdbZf8SjulPEQxJxjEsv8yMVKmW/Htergn
L1ZAYVRH/zZAn9ikh9YwGOylw9Ft/cPc63p49LRWGO30EARWmhuTPjPmOW/w5tG91wqvJ/Ley6MA
M45OO0yEUkmOmL8B4E5q9JreNaNIr0IN/9gMLohJyPCCvORJGaHSQHYCU8fHZsuPt/6FSmm0Fqfa
AiMH0QO2g741COrjqX1BlujwppM9KVjhGuHbnR2bUbE7wlVYCJP2mGM2XRGRDNN0nTDSGCvMNC64
dEP+WILUr+wWXcw3fUFCPr0FHA2SeQyNKh9dUmcph+5oULINTsVy0NMvVlijgnPQhWZlbCx3gF+M
t+R9E/sWWCuZHAuq3WzKcQDX7UjEx7Hf8kaHBWj7/6cknERNbUc0aSvuFkP2j2Ho6QCoXRQtYdoS
HOZDQR/x+4A/gWcvLJVmyhBCVWtiZVCINQY46xes/UyjaFKnEqG6Qhq6/9IUAp3wPTuaXjhWxzna
JOSm4aW96oIqTj28hWE5GS5gjn0dgCrnHkq03wALDdYROig4jJYKGDkw38gZLO0TeViqW2gETvRz
ER0/sfQSTKn88jxu4vAbwJJGgSRGqGc2JLJjBXGklZUODNJ/w0NAcaoYh+pKo8jOil1CcFLxUrMI
5ohLCmbEnRmEffPtyKWGIkb+6onAeKiu9sUNebj5bwJz4bjuZXP8BUNfJlI5L+z+6hSED2gtva72
HRqYQrcJVf1pfEtiTVDCFf2+BpUEL9oLoQ04V91ISYZ8gqBzIl8KPw5To4BsDwQG0qlOf64seaIQ
dQqZZJOYuVWYP/BWuKvlsZPDaGBzDb+okVaYl1hu8e4prWNDmGLlK/RdQELv6n/Ts7XTMa7IeAKT
Gc32w1Rne0XpkOneLw1Olbwd+fGtSvE7QQoQ2nlCETA6LuGSXJwWyJPx546c2cKopbntgcCyquS7
dwh66CnLJVcyiqDO5SR9+SqUtVrkgwiq9CGYy4jqn2PxmGnrODWh7g9iBts9xYknzz2gZQpu5Z5U
POxX7j6/S7W1yLEFw1CelurmiQjUuKdLcZEDXOdkVgemwa0Bdw0Vt7rlRdecOpQL9d/frUhzYvDe
XHCMittUSefr0+ExghBTn7pf58iA79B6G4jocZdYWhqnMHSh9MOLakfvtnuEx3YgWtSa/xc0QpbI
XJJdctf7YlVWDdr+Nxs8VPa1tsHti87NSYAioF7MRMco7uA9rWqcjXhGDu9p2Ogvig4Ka6FwRHFe
wgu90J7NAcQsaJ1o7bKDsLextDYSqPH5k1h1OBTMqqhloQmW5TbHlK1PB/SK+0Rgj7jhJsHjE5eB
9OHWOta7Tl7e4LA6jsJmQCHGmUhEJ9P1NOMZADU8V25Gl4WY3aH5SzDe59C4VZ+8WWGNigTBQkVY
jnrD0Q9eB6w/N+Up5oPhhAExvOEsszK2iwaZBpHZgNqF06QXamR4OrtQlPcmOVkEEIQvX+xzoLNd
GFjkXmuTyVlCD/aOYp/70Pm/mxH5jl1x7nNK4/PVKhZKL9TFwResGTiKPmu9lQ18Zg6BMgUfFYOt
0SZsUVVUbaxJIwuclo89LUlzzLIgI08sFfTKa6oY66DZjwS1K9GkjTYnpG9YF4DNFX7FLfyKhxJA
/CJ2SslZjXb6/YsTHPzuKS7jmq3sCBVm9I925LKGz/GyM75LGwZUTz5FEa4O0+V+QCQ71vNLOMii
RJFN2vcThJOHiOHbJh95tcUlts8Mv8loRJJQwhJASBJNPGbky4V5+l0NQ7ve8N88XoaqiN+h1LOb
5SrVs/EDV1AAX60Bjv93qiKUkL7Oz7NzJlro7F9C3UW82LGexqCq1fc7zEmb42B934bC2NSXqAIt
KEfkwVfetj7q3mjSrsfdH7Ug6kJ7ZptmwMu+C2yyFSKkd2NN3WRGDuGnJHSn7noP66PxMsphpRSW
f1PrXB4r9HZ783b6iPWZ9mkeIGPQplhs8L+svkjd09kwreoIVGPfOD9ZyPwDSeaqyDBu81V4fMBX
N89lOR8Vadu/TA7Y5omiNcLPvP/qyMsZE4wNpmggZyeDAaxOaN+Cr2ze8bKmW3h0mXojfGZVpHgJ
shDd5BJrAnSucBUbh2WBnm8N2RrXXB3iKqqCrdOLGb32HkWvkjgHg0FG4/ostlaeRFFG2gRtqS5U
Abhs7WX2KuoiyBWNrIv/nXiMFXETnPNgrbAOss01dcWcqBjelKgfezFDeTL/47fomAfvAx3MwXim
oiJtkC8s19bX9XZpBmRmsWatUtz0aM13Fbb6W2dy681BOl2qgolvos2wrLzS2MTePYhNjmYFDsjO
DZ0OxAgX9iCg2lOcxb+Xz7x5l6SlFIEEMQq+DljGFHzzPKy9n3kdU/iBU38A/YTqWr92thTxsk8s
UnfM8Jx8aog68ReHTPu66LraiTW7u8PH1ba3hB7Xj8Ikf9RuVnltGe6FMGFCv2x0AwkqinTTvuub
A+aom58snTHpY8KxxFIyCKdnBrKI33uOGqX99sD/5eLpjOzEADlRjSdjqRZ97120oUsYE0vvhBA2
elPIxE1wC7ZhUj8TrJgoXc1EPHC/HJoca3BYvomWnfG8lyJsPJNH6WatER0IpFPLW3WpVsZFvEJI
uXNdRWYmgJ+wzF7f/3CYH0AXkuDI7ynPnheDKs2qxh7Br9ShSD+jrpVt0G7DeK05I+wuwTuxQKCZ
oy+Za0T4DBnJRmso1kSUO5Fm9Ou84UP3R5jrHmsSyMKHbl9ljmw4w52kRYlmoM1VuAhU+KqbzjI0
I6W9t2R4f75wgsGvsvzJOqpsBUC9/GNhzefEw7+y4V4aiGorum2hAAdqV6Arn2THsDMXzQYQhbII
m/CL/O3mR1Ze2wy1hoTxKo6d++yG0DSI+x9BJlPZQ7T0r2+sMIOLg7RHtKEE7A/r6eK5iPofRdMv
arWxARiMQIG8qmILsFRCIDtqDR2JBlCoretndNR7S6Mv7ISlNcoNqIYOKIKoB5g85Vu7l7TGnias
Lj+38kEeimPt4KZxhu211mvFaAGqwXzGLf4cFjKwUxvwBoNyKoghYNAl0G2HCqP6a6XAwLyMhOcM
jghggCXk/Cn1DhH5s6OaCE14KN1d28aV2pOqGIOtkvDCYkYla6XEAkeevXHr2hvr38q2oQLjXfUK
jCyFIGwzKM0SITrXAX/iPO0tYDHkFWjNG3hKqIkzbIhUi0OVCBNMIbjmTIJRNCJ8r0LBUNaQi/c0
x8gdeRXcacXh4jpPDkTmtVLssXGOzhkPTmZEDPgzGE5J4AdSLjjftaMPIeCqdr4wTPfATmvdTLLD
KFQ/M1OAO6td1dcVZSfRRAOSUAHzVprRHbYTr0FIqxKzVN0c8Ie7HG5lb4m8sjS3MtkJQZCQuSDS
9NxydFEkwPchuXMD0b+aag0PB44Qg2r2Df7BMXvULxjanikXyPkQatCQW/ce+L0s08aMa1Uh4AWh
IG6RfABwPngLQex/f/DexO5d5nrzdCp/Z48n9xA+goGGSEzv5T3uSckow2zIHjlEIjbjQs2EmkBL
cqg0veYn47MLRhcs6o1n0KzDO0ValQX2RFLNqYrdZHoh5bOX1xS8N7XtfN0ve/ozMgfxoyhRwAXJ
Ead8xNZazwHLb4oX+VWB9Pd2TLyKx+JbqWypEhiNkrx0O2PQBfhTxBh3VVPnVeqDG7xd7iMKTpIb
iE6oRzOc0miKyaAwrEOPUQfG0IgscTBB6HFSO8Ng/B+Dgb3hETIhTCSGrS9SQ5Wj7iWPZ7tdizGg
uVY7MAqSERiMsEzei3UOX2H05nMRzQn42iU18j/FQ6S+7llpzZdJ0NZcyjJGMh76f7FtZlvvM3un
obDIomUaP3ILU5CbM+avtuSPeVOF71fA1+4Hf7oXnT5fuwZeOegodSJOpePP3g/0LmPxHBQkmS2X
8v9aPKWn66xmn0fqSh3DBxvHPS6/XTl+HBmjeYFj9zYRpQy48vgNmMS2bVo09zjHGRKXiyBRVmfi
umagbTNbHUzLF58QnyHDcUEraGuBLoSO6FC2J828fxtHGNDypBXnfgQDcZXLnOQA8rc47H+GVPuh
VLgro+3KK9VsZkKwr4na3oCriUQ1HrHfB0SRZs43LoOLA9ByFUEQiwjuJpF8N2mlw3/iy8V4r8sX
P/Kyj4BBgyv6OjakeYM8EW4jPmYrfxmglD6tSR5IkYB69qkDHjMy9WaRUJfh9515ygXNPLUGJbM1
3NAhUoCGN4jY9cey2gnd8GC542I1h6oN36Ii1RCn/VK8z7Y6hytF2XsCV7gl27AFPTvGTnwJpA0V
G25kZGejRWKCwOXdVCoZ/PICQlymKTcdLPO0EgXynTFUqE2bdl8yCHncvuGiT1A1NfthaNaKnJWv
7gQTCcqXNQ/9fHaK3TCsw8sSIOjQxN75pVDwfCOxkLeml0F1b+IAUo2dKADwntEb7AzcvAwevncD
2xUng1o+R5SJ9ONogQwgYwcvgGAO7q+SqcCLDv5TM+XDYJZNMyosH6kVrpHTdY+YK/S6pBRZnaCa
LSYKWYphCD1wGyi585sQN3s/PBACVW3qt9V30Cc/4WIpVxvnhyQTTV4Nlzly7HEhMsUYsxZmzER4
4M1yRMWe2YgxUs+96xc277NEj4Q/nf2HoBZsZOyuHZmpeKHPZXsy8e9hHAP/8yM/AZpQYXZ+JPif
l8xBpcpm8x6YtNH1U1p/7h9819cGU7a+5LDnLO81e7s4em/cVJUpVUPJxFNja2r3YYBAvf3yRIv5
n7D4FZGgpW/Fr/GMmIWX/wFBGgX38NA5P0txU6awemr7OCoahTit1NUsS/6GWnFbz90gZKV2K6zb
r7OBqH35ZN2BRNBmGo2eYNuMkfThXo4acOpfxcJENKTOoeBBI+kMIFoegD+HSSt2oIUHdasQvfF8
sxUhOA7Y8BuqNovifoUBsKeqOXZwY3IF8tymlo4vSimg/JD5/N3a7RC3JGZDp15hrfiQ4D7AlzsT
QhfRTKrCeTsZSd5QPeOXBPgwz9zawcsiBIV/0UbXvQVg945GtP6Q9wQAwufwvJ/IJiKANXXAEML7
MsS5ekc/GweTFJyp3bT5Qqp1b/AGhJ7U8Pi4LHFliFG5GOpB4J3g4loneKiCsZRaDm8TLO48Lrl+
32Za0a9dxynzNQgLZtxT1l9JMxFF3Ibu83xUcrxYP75o6OcjKlYO45V/AChrDYfyMO4j2n0NvaMK
ke5nFFkdrCZd0eGB6emJPnDNy7pv9ZC6T4Bm3q17qQ6Hf2Q3FSY5UobE7VW8EvVgc+emYM1nxQRr
zV6B+q0jkBTyENh8XGu9+0ROFdOyl8MvOV0c8ma/EwGfEca2iiEGZbDLlntBTUUb1FNurdA3tmzI
xGWX8QqSgE56yWULO/woT7ANky9salFQhOd0WJdZgRWuGO/j9IfIq3fql6CTkdDbYfwmaxhYuiv2
6IIhLjtoKnG4z3GtcnM8ZT+1KyJzdmvZON74pG1PT6uvBbnGvKv73ECfIAxwkUf3Bpfe029P51Rv
vy+ZcC8eTWxEOd/3eyk3G0BjOvXz+rmcSlAkapnVhbV1ViM23WNoIYOEl9G+qy/FjpWhKs2zUndP
enI0ts2u3Yj2hrUyGDlYuiUm6CFIlXliz6Wq/7ldqERWmcxamp3fNFVWmKgElhYQHs4QVlM3vIZY
SJ2ea1hf/GBGkMR3jmE3KO3PoFsqusd5hle84XvxZP+ZbohgzBx7i2mfXCDsiR+ujFOYTp1WoyEB
FN/yYBw4x/KR+2WG5eowMAPxxRHdaj+t5sZgoUKXoE49qpml2lTzIRyvqAGQth/v6W0GaHurgrUe
jYvyhWqAdw6XXspvMT7kk3JzoYKsymxRq5BC/2/hCPik5srQsQdH06a+8nzbuRGSQJWi9J28CObc
QJg+vqC010bn+gavD9h1BnLDwLu1Bc8DI/TQ9bLcLh3Q9Faz0AKt90rvQlZdqozWLDTABVL7FpwL
KKVJPuRvwgS69QZSF1nPs9rBtvdsP03+dhAM7wn0Uqy/oNh9KGbeQBzsQ/9DXY1X4zulwjEwHH5v
3/L/5AK806Wz8mw/UBvtINOB/TM02QPFrpSyFd0CtI/omvd5uSQtsTGg/BvcBUrlgcO9MvaDlGx3
su/jh0LvVpz3xFG5RBBwFyVD+mwsNmmvc6l4JXRHdYzcy85j4TIrY6DwEj/NehFdEqFFSFJCLro/
jVt7evJClTgRF6Eej0JQKiNvf9tfKZOJy9jDfkA0z8C8K+xf+MmVHD+/yLmKMmw3zSaj1whezreh
nN1Rcb8EpUTt8aGm3MQPW9+6INC9F+9QvIPqeF0vie4nkD6ts9HIA1WOuBInJhFy4rBe8LtRDqSN
jwGt8lzhR7Vyz/zKO4hSE6vWsCaXsOWHxB7LS7s1u2bEiUqBy4FqNkNzRXcES+vpyguqPfsK23HS
LJkUlHx8Xs+BJVaDBQkB57TEAXD3sY7g4ns174o5BUQdlW1R8UMXQIEdnqDcsUvv2258vVrjbCUJ
6zZvp3XY+xHoMSO4qJ4gnYy5G5IOJNO0ws9cYCimZWb4B4YM+sHilohLBbplE6i344eGD1gWk0iw
Jx1txYc9f3B7/Ye+RKo4bKtklveikBHCgEFGy9tXLCc1U9nJzpaWWIZAQwAAdNr/ZnpYuReYotb0
O8PlusAmcPJ1pdEzJbsr2817GbBIp8TNS0Dwt8xM994Qc+Cy0AfmRYUKvCeo+wT2qq4CgtscQatC
5wih9b8wjmB5Nhnkd6h42wGipWxxNPdEjeI+EVikH+ete+LimNUXECRR77nkU1QeNOqO30lVXFkh
D5sDcnhMtyMztipPIovS5PM2ZkIZ2jV0c5bTy4G3ZYGI03Fsil854Y7gqL6z796lSlBIw3TWnbUJ
M8brADhm6QPf1UbbHpL4jSpuKVizRBAYIrzCj7EPFjwiuiGnWh/mpPLoKvEPHaqgau0eNxc2bEIb
Fv0wC+XGwZQk756WB01UiSQ5jdNDadn81lCMyF6a8GGUlg7pEDNYbNMv3lZQ8UoWuTRPy4iGLLWm
NTWrIfGy6r6sllhwUTSWbMVHSlO+qYwd6XHJ7eN/CBn0ipj8bo7NDU5Uh7D+u9i+IEz8yYFjRXRA
zC0vMdvrxZ4nKIGgr4EHOLjp7lqE6G2kaKlowI5uvTo2zX8sYZlbpHEcXEva0tnywOUigzFzXVi5
GzViEPpJb5MfUwzkb/ydAkGGe2jrFMSQoV18wzlU2qR8wQfkpbWfQrHMgw/XDR1suqr5abvaid87
Knn1Lt0k3UqCvJq/j/l1HZeP232xaGW/ubNFN4DJ4o/jkQ4c1g1UeIeuhXh/0MyPEXusMF8PyFez
1Ir4ruBf1dImXCChu/HmkMvuJ/6YE/0e60icEJjuMgaiCP4abJ9UO1K9YabkPcPFeFRnXBtubWE+
pr//bZLsH7/fe8NdXwzm1egRFZmHTuneikvltBBsBilvrfW4t99NLQUnz2o2IrpTrabHp4anDk5b
FghSkPk9M3y7PyU1GkpcAGo4iqSSFUhXvw+IrLHXSBweDBud/layTyhaJlUKjNVWbyzkH4NN41bq
ASIR/RdV87faUEoDEKMJrF3ID2OFgNXQKNrCNPNaXg51TUHDkAHvIBhrldfJW5l8oLHEL5KTW1LB
IPwm7aZGYXvGDNzVod7clf1A0qQr4d71rw46WFdGHvknNFN88ciBuU1chT0KdWiZEcmuxGgnhQPB
9MRl4u2TpX9ocovPiNgi/ykftx3OSkvqGgZfH682nTGi+yPWYayBRImE2zsLXV0neV5vDSwQeQ6y
bEgS8BMxxmOdHv2xeeBzaxNxivRy8iZTUYV32iiRBiVGmPLuPp31uo0RD/7i5k79A2vXBvJ0Jqz/
ZUbK1bV1+wSUHA0i9WcJvVzCzmXEarOH7r/KViM4VaVNmniTBAP+O0X5DyWSB6hXbmOJOI4lpZLh
QwMK5+cwkZZ81GtHGrICq0AkhwEoNRVWiKzMVYi0fvehVhES6yMX7SbqyB00ED8onxtFZYUIIJi4
2wpD53TJEkDOe52tTxVpLNS2An3LTkridx5vqSZJPWr4Pzzz3Ma4f75/GVGbIiuO9fwCk43WTKr6
7eNDkQJTz+5WAryOxZi6Di7IeNKY0/DF9/T777t4Co5FLfV/H1XSu1tIlXD2ZYiznanj2z4BGq71
xOvUdxc7HyFQFpsdSEfOIG8lnsa+WxIFl7tMfcOi1FV1NBDIJPbkRTufx6XqXr8/VhFcCc9HgOnm
7ZWUIkoQjkGr9nLjz11FakvsZtsxvWZI2CVD8nb87WlCyP8et9G7BNd1hOjnttosVbVyxR3j6IV2
SGPOwea623sLyrOJoIvVUG6YnH4RQcA3yD4KvFOoBONpKiqPrrPYLRZICMjKe75r3yBGoIM+cyJq
NbKf0sfFXcUc6nKdRETsT9Zjpenm1oozrSRpBbAXpr+56N7PwIi1uSOTkTkgm/6q2SFH835SeD1n
y1KFgZxU4AshTCY4FJiuYEAj2k/XzqgSgm7TiyiBBR/lU2I2+6PlasjTrcfUP9a0ICJzvLUBVDCU
rNd7nbkWpM6HG+y8hyBA/FoZxyJFvrHrMaFFp+htFrW2kO/5/SsKON2SAnfxQcpnxQCsQxM5ks5L
wCJ0/FMoyFr48nIuAxJoGXLrgI95R9tSA6qgju0qnrETUfiKf9lhbUq0SObzH5uFVaNLev3I74uu
bibut3nAW8SEkupWi0AqQFv3Bwnv3N6JodoE/vC7Njs1CCdMHgU5UdOJXMQJzouvwOf589w9JRNB
QrBmuKuppcCsR0ggPvnEYUpEBVqJdqkKEIPgQFBDbOQCJ5JHgcW0HKf7JguY+aIJB6ODTJDDexhU
P3sOGhMe/kjdMXqBgHoXm4q9Eyn+z9xnmHLr3zqT9tZ+D4ZnT/EhSi1c21UJzhG+Nmf9WA1h7k8B
3/Yf7iyF1Od9UtJD0m/+5Nn6u1f2mxTc0y4hqP3nn8sGTVFBtbdnpVLkICIxrAuPHc2M2AZdB3GI
sOvU+G2ATNE+KVkqS6hlW6Oz6JfA2QUe9ITnjTY9QniMQX+7fd1B7mPIoeuOOKn1pdaZN2PrjnVg
jktbnxpjCJh7iOqckEzZS+tdQtL6EBk+yZfc2kEqltCep/UYzUw6fp9xBj2ufBtO9vIDy0pyFyF9
ugiO7B6emRqBp8phoRdMa6uC20L4ts7VyW1hG7xNvJG/uqFvxr8mi4PpRVofzPh6oZsGTAvKXPn3
4tvzcfnlfPtiZQUZhENPwlzNCBLABK3N6dvrkm6KlzBx6jCT5m8H3E6O6ubBqdn1uoKuWobe31QW
wiopFqlG+/XGdkCxkav1/zixTUdw04g6IAWb1R0AUFt/dDrORNa9iEyf3FUEy1HcZpH4hY+9nbHs
3wzOl9ghlrEB7I8JXZ/xoNlAI+Fvfc3SsSalqJAPEYR3acZ1MZ1SsyMPdPBQ/UuZwAILb2AftoB7
FgmFP8p+/PFQQYrPBa6A/AhDtgoFEpYBBkoo6u3VvgKElzTimFF/kiEmUOAJ9bQp7McEMRhlceCk
KY513zkeVPmsDn/kbpM8pksJ0p0THSing+VkWnjYZmZKmorU8eUzHBL38nNlij6LypTIvQckcxrk
d3//INsuyhRhiXJpoheYGuXazKhyYT/zLZj+aY4c2r6PqfowB+hs3GGcLqHd8MmfkDPLYfJFjfQK
jrOXDDgnJBsU5jL+HM+xFFWNnSbRfuIbqlrRcLsc0dLQ9lVezcVE1lyljqgFX1lY01OlobTXgW8q
Tm8BxRNgjBm3TA4vDCWCpQlcJ60dRjwdGLxW8aLoNdDD99z/NIJHUxXPU9QrkrK2045JIChKk10J
vMhwhINC3E2i/1p+PrkoKSeowWSNuImiDtz/ErJUdyHvZI0jnmqDWAdY24rDTDRmOtuKRP+Gd1DP
LKbAuNVbIfK4gx7fFj4NhunHDQKg4X/ibXj+xAcJnXTbt46zL7DL2XHRKi8z7SOS1zNj6SWxAWed
BD0VxgSXrMs4D6Z9hm7WAUcBPjSzGqMYEXSWyLiDzh+p0QRIKVEJCwdJm2nHVg3yMPn3QeMPMNgk
URag3r11lzg5p+//v/CPVgLxzE+ewq3IKD1aCxbkV/n5y0YYtX8LqxTGA7zfW5StXm6ufn4FDY1j
fESSzy7My4aEDRV3vKCk+JXnpsKLj1fw60bv6kGPufw9bXKCt9vfNkw1EVUfyMjKFUOjSs2epyjE
93bO0Of+dBELXO0UUwY5JL6VZw2ap+8bQh+FAslf+J7tUz531PAacsHb5x9d92IjHocvdnSjA4QP
luWPTtvfzM59b0vuKkBzyMXVH7c9gVla7fgIjPw5XMg+vHmnFdti5kguySKgdoc+qxCK3RN0n58h
Vw5f5r+JGsjfy89eqMfYJnwdoYqeVF+jvJb+YWgEHASvIJ5b2+ybddfoouykWCx1j0hdA9OBQ2Ip
ZkZnQBUnRJod75fxqXURnSEbwobgYbtUG3Reva2FInAyODlhys5sKsli6TtnXXUvlCWqKvb1QBa4
7g3GO3hZ4vefYWieYuNFp/OpwPj3ril1TlKOBd9KP8PkhPSA0ldH7E7bOIw4M0Xt7zb5qfxLEPaG
NwHKSkB5Z0lxC3bn9Uk80e2YrGtq7VnsKY6YcIZ/jl5b3Y4VKK7wW3usE+23bVLjjVehs1Xnkxn1
BQVAV3Qf4dDu7ZVczFaZ+mURxjPR0uEPwWuL7LzUUtE6SElm5L12VToJMFStFr12MybT7XWYekxp
dLXvarOCcBy0H73qmZNvoAeaiB4DcLor32qquGTYAPK99aiMo+5cGUyPk0j8fD5FPpi2d0yQSI5/
DT1Jg1n3Y34l5Y3bsbrS2OgcZgimIp6Jdy1G1nz98A5uP7mon3rTKmdla3sm/h5sgWLJZF6JtIYM
VHk/klyvi6+1rfCOm722OJokLrh9Q6Ohl7clZwd7qw9lAJReeUjVvSfTqo3ZgZwFZE/JA3XypPxz
ym/hRvQtKD/AzqkPaFGOLDxbiA6avl3ABjYZ88nvCnt8uuRP35rQTHLd9A7L0YBFKTfqekIUavlV
XDLdteX2nR0iufNS3+XsyzFEOkDb9DflOGKWLb6ulxdYEwQcNpiKcb2ki3yE1S/GXiPSz2bftgsy
LHw40VToo4EJrKYCDuC9/lOh1JzPr1zWSrgpLxeA7YZaNg0OM/bA5gbdkouR1dRFOYwLTkTdV09X
GbJDlXOXGy/YF0Idx50s5vbsd7M2T3FU/spyUKqbDzTp09ebdV5PJof63zlqkMrBMfL+XEdx9Zyk
uhHajuzVIrV50nWBtBQJjslUpCapT2vRGJoKnTJVRlhL2pQNXFrPUGO9t69LTuSRS3ih9Ewn/BBM
ZyR915LlBgx4l9pj1S33WpaQdknfbs7eVpvFqEXejEWrVwzjEOeT3aJype66k8/yik/DzsuOsY6d
WNZwp2SjJPSK9nCBdRxiSBBEfmUZuAIQT3onmNqh+hWyIdzSKMuvxC/vqYtqXPOqzCjHXn3osAUM
MzmbpqnDbRl5YmqaKVb7JC2bR5nzeO95OqMey8ZimOaf+le5vv8jMIBii8BvITD2WAdQ7ZBt5520
YlTcjVBMLLYLNwG0lNPJ+FBzHRgNHDM8JE++mxRCAW152wW1jav9+h3tzLD7Olo3htYRYvLRH5MP
DRfjbMq1UNMNli19iWIC4RtbbZBgW7VyhAs23EnQVR8tMlNhhGhJbN3acnHv2PkYAjGiFfHn35u3
SE3Vr2A1gVkPexR9fMB01tB+OwVi7fvHXlZhF5QVL9d8JkpNQNnu4FI1RIC4dZOmhKAdcYP1DskK
+72UMqH5GmrH+w6wtMF1Vr8CvmEfA5Ewe2S07E80TXIHLD3o9Aeo0XUQZ2xAakhEoibjIrVENRYF
CHRY3v4iTa08kBPxuIlwIJu5h9VHew25hJyhWpAM3BmrU9ghRo4CZ2qWk7ODpq6G9Jv6SC6b6LZv
D5GtmiY7QBGD7cRw0MS7KAIz9+tCXdHLFhTjVPcsd5eQgugKQES5imdNuj9goeDtaBQ1ql7v0V0T
AibIxHipFdvTKAr5ok7gkyFPHxDZvq20KPKDkhqKhwcbx4GocojpQ8e5Vx47Dyz9hkb4a/3Yp8HJ
xSqR7jckFUtvAdbkBtCTjtMEuGtpwsnRgw6Obaq6584HuPX7qwwvgdzIOqL59Y4bcbgDhvx/Yf1M
HH6s2ol1XReDuPS1LobG48Uf9Jn8fj73lEdEqNW0SiD/uiWEOSUGErt9zRjfPH2aYhioxZA0QTjs
NfKvf/u9yJbIwkphwp/K34fetz/E3Td0Oo/zYFIrH14VsJtWeFPE8QH7TmmiNb/JF3tmL87FzisB
IXD/TeEvrtOfnnQ/bMwg92rZyD2b7u+PmyubOB/4mTjHBYx8ZMfG28i/ywVLgK+XaDPhuPa9yefs
F1hxMpcdWCQUmnF71Yyq2Vsn6fvJe5eBnaD7WTsuPwYFa+HYktCK1nljAkDJtMpydipFizP+6wSD
Ec5DH3yNi7ei8Bt+azBSe4yU/C1u8u/hQrqYm8nXhSFPWmny8O94e/2lKBh1T+pl4DTPW5nVZfJL
ZbwlUDiz3fyV9kotTRslmksYbDh7RClm10KYzSSX+7czLCKVglGZWkbZYCuXvnKwgWifjIlhOSG3
RmuVlYh+p775viRf69/dtW4WKjvtvpu6Wqea0JcJR74jNSAh1FrbbAvrGCmjbC2fxQKqQETtzoG9
lQT7sEssZvgxtAYExA7I+cl5NcDBFgJNFglyC5D/5k4ZEKxoota4I1s6eQCFSc530gFF4WG/2ff2
GOdwuFBKqRnUyiKIF/N7o3aTaHnsK4XsIoccEjDqQTUoc91XQC+4D0syxeZ5ojFsGa4/VGmgwDgy
m2Ue0QSID4LlC1U8UFzUPjhHMWpXLqcLH0oZpa1P3SmFRL2YFMNsrb/pIrbOe6StAoT29l8iNTpC
zZIm0BMjoNNx6kbLOaxvfu96CHCOZXo0GB6vFsydvuhnRogGOQu7Rbigxj2nGv4C/aGWtv4mYrn5
ZdsofbI2YKwtqIYHuQSv2drtKHDwGxBwsuyNQYUSkI2FQvj5HgjkRVYkPql/ZtZYfpGEL1zYaF0+
SL5JoDEUjOQPsJP13vbfr4gevaxXcAafoE6/AfsL0K8p2tSYdxt0z4rRj/eOqkg9ZGaWxSujaSbe
VuIRbdyL/pzdZ4YjcoNmHuVobZFkNmoBwWZ3npBbYVmfyhx/TB/RWX+BZGM8efXZHIFrdfD0V3Wl
jkCHsaZJ1CTZortCFz94KB8qZCpPWiLOwQrT8O+1xDEsjn+mPtNGSXW0LDRErmaFW0JrZRGlcKmm
qn/5UiKr95+uuPHc4qGjaWlxFgEVzkfnmkaTEoUe6al1UE2sv0CWMeko307K56Rv+E+YLafucsb2
FRimhvTrjW/9eDD5TwTIBNli1KUKtRthK7e/AQQQgeimqmEY1MhhgFFG8ANAeQqq0wI2i2f9qPYH
P5doUcULNebDlogqhFiw1KTnAeFS/sa51U62I6rh2jg/AFgTl1dHpyrFrh0bK/pKBKtCZWGvPNt8
TFcss9NNn5B8Lkycd/AiCaaYtxMkbyjyL4bRR+5/WFdbPz8f7ufnYCIaUZl1TNVvdxOBMIUvkBrX
wTvrATktzBeqZ7as/5wp9Yl1onyFeT5gc9yOYw2YDYAJyjCfHSlT3bCqYIa/l5w49OCHZedHYPmC
VVDf0oY4CioZhEYiOE8b+ULtcnBayfDIHwbClTnjpxwOyZ0Ir5Z7EclfoRDH64XfFvO2I+IaJKuB
MU/au9LOxE1tyj8TBYwgaFxC+pY22jRany633f73BdKwy/uFROqfO6WUWjBKnqmmkL8M1vb6eGJV
KZairBombhSFYvKnXVePVWEZUIVT/OquKrvncS96Lvq8OVLzYrVKI6NLUHHrS4W9MZTNDkXdg/Ox
QYkQKGpqk1a2WsMvNQ4QUVr5uByUFEhu6WPJGmzOMQmyhKrB7OwH8fS4P2i4nYjkK9vr/Q59Racn
TI15IIa+euX4yU707XN6PWy4h8fmedXD5DxihrppHMHLzg5XDTtnH7qfOGJZNYkMVIF2U5O+83XO
R2sy0iI/+mZZKrdi97guvCnXTZgSoaI+yvZ7X1VnxSSQGIX6muo0uBKl2jA2RKdllvTwUv5rlFdC
IoAZc+SlkzMhoW+jQ4FCnFHQQZOEt5QEE+y23pufsFFT0trkOTY9Itb1tlVnLxtHCZONCCM4ed60
PnkAmSxQ6WUiW6p8FtgYCUeED2PkEI6B13MyuCzVO809a3EsfMzx+lahcAlheajPklOfFe6alJ4B
Ou+Omq/vM4UsZHmgeH7j4HmRB+o+YxTP818m8oWk9GQ7Fbo3hlbm6aNrGUeQVMYQ/1+S7KoCbo7f
awWKM/UV2xGmv0Oh6qh29QqFRGH6NmpDFas8AFXDNgq4cGA2+gwaqopaXnOzR48oHXvUTw7Bffin
Msho5So+szcSKcp9kqWPDcBkN80y+bqG4x0OoG2woJ61JzGtCfxX3Eozi82alYoAcF9ocBKmTha9
WeMQdBm8tujmLaepXuxyEIFKv1jG0eR6zeVN+055yV9nmUrw6bbQaK0o0URd20flfP/15YVF85Tb
c4sBWsDZExrBurCtNgOxrbtigzKrCU35Ms+AFpkt2rHwXpXQaHBr/nFcSijxcqpeyTT+YaT013Nl
ch2zETnwmdnkiBHv2NQpjnPDh2mDD472k93YLoXZk+jo9WDag5ylm2bAW0VGoZgN0+lyLBtldjmr
WE++c4IMRY6dFH7ckdMulumc4dbBVW+cU9gWg459z5uYhwsiY9QKyq5rSSE158ZI1iREedEjEGJY
xCMlU5+1BX2O3dWXmcYwVIHUMWZa/KfW3bdh6E3feN71uMfkQV1xRXrISWgF/Xo0II/PShvQDqkL
XyBjmSI2lAbXgnlApQlPsZGeEL20o4kde6zWYp4ubUYf0ZBmNkeF4WLKPspw0bRx11L5ak6XVO81
/kPp4tOqEcZqpvq0CYWavutFNhAITTK72lSRPLwhcoTH6VZAreCCJU91NHxxsNaa4SVw/oycjPEp
HMAqijjVng9x8WYzvm+5VjAzbeNThVLQb6nfGbPIil2Kx2bWVe3eVVaacRM7tSxS8P/1W8sIT/sk
OPTOvZIOPXOjhh2dHxHFnOiGEweXGjpJ6W8QA+2SUvOU5dY1Wfslj+jVHwBH5vr8cpyQ+jFZKhlC
4Dc00agK/guLKbI/dAXPACGbPGFrLrWAOwUw4ALwobuVgPJ+mrSVKbhoUeZ7+8qaHEzNWdrNDoaf
hcd3c9J7Z82N8xO1Wd+/AfXDiEPbQkpwzCipLHWoa5IQQ3WU5j+bNk3NpvKUDEFkRwxnUyTbJcUE
DkfhdP/AXFJ5r9tWUt+O3xjfQskO3LnLpPd3LGan1eiWodp82hV0WOnUxMWGLts9jlKtwBhzxt0B
Kq1D0cU15lKwDIIuGlVj3Z+Q1StojF0QLDNG/pz2K4gw6Nqy7hQEzKNEjoum++dPkem9mO9RU5UN
LgSPpMp+59llFs4cmmQ16Ve2K8GJvUZW6nTmeZ0ZM5uXjOn0LnZJDw3Erz3ZUHActkv9eoIG4Pbb
3m4gyCMEZLYsLNldhj74BqwJm5VL6HtZ07sipnfRDsYe8Ndw1yNy+BmSHd1UYv5iXsK7HNgTI0n8
6Az78PM5MnJ5ptGslPCy1MQmOB8PMss9de12zq/tlDS1HEhQo4vI+T/+WaiJtacYEAFrojPDDvCo
4lFBGxt6Pz4vVGdOYPw8Wj47mv+eLxOP7SafwcKUMi3Yn3Ir0BxLPPceItKYr/d4FZC+Tb22K4xT
lW4JZkTiKoLO7va/vGjv3N7I2v2ZoCjKPfb+gC8+dNXgsyH6zLg4tjbU6S6ZbPiL4T28BTKfg2x+
rYRpQx9wDMXk5+5VPB7gEF2Dk4U/pR78OFPRenfVRxFKVvHdOm1n8bBYObns7KBH/0VZ+FqQMm2x
CKr2czUwGRA6qiEGNdkG7sk2WJB9621Aykl6IutHEWB2QBAiWelIpWs4PNUcYHqRQac7M+ej3KWk
+JxrfDSKjl/dQx4b3hRPOcGpyb3AEK7M+iArmOdpGPCteuvNKyXmcbT1h3vGI+5ztSSichu4IUUN
U1BXwPiV4QKejyu5aYcrc67c/pYuG96R1JG2oUsLhySBmAtaSVy42MNq8OerOMJwvv6ZL9IW9aC3
m/gZTYLem0rD8QsbjYzYh7Ybl3FNMDTGUHumGryu3b7dl8Ej6CY3XcgWa+1bQHc11MR/9TNUBXVA
cOVYNn4h/ysvsRhm6yFJtjUD7YFxbPqYSITHiu6UOgMAZc8AwrLLwWC/FtEMg17yWWN1/bItQ3CV
6TO8Ae7ost4mWodKPBJYtoAL2eg6d7xjYq0H6OdOsTjgjinDbKqLftEgiGf7kMWkEpaR8GYRl7/M
4+R7yGuDDA8MRtqUZi4WokUxHoP9pKnouy5AGV4+nTb6kP8r8MwNThm9jWF5JgRLB2R6jzV/nch4
4kuMt6otdjszoRQ3cJFIFq7prdqkSBvtEhdmDRrO6ZQ+AdOyT2cZAQyfgynVQNr8K4fmiTIOFuJ3
8dY+me1OGoQKMmPFRHhUzzFmY2EsgrhpW/1XxP76XpGFmoNGyRLxJ72eY1jDaAPHF5qG663bKYfZ
CBvbuy2DKAFmj4u9hYLtNrB6sHL44FWbZnl4Q7m9pw21h7vD2+5DzSbMI9BhItCwQeZJTqA4lZfG
ArL2iTUg+2qTjixFCzzRQZn5CpAJJ9+itVg1zraBJoFQ4u1U4Zexqtc4hP0FYJIMvZuk1zzMKdTG
uEmCLp/wmHGFoPeZfk9qYzumgk0P4pYlypW1WBDC8J8tYQtgkg9fwe+n8Fcls/03WsEF9OEDqArH
15kWxMtlZvtX7ZNh9XQBLTQT3ZUN64b02fx/rzxk4O+xktzwaZuSWAw/C9T+7+9uUyRkTju2wABp
Tlj3AqUh7giz7WrYz6HFE3KBWb6vowXbRs4mqTA3Wvlx5Qk6DQRitHKokGKbbTFSzul/EQo9igzp
yqLEhadUtDZAtt6krGiIDsRMaPY3yHsxwo+mgErUceZCa9dytslRVzShRI9vLhc+p7TDSKFK10Ca
jj1Io6fvyNPGiRJGR3GeBcG1ZAY61xac6QO2sP3Dmx0CkkixI2a+cUXrNU/RHdDSmOzp7vjWrJPf
I5Ysgt0NT8ZWDFuq3jZQCeSzqpeHO/M1q3G4JeDxyolsJuTiCCcoDRhu0JzEfTCr5EK3HZjWv5dg
QfFk/gzVx4xyj1vz+x2D0rJPSw3dR0qwWsZz1NRRQXZcuGslRkf+1ymOkhxYtEDufhezFqbdycAm
frMiIPFVWndQmXb/+Vnt9r3m2KlgV0yGzTpPCW2aOzm0WKTkBPAY5+u8H9PxX8PvnCxCHHLO6nRE
IFLlveYej/DMUbNy5m4vtF5AUPCLEjVWzcKO7p5sSePCLssMFLJm38BZtflmeAM9QkZc1aGrcrsd
hTWOEpmbP8b2dvwXkIcjijQ8PQPLMsrNiEey5afuwAGSvY8sL5WbXC9lHAuKP0Cb4sXC8VWKmGh1
yO8rvO1AiU5Fwm8Sx970LicdnyGu4aQAs8DTlb60YXE+7tSSFYUigMQAvAdvYPOijcZlzJU6/5fx
huPXSgWERroYvrcyf2CRjIvpT0G9jk482B+dns6OwKdR7+t2I4v8XNaJQYB9qmOapiK43Z/RJp8v
MfSBI77C0At1hyzvJiBKUvwZRYonyZkfVU9Hzb8WBzOCK11cQJzl1jUFBJDgfXrWfiSipqxqyiug
xzf4FhFi7EogZiNuRSORRjR+mf4PR/bEdERP0L63rSu6dExDP6VEfedKgLr9yc2sTnpz+7g2g7TW
rupI6/7FgOAuzjw+vLVf/4bdw0mIy84BE+YUHMNq2EeGFarm2tPFkAXUWKKgi1ZQQoC77wX9X3ce
CV/QdOM5N0hO4faQrS+XdpSJlsWlShTO30BVVr4j94VJyKuuzKdr2+FyCGNbG/uqAyR1XnaqRxyF
mXhEy1Obx6Vra7O2YA/VmMDH9VVL9lp61A3Wn1nMrqcYqJDuUwpKx/tFSk/A9wbukZQBicaRpt6i
HgvpXal1WOmOvtwcoG2BulW4Ajm9vUXyjGvc7f2qbzIFcLcEJyVCFoo3x+x7xpkxQ43jYEVkCyhO
eain8XU5L4ZArGsxMwQk7NWYp4blLbCFMdtettl0x3cLySkeRxtX8dTQLKt2ycd1HvhSSF2FiJXq
/Nx+MMuHYfT3BGOB+qT9+NmyeCCvqhrAWkgLP6y41KV5dh81ODNl96i6b3voM51ybeqAFfPa+Tws
sBFY9fXH4B7ued4NiMouwl9RH6Wx7BdQbD/MN7HqWaidLZdxiZqbdqI+VsLkbil3LI96qMz6bJKo
7t3Ku/PEUlvWiPj1u3JxdE0hdIWIHMwhniq9MlUHWagNo1gxV84B3R+op+zDFSTe2Y36RbMHqSGU
TFFAPIPHfdTEcjmKoJfta/V98+DVDrEbuXMjeRwirBIEdZr6KhVpuBRyIBpO66AA5lDLBhuGA+0t
8xs+Sj6jTXMzn1K23fbD27gKLPRQBdY6B1JrV+l/m3+BcCHx4ft2gX0laAf9Tepo2YpBV8x24DV0
r85IWS/zyF7fwFGEd3WFfy7q4UsBvZAeholbwby9n/UO+68xSEpDRnopT9addz1bXI4GQizlVsjj
vJNeI5xmmsm5VP5GZPbBh8HNHx84By7Ri1bCl1fygg7Z/VLiSAdyvDxH/BydtgUGL7UfAEhULglF
XS8zUofYaIxrY0QSIk6xPBJTRYER8PVW96ugh3+vuOskbdkDA0ewVmzkEXFbsv8nmJNUsa2YIotM
O+nsibKxqku4zzMN0N/sB8bWapgA5jzBn6szakikaNoyOUesC++atxmWjCwG6fl82TYlWaDuZJtl
OXc8uYFale4K4qI+PufWEJ/Z1JMb/Tomq1YZR7ZIDMqxdWDGUimYz8od0QC8gSlvoGT8PY6pPfYq
vZjyeK6UEYw4OjSGTUYyZwax5+bg5bEXun6Mvit161IfIsxLn+0ZZI2vtLcXP5eklKWkvVLITzf0
umNJVafPeF/Ar9u5/j49vxbzflETbFqVG1RSTYvyVf/Qy1ig3vTHDg/CYY5ecMvHdi2khC2xaiSx
966CIXJaYmhwJ9D5acfSWGU3xcHZFx8of3gIS7xqGte4CDo7PwG1v3lOE9GvDo2Lzx9rDYrkW4jK
fwPRX45tGJCIKZexFMSzldO3dobYQqT/9PQxnlW1eoB7K0lXIUcpP0RDKBKFzVpEKVVO4NsFXkDS
fIqazHz1hS2CafAndXxMTwMHzPqxWHcGWDhEf6s2Bgyj1u/cyWeYMj3wir+51rbqqR48BdA7wPHS
PVTYePygFyp/cdWQlQlVgfnMRDYzBAIzkjrE/h9igDYlT3qOkW5s3cPNPYmGD6Depe1524yDD6/z
vK1TQt2/hAg45AsShM7ba7pLL7jrNjj0uXhr3tjaOufuviJDzyiXo8htMJ1EbsFZSbNuBkBvCc2C
ZjZJlaSJYQmRpJ6tcm+TjJZUBP0RQSGmTXjvXMUrHtRhtffxfWrStcTomUp2TMfJevKogNYpg5DH
ulzt+kzOLjsCPC/klXYJLl3mIz/M8WCPsktegF/wiCkW4Esg4adjoA5PEJHms7Zh/2JuNGkVe4QB
PIG+qdfkZNFjZ10nQaIEAoHv8fwK+tpv5i7OWFgMzkT02mH2qha5/l94wu7a58SOu1NVoIgO1qm0
IAC/Fvvv0QsH5Y09yPV3S81+1JIiDtqciNFP3gwZz+mKt9F82YCj9e6BquXJln5JsM05pbEKfdqv
GFrVuQGWcyMMJun4IxY/xeM16/pwyVteSQKnYGi38sNl9l7K3pnwiu+TW8lDDeOSV45GNqHJoy0j
Wokp30AASENdOXIYkNOIvLUqGOcUYGbkrHndzJbfyS8hK4TSP7XYzLrcIZYkRZU/82Q0TX6bOLLP
xvxOVaGq/p37l4l+k2PVitu/DAVIBgxBY0gPby2Gzbxl7W5eTsKgNajiFzQ8U5gbyWbVcZj+hq/k
ihp37lk6C2M1gfwkOZ/I0m5x+YPGMCsN0uw05qNJyRXm7TYZxt59iNnwlvCVDI+FeC4BavAn/uFv
pM8XAWrcGlX9HjuH1Oig4sacXa4YqPu9XSND6hIjGWn8wehKlsAgwQV9Hp8WPuJyHv/XrYwuGurc
2rzVHoff8kPoUJu0YbL1c7JDBRXfot2CSY8Ic+fMtUuaZZhPBt4SfdAmj+9rrO0r+x0Q6DnXCjot
PnnqldMVMsDOiUYG4Nx3KT+D9Xtc2N61eEhzz5tsF90BULRnhW0OkW6DhHHzWGARGqlx28Tkxtcz
lmma7NRDE6sjVG9mhUN4lImGVlwC+2+NM64Fsg/1euEmTN+y9dnwE7XP8Z1JOVLlZrgMGyzOWCuR
J/KaXmEcwXktUqL6wT+f7XB3GW6mIb/qr76LXfVH+4Gu928vxEakCE3CFs3mCsqXaAe6lb1W2vVC
k7SMbFOiL0UCuhtPvGL6XwGIAF/rWc7NguMDs8lWZYBqlch//UM1iEyglYH1FIt825O6LXnx49qt
n5Tyo9UNmY6Jj/FR6hhpzRaZ2XTE2+n4s8phhIrNOfmO0TUwslliz3+HBhr9NEwCKU2VTMOf47Ux
6dPwEAMd2eVmNNZvBzH90AKuaA19COB/rmSte46P4RF7D3Ic+n1XRDqPeAWQbSRk/HnNi69+d0qD
vOu+IoySBuofMuTt0vz0/J87+1wdsCAp/2+cJI/6k7sx+V59dXgvYhwhvl0G6kA18Xv3YsoCAeh8
/44Gf6RYyrMuWNhqYnRcFVYZWaqORygLrFlR+zqCPAn1yZC3s8+NpFTh3AHkiOaW0/LDrFxiDW9k
1T+fqXUDCmACuANE25QiCL5sZqtthiHJDpGVKAyQllCF5vn79FA1PYXJxP3yKOphCHe/Mbieey57
ExLJJlGNqH62mtKD37lr0iS7Ld2dYWZideL6GVfut5lkIMPo4d3rcx2dCpbkL2r/eBGizIhRxIOf
iOzBwr6IRXbnAaii9ze73VC5cv/7+hY6XgbqvpZMa4f8UiLKKo3TAcBd/16vNDR/UYciCXi+KaFh
oC51IuBWzoW1rL0CDjJ7KbUjgssrkM8QJQh7N/SK2eGrTysUJA+CYUqMplz9c2eF/avm3moOl0x7
cb8RWXIB1T5yhw5lX7QZt0UoQpcUl9AA+u8tLJU38o83TsqBzjBBYr38axGQsi8UumcoEtjQkET2
MN8ysLPICXLRmNjv24WbsgOJjvEHyIs2Xagz7PpSFg12sBw2MbxzsFrGAGHw3/IiV04XKqPBftcl
sY2XaGCvTF568sX5pP5HMT2NG/knJgTz7s5P6T6+0hNBF7sS85zzI6ntMBvgXxoHEZ1UIWCMIKN6
Gkq5tKtzaTxYzGBv9B9NRCsY3QY23gEr/1XpCpWSIwOSl9XoLe/BpH9JFdqG6mouQZ5ZOky2lZFt
+nL+43WoRIAsktYmC1HJXsPm4lCx+fQIOE558v5tOfNBg0ogBaxyxHd7QoRbXrq8filUjRg1IGwo
BDumtuJ2lFPFJ0n8R3pMyb041/MULZCse10mlpr2cNGucSsETV1LtKSVx3WaqZuzKuKALTVYyDY8
ZPp880FJHOmLAC7lfm+t6WzZAQt0leGM57qPcNNdbFpDdy40+C1BfJI6YGZwsDx57WqFTMBwxV2D
6pR3NPrx2dXjZZVZycnsR3pDFIHynPfCzah2F0UpS0IfDvOEbJbAc/U8vO+OcJrWsjSUqZcpzg9g
lM9iZKV/lZgCZ0fSuicCSIzKdKbSbKLRbC2bdX3u/u8bUTwHAaKfjIBUq90n8tr+vOJMj0IB7auX
2Y3Cp/DiMf/ETVw2PD6eMRxz4MZKyYwH2ApnjerBUD5NNWaetsGh+FN+WHzvfFttLdI78orZcmN/
VSpDEMao2GvN+8umKqXM5cQxxU16gji+ASEj2zIDBCzpG3Zr6vkyFOte6n64oXKPC0ZF7P5lvuDS
UKiAIImSzg8hdMzXddICVnghQ3MiVrJAhcyunckGeIpa0Op4I6VeAecstHhCXb/p2bHWOUWT5dBi
WXC6uWn/tvWnQbsvZBcBhj9aXuV5HEsTvdlCCJRMTEmaKYg5r2Oe6+tKXfw1vTFB/PjK5CSdiT+g
2uWm/ioxW6cM4Kz+wc/Hu4ULwLbyAJoLbe13FqOl2Qhq1paE8jFsJeQaJoyYP6m6M1mhguK1fyw3
1rDF1Tq2aPZy6AhyBjXOzgmP2o8yioPXUf+oNUNqmZjmKZM7/WzlPOnm0wTfqYz001Aj0O0B0WPW
KDRXT13Z7FXPzCyzsbjPqQkxcKqCBoqkFpw7cARvukeS73jSxkkeZiMViIpFLTYJdC8yFFLOtkLD
rwiACcOH/Cb6Gl1o/m2vQUClZDjdwsU+sbJjGM13D3lj1dYoi+i1D6ifw7nDQ6dEn5bJIfh7vHmL
If8RGtKOyk0j8SjkSpYZh/WxCSp6itonkXNSXFJaCyqkQQ+utYQ2GkGumkUuSprBZzf/mdw2ep4Z
nwcUfXAT2ZE0BvnT1jq/XQr7OBKS7ox4WLn98wTeagMTCTQqcKq2UxsgZwWMaN1xez9rCFoNSJ1Q
AzXKZsjPFm4badmOd9BQRO/ukvXp0FKkxHgE+eiFVKHf29w6n0e59nX/pkP+AI0sLy0mc3eQM5g1
Xyb5420M36raLlg8S9fSYVVPcYnMnNV3wdTkszWEqKb0K8POMOjSxzWsJ2i54SD47xM2wb+0o9J0
fdfgCvL8eC5cwx14C8rUmOrjfNAA0KQMoKjJvxSGRFEUEypa70GwWlKcOBKI979TR2bFGjf2zhqN
317xPjIPWfHkhGgwOTxsLUiqIebL3vzsrymOmQfyiXEJOcJ0bVTzzUZskxhgAg4cEkVfRnANWTNh
M1Zn+SQBYmlo6xE6ZvtyQtajL/fbUKRjJdifAK6yk/eDJZI7aD8jueAbXw2AXA/CybfjYAxsVqSM
ByeZAami/5tWi9Y1OlxSxagzo7FFPzAYcClNYQiP5f3lc6SMagpi9GMNmze2fkSBSvAGSZrO8C2r
oN8jpjtBFBCBzJWmnbsRCErYO9wVqCq6IQLmVkkX5gOho4rG8GVXYHBjs1Fka4q2MTptIdrgSdIq
4RCNhP3l2wUN0iARCz3vDkxXWVNfDhFCtd80j5+iUBV87Q0YPextswxN3xfnz7URgUm/G11d+SSv
22FPocvRN4dn+Ntey3o/T0GHm6xsCdDtshK9tXYqrzhk4ATaFrjwr67qNzCUjHzZ81jS85V4dUBv
c6GUvwEl/DyO8NUfRWRz6pYiV7vgo0iimfRchHEaM9GApKgpUSM8Ky+bS+9ownSA9MgFynijfGg9
Hn0MsCgd7Q0yrFJGy17XkSw5OVky8Gp7/A1drwZ1muxsVw7MZ7JR0yqgd5EEdbVK95OvFsfvaR/2
AXI3JUioWAkcgG01a+IN31pIlgMwV/3EWiOT75nwvWgQzqygAfiLjssHfyluXtCkjTm5GPnLITMn
p2zRDHowJ2LKjz4A3XJ1VIlFdhYqQcMk1gMSZlJ1PctrsGgx2j4DM2VmehJSmd0gozhMzY5CjQRu
UikGel3E6lglm2PO0wz6ALDrA4iyutdQBHC/ey3Dz9uj96NE0+cCn8fPNjYZMO0kIcJdmISkEbw2
+7+tt1Gkgf+hfpYGtqJeAlzDvSqRKyenvIicGjP88ySnMAloTg5G9iCKblDDUHgxqrg9/5SSGSa4
ljqhhH/v8ykLu/ghwjNmpbyhxoFrVZFTAjh3zk8AkM2euETWFy5KWDobjU3ebdG19CA9GCNfIFhy
hqHFNmD3TgEzjdhOUh0VH2trbuIqrDn/djRTyrNrqK2r5uuwbT64OQIJJJkkRjchjY30acdhobmc
iAUYrSnzyJUU//V3HhUGUiOgD1JfamM5ChDiUtd8fm3aoFaXYwucSLiaC0SWs6et10AgjqHrEP0x
C4M4HBNXD7TfTd/pY0V1QujsYZhEWY+H0UCevhFifAr4XABtcK2dHO+/5+7EANhUyn+ydgSlTdGD
vlnVQKsHS+VezSuEFot882EXJyE5HkaK0wBtPyzc72gIgSYVYP+69Dlk1EXq6FST7j70aca2upp1
b+bzWxr4CRb7yt92OU5SVxo9/r4xZUZ+4qkoE3R8irqI2wbbaFrWKH5IlhXGb38EYf2kLOsVg81p
VGNoYQy4lfz1mNymj44ysXeI3D9UEr/bXRa4UsHwkEEb5KpzhDLYkXtyM4flcrOTB8WDrcSd02xF
HEGubpbthX/YgYo7uZRpZ2PUWKTlgs7obPDhb2kRk5dkUQ28dlTP7W2qGCT+b3yPptOOITs20IBG
SN20BgNw95uJ+krsoI5FJ5IsSbtXXHbXkDYG+fgGRJgXri6h9vq6xjzj5wLCBjNcY5HQIKNCcKa9
4KBbGI2NnXkT42LzSmxT63Whw8hf01HIIU1fABm1RBePhdxdd95NQPyrBKp7Qq4vU2q7cUGR3dPv
U9yZnzdJJfAjqfncU7eRtg8QgiPktLCJtUVlW54dV4YLM3TF74VagbkrLriD55EkpjqAUUex1dJh
Zj1C3xS7K/mI6rxevJsezZhyW2ICirtzKPK3VAuuNUbKc4bCqy6N1tvBL6n2uUWtRAzxPZqPqKB/
K1zvFY4beKBnqp3MczybOzDC/XDlRJBn4VrLWVNMrAWIeuTtM6YhpHtIR2DXjen7XC+TXZ/IpbEE
++6RD30jEg2QbW0VDVoos2EvA17ne4iMhlA5GEfB7fueko5Euh6PcaU7KAieAP25vwvese0MFgWu
o0Qx3Fli0UVn/iHLvGAXWf72kjtSPuxeCjNGj7xE0eSVgU/ALSr11GVlzmglA6RHrhyjLG5c6c3E
g9L6d2kIQxi/BnkD3LgT943eEEPI7P1rQswbnReMjfEBh9zOuHHmUp5e+zOMDYFS06tjxiMkEC4h
w6spKoZq8FunGd/YtNhLfsCCY42z6yNOTLZ7wITuGH/7yqwssbhZ/bh1K0sgvPzmKEeUiEbmGUfW
/ZGtmLVSlKpkQ/b2hPssFkWoRyKs/3EVVu6En+4OJY4NZqjX6M6EqfZcg5q2AB1nrE8AASxWiVJr
z276Dz+FDGUeOFXXQY+UIwOY5zO1e3t0dFY8ljp4JZSyEuD0/bwxO+Lg7iW3IfEnLOv0qtgWpGiK
gGLiiSweqlAWTph1fj9hE1L2AIker54AIz9OlUoEGSm8R0Jtv1c5hGQTR3k1b6o4ANWJzyJ6ffK6
FryOhzZ4t/xBWCfo2Sb3FLQsqmEdBysq+aMRHVbZUTguuKvoSD9S8+v17JzjkIiP+a3eYnnvKt1J
F18pCT4qzs1wZosMl6t83Xg7vKAMLIepgyE/JIGXpJiG9Zph7wRtNHi2SrETf9N8VgcOnt01LSDL
sBGa7KOyT6VMYAnIJMunDbMZn3S54L1I0hCcrOr8Qym/vCIzwjk0fNeuHIEFV9xtxL4mLyQrT7mk
g0CnFFsc1ySTxoHGuqwQxYfASafjhYPMjW/YokYJIld6DgFb//oBfkK3oXNEoxlLs8uzelXReUio
0YkixHODwYscI+3JJx+Ta5aV4xRqmXcS38qSnzNIXXty74CwqPuFw0DvIwy6q4fG5R5oVm655KU5
aV9e3DonmuaDsB44vC512c7fapkNDpdIaUdsgda9Qm21R873UIhEPoAKvDjsh1a6NoFPWsh/HxfW
2HU533/I4lcPUyMvTe+KDHQohLP1WzpGIzf4TKmCvDL2XeWZGnth0K0/Z+JPa6y0K76uDxazrpuL
rHIAtsm2PGVC2Tw7tDPef4HYoe/C6FInkTrPPhXHZt74mRaQUIi2ufVS/AP5iYJ0N+QivnNMqrrC
TXzkD15jo9k0hltnnNzkL56wJXbdwUm+BDJO/Zp7s/visc60cZrgy7E+R3D9bdbEKzPT6iGOiLsW
1RCm2LS4bravQU2Zjq3B7W2b2QQjplj4RwUMwdZKGqt7Ipyt43S9XgU0x0hPCvogI/ZaQHFJNEJ2
g3G5JAHWbpx2cByb1YUEG+te3dMHnjsivMP6slFwKsjGtLTwRVI76ql1z/N6RKeVoUTsbhdBwV3Y
VKF1I7Cpvf1PzS5ceofk65Umme/kfXczuLJrEkprRZM5a7X9XvQFho95sAXPzbkg+cuiM76yOnMZ
nHiucTnqCj5ute4owAldS+/0iCV03W9z8HUlkRipEPYFVMOD2sGcFQB9+NYqnRgQEvjzhu0atk8M
VfaZS5bymJ55qkEuX6Z09CyHP1r37aNOlcKFiSxw3pA/oYmN5zylsQDo5+W331ZKPgHBLyuoIiyU
4C2Dv/7MxL7hO7rXvb866Jb76ttLGNZQd6cO9bwFvj0XRPsocZYHg8fonN5oH6DiyLamQ9C2s1sd
CwK/bV9eCkU/m7S/SbvZjg9wyr98oLAJIg4LgXH8eo4ltElm5dcf4gxzeqQzJSMtKrRTDTFmxGqQ
5Q8XYj4FYSzI1Z5htx0XNH/vV7PUSURe52He1hl01t/Va90B34WB4k5YRFOJzhLGFR5T5II8cOV+
9fdnlqWM8JVvDHaHG3i4jV54DUTKFrAFnFyG+02JeOSwO7lU/GInB/7tjnY7hWHOzhzvcxIWN5k/
qUMSxgjo1Ea+yx1SyVKeNSXryCA7OhxjfssBZc5nWtOy2t9sg9VzxyLN7udjkhQlGp87Y4aPTlte
JVUbmPkP8LM2hjhBzIHCUHAlq0Am3FAF4rnhXxhxolGN4k6OAz0p1e68+Kj9AQ7B31OdKwFxBi15
lZEk9FO5vHjgffs0TZ3heGUJOR8hJWdpayLj9YzZmyIrSW0DsRYIVSYvqvCh4lkfqrdVR1+lHsFh
siYHd8YEcPQVKTdchiF6BFouC1yvePtVuyBZ7+1SwmRtLjoSZSMG1DC9L9vbhY2HGrBpoBHdCiqC
EzFQu8ltQCiMl7Vku/gpe0i9HBzN0Aj3XuS15gEV4fXqMQ55/kU9gT7IqOeDquhD6VdeHqFnKRsp
oc8sG8FTS+Y889EsRwaQuE/Zu0O6gDWDKbJKuthixsrq0YnEyjY5pWM2/tPkVbj3+eWw1ppWUJQL
6y7iX5bOX9OhU0RMBpOg4QGGT7Uq0v8WEQxXG8NThqaREhqojZatSyFbmJ7/xwXqEjeP1Fl/Z6Jb
LsnMKkmbby4VWMidBhEAdOaakfN7J7Hw7gFOf7NyjVFo7pnTXFimUIj1NBerrx4YTp2zAX3nhrAx
nn1SgHr9ztfQ/x8PJlzlj5dMIm6MbmA11rUfr2dREPqSk+5nto0uXJiZZDgDtCyfmaJ9jsUNAoBD
tUqepBiKAJ2UF8aBbnqWjM+toTOxemAJBN/oM49mjuWGtMnlHOOB1y2HVVZ8tKTeBoDnoICzV4Fw
lBc9jKWNUpJBc5YXZ7JO/gqt8FxISY9OfPxTxi4qjed5prH2ks8D1B93N1mVvblevyzC7oaHggiU
E/A900o9sEfld3wuqzXyb1zic34ZNpee2K1WakpbHjX6+wAfvj+e/Byyn8v75c1gHAJvrAYBjgRU
XzLnLJ8tas4ubuNDdyeri4qjTWMkf+M/8L30V/tt8jBmdnK7lCXWf5JdlOtyX0MOr+RKkFrWQjso
iMJW5HmVpr/Wf94Sh2RHZgizlt//oIAVRbsaAG41CWp7EUdYlbb96kWjeLuy03vR7eCLu/UVIHoF
kvL0oaHy29l6ebnQYYnlNlmRQTEIM2NJ/Fcwif6MzudG8Y3xrUHTidAcnL91iU0IvwG0U0wTMB1u
sfUAg3mjwslxWPsqTyePZBPSyBoe549/lYkFliMMVGYXaJh07MbbXuTs2fmgtocXhKxJ0Sl4ruIt
6FtfGjayeq5235g4jDfdTL6nLuThsyBKyMzf8Rol7WcvqumURZwZbAJJDhAztqozjAjz9WaQwkod
UFaHrYeCIMi3cGMWQdSz4kn7w1RyMjPYqtJ7f6VMlU+5PNYyEq/cOTLSaMaI711A/isKk9ajgZ8n
cyZOtHm/ybyVkQHUExLAgOz99Box221Q9ecZq4BefiNt7NyvFQnZDMMgnfKsiI3t9dlIp6QsMjUC
rKt2iG1KOXi20iLDg8/q5QQLFkXYlpVgPUt/lo8iFtyW6rUuj5q42W/LRfGf/pgeTyUaCBQ01SXF
A1QsJIa5P1QckHQ+B581r9JqW5dTdRB8zwLpphIIXXdt65ImKb3B+aYn8+UVdyi9Eqam7D9NTdqA
kPZ7T8B1Mb7wL/444vvldGInkr9BrhX98uU+2CP/ciNPBzcRQHu4oaqk2BDYb+midfPAz2C1OQn+
wrsXuS4P/1UyhNUNN5A1xLVIiZyTk+2jB5eAXjaTtwkHfL+lH1zzZi+s5GgltdYaYKVqWtgeF/7Y
LPXoFiLoujlXVcaxzo8nJVlEkbw2gpQJVAfzExQue6SInu+aZJ6HA1nY5rIRskDmUhIh/6fFu4g4
Dgw199aa/oP7QHRvYqub/zxpsZ+kEJ37G8ZOQGDXAmHCYVnK16hCEldDijWqwLnqHuZX5K4780Dv
NNs9UKUs5Y8LAXjinHKOzp+8/qTQoG5BCfeICquroQUbC/cKpr6BNhydazCm3Py4ucHducmGZOfX
E3rdpxG1hF9BqR2quySIH4O8vUSXVh4wDKZK5M3qq+kAfqqk/1hJY1d1ovreyc0d/ofzHZDBrVor
Oue6n4oa3BRuuVeIWSbNLc3vakkUoH8k0RsCIVPb6M7qO+M978kwwoo9qFcxT+4E+GrqXM9PjcBv
RNuxjutm3+gL16aZzCU0E+YtDandcGFM/TJvlz7B9PpLK0S+knBXlb7gKrFaIbh1QWgRKQDeyqPb
xgR9Hf9PEqorlFDChmE+Hm1L521HmG8RbjbbyEcEZfStjgN6JM/AtG7JFb9u7ZBI70Yurid/jQsQ
r3hIC6x4L7QAe2Ssh/qjohi5zA2EkmhhaluNVaxwpskEkyHlDePH+t0u9TIBqWtTtGnPbED7T7DL
NxPZAkz7je97RUmMz4BMIe1rElPEK9ZruDD/AodDiql7NIxcdBxm6vUzkoQoZIlFHNePlO2VUNoC
korpX962qIqx9ZTPFx8NuM/gV7+U5lduNgDlUZmjCC3LVkchQqFP/+Vwq+pfpgwJDYcKB+aze2Oa
HM+V+73db/52C57ljrbUgManq3NiPmVYqfpn4NXptpFb5D1IAvw6Amqkh84+37GJSJ9TvCHn9Twk
KKNu3kDgf9ubOelxDF28ylAz7vpJzJySt5nOnnxAxMUDZaGeSWpXUga1h7QmrNDTZxTgTGHxFmh3
vioHzAO9T4igU+oFDBd6+c3aNF+hTHQzzlPOxRnT52nV0Klsw/IBGWovzXoyoV8C+2LoT4NE6ff8
cptF/tcH2ZW/cfD/QfmspzTMTgNHSYrFWXgEr/SnIMz4wo8JU0RECdCvjNxPmh7SCyYlsrhg/7Xh
RP6jdxf8qgIu4EvPWcUbEcUmp1RcjJP92vdU1Jt6Dcj+a2lfDkkY00a/EftcKaYdEhXr62siIFBP
7ELHJRviOtu/bmlSEZRQfmpN+ODhLv/Y4OtWvpTsTYnl08WkPG7Jz7WsV6ej0dhNPKsDkONeU/Gh
e+s635BufBhTBr6ddSt6dJShMipYvUk/s3aIMN4TpHOOmQrWXLpXrlduHKh66jSvc5TNQ+Hx7N2W
CyVUFQVMkHWpIm5WKw5o8Xcn1d8rYqVDyK/RvZW+XAn9DskBqfMMZaS3RgKvIJeC0uD6REoFU5DS
YBFPGRLQWnS/++WgjcQNaPGO6ThmR3E0CmFY9FuEgyQMztzx8NckYYllLuL3B9f482QjJkg/cym/
ZlO7v2EpRrVbyyBcZi2hlk+6HUctC9FJkwYBhB6fmfzqsFgdKwGb4HfeOHpxnkcKbo4YmCdfSvOy
9wPV8lo8YxGcfIjSD4gdaEhl3aUqQjvvVyHxR+muyJgWIjEPPB95yWPNH68pGJlq0U5ol3RmCpWq
oQD14mpGPINYdZ4NkkPT+aGJpah0Ur2w+YXKbr/yCgaRN8wK29adHIVaLzrzT5HAt+ffDQYoofem
OK49/yl5ftQDGZ2x8RBlgD1hAkWkX1g3PFnuDefYweRUbtjR+pO12Kol7wPIO3XsTHfC9aaL1Ccq
PriQ5HJ+hW9OqIxIcfuEiAJW2Gr47LGwlA44nTp6Kfcu+9HMlsfM+oPUYGBNqo4AGtc4ft3yMxp7
AnX8YaInvYPn1ylI0OsbpfsUw8m8jwsL7BXs+t7OZlj7XnSMfSxCdAE4lpMwzmQWwKnWZbiSxHm6
+TYPdjwwHTfmOvkkzddIdPXy77vmWQJQ4KnO9Q8vwyVk9S6ogCdsJL2DiinOLrtD9En6MmuA5ywl
jDToqMXCg5J+uYSQQiwHu/mXJa9RpK04ijCiDTZPylR/wtU2UED73PwEwsSh0tKY+NYOYnPmM5A+
WEOVuvkDAX4ceJyMf54fCUkmogY3u52s307sFQQFktql1KZ11goYacdhYItx7OoyFh8qsp8EMRfX
ijw4dQGVnb0/FHLwCFg6zXPcmoE5a0gxYWQeGlIZBW07HPloid4Tf8ZPIsUtXZfBdB6n+VlqWHo7
Te2KgZcbUtX8g7mjl/ZZ17gBV44Y3Eqag0RqpeCc0gjNT3chlgpkVRTEJXOpPxqDYhI5jAm6h0xG
yFo93/WrImK3nKnYMc5UdbQProyskRC3zj1L32IlaRHyAFDhpuCRZ0NY8DXpgzgsVTS9JeYvpmjU
11cCbuN+enLn+ohBG0RoWMSK7gxBxd4LVZ8dSAnMzoLfrIavsLaPz3Lqu7ktPmCE9S/++0uCOwwe
0v6AQienDVEDHKGAn6/jbyrWcaWD+iWF7832ockTp9LhAaryJ4ZmHZJiXDaEksYPOJrSzGdZ4vYe
uqlx2oluAKWWeEScPfl0maE0sYzL/VEEQaidMnbAVPZ2kNyqj+SS8ySM703pWvZR0p/piML4+Nee
QE/vvoa0kkWGHpq31N5PZl3L8OG77aEFtu+PzY4uOh5uxx/FhqMDjHB78J09XEuCrrH3cacG+vel
Fn5y35DCFhJ28vAwPyQItNaTo3tND21uP5VJkiQcTFohCQMEz6L7gRBj7Jf0gCnph6p5ytl2qG2Y
jhegpjDBeH2tCB/mzMUZtVZsNGlE0Yk9QwP0X4yP+PBRASGz00IoH7WgtOWMREqSLiikka4HGOUD
XgiqrRE01HmAEVAbHFuYu2WGXPj6iPYJ3egIZ7M341txYhpkBZIyF9MS2t74o/Jdof038yHFTjrl
rgmLXbubDnnHKQgTcaVT8A7vJ2ATLf0e3svRfGRu2khDy7z9DWn2kyIVQgKS1h4pOZsH6aEoQwgt
OBCAv0cta7dyy0TMTCxD3V4MuSZxm5M5lDuTJJJd0DgN5ghhwBhOV7oa0UftK8HOTrjBdXd5mYmX
+/6rhl1C/rPqZqdVCCxBbRRnU78m2Ro0KxqLizarnG46QwHz+QNCj3mFULhoqY9BHp7eTfhVQyVu
o5lGJ48340IJaCri88m88DfDpVb/lOpHAkeLbtWmNxYTsfWCYyhD0QZ6L/lRvJEV2WO0JjZongsp
bm5FBQhHHHFiiXVTCWP3sf7Z4nMNUr6aeJcaZ+2EEsR3CpgjJ+hFDIxJtpwLlmoU/fhGUE2YgT7l
2xjZIPLlbyTHCqVpuH6Y0ppcpTb5mKUY3aI7zpN/jSYzI6f8a4s0hijBfC7O0uQBHqLAT+tRkhNd
Y3Xrp1t75SlZlCb0aNPaK8DzsVp0ftyxnT6uHyDAzkE2tLH9fKvFfVqj3NbEKDhJvC05FEe+fk1Q
7/a+44yYvAgk8/aNoZcCDDXAyqZ5b3oGs26/sUHNHLzgdCt2E+Ca5ZRTB8akmKuheqSkRkPXcriT
+VPuLwsDGvYQZduv6j8ZZQtzCEs75sosFMNutLdnUe0GD1w44Us3mp0OVXh/sgX0Cg2C1CwgkyFm
zP88DUiwuUI4Sw0bfkOGoLi/YcDLWAVdjZxnbXbqBmb9JaU8zA8pzhUcCSAMKXosKAONsi48noQX
TtB/5aELtdnT7NMTN9xNJHIWkw5JlgBxMmIRn3b6cPu6F2nZaTCJ4SEnN9/E4qsEvqb6TpCgoKiO
7wAqOFVz/47u5E1CL6d4qhhcdxf13jbz3A01SURNKhwEWg1Vrwh++7TaSWyAVS8nSL6Y+i4gAJJy
tdkVaBthKt4g4JRIY4zwH3nd1wAyuFrXNSRAgICMGYL4t50bwxhoSI3/Gj8NhJ+zFZe+dn5NW4X7
L6fn0IZ3fhuUMQuXTTTL1Y0nGaSde0PK6AA1ySk1oxhk3NgnUFVbpyW2ePChZqUH0URWBWhtHpeI
K9sdl5cHADSTCnVWcGTKBBJU9M4naWq2Ha+pAliXSOA2H3RDxX0dfHgQMoeoZpFyYWkZJm2CbKAA
Gsd6JznujtjJyZu+al0uM52q0bXke7Yxddd3mLxRUsZvbu1Zz7fnO2ZFjyQuPHbjBSpAlqb5QTFM
kskWDe1ja/SLlcJ9pEYYSaEZdRj+o4Lkt7NCfsD91OsHGPXwVD8yqKCnHeXHZckB0vL/IhUhDjoB
NRiqETbyGopdUM4n8SDq7PcgS/EajqDo7IekrxCHCU5NlE5uf29HwNJ829iDBVHiDyPUaKcvazDG
DueqOloWHFRPZ6ut1hH327l9HsP4e1NJypYlJoljt5NvfIfq/qYZulJdP36UFT95LbBOzwrsbbIj
4JBwYVbuy/lunvqNONajB+XTiyV87Xw+L9cyNkaGUF6WQXlGhcRYed+oC9W1aSelwIkCVSBZyPhu
vD76fUprgfJPXn0UNEvWNqE183rNXds51YBVZG6XBDfiF37KG8/6ANy/94s5omLAAnoDFChY153K
DocE4riyaDCa9chG/RegFUg5WB4mrE6j7H/MWAXUMi1p1PivfNBUSTiz2wrsnt1FSspKp5jxmj3x
9M1rQLfihaUn7utoNVTQqeb6dZCyKht4OKx5/X2v0r17wVqT+DpKAq15ZUS5H1U5uLWkLfsCPO2o
Vq9OrGt0zGbcFfyXa1UsX+UELEZEv7be4R3mvn9xTg3uGEZQoLdfgaEmxAn9M/6tJkmN4Vw7enAY
uZsq1i5/IICBsrX93VHlXSH4HWxW3dElT0sqPooctYZqUR8ULafDMgccaeQ30pUF/ByDxV62+mQW
xPYqB92GtWAsuOqj8QocdRIwBVVPNsB7loYRH5aCPMez/+VhhiNQy9W/G+U+3EZ1n/8Cm9JhX9Lc
qVIzom8KwoKa7zzvZK+duYSMD1hY67jLYk0iVlwZhIXQrepCpkl3RSjpi75erdXlcppDIyIwhAiv
+ADhT74q7Eafuln1kue7LXmJp6QvhEBnh6gjxcDWOn0M/+dT7Ucy/Bt5N1UerjAZCQZJjPw9GInU
IPeERvY6pjatVmpQAA+47w8IvRoaXHUhvz6u6oRNcYVqzc97Zs+JL3TG3S8V5b7UJGnSaoEUSWo7
m+oZ8pJ4PoijkryywL+cbCa9xzEwolXXp2r+rCtb+/bOR8uGb+8beLZaAYYG8ESTIOgQCZm0th17
HfvzKTcl+dI6GjC7WQg7ZYx23NJZnlQiUldzHMmn2irMIMqHtNqWvBl+2KAtroVfDwyHPMmkMtXy
mYsMbCb6dV6PAuqZpVzJH6DRiwyG2C07svVGL1ikexIYuC0VVNNATW+1erXu7gSr67+Yt3cXuIcf
RFnVmxkMez9xDl35jrbUqI5I5dBY9Jia7K9OGQB0Kc+aBoc6HcBB22uRANH1TDGWNSDBwuBchHOZ
KhTzaz/+OjTVe9tosmmWUpTwcojtz4H+OiMjdX01QhEGl0Z4VDyBt8wMF45dS1L7Y5NGggJWVvwn
GqrSDrt0kyatzqNlhXNy1E21e0uaGbTYZ0OzjPKrVcU0SwmuYN/4/lp2aUXO9+We7IcDVq/to+pQ
165L6cypjwO2tLX53nJ7c2PGtYKgy/y8S+EnswEZW/MlHuhmYv4zvbuzugTUfkWpAz40WXqweiFr
YxrVtPey8eQhikNuXW5aOuB0gqJA0LczJHHIAPZPO2SauCxdNJSlWrDSCHuao9yRQ5LY+WM0VGoY
rI1ZpaFHAwhhiicINTqqWlFsJeMv1qv6hJM3qMJIPOuq/XBJhddlvlnY8TDRzxXZE/7sa/TTEGhV
JbGHbXD1gVMz80/S/g60BEzN7cjpshWxgdwXd120jIuwXmgex0d6Pr8WYAlZEppkJUbegojNkR6W
/ef+QRQPgQM7lVGwqrKVhpGYGuRDgVlQrwdWbAQ3pGVN+i5GBSXiPqFZ/9gZYe4kF0ZQAXQl9mHq
UWtZQZVahWXnMNkfA3liT3zifIerGyANwfYeNylFG2y/+aPDQzMNMyJMfeCFuOEPZuwVulWiDf0F
N/vl7C0N8ykJv88Ye1bKn0+RFYdPcK3vQPpfef+fErcV0m5aNr+K8pVUOoo1fNC/v1L/9e2YjXU6
p+hIfHlDN4T7rYohtlFzHHNIEDPv+dpoFa55kkRSU09ePRRuESwipbqZucd4bcqVL9wR88dKGqME
jYrbBzKvgZbw6IGMD3wx1f3yDgIcs5HJ+B8VmtFSl+O6vfTiuYNR/OjpAADtQITsksLaLFqGXhUB
1gjKyWkpUEZAIqp758+0slDn9mOGZOg/Jdhh5qBlk9FxAxJYDJh5ewGbo/rT8ZUXpMTbIsesDMcL
+9zae37HQyHhgzo2vgHHXRFpfFMVRqJsw2sm2NTCaX3oTiKV2W5rIGl3b4sxEXIbjcWpUXmqkNzh
4gKGo1+HEtmEb9tZFs8PWDwUFuNI4gfCp9GhisGvHv8qF8HiknC22AQWUFB5n6OgOHgSPicGESsj
dII03WMmayGGpA8in8gpWKFi0xUucJvwrIGBH4OJasgXQBC/4GBZA/h0+VFpAdLr6LXtH2Q18ok5
RB/7bzy8TYzLC2teMaiVD7FvtuxGiaoFcVrwcMHk+tv59YgFeFehKusBB2m6jtuSA2v//uz9hFBS
bdZCz+YKxxzskpsh8Cf30v9DWcoojpR3h2g+OuyXQRfFtC1DzcRvRIayOUvWGjtT1MwxmW3hXeJF
fPoeIElCrCF/PaDgtwjwlCzasTc2VoeyWglhm9a79R4IgEK3/be9tXe68SiqO2Nb2sGTufJdOwnr
6ixy6ClGHJ+cE9xh+TN3FMAgrh0SYeN+xka94YDBN0gwJdHZp8E7oJhtlDcflBx7f6vJjCJM85wn
3ZxBv3g6aJi+8TyweCw/04A4FKPXn0R6038H4DrOEXo6dblTE9Cf3BG6/okpZmb+Y+SjfUOFAMhy
I2rRAmS0Z9tt/Ekgjoh68f0HThNhsNxvdja9fKiBOSxwQyMfp4Wo8tG1C1Ktw2/PRTj6HfiH0wkc
CnHUdYVGkJEpkHAYMsheym3+zroRiDu1TOFPj0b2IzhqXcoTRyVdTT7eLos44BMWu7MjreurSXkV
P9qo1LNWPABS+r6kiUY/+SRz70BBWerg5ctKUj82Ro7OQWS22dqaAnO5eX8Ijx9IwXDnfJ/ae0rV
S6KPSa7lzBlAzWdvpppD1z48vLHvCsiaObcSK7TBhJ10dvCqGyfrTMfm/5Me1uTIliQo/KtsTOp5
uAtpqQ6KzuyS6B8i3dtKVk2/dVUqPefhc0Ss7d6LogxJ+RyWQdsRSbZIn/sJWVpYUZW0Kad57rv2
RL5YwxFzhsWiRmF9AY/5ck0Uaqs3FUDYXn0dfEjIu3f13oxBbtFTZ/Ea4OJXJ1eNAbMGqoss8nR9
Ztzg2lgNKCpwRqwMYzIuMcheoaZXZTVmnOKeivWEsrDhy2Tl7Ey053hT0OdGvYZDGVLjk0bRxmHr
v+kRsuuy3J21nj8Yf5GBf5wzHjCtphbIG+w8DSQkGdZOBg4cv7mwqIIjBXZVCZ8E2i6W9qPoq3rw
wo/G8qLGWOaox48VquwX/Lb4zIErlKtXs8oCygF7n8SvBO/zKeXDbxttRQn0Wezfn5bzr2UY6+jx
ESjkL4u1Y/gKkkH3G+BQR6e0oW2wz5dKB28BloSG+J6CIqFs4zpqa+yaqeVYSMLo87QcgenZUK1X
/VEjDAjMXcrW/EIWnlnV2A7keGRZFUJVjtayMFfmhy+6slsHvLKhZAMXEkJDCZKP1Lx8S/dKmPzI
xt+NfOzRvc9E5jWTdxhHFODMOUz3C4Ubug9wzP89ir8VFCIgOIIuJtYWBpO0SlE2luFROlHCzlkV
qj5pP3QZX2k7Xn4d+rZ2w3P0BLSZuIqYgAe6rceGUUdOX0RBVTUXZ1zrvovAo8lESxRe4Waz+FDx
iVVEojc8c6cFHjY5fpBoZfsCvFZWaLnilHOX2MXXHE4dfFLrWUQ76JylO0HyMNwlszanm2wA4l9H
3E08U0cJY0a/CDQqRD3R0U81RPTdJ45de3R6PiTxgnLE45I4umoKH2j2lU2qiBkfZu8/yhGziA/J
3dkh3VDHunGnNgpfCvGa4e+R/uGdXg6wwE8ULCcvsBUWQkq+yGhZ3whS3s9KWqvSShOJvA0fB3Ho
cxDRctRbqUNUmu813yox13L9utvykpcrTrA/EHwHUEE58qQlz/6Dxf2QOssmd0kY9ynbkJc356hC
c3F6FZvIXZDgp1DWlsNzqaKWpEKX6Ko7tXWs10fE+iBl6j+Pj7t2FQBbNzx6DsO8cappuFLuxyjD
H3AJPRVV3WRH68onpetp0wYDEL0WWLdi+02coe6NwvWs44B4uZpilvhJLZqGdyndFZtdwvEgpxFK
KE8PhtWHsC15AmjTyIIJ3FM/gLXC09OiYpqqyv6AzWQ7TM2ionTNUSf4IVdi90qExHo6sPSrj+5w
Dycm3rmVOZJHBlTOtD/gQyPAv9LKvNQc7DT5WCRYf/b1aZ9pRL38jlbm76BHmNeoneD+fbA9HOeA
h64pU8cwoApZxRUpHR983E/PIz/dc6W17303koBUzwlS9tMvOTb3E+IBLVKNWnWHIDmO6KnUu8zn
a0LgqLdBRVUFtYPCnv6QN4muSnusy9rLUa8DB95d+PRsKGeLT0iH7dpjKwxzQmzCl6CA/W28XcWP
xWrE7BMp5HjvbMraYp1HdKVTtVI2U7X61M+zD8a5l1LXHi5JEIT7jOtTqVopScBFquDDJlHe3Cg0
4TepUurCQEEJwuUrOGwT3V3BwLslBm6XRQ6SexTrtdHXPIxVSGcma32X2yPQHpe2JLIenbtUOq7K
9CxQHXEDeydCy6lRCFEaXPLxLpr66yJDPB44sYHngwxkgRjEmFyueg9sVAv+KmwVrNXcSWV3QxJ1
/hLdENrxT5Dw88FbD6hRSw55vvq8zQzjHwPE3HvnSJ3oeD7ZEIP/fsrKhmaHi02PBD7HGL8cSrUB
D8XQr/KR/EMf40xJIlI7Q4oKbJxiqsFHCVVDTF4fJ/i5qGguonNpipY+zaIyjZRyR/OyhIDJjaBn
+LXUH8yJfXVjzurEThsqa3DlN8kUbvOcCxFlpAHvLXfUV4jgH7NrnR+9rb36ChqxAPTdG+I2AarP
aJXErELo/tYhQB5RTwXmUod4Wc1+0osiB2wQdf4Zo3/BDQ1SymfdyqKbx7oaP9kLCidGw0AwimFQ
S/Pq3LnExMe0Fk/VQ0rVhDibPDyXZhzG/h1D9ozACjXc5Jh/kpj4SCvJvUNT5QPW151XhrPP/0Ar
g7WJTHXZ2yajI7DqtsA69HEuvV6uDV9QJ1+n94HReI1hIKhCY82BJJovqheyqndvdTuJOA+MXG9P
iR1ysg/ug8VOSjC/ZafNkfKpt4VNWHLCoA+L3Wy/dmtUUqyFoLUjCuuFZRUYmtxcFq9yhy3qUl/D
D/0T1UWyxKUZxiPa1AVIx5lqz9ZqeRQAVxTpt6dkkm1fInvFINqL8GcjiKcdeNJqxPeZKboodysr
b1TnzgiuLRifsUkynRjMUdN0ofVURn0NJK4UqsHxhr4XrzGRWFGx9GQ6NQlb2nPxlfFw9V+CaZxu
nxqru0b+b9Wi7srAb3l0vOLSXT3TTog0MMJZK11X/w+OLHgb3IYsTXuU803a2X0If18cPPUHit5E
1Hz7iOwa2Hvu+pfQieyRcUhRHEedoiY/1pj833vzolKGd1uT/KVxYAa17n6HWtUScSp9Frhm2lw6
vxrE/dt4nJAbBlDKrssXWH4s4JI8MbMoJI+0HHn4WMKiZwiLjzB1l2YpL0uWK8NUfPvOaC9ohJp5
1WXAbJoMH/nGB2Q1pXCmmhrGbfe4wFBnoXz59XK5q0tr00zJsBrJ+sm27YQ0I4iPjgiNm4zShOip
uDJONGQ80Jh5+5SOXqf8mRf21RlXil0aQYkapS7f0LEueyHfJsVo1gHDk4L7QC2kZPC91q15brCE
pvkMxaSmauQd5MWtyktKlVQcrR1DMmmJ/GrF+JxeLii+HzMMBz07B8OT6dsJ39Ap7fAmpJuX1slV
XmE8w2XFMo05MmWnDc2GTF228lzPuG6uKmkSiwkbhTDFgwktFCvHEIsCOU/ZFhIxYEvhR/CGkr1J
6TXm4XDScA0CYUSco2lIH6kZyjbAPb7328kq9NNS03W+FFubYpbwMfklvRUImNs34h6W9pl5fs+K
+m9e11yM5shXqCQN2yGYTqygPsPQ6i3Z6zLWnosWStSDWTXtdBHOon5n1XtIqbx3J9f+OWdWJTYs
ExHWYVxCaC/AQweJikgErCreBhjuUfwIQiqwh8HdI+qjs4qM2OrE0Fcdb/AivrXju7lzWZP2kGjc
uJbhUiWcso7LsPwJTu6ZrluzMXp2m6fcBrS4OYR6XOSTOID/FkFYZZSLKlf9pE4l1MKZ4FYlbCzk
RbFvQMtrrIPaUuTbq0oLPEew42+k+GKVabyxCT5hqcapzwyAk9l3+Fpc5YKL2pNPLRDI3p7x8RNF
ogfQEh/c6W447w1Y+XH5E9U3q+Liej0ffjSq3plTcnaMk0FnDoyUGbbjKm6eXhvkzd5BRiGhd8x4
Ik0trDf1NtX+Yctvr2JYBbEzI1p5yE/vY4WxfM5APPgify6P398vaHoti1l9F5wOWSlUEJtS8sYu
l51oNpgrKoCd/YWYwA5mWNcLWiN/l1vmJPIRWfGhuF8e/kCfsJAo5kHfM7gPNhr3EMMxWHQMtxLA
Xvn++8UJbcPxEvnXeMKyEdFoxll8JbcN+MRUFJEgS6kyrnzj/nFsLLVaw6pqjWy0x+lqG+6XWfUJ
BCfutxHMcgcJtM67kHlcBTfeg0RsaGQcP4MmeTzPoUN322+OfVVL12/W5P03m35QS1VpzaF04V8w
IYuB5kMd9MARHT7M1y9NxMXiRa6YWXuSv0nPR2yD+epKWHybK7k2DB0cR/1M1cg/YOVNUp9SxlaG
+MbZqR/Llw2HIIVhmbayXfp43CyNhOppbupnPeD91Hd6oWsm8LXz02zmI8sqQiscRmT9gDkEGsG6
LddQtnkLbaW4NOoIscEfIm7ZlEJ768+r3cwLknuDwgnOjv+OaZWLfjC4/k9WUAXIvE+EwTtxCxGH
DT6OV5+eYjwRPnouOfDnonl26X++Q/KqhxAL2YYPLvaJ2atsolEW44XI7rJP4wC/AYpA9Pp5yIMD
rcEj/hx8npQtjHUs/A3neGlDzD9Gt+/eqQpVZdAsU4KTtbiVx9v4xfKGgOioayWoS/1khNPoUI8l
042+RCaGHQyPFu8XAjA/OX5xQrY+zreyx9FEhZNM8mEt4neOSLUAopPUYpVlGX/eBFPcOLdSxUnJ
d7E2OzL8McjRRs6x+KvPKtBMN2giRwkMiMJhRj/Ocn11tmLbH1CvVI7lb9myG2+4s1nmrjnTRjFV
72pyKknLLV9OtS334AadfTtPhXUmxp2tcGY6Ux6xY5ocyL8806u+Z6DdhWVOP9a7YWJqEJWcl2Gf
XD1WxWhWcaxzCyFFvhSsMPk+Z9TQISkckjewjwIrvUUDETUJskjp1CJbq1wyHEEhXZeyTo2KYIIx
XDyLqf+aaUQM9QuV2DsZQ6nZ92NG8cyVosBObjVXP6ya5jDkxxMxvjrbNYlMxW096e+xbAepKVcQ
Li6lX857s8T4TMn6ZBqytvkjwvuT7nXOj+EgdTW1PBlhXWs/VH09Hcz/TVIq7k/IqnpcLasKjTGu
3RbksHiEHu7/HHVjj6vzngvPcB4kadnmT47mR4QMMWX/++IRerBJehrlGmiKKHVaDerNo+K/1VxJ
FUeJ13d/LUz/5TFF41xH7K3mxGu5m7K3e5qAkaO0+M+lPuwDDB0WvF1RH7xmQ5uv2QkecHxSsJZv
PMrlL56XwUTnWKvx/cTXNCwKgZqS69MgvezTwEllu/ksi/P4CSrhttT3W66Sshbfg7eBTCjZ/ws6
FVBaoK/J+c8hDqRntRt5gDnEkrdRCNV7KoJkp4dOUStJML6Jh5UPPtVDAbb6oZNoeporcEEeumQt
EOyhkHcI1qfcONXsVWqWzbCzyu2FkYQhxJe1JvawVq+5tz61UKlxcEx7S2No8lHLZiYMcnI3sZ4a
as+afq3G+KDzmcQQtZ+G7awEdPB/gZ7miJrucFvKqqZUqxCLAQPf+LfITQRC3drLtFwpBwI6yFl5
yHN8pPjpxLeXMThfxqkAO1ygumaKT01wcfyXlGf1UfOthg207f5vsGT3BkK+IWzJjPQ5gp9bTTYF
+ct+B6WmKRvK6nRhLXCChEYFcrVXrQEdc8fQ/LGBKDRKrndiql8xtmV57NedE8jMXAC7pre2gLm5
GdtinYw+A4YnaSXdmUYp+rNlZHEM9M9yFbyY7Wje4WwFSf8BqriQdQg571TrNDGWry6GzdDdAZfY
cfUxBqYDAqCe4evVqUh53daHnSz01amKiTejeblkVVx7X454tBg+QmSKzOUT58zci+WnozGL2lL4
nCr9brqKHlYdqx1rxsgJGPxFp+4C1v+hK4KlvSQgQp/VkzLmDLsqWEzhDm9vhePLCmKw+ToRbIwf
3j2b0xCC/gYN8L0Exrvx1GaUHJJ3A0QZ7Xe0Vsd2WtCwh0HR99IVYTK+f3uRaT5Aqeeh/6tbeQlC
ZLTrfULjswN6a4TFwmW6Uhrvfso7RBcSrP+UQe0CQ3a4XLYYPrGWgIxK6RpeHswZXXwFCXFA/wSM
P1m6/5H1Rh7t/H/BaKswJ74+EnEKM/bn7iBYV93EkJK2bRF919bzpIdXz9WgpN1E4Tl6OX7Z8jjC
f/lOM4YLNk5br+q4GkGGx7zMjya/osdbe2BDAn7bH5O9wIQVu1w1iZE2UpRsT6sJQekeZHI5Si5Y
pcX1vhGJnLwCWm9ik+Ez9VFiYGXKW42lXEl5k+oZNhUVGuc2M7LoA7zFo/eBiD1Yv7A5z2iV09oD
5IQtGoaJKSGGyfgnOQrfW0U6A+g9xv/xmw9A400ovEsHjYNmtpUp6ewBsWMf60+9axwnIN6UTj2T
Jaf+buQGFpypKSUSPECU5DcCrJQcNM1zrtIKe5sVzpYsDJflrQKsuTW7nS7kVvoDMP3y3DQ5P8iO
yeY6sH3cXq+AV94Xogjry+JPHV6ZunsNV8hjp5vnXNmf7avyXi5qeLxve+/U6WCzuk5J1mHHlrmE
SuKRR0KnLNFjAAXPDa3GhDTdCj/53kdhyRRCdFWiDOc78TIx7dE2AOXzDP9BxKwDXTDPe9Etjp0Z
+KZH9cBxHqNaPg38e3tR5c3cHs7Pi9QvN4WMTnCQhGrZ2aQjOkKcSfIXjjJV8pr7L+4WOlIRBTtR
pOFSXXdXe8uX5/E4pU1wLVPot4L6DtXvFuVuYO6ZwONm5MNLsYBK9NhdraVxzyaqSBLyQPwIPdG0
oEvSR1GvV50x5EwfiRLKWvLL1DIId7ZLjlvXRIP4vlqQ9R8g4N7x5Oln4g4raJ01pLPbjw0ggOnZ
0C1ITRmToKYs2eetwnbhsgykw15LnyHGwD4pmu+YfcvEcp/cS4IDu+nX0x4w06aKwxr5wwYqpbtg
hl9Gkvv8iavTe2UeZn0kOYcyKYYJdl2H+sxGM1nFPLKPXvWvEwBSqZTZiKWad+Y3FLJxiR1a6Y3S
yNcq6zb6wxjjpyWfcDvG1OtRLkQJ+5xNxl8TKPcRIk/FeWu9jk4W+x/Y49f5TdJ2vtBxO0HBFkfR
WarBwQlbkQE2YSIK4AjzFs1c14CVp4cD/vlNB/49U3sJ95fj3JdJJpwqyvGo7wG0FtM4kvbLRxqj
7FDgJ+tZYTQ5Md931MZylUgiiq8VnbGHdkbH0LkqOWBVCFMNquzpZzraME+Gpx4dL1Qa4GdxWaw7
pAquYgwm1qfg+1ExcKJOzHxEmDkMktpT1RR7zsD44d2KiW7Ydbt5eHe6PzoZKkjOw0kYSZuYGvSR
bzJZGpakQff2H+bymt+SNInECMeZ3Fgk8EHM02wl7z5SCQXXBnEZvPs2uiO0xonOxW/9M6/5ROMJ
62Qh/zJI9clz7lSiP/FclXjY1wx5fi3VvV0df+w1xLijEG2xq+Y/X0R8CVUN9ETa/qzL8aA3lJbg
WKeqKHC6ZToGrmD73W3CpuFi7yQKbS+E+S/+HEi1MsKIU/dWXdUMIA59+xjAlXA8TFzH1cM0HZOg
oUtP0QAvDtj5db2jcSkvp1GC3psZgVNUMlurD9t6Q6kY0DXV9Rv4FWGnpS8dIoEf/fM34e0ICslz
CXdEa9+puFX84j7rP4ARQwBtGUARAxJ6DUR9jPvddZjq+uEHUZlbjjQc3oPP2NUyvXCSVYzMJZSJ
+p80u8mumyUS59kbGEFQVrt/QPGrXyCmz9ZAhvRJZ2UC27N3CoOg94rOa1d9SUKcoud69Dtqbwlc
FHgPlka0oAkrZW51QlCnKf1iC4L3C3Y+liXqq2LrkLFnivoY6BtIxHlrXiDwN4JqSaJhSUgNPtXM
dWWzEhO1ocSNEe3kej5MS+Qtb7aLhOR8mFXB5kE7+z1fguHVGD5byDsH/mZuMpdzAKYMmI69/4F6
MPr+v3MVx0xxRwx7UPzBhwj+kUa/ib66s4MyYv3JXdfQsjLT45cIqNP0wsPdW+L8TwonrrEaOWYc
gL9eM7/++VYpYt4OQl8N+RenV0SggmE0dsLa4WvIUEs34It4s7rSmSMX/ic/4RAp1z4I/naKjHvq
1Kc578ymv01H5aeQFUH43vwogIRVMOyinL/EOQv6Ws660XZ6sPHZl5E0ztyIweJIUQgWG2CRhItH
uSzWd+8UwabZu01DHV8DaXf4bG+cGfW8cUiBgarQv1/fk+HV5C8ifwWXDCZFORPk96F8scnuik9o
OhIpx74Gf2KOHaLGpPJXcdERiA0MyjRo0fT4VDtl8qY7r8TTWaU12RDa3/qpw3zUA+ISmU55a1H1
iQdYSb/xSG5iL7q5319UZUs3ZbfEC/d2W5jgCNUYNUY4bbZTEJiLaaeogRwS4gCygvha2ifOycnr
St5kAAH8rmyE78B2g0jBhOc8r+KiQ1jnRJh2Ym14QfpEiptJVgoC4S0gUXAwRXVCC8wmaEyEwq/K
P3gBOaeVgLQmxkNrl2falvr/Z6gLsywYKY8+GFnCytD2LkkLUyjV3bN84K1Uz+tPWV8IMKVadG/k
Ht4k1YWikVVDQidXeVQrP01KozNRd9l1HGPAA20M3U+47jbbecqrTPMzFNqlYS3EYgKtBQ7iqT2T
W42tvPAHYkumiK3CReS8coETQxYeIXbkqsOLtgk5q63NgsXQkd1OSQOhh4/ms5I8JrVz3Mq8de3L
cE3PTY7eCxr09AizzUf2uP8wyw3SSK2eU3fgn7797z6tjuJOR15VO19W1v/LVCh/1GMhVkDCKWjS
rao/zJB/0xV6boV6XRE5SITcBVoId4IsYZvv8RgKvXdDkj7XAObIEgCPvtRG4j2X3kUt59oj6ybR
LHx5d4fe5zlvJKEeQ2Ha5sx1hdusCM622sgl7rwGBIVa0arQyf+Krjdy5MfkYfGeTGW/1kZQFfEz
inD8+bO3GWbeYq/rvkrNMAyZoG6Kn/nuVC5Csc/5AxRkEb3mD2DjuiakH9PxBvUT7fGd3eLpS+z/
V7JyoBkbVUXwEfbNUOkylGqEjHtmJ41nnRVTFYT5qghoYrAyJplQ+HhGI7Tth/w5cfWT6lIwNmhT
50PlAeHTREHxdDyXAPX9xtIlu6diQSJqNsgCTChXleJLYqOUjB3jin/nLGuRQ2E2czw45zuMsDk8
89uLlDBvgFUt1+HZWnoHkbahWiDr5hMO84r2vG6zXZkvNBv3nxcUvbhrHug/xbOj4fbBRWvQxpT4
ld1IUkXMZAtyLKPEvn/SdsUxma+RcwcbkmHtk3uXufNaSnYA4h35jOJShkglV6V+0GPna/2Bwg8B
YDN76vNDe09T3QhpV4/spa73K68Iw3Ys7VroKwwukOOUmURZ/xRQuqjoEh2qelHLjPF/dZDxH3/l
XBKHOrvW2kIRsSLezSIAxYjWpNxk3JsIOPQmEUl5J444IZbxHzjV5KQbv0IRhEE+YXFoGs6zaAwB
IUdnXjw6pEMe/leRhcC9ZUaEmivW1h0A0I9I7bJGn0iCrdSrbJ7ZhKeWTN73ABgzOAEVf7KKERDi
RrdOlQ69m06THu1YeRo1XQUoCHVQDGRXlAbULAUUTtlIVMUyhisuNPq/aHiC1pYu1veGZ9CqP6j9
vTtNOjoSK6wO8yc4GiCq4s5PN+z75bbm1hvIYpYsJ7OMgaf506oEjEmjOEIwxNUJGViLgIHcb67g
C7stMQ7xzjY01txmbtQ864UwpIPflOpO2QADHznxi5gOUEyyB9OaP8TyuFgHV9VAvuDrGtWIvcYi
rr16m723dafErJCKb+U8OCMPJGOJELI51KFDqmhrTzxAPN3xXh8JBVR3DzvWbdR15NK3V6UHuoF4
Gm4arrLA5RIweJEQOcruiPAqceCgHAyj/A87R2fvpe5F9otsYgVCjzp2G+Ona52ZGxK4MzbbIhj8
0l8aWqEP76qnGuOEN5vXtmf1V03OxlNAn/lCgdm+iWr5mcrhTm4ytpwBzYSWClxCbEJ/0S2fvcC2
J7SwVNt6ZtHukNOXyRQIfg5AvKsQsLScAR1Jyje0wIh/7ZcDl40jVvF+MMPez2k9Rbor7RnDD/bk
uaWc29+DlGIrprgdl6/ovTAAFrRNe+txJ9Nb2aEYEMzrGOdtTF6C6DM5BQlxJPaKdAXGJtiKUsR9
FQBYZMqLI/6bmFBuQvZkDI2th0zwGrLa/s7NSk9Z3OE3eZhkQfdy4PKP+thj91Votjlaic0ZxpJC
Wmhu7kC6GyQwGprMH8pIGYXSoR8dG7xD7jYOSa1rDCpAj++DRDMs46/Q4pktTTO6D3qjFmMZJYfr
ASbdsowjv91xYP/a/wWeC9+LqRnd0386MNcBM5Oip8rrxw1n60UHVyVTCjSWx1/4xWsi4GB6VDTo
AUu1GSUQ8dIEFQgVbr7XCRscdQRDMF4d3k0qes81JbBYDXpz5DG4Gkoc3Sjrj90PccJ/UBfXYCZY
7So1VudLb0ZIeEOw+6vMOtNVhseijYItsdn2ZQbH4JXgd3dEasCL8vHpe6oMoZihXkw9434lSK4F
AgYyxbEp7yZ4gbEZRJL3q0wUPudasUFw5QGbeA13061CNLgCOZYP4upcd/wjK3FJEDv64T1Qu/NF
uHkgOYPHeClZpIt/5PDb4ehaCGsRdqeB+x/b473MMJ4S2dAkh5PpRkRF9JG9/w7gZrd68X1Zq9rV
mCul7pGVMZY21z0lc8kulbxFx77kCgzUX2/r55+B+Mno2dkrPVmOr81gdOFu2r5rFf4HwU1cDajg
cjHW2Mp5xagqHpCcdrxk0YmFV6Bu7EuRPFsNC5nNgtOG7iZKJ8uO92DG8spoujwkrmJ2E9mZKZZr
3iiaRrYwCnb7IgYC++ySjX43PrJygJnh6i4AVVDV28+gpSx02A5p2Y+7TFkxn16B2RwpNAj2074D
Si/a5ewLKooTHqt1EdCopTwViNUqXVQR0tSy4vR8sN2D/tR9QLLfjgjRnAGvDvUmDrdYpFL9WVR4
Wj+H2Odm3yr3RMuNxrJ5LvBZ6Qou34bW1IzX07AAxawY9sqFATgcFCUUiw+dZxNjzL6uIMhe5+SH
28tIWgVKYfuZCiTCiuPvsiaMBn7uMj2AOEhe7Rqa8w6ERUvP/N/mTvJJNDo0SF2sG2MB6z68fmP0
Sz+txeNgih3pBy/iKwYmuSmZAHixe8Ub0/n/XjngTSbYPmFupDon6Lk5ct65ASY8zdbMU7ifm6aX
rqSMHuI0lJFJ72Y5UWftZcM4DE1kMOnpHHtNX4ReRmhu/AmTXKLgHRYa9D+HtaB/biaacStKKLoH
BpuGHjn3HVVAiI5kJNgkaRLvBTC+y9kCpw0ZhuB2idHy7Dfo1pmN+WZWOfdeg1b+IV3gNjwlrqxQ
7b/OjC3sOHSyWmLacK9lq7uoS1HX03T66gV6NtEor4fmSMe+vngrv0IaEZLz4eR5ia9WnnRV63IC
pxAZb6eo2LigpDIQ+PpcJop7h6lC1lE9Jkz+n/pF8PvKFq9PuZPulthLONfkm9J6P8XsdjfNj/cv
5cQgOL7mzj23Pa2ugIpR7oV+Y/l0VH7+eNvrFEhf/Q1iNdkfqlCfbm8Yf/GnJyDgIPBsyeImUfa3
uxlCT5EyXQDbN9v/COWnAONrl/KeJ3kXbAmaOxs4V8V+Vco4EYTAWh1kRS9W1OOzI6Sy1wKIyde+
qh3qoAsgeUfwVCBWYZ3mJSwHOWjhqSW1tq5QASH5qAtmK9SClWoUwnx2JNhZialceDrLkST1Lwbk
6RHZ4CS63fG3t0y5Te6/tXlxh90viKRFO5tyX9awpby1F51EhPU/hkSejAdc+l0l0ITxNC9RRRW/
0EX9xfuGaDC2lliT7v+lXSve35MtnaHJSKGwnv0077FzJJ128aIS/2yhMJfevoezmx4OJU20NdF3
kuHps7WTPoQb3Pdl+5YAT0YZvdNt5DTpxqeEmYA9snT8E/+33cXtHgpAs+p3C2KvdwuOPyYr7oMJ
del0CHGGGhAXuRp9EnhrfpMb65ZqfjNsF90noxLDFy9JmftSusXdVUr9mpZTJGPUSEAYT/9GjAIl
uEGkMapv0tHfro0mzxSTwsas+YeOj9UMAHq1J5OGVYG/aNZalT0gNkzkbtaydn8kddILCqJpXReY
2gg3CiBvnPU3/a92jPWhziarCBveg5CgdmwnrbJ9W1eTL0wPaT+viQwj2qgtdvoa3AB5IH2sct/J
aJqFV6NpWu9cXKd/Hw/fv8XF/x4F+f38/NFxIiZU/uw6XzLwKDLLwM+M/7JbvCfQR0GCRKZXzpvj
UCDZITQkfF5g9I7OjxTzdQOjUMEMAIpXlyAkT4SGW8XK69/umoU6hFKIUpFb/Cnt9sL5Hft141Ey
qkMJoNvyUdNRB12HfaoOUNApi2/rnAqTnxtz6QlPbSiHrhDZcYPJSXV7hQIMDLqy32EYvNtNr7F4
SMeHwnxluLl2tbCPTGDro6vurs06WHsT8v4xp7tBWZROjOWI/OjnGsqS75YMd7oz2yLHTx4NEutd
CgIUyFiioKETRc4nyFHbAi5dQ6/Z0On5wuC2vMuwk5qB/rtP11DkzPEbmtDE68WYwoNjGBzp4+x3
SzGyckPxAVW+Asitw9UNmOlGnPB3DAg7knfvQENTSBfqUF9kSjZgB1pLwFPEce9Kb+oPcBITYQOJ
/PzazVUU8xayLRk3SDjUrJeXcfPbgJM0hZ1aHXwF6xxZPkDZNwQ982JWWK2Kbh98TfofvomIrFkV
q3W42PcI2mKKVKaEu2Li1spUrVI7mzhcwGIMFTm2zZjOgXWCLxsGdgIrc0bwl5T8gW1dmN7n4v1M
RQCAMgKioBfmp+ax1d7ucMTPJb2t0IrI3kedM4swZEaeE8cd3kvDM4pjpGnkRgVX6/TT6kQRRW7V
olqbq0NXUxbtF45zWL7apYsFDXThyWOiT4vzly3aGBUTIYo5uxFVR9GPNuAgLPuINjAmki7uWTpC
g53nuBnqhfKUxOlKRDmhvV7qBel2JReIp4LTxai99szfSM2/R3z9L26GWlWk4YkOfEoK2VY9q2AV
ILWYu9hKuzH/STFbyapETZVzf7TixMg0N1/NexDJpX/6zwBSWmpIWMqXMgJ67To7lWOsc6qsXtaS
H9xkhJUKNCuLneKo1FNNXogDhbTsQOssjYFg1exf5uGZTuktSVFx2vs5wdLcyi55jdb0EVKYS4eM
R2X4AozvKKAtqJ17+GfIlKker5T/0xP7tfEppm1R3rF5YsuuxICnJeehR3g8uEQuY6YWZQWVxjI+
Izh1WXv39aD/EIa0mVe++4fc0hY6WD6np48e1lGvliltwvMG/DbqT1MPd7wv8MTaUBc3T7cZ6kiG
Xt8zUj0ZC9YUaycppbCz5HIwdnPRp0IfqTZ8ZnrMbTixY5h2qUI/bXrYAly5HrbR4ztRnqqe73ix
BDoPCNbMYehAtt32e825HGVOZYW8bDhH6NPd6Y7IT3+ySwBBsWizQ97jW9qTibylkZYx+DC52qMe
Q41MR/f4HrQv0VcguObqaWYeoZ/HtXvs/HCR6AXYlB+ybG8r8TsKsY1VQy1AM/ob4zFGgF4B8FkF
jNYTVSBb38b0ecxFjCGKNrPjDsRKeOqNjt083CkeK0JopY/RVEIgaf8cRP/WDgqRsNXSGQb/6ISn
jmGg4akQaADke4ytH8UPST5hHMgH4OF37NEo5b8pvAw989TDD4yGyiPShQOABdkPH+WTS4AP2VLT
psFEO//RWXn7KJbntxmugW0rSWCupkpPssChMQAR91mQgZJhjoDmyhVsE2Ez68tZaNoB8lxgty5/
a9w+ltLC3RFt1Tj8+srhSkKdvjFSvijg50Ixay+1C9kcNlGbyyTtGF49qHG5bzW7/lgoteFc8E4U
5V01FQSUshng7ZRN/vxpCazgLLmvhnEe2JiliPen9XNugKYjpbAgdJY/rntVS44HTsMGlAMLMayB
76XeoKnkkPxsYfpPpT/i+4meVl3IL58rLppJ3X6l+OQWxVU+yYczDZif3jRzBaa+1+Xv6SO876bN
EYjKvj8QpmTuVKuuAANDC0j2svyM4W4srRb07U6f7kmc7IaalG/TX3noEHhQ90Dhvl6KOimBl2Y3
FKOnYkupU+5gik6CdyufCd5TNmnHenUpMINcGjEtvM4xWz+GZPovoG0DG6E785qShE2o8bySJWCg
z70gnzWocVsTdGPgo0VstEQR54fqjL8sl1JJV1JY56ngyse7XJ3X3G/QLnAK48SwtoODJvQc55ad
qvzkdr1GcywifqFW158zW6CS2QD1PAJEc7d/1EthJ/5GEpP+mTpES93Apm9ZrDVU8rfRr3U/l8Pu
iJ+JrSmB/IcnNPkpV+W1tdh858IsT+GU4DbAMblSLNbtg1n+MjR5ZbNBQ0X66lmn7LwMD3A4kxAU
40tGkpZw+0dqdL6O5uXlSHS6ZsOspEuyqf2rwxIAwGPnNnZaRCtVbRPEYMRLK5GV58Fs93xcdSF9
G/xpeBHEtimKOuyyNjnV7QfYVdSedjyNmVNjCcD1ygRdqCtyJL+QUuGJdR5qFmKJ3BWgYi6CgJhF
xUKq9lwE2u87j/NYoH0uZyYBwE6bDZfBse53INvjS+qLivKTeNGD6p4SlrPxWwTzjB5OBKsX101+
OLUc8SeY4vodm8DSLuPmt3YnZ6QC8P8mhEhOl2Jbtre1abaJy8pTdj0scLPza8lqgGtp0zDO2TeS
UOP0nV7CZe6xQoy7d7BkltSVvN5L8YolFq/r7IRYGzGIZ5rbIL6ozWd/5rxS75/IS72gPUe0XWxP
S4eAIWfqV6pXi6suiwY750lCeSBGyczGSHhZ3XFbqn7KfUSQnA5ExJ6LDIV0DyzRAFMcBSscDYa5
aXDMDOEhGAGKuR6y2W5pS513yK79QGUewxl6n9hmvWlZTTNJv6ir7UjhdfLtmazOdCe7J/w0MNYJ
jqlKC7D+P7lDH3z1sF2ZtYpZn3eJYHHOXf3Zl5k82abYAPc0yYljxdwCp9t+9LMD4mibjqlU4213
cV9rqUgOibHrYs4ab8M7yhJds1i75PzBenPyZ54wfSZz+wknskxULVCKxsZObjocL9k0EGMKChv1
D5bmfQCrdTX8g9ijApcxIxLzohNujsl1tPA93QSqsYgcHFcPUjszA2TnXgHDM1Ycr+hKBd9jVeR3
YgLa02zdb8Mu8AI0Wq8iQzle3D75WRk/gouoLfbganxgVkA46+K3fHAzSFHoi/+9fh2vEGR1xTr+
tolV6Ml4cD+aaQ5Rpu7m5vRcQ8F7aaHAd/MQkvXAFpmao6Wn/dUzMJOMH7VWQCyP+QCbMySVy+3+
Io/s8AeRPdrEGfDGYe1qvAe15xZ2XprWaIlhBAANCDItGKH6xgN7DPRC5RxtJQJ0Ctg/f1w/M7YG
dDUOVsPWZksXXpTtzdQj9MB90Fblnwm9XB/lRzGIsUTAUykWlzjdn3KX9H6vWp2ch4mI2CiRDf0H
/rbASiXamzcxMvYUTbMSy9b38tEASgoUw/Izt1atcHaaEGM/0DfQLJd8EZ/MZ9eyVLrIZDq40iPS
WHjT03UpiOlkmZXMJUoeQ1391N1gaN6yF1d7rXwavp+zgSYWJmFRf0KzeKrXGtyDtomm06041E93
rDAGusOGvV/HRUz07B+WnelPVkgL5M84VndDVxPbxYBZWGk25S/SriIr2gclYlTzONrHD8OSMUJZ
pqvRzLdXUC5lM/dnPoSJcYKR/boUIltVqX8Or+XGg8kidcA53hekNEMqxfjX9C3cdW2RDExvjmZ6
sZ88QBhAOwpj7GQCK3Kkj0GXJyIW+2hmVLxjCpgyihU3Ff/ZfgoKR+PmsHDk1PW2cLn9gDgrBmGb
AOE+qexIUCBj/3sqprRMO3UbNw3tFeEadjAO3R4WbS3tsfpde5YImclnj97XKSPN0+pgZVfroILJ
uwbXwmBnpkWe/hyDWVxWYME8cJSbrAtnLldtml0MgEdfVrU34x5WIm5p3IUewQWelLHa4g3eAy8u
+ymTYlDVSCl8fNcs5vCJbeNfenLMZGGGWoQLiEkLUMNLE5CZKMIflXdofr8pKZW95dmiTnZtKFhQ
NNyZeN5hjieGfLnhPIFUVGmSTyTYAorEFoFpffbpZ0rMz6pdlP20Nj+XvXZ2VqPeQ9kkl6a/6X2B
rkT6hSycKKdVYjw+3ifKEeDUPmU5HoegOwAx3HyUGYil11VZGGLWAE16WSdsuWu7areO5EvMkqcZ
p//Pad/P9/EQhmfrdJ/kFIr2NY8PwIYdRUTmulE8i8L2WbYw33OTcOdG2Ti/p4xxIaMlHAS2qBkI
dObp/SKpd2MdbtDa+3O8QcJguQXawzm6ADNj/tS4LfpszuhgIY+hPvtIIW7oHcM+vCxFsWb2SOnR
ARSSk7OYdyNiuWp8yKkdM3NcUvpMdEhRXhJ1aiKuTiCvjFhB9MmRmsQsywFVoYEKZL2YKUK7QuWm
dte/1KJFY96FP1vd0udarRj9deZjs4/NcI4FsNfD1gDgJF70SQ1FRqB3MshFiAzEObpbfraq0lb+
6DxipXKDSjfc9ierQZNs79Th1N4tlYJiiERT7leO34R6vZcKbF3wtii0joGU2I5QQ5jGt1yfDZQO
l45evCAx6vR1SmpaAXAomE8S2aMY7ePMkaM0LPnfQeStKsrviWnsiGbR8+d6aM0Xu5tjzVTdLsqe
C2rN5D+n6ACW68PeU93pBUZ3U5js+1OnQewLUDr5nmJCUaXjvdwiwcLgL+AzdzWcXYSPLNc8rhsO
b30r0ElTHr0AAF0HNuDRI72aueXpPtrUW14TwxGuHoJnjPNHOzHrjQegc6pHVzKx2ogfaNRc00z3
KPdfy3UlVCqpOxPRyZcxiGlDheytsXgWfTNZ+GuCXYZ1Wa5sB0vwdHp6hRU49ndJCkY9W2Z/wsR4
Eh/iPcoxTc5V1Pb2o2cF/JQh8KmmKJhOU30tmbwfG4WNv4l0K10s+6XSFCVY5L3LTY+XINDa5BsK
mzK0+WNZR9a//UfsQklxPD1RPjZl/Z15wEKBZPNAvZFvzVtjyEzzXxqhnoALpDHRPlCaV8IbePgO
HCMGs3Wkn5y9a8tU33B9xZ5N4H0tw5ccdC2dAViFLphdJhMBqq5mM03gGl0LypXPQGrgvFaenqtX
30brF6lQC16ZW7xd5GyfIroKtzh1/pRY5FcQuFCvMk2lpkrjFaAvCu5zpQ14Z8F1560L4mltVj3l
WH5We4Zo5gM3cw5Sb3k33eIVpLDYJ7PSfYimQppyBFYAdhPy5DXrQbH1rOJmPwDyglTSsDqApAwP
SE5ssMe+K4zskQjcPaNcHSwlrSti4RZ6Ut68Obc94j89IQgvIYNDnjtPc0plmta8AtRBykl1S0i1
2ErDD8+4fc5dOD3ihiyM8IFhSYZ0mjdaHQxtISOr77ffepaF7iBM+B5AgDGRKKXVWdkWVIlvcMit
ZFigASo3WP+fklcwJvoeJyVYUTqwFKzOUq6Xia4RB0YLCJ8j8eLoTqL9RjDub5x3Dkgc9tdKDxcX
ADkOFI1bWGl1rSrQoZgKQ1szC1BAWEu0hBj5MNalK894ZOqiHV7gdjjPWBYDtlVlFQkI1NqqR1ij
vaf8RWiGQLrmOW5F483cqE/jFAbqXx+0dWfffMZbWEgIcisLErqGTmOVXxM7oqFMELrVsYbLmv0A
NQ7l2CN8r63L92znRoELLccVd6ahPX1YX5fY9Ut8IEQFHkzQ1U37XpVPsk8XAmCze++XIHXR5D4I
/X8c+1L+qL8I6CxYK2Hvcrhtplx2ykYVseBMzjdtCYg53musBvigpWVRUCXB2o+G+axwAaPbmkpT
G3QjuMJ48xzGI2LD1qUYoI7RWY+svYopIJY8FeVaif9rqm4odNh/4szESXWCnJyGXJ16ZYUXn0Dr
wfEJ4KWSv2+C7Al2+Ll5T7tNRnZsEFQomriQF5HmI69v2s7+hsYFR7MG0A/Ga1qzGqlTbbQH0JW0
nh5tysYJb2GwF3Q0+OF47iULKHLdk0XLwj/g36rhst47eMnJZjySmEYzgJ3wNKdB7Km2mFJM6Lgq
ugSI3BbcHg55maVoy2J4zbnTctb04OzDZb0qOmTOQ1xG3UDTJxxR33tB+gnW49b4bqyMqiSz83si
KSui8M/yhQy7BeywBOarOj52FpwPyQ/0zAnOsNNxgNj/be13ieZlzq+y3W2SnUva1M8uTTL6JNT6
dUZNcqeGEYGnFUxyqlw6uDIBx2M+UBVa9kiQFMkiDJ2v1sQpi36erA7TtXtbZpDtfzAvZnnHJbE5
U0deJUbPrIuLUxUnGLWxfQ2OHx/WX5X7IfWGZO8e/aAGYNy7ku9JZxcXbLoeS7rBdRvw7EcCpKUM
N40bdYT//6PBJWEAU9uJSlFKf3DtSWFzAtdd8l/QFB2LqzewJFlNvO9QIpkdcbVN2UefRCTzCjZO
dQrYKqyIsT5a799Gm7CEEjUj3JyOrjLbK3BMnbjJ+xfjPfuhx709VZ5FhWi+JdHEQ3s3LVtpngmU
MHiuMadeNdbLHSNTf3Vnq4HAHHJ/4NFQlX8LMKuCOnqc1REtynkAUoIppVWo2BoCsUTZVzROJs74
wJRvpXCYSihRn/b6qfvwGZJukLSRuCx2ySdjYBDo4f3vF6k5kK7UsVGuOVQgFjT9tZNPLKKX8A0i
N27OD3XKzqQDXySVIcGmngEu4L8wkegZLUZj05ceYBbHdzDgES+9oBLb6qF7Wzks85XtYSh9RfDg
FbKU7ZGOqTCB5ePCe9VWlLjQn96c4cxtJxBy4Nb9BwGodPQNjLhHj+GscZLT4uy4aVRfPfINjQzz
OmQ0wEKCxDhsScLVR2y2tp+/RDwuy4izdfzOKs/58aictZqBJ3AfIvCQZG2b4BJ3a36Jv6orxKNT
/MzjQL5AxqpC/ikTSs5cKwLlNwZoGh8beJYiD0fWhYT1SUh8pGMNNKHN7iPeYTKQUUdRB4/EZnb1
emuz2irOOnZhQEG8jvK6UOaWDZmyeo3xZMHbqwID39067rZYQHAT/EuQyatPwyxor4yD4cjtwEPI
nQudxR6ZnYhvRi7t/yjrPwL1/mKvDsM0cWetMGFJS2jkXwo2mMGZpRDjukGiMnY4CwntfUvpIiUV
ISiv6Iya6YSzgf87eP5H4uFfrh+9Mnpgx4pgkJk4mbV3XutGUEamqmWcnnvlHs5p8Wt/s11eJcpE
+dwyM2LTl+xVFovs4bHJJAFFl9NRSYRnGeqK+pdu3l9UI1yZe0nkCngS1rmIQWn2mwJ2YwpK/QUZ
/ftUYblATHVnRe+yjCSzYXG+fK+Be3EOMJ3K3RA7mF1TULOY8RzTNmNerpUqyQjHCBQ5odkXLz45
1aWqrlaaCk9Wvinz763tKKUFwruXb7muGWMi6IcaD69GMmfCcnCbKsNr7s7OESVoQpeDTyH/MR/y
YMHwxI8zNvi5KrhCFAzggLudGYc2g3AiFq1mLTxCFs41b7+q4gs6d6d+rOh2FX19EJh8M7zTw4bq
J3OJuI5iRieNT3zcxFDzHhw+Bpc6dIQe4EfxJqkezuXHRilCGvD9h/NXt4zu8WNQ5RS3YXiP0YZ9
LtQE5+uTeAG8FJNTqTQb7oBMZo9ejEsvm4IGt6rPxkixTRzmhQyP2uiC7CNnQ0fBF1+hLytt18d/
Ro9URwV6bMz1hDkvp538ez1Cqcp0dePGB6ZT9cv8PextJy5KPULqTKL4xNxqHUk8VVSAT1Mco6rj
FbC35VdlxdrCjafV+22FkhBcCAn+k23IvprKNHm3TGTB+Qr7gUNVCzHERr7CT6oI/28JXArcAAwT
orEHh6y9Pd/7HCjpbPYeKpZ0HMbx9DfsGEBtuH5XwuFWEsAqr5UhSvM0PlAu4TmQqxU2VX7p3TGg
9kQO3w6cIHVrLSFpT/FK+4PfPVHVnBtC43rcqAJNTksVA7VrW0wKIcGBNLq+FhOgMq8PbrLt8pTd
QDm4oZbA4UCONQZ0qsV61qXpabdKVoP/5PfZM9cerxle1eiDGpkamQOgzcnkHBo4mHKEmqVyP/O5
fUEhxJdfL3nven8O584jDcwFJRzoaVwkuia9cu2l5MqjU8nDSRH3Ne8fpC0+uONQDinxDP1oOpEe
hoDEazr69H27s1O6MhKUY1yUe/JFrGofI3E8Bn19g2bRdf0UbFgbNAh7G2ee6vs9Gba0aRWrFbSG
je+oY2MTWmr1m2E3Nep2Yh7+enM41Tr3lO8eupDMecFDPfuFDTPUKriwef+/5XoajXeG0K4KuOb6
lyPBkD8B6SQCQgD5S6dWMODwgiig0/ljZSzV/O9GftEtK8DRnl+IMcX1JiExBqtAaIDkd/wAbRPo
5kpOdgu69a2XNTModpu5TZC4cuZHuDeEQkDB81yLOcmK36Qe/O15HfRZqspXvcXnOzpTsimi3nBS
n+YePChF0OuXQ4QqY4Sc8G0FZy0v7i+P1LgO18KQ3osaHIsp8LnGo91Xy2FWCY90pKWPBW/N3PyY
SR0YVla8/Nk3fNwnetVkSiQviM68m+CL/+173n0D63Fsl5gX130C7XYfnahgwEuABkb6U/kRLnkD
JZAmPXli4P/DXNtHQZe+K2wxzSMTeo4P3HOwfiCaWiIZGGsVEfR4Dl12jHlv8wlQ5QiGRO+56oKt
nvRYbUuY4fC5/b6WmnRuhI6aU+i69yfoO1cuyXdNDApXNO5OZKLj8rItwPP6rEF6g+GUAVRphi5X
TEaFZeAs82GR132KoL0Nh+11eu7WmGQFpRpuLWSuFC0oeXCYjdADWaaWAMaK4Bz+kKqbwiaV05/d
R5uaxfLWgOqCl0Qd4Uz86r0BvcuTSoDaOFiVXVy6eopqBZMGoBcvJ/UHraQ4B+eZPwdYIYyJCwfc
wGhxwEAgRMsFiLVM9+sMp3/Iaebp9lYG4yzY6HwlA49kIhvnwNgOOPSAdxo0dd90hgJd1WcnkxWD
lxVfvQGo5HVb4IYXgWJVj3NAFWCy067Nr56MeHUP9oAneziIh0mNdX6cGuDInHtu0j/TYSyMn7RB
86vLgGsxYmLqTmWec8BClVuvi375SzSDJjFT0nxG49FLDsEstNoJ7vXruuC1GOUuzOEIw2MfzTdN
5kmjDpXsa0XvgZnoJ3ieuvRudA4X2tCNW+X1jOlAb2uA+ZDQU+AOTDevbGmayYGWAfL1QfUofDyP
92/i4DDNp3H4e4f6MhNbMjnPJeICE80EZ1JjxopclOclkyhOOOJC18NHuRSQ96tLrR6bkjzAzLVW
yB+2nJFAaQvOaFhTTyirKZ4g+bz6XbWYQc5tepbKRx45FQ5oIaENek+lWaI4d/0Zb0BtNzZ3eH++
2jPG+JKEhp26SxGESU5vq86vrvRBb2swt5pO71hOT0ay3LHE1Px70Id/J8iGZrdjtnT5sdKwm1Eq
RX8AGOTZYaxfjSD9gCAm2PoDz1GM1sgVUDnGwYUYnCptytzZykgRlm3s0wDU6h/qS7tTtXu8w68d
fGwt919JkuWsC7PjsthVG9javA8n4mBU4CtGjoQBzijd7SY2V3iOqZx7QmLbZKzZYX6yzWBBa00a
e17D/5H3qFnRWL94Ubc5twMme0NAzcQac53cAfMDh3/iEnNVuNKTq3OTIlb+zNK2qToLYMqq4p2N
OsOvBJ5pwtOTiHUfJL1k9/esW10MjQnPiNlPCmqIADhZiqr4bIvGPrF9atrUh8DrJoWJFHeLrbvl
JuEwJIZtFpOTpoaw1x6FuV/BFzglm+iQbR/1ezvSwemj9p7Yx1TPgyLWRkiUzVD2BvC7PIJel59M
ka/goJ25sm6Wakz/raf7ajJe1dHrse3ulwqw6gHzJLGI58EZETMnki9VGHxNFeRHxUShX9o3a3Tc
ckZJwx1BN/EfWFwksALp7Oc2HvX/D3LkDi3BAE6WY8FrRv7re0p9+ZNukEo+jNYRR6p2kwQpGxrg
b9sG7aKOHclWC4lx/ddrF8p4eF3PioGKh7qvVn1iSQKsRZERJNdb7JDElI2dpRGGtoqeqE1lREoL
JIx8x+dwVbjhHS9lLgKpRtFkDTzzbJMRPlIKINPqpwHPBVTDpyeMMFngi7hjtkxvASmx+gVA17/B
Nyg+vdSF8GAEZ6jLiNuV9xkGpVRn3rtIPr7J83xUmyIByUg5m0Rz7gBKxefzCHhPKywLwwx9Hwxr
hgNZlALgC2Aps0GfIKl2HRCUvuQjXEYWXjZWDfed2Z6qVtLJi8TnBQ9v9F2e86SN77/Cq+u71rkQ
BrBNSr0vn3Zkn5bSOhkMosiO0k5Mn+pw7KskU/olkMjQXL+Ykk9QGe1r7C+eVFXZboXg2XRwFMpV
VT0+l3YKm9f60swiOiUquLvPHtRtesEjR7f6ejnRogyxby9GOspjpYrjRlPsTyeMPQQQ2jNkQoid
1xJraqfB7EwSrfrntzPa8iIRoT5GO3R6jaVtWiqjXckeE5pbcIOFp4lCataLdRBXWu81ICaGHpNm
1EuAboQ/7V/psq9Ez3z/EQKILqmlZDMbC0QbUFgkamRa/iUembfkvcLezavpoKmcdySWYtXwc6Bm
rc0XgZR6esmbbcZDnQqVCzMAF2DvDd5zlOlSXR32GvyiCLanC6pKlNfUmilFd1eo7CYhBDMs0TaX
nA/TwEFkmO12eUyz3nnxwksF9KVKgO2GcKXWy8N7vsLTZb8eLSBl9vyqbyLsW4BcXvYgRKNvmFIE
fmjxyjp10b+k88arbxRKHfhRyWakJE7XkW1NC5/MfGESIezd4kxLDBv984wAsFJLDw7jsvlyaNVx
14ZQJzBzjWuAywtcTTlpAF2Ssk5enbfi/8f0gBk+A6f8NQTt8JrvJFlmyRh3/HzWO+EnZHR7vCVX
u0i9hS/x52UjEh4l9PaubtUbE+s0+KY3p5utZN1r6SBPw4gMvOgp8nPAz4gUrMRs+gf7eXy34hby
gTCfVtbA44DA3CzFxg/jpYGUH+96gZBih/anyapjJ91bKXJgYahmOm5xRbcuX6QpFMFbWc+gvGjn
BxlBR3nrd1nHgm+0LKnwDxsKzKewDROrRqI8vWXAlSJcN6/Wj13JJ6bhxpje+6wUc0AD4Lac9ALx
cKAkwBBm/8S/rG30+hp5oyzf/GxdLqshBdrioHAcvQXvZf1GJYb0QaXNWrWICpQOMVrEwalTmhvL
JwQvi4OzkLAjU/ce7wmjzjGUnJNcThgTwJwlX6iJ0oYnkMK6TQRfJMeB1myCS+FXYoBswadoEqNw
ire/pCA2njPenQCv0Zx9RCvW/k5Qfawa4gQymHRJrL0qtplfqWArvAWc/41gSfMY7aXh4YWio+Re
ZIxVEb2fWvCG/uFrfv0byFopnMTGBf1KJckFy72Vgr4ispwYu5GqABLkbxpjwMWGl2ShVSxdfxHs
bIh7fE2of80SAdkvLh8iKUKJeqjSar7couamu/c9affw0aXF+vIiDSRhN7Qp1QTYgoLQf16x2LFo
iWP6nzJokH9rggr4N2OA9o3oqNqJG3f6QRmM0Df//I6sHo+ARg+1wlkj/UaNIIlp8ud1JDQ1p5pf
Dq45n+gT6FK5awsfa0dVM2N2WTC9ApUHs4aNwmFCTjagt558rSUIZcX44xt714EeT2dWeN+5l/x1
o6k9VC8Y42EqePTog9clfyP4x0ZjSVGGGHD6aNZEycxg96noiwbiOHMuUtj8et1ollUubyxa9+ys
meALZCjxTmwvADLAakwhzPy07HKMCv/uNY3kVP1V4pGWdKmTtmmkrnsJKUCFi2Z5VhGa3Tsba33S
KlVkwTyYLIfrbR3iqgnAsmk9QMp4/EXx+dsggY/kMRHveaYhbbsCZ/GMByJIAaP1GhYakHtaINGY
tADEgrOFMYZIeP6Y/YQZw/DdVRss/41Ut0VL6GXLXIIZvo7YR9j11PPFFI4m0NLYwDcMFFxmEZo/
azvLpF+QMN7SQGKXJSlHnL5rdpEFQ4O22VWp6g60BVoBnQ0Eig/UcQJP97JrDAhmeeEShpQMlXCT
VTSSRSvoG+W2LK/895bO//9iGh7lwc7yn1Vt9PyVx7ye2eHqdL1v9JRurqll7cGGVXyUhdwVPKCg
kAYsfuJ0lOuC0dwNssaZeV1tDKIZGHy7HhNhX43HWzXRzZl4WXf0/F0jOdMAGVyZZF2b2SKt41bq
5nI8G/xWKQfFpHjgqR5ti6zKDYBLt2R3wemuYXUgPUJqSh6CPRCicOSbr7Ak3sWRw317JbEWHvOT
y70vRjMk90+E++b5QNFwbvvdodT98fLt6aigHDYCy0VV/W+Cl+RVP8Dx4MYfExCGEX7RE9hed4bh
AEvhcKZKzjk1exafyyFPAp+aIRkXdFQGpHdTrbner7hHJiK+9UELwErbPndfWMhw2C2MREipdQXy
J++CxEaNdcsYG1jd8Dd8MU22rTCvO9VbM3IId9X85yiyqlkY7YD9IzKSOGzYM5416klFLHxe/FuN
2n6xD0tT8y5shyXNqke4O8b0LDxb/iNA3fhumTzXPAjeq12g42Ef4NkmE46XCLMU3MZARe3xHG6L
lSEQkDy6Nl45sm6IWbqy0OU/wTNxKDb06XA5ADTs1pzKoJ2mhzfTTeGgpOyfwJc8bv8UxzI9L48K
pH+fKi7ir5geuWCfKl+Gkg/r0QLZJs9NEBf+odKexfufJMuqGGI0FYVjoTDxI3I1XRowVfygk8D0
rA5H+IGWvD5bhtUDy7idS5B9Rie2FZ4Ss1uB23kttztQBsSDKEVrbgae5br6Pb2rmYnjW3gXFLsW
mKbr01ubjSKFMVL85K44jcQA8K5AQoZalRF1zVNod8p2OEtKKPDRMqBFb+rDb+BWF0Q86rdMYiIa
W12fXn4cDHU4aWRtjZ+03Wv+LOyTPyoKNaH5B4Rp+nX4E/9MuSQCXqhqN6CSfHhVr5z4hBcc/oNY
j8YsVh//RIizGaeNtYBtWRZkcPWpmmfTX5nDrR66B9AlYrXnutW+J/p+LPtQO/hkI0XSQu8F+3Wf
yyEd3hCS0x9rnp8m7O9p2Nf4EYdp8S+wr/g1bfe+/UFLK8zb62t1W8wZkhHKVN8WwJXI41ANprlT
ixCVsk8MNq+uaRJxpxrq3ygPUaTgO0K8qdMcmDO/KgwNnKsocqxuJBADWGInOCfWOJoq+EEo1Hix
93ZB8l93qV67r/xRj3Yr6nVLiJ+Pw2D54U8mUlAIAoH9dBYMcQm4drBmaHLNEVVNOigzLiHPcLsD
ej/D3YtftooJcDu9yBxeOR4a7vC7nXdxz54FKlgeaEWHHyyYKnJ5Hx1J9JGfsvyGlO4EmOcYlGeV
4yDtcR1nDJQA7i7oMNhJMVlU2NFnQQ6d67430D6rQYIdN5yhvdyQ5cmxz0FCU+BrE8sosTMfVbB8
dPwzZaqTa30c266ZCERu05i8HQ80E9EdJ1kpOVecdydi3109NBfJ9goPOZSR6sw9ebs0nW4iWkSi
nmsMCohbolgWZ/RiUGbSsU4qoxnuAR52yyrKmI5XPdstb4teZhoADSyQqgfw6fzEIp8zq2vlDits
u7EEA7e+ajdbD5dw/zzGKJUNa2DaAFhivzW8EQXyp1bhIF6qw5SDkmtbNMQh/u8Gi53w39mauB4L
Tsdsa/il2OJq/9BMHGSBHSbYz/DKfFGiQuHPxhNcqhpAS2qw5PRRWk29QUfg1WssiuJtdUghzIPo
/E/PiiMScmGENZyVp50qItr+Vsavf2kL8XqxVBmRynttypSEYAQl/Bgl4tZ/nkFOGyUBIG90hFD0
SwY/O4QJ5KZxG91w9O9Z/bKuxyn2nQce11wHimsk1r5TzNd2be0gHaPurhGDwxUv7WVTVJ5nCIiZ
5LUNavRmFGamxpv+xOVAw7N454Pw3I6kmJuSpu6N/nEXtoJ5TM8JesEdU3/Ry1ojswSgctwrkV7x
OuIq4dkqt6lEz5AZ+/tz3COGOLtyS3i96h7dBHDnalOapyeFM0ZlR1oLOOJyqGdSe9plGE4DIY5G
ozNentlSH/YCrZQXYfuuOcZ+Z4c9y+N3TxQMdxGOMgb3ui8+womxr2t8Luqg1d8bxpqnPSDk1BSz
V8Jjgh3cGaEWOuyAKuM/sUSKDqTNtjhS/Y+r+E0IEUSsgwfXS2T5VRZQ8J2JAhX1Fsb9GTztgQNH
FQVrxbhoK4innZJfb3ocsWEdgag7mWhps86y+5B3CSLwK/jtsa/aF/E65rNOFXvz7wSypPnQNKPf
DYZDBvChfGnp3Vxi8i41Vce3klP0AZScWnNpRfRQzEzNsN/ejE613eF8l9Ef2UY0vfmsCMbjocR8
Q/73iXKUWG9UzE8AGz+989wYW7NJZSOJDPsoqRvTClHDjODpUA5mgJBKM7LfyMS4iV5vLFfPI1/J
B+u4PQQZBbzI/TkMf6ZjDVGRCOse0J/3zH20eCYfyFTmxuPtG80pOuNO9Tr9G0e8wA/ndNDwhTET
Bvchhb66tun/mFKmiHom/wrGUUBWGLkYXy1d9JnV+hawivhl5LV3a7qTW35gw1omdwFfmvD5Iugn
eQtz/RGpVLS+iRRzYnUgm7mWjoptCSB/mUBMKXUYWaJK+Wq03OkcD0TP8ZKItA/JbzQBAAp7zXwF
csQZR/70bjM6XeBngm/kVQ1KLQoKV2GC/C/vklRTUd+fxb3TZZzXrkkbjXcANH0SdHJD5JZsAZaT
MnSJyYMMMYo+VReF8h12DK1fOd8ZEPN7JHdR06NqE4/1XkCD+6MGuB1iGNaL7FOInFiLTdPDft9R
Q0jViKA04PezRXAuqBpTzeQdnBRL5vTpgepSC+J4IU6P6/USFgU2XxweDk6148hwzwJMZwewa45i
AEfNBzqnj2yL52FX7TQD17RHsP4POY0drwTb1szmx4cTejl87cWzmqUp5MAhDOWCbM/lzPBXbRP/
1S22QtUGIk7hXSEFSV0nI9oqC+ATmWMUyrzcegNI5fBQXWgPzQDEpgnsSDEisMH6StefYKW2hlmp
kRjtSchFLD29R7ir9ksEFZ/GCGLY04NivHnXHzVZFQBTZZct5XrAEMCSTLG1tEDP/hjLw2RGvHIU
CThvgwZbXradCsCLxzLQChMgVsaO9subi+R9+1iypqulnNmVma8fvFA7qF4+Py2trZFgaXiDxB90
U9MJpWQZ4hnmAYj1MjcN6Zts+fn8U6CgU3P0S6/LSUX7shXwX89zR67TiJl2FgW0Hxn5Rw3qj1Wd
kCPQKof/M0HEoU65n9N0bw/e/PwoQ0490QGWIZNpxO1ueRA4peTd16bdDOK1pwYLFmBNmskoiQDn
vNdWD95TDBdTHESjR4L1s/do1ke0V89M+umi1x2QoMbo5HZGnAeL9gedRlTGty3oAzM7rqPTFDD+
wSqiHUj+DrBUy0mLgu9B84xV/IpSy88CiXJbwTTVIJbi+yPKrN5OoR/CuzE232Szo+AmsPg/sEI6
Ar5LX0Zh9bq6PkHaxi9wd9Yq13v5NI/s1tgiZnRuXhw588hrS8eXsaFpaB0aq/bN6EGfC97P6rdu
s9lUASiwIfRcf2nWHQQYmOdkdQNGg8STkU4anNsgfDlNSEe9CdnvEUJJ+avZWlvQyok6a10xpFID
CxQewV3Qd+N6/Dfaqh8XIEogx28AJvb9BNoDWwgJypiPGSPXOFxcws/jnN4XVyIeaFBjTBk9vmJ8
XkwvGtIjk96AmRKNWst+az5qi5yeqeeTtbR17WWx2EowL8B4X+wq3J5e00QwnGP3BaBJVEqeBYmT
mdIMN6tUK5CbktR92frO4JilpQYfNyXiYppU5vzXvA6ELow3X65SIHig3jh2435/vIFZRHb0AiRR
chHbRjfmtKJqjNcvGRq5UYGi72kpr6rn+dqBH7JxcBG2V5EBBBiN1nycTx2UVWFr6pxiOf8+SA4k
bU9CIPCohVUKK7/7Wv2UCzky3Imd37ewTD1tTh46Z2HaETGNZOtD5mRJIc8+pKYm7Q7vZBD8/kuf
9rxAd+fY2JQNFsCezB8UuRuNjG7GtqjCpXC9hJuKh6siB4fOnlNicoFk1dxO9asP32VKlE0i0RBP
PmH4evqvdeyged09yBPkdStP981mqlq+5BM6zpE8Y5ZehqHId/VR/wEdUGTQMKSTeYD4FTGt3Ucx
HjiNsOLcvn40W3IYtfBW80ujf7Z4QYFrOwItey9I3SboDRpmXIh88HkvUeAS2uSocxB55rWuan1V
Hi8oDS4EYbFbMJu4JPQU5bM+WIaoGTAME3+kuOtT+S5iz5bHlTaoap202bX5HKO4iBMSfgbWuBHL
ViNS0qY63+YlF4/VhKIZYLCobYHyV5QPQA2Oh/2dkHnyYKgNAt26ql+g8Ocu7/wKdPvOZD9HFsJ3
W0crVcXcd263sDRGOOZO10OOy2OTSM11/Szy+hFgwF0NByA9IZHDUyLH6WFzBGobFM08uOxc2wPe
wDxw/NV9LBeW8ykCemBajXAwRi4077XXrRd2Pq+QvTc4J7ojZ+ItSBC1DBdgHnjYurTEchFC3u7Z
tlJQzepTvZnKAUHZFcJAxNQUS/W6jJiv7zJeFQrQuFHve7SNF0sU+dLEFt0+aX68SJRg3nkItMVY
vM+jqNj+/6sGd3boaFzhlM3E/23zuX2kv7dfDGl4P8ZolYzAhLxX4efIBfvI1N8os2EWTSIqXGcG
cx8Tlu6mQTzvQAiL46b26GExVJClFdtNTdTzyXMFxntQaPWVPMk0laZFbS7rmG3a+vhBtumSBVW3
aowyRxBfwYpRs9cxnc3bcf1yaV5bRG4PDwAczMlP6UXXZBXPRgIcGlZnh9knbuN5UZAvVQcDmxqB
TxtWPIdVrXqnPxtMko1YFO2kf7c6imsvSEuut8xa8qF3nB31KSfPb2hi0ERA2bn9601oecUsx7cH
/f8g5QUNORwAcWbF8oRVQZ3hLoAbhOY7pKCskYo58cygvZKsO9/V5JMBN1I+FIWWyjv0OFRehgkl
mfEVkR+rc3fupskZkMf12AnTYUY6oSJOk6vnoGlEm6GzPTAl0TC8qoYxSUQxvvCPX3KYDpYnqZe2
BRnz/DzPJL6i+ivnz6S2X3r6HNGDuONW1gsNmG+vjUZkxcC7h8pYWlZKzXVC8oN/Lv26M+RRtLrU
q7AEK/ZpX18x9IJ24gAPagtp7ZCTjsP6UTElS+8VHYf0IJFdQNh3SVXB9GkQFjVCwady1GNcf5e+
LaTiOOmyV3KXZEzA+TCjTAdiUXPfIiqnGTJSMkHMcHpSnrJ4Tpj2MvoL7szjcnu7F8EIrFbI9rdY
wAOxcwGLvBRSv8O/UEj87inQLZqr70U84ykTuNJhDprp4LsfxyD/mRBEO+WN84EY9afKBs3Z2uV3
mPadqQHWGl7VZCh5RiT27GczX0GJmbs/Z3uhlchFQ7Jqf36dMz+ZHk0gCZ3KNmNcjs9QUDCYFap7
l8dT3ZEs0FLdcj0ofJ0kMiaQMrQhlCn5NqlUsDWD9XP0mu63g4sEKLsebLpalrPwhGR6ipVTvbpL
z5BdXxExEDbSIDucWhkLzd+zKbxS+JgSE9gOlqUeO6cwF/3uZ80WmlYPeSrfcizbkLboIYhweTC4
k57rguKZwZS6rJp6u4GZPJ7LGWbo8HJRY1AsBUXrn0yZUvVQKHbC1/jOe3PsHP70vX0T1z0Rcq0s
NfT1lm1muGp7Zw+fC1nTBZFEvwNaJ8CyTXgDf6Haip4DvjDCr2N3Rnx0cSGXcq92LBGKd18+eN+s
NGuoM/fedDn3vzxcDYY//DnGqb9LMbgsylUwkoAKNnSgPvYOO6H69llkp9K1tk4gNYp2jYhjOD6E
GJTN+xA8/bcHnWivL04+Q8//YFVEsARJkrvp8SVCdA8JsXRrE7EmLiDCYYId7uWlX7LSMWD/GW4Z
rLKxQLXUwPwzjFJFAtbAoG+fpsVzGrlEbNAfizqqXOi2KLQviU5v6NSyuUtJmeA8/VS/ybWzDwGB
BLVaewac0kTJnVCiDwbDIdlMAHawrP1X3KczYSAdz7ZMS3e7KAlsZAsDQUSB1KFfnHZzlX1vJKds
FQXuA7bu4HlKZzltdFGAfP0m4oanJfRXtMNFq8KnaGlRvnokqthosMCPuFIGlDqs52WI/wVbW71p
dpXCMNZoTvWGn5FWRM8M1vsDEWK7V3oY1zKeV8nGU0X52GM/sPXwaxnlqku9KX3rQleECYPdZcX0
FWq81+aFFZrqX3sN0eK1uX6kkzhCqUJMWHnk5UQc+3ZoSi3MBrUPoFsWstW394dvRcF6JYzCa2vN
N6dnVRFE1dpf6OGlfs7LHUGnNSsZotKrc09Q3OfvinxK+aCKgJr9JVXqrC2PbcULlzbAVPo1gGOO
JcFI9SrnOL3TZTVzhgSN1rTaCoiybkkOdQxHQTyFt+ijqoRnJUyXwMckkSGO3E4f7j4+KS1P3F2E
eYx1fNdSkRDa13RF7xEwrhM/XWKF5v6W47m2+jMFGAfcT7hMRqvl8hfipHSLJbXrNc2xkM1elCK2
FTZieEwzzt5dxqxLpVja5Tv+g0O4Wfk7OHeO86vAZOEFyXGWw13Nn2Gtvr8GtFsd/AfxIXQmOdTb
2I0Z+qstwoesiEj9sATFDdOeFPadGAX9Xrcy4hSkW6pGgwEEIIbUpTtHnQgg0gM8qBJsCvmu0hss
dLkSBcLxkFDOtRSuY437OiOeLXRg7VHjMV+Qge32RUUTTA0RKPlytOoq6Vgeq343Al0gPxej0xX/
0gE3h9zNT3/T/w/8gnho/Kf4W3l8B6W7I1jz0WUMHdu7oGm/gXDSdDq+Ycd9RCODGdUHbDZcbNh9
LeVfNiUfSPXcnR1TLGBpJ+mIHB+caBKwQWvSNLvUiTj5+Zi1eRXYN6oixsjzkCIbTNuqXm6i8tzM
JJwxJgaDK30Ph9/kTgkIecdcet8dtULgerdU9Ug8u9Uc4P/HDzSbQUHVr41g3ERZrgDwV3HqjzYR
jM4ZQk80zuiEOLM8s4KEdXoJMXkbejUVoNerUyk3WogSGo10JfO9zomf9pL+UMi4gjdZyZrnfvN+
vpWOaIN8hUjXvcqiIqLacbSYuc2K9peC52vCQdwprKzcV6LR5DgybGheleU1sUgL1t5kFluLymdS
CwnJQi3/odlijSW13r/aoqyDSBX0SEbkL1RePdnSsD/pirUzqtzp1dlOQDokzij8FuLPvVoAcQ/a
rks1uNWUM84bXOXrLC+mtqBSlUFRB32oyQdcSvP6i2zr9jQL6F/zT/0ltL4ctaJrN36WZMhEe0d1
XlxxRocQHlDf1R2o+IfCG0i01+5WmBoecy2p42vN7WBlCxYkKQNA8SXxBiFX47WviJ37w8Pak97B
+f970BWr10DfrXNslsoXtjv4kiV4Af6o7d9MQ1k71qmmLjbpMm9z0enypixX/8fOjPdxKMzacTby
a45qIj5VwEbG9VhaeGOEjJRwe3ZVLvjNNwoDC0bofUn6mp6RVpY37cuwOZr49eQwAjw/p6wcutO4
j9fDeCXk2dWwgOBrHs39884WWkLhlnElSkoKhwqXK0W57h2t2spW0wZdri7c+Gfi2WGxkHtr+Bi3
aaefp/yOVAYeSgiTRckcUK00mLwWG8JsHRyOusHSAYPPeomtDB3uWYhQxwwv24lWiu3oiVXWSoHK
+LMRfkcdBm7zazJzFAA3wM27/AQGiKOUO2xpNZaPOoyVL1PB1IVm4dq3hjUFWMpGfRlf8kgUyy2Y
tIR7oZkVbnEL/1bvqdoLIh0MGiWJeZLZTtRSmsoUP/wo0WjweiJFlFolfd+5Ha9BZT8DEvVMEO8N
Mu0Gw19axEnlzO2gDXEO4UZVbi5RjMAK3rqUBkLNXMLlKbX65FYr5t1nVzhdfrgtvH2J0MfAMDw3
1WBEbFE+7lEyMylcG8YzrrZa/T1qAMPRvuoQ9JUPTRa+hkYVgpPk8Yja1jJ3adhhq5bPt15pZShA
ZjtM6QM3cKXUY2TQvXYQyuomwq5JJstkFV32ZeXZP9aSX0xImg2zee0TOpgjBs1tbLClFDIsdTP2
1jsURwz+lgM1uuQpJbfpvfCEwaoGMMrwYRu1NGLxxGwq8FIPhuKuTdewUmYypaPP2UwX/x/5ImEa
72SewP4LJumO7OeAuqT45gGnDY3GbSL0NnMfHhb2Tqg9WLHjoKhHi+/5roS3I+m0UnXnR3zV0dxn
i/Ke/6GEBVwjdAae68YM0V5jdipi2XwMiHmxj/xp8Qc00LuPbGRqLtmLgyV4jM5clJyS17geNXdi
eG230vPiHI3075YI+GAnbycnpTTGkAn34ctOJxndb24gD9eIBuMdQdl1TgtfLCCGdiJpeSxeqsf/
VbJlDn6Pnz6HD4IbAgpJZys8edAenJH89j6TDlagIurN3FHAVMmWOXB2KInqf162djFXyPu8bnUU
44qSMlVnQE07bbPobHdA9ezmSdwkXHoZIU9n8KVuR/zsR5DH4SJwdD0Ui7k05SkPS7skGQHW+ggR
yKi8AMJtXIxjhUU/ziEewkor5J9CU43boW1y3xatDziD89qCDultaXMgU/0v44g1NqlolZZj5y+z
DhZpV9eRj+g21wCFkXgEs2LDUvgjLUHxUlxmM6baWNgDT45DJnhz4zrQBpny2IYFwIZZsgIZmKZ3
+jEQQo9j0ZD7gKb4buezGvLEGDmk9ypVuqqIUbrNcLJv9xDhAK1DIG4dRlvCdfOVCXMs7gzZEPPL
1V+QVFWj3F1nNJouQfgMpkrCrBNUQG4SxB5QHn0Nf21PK/sf1IgKL1x8ZQPH+xG4rAQlNVXuygXQ
5HjenP9Dm1PcPk2ada9Yuo+Hub5epXhi0cnxvfAvrv9Qje70Sr+KOIQfAjq4kTDzCgC2if2LWSZt
HQIiJgKBH54Kco5aBrXpA+JgodXpW7OM0Sc8BPmdUfpr+HW+4UAJmXdmfeg/2+5a2k5T7gPRs2Dw
viD6y9R5IugPmNAArjOUeQciEPbvpVKnREeRpBoNI2GiCxDwf9QOEp2evj7JMdCV2aPOFsPwS2ug
gxt6EdZO7PmNmNlGWDi/jAANwK/mhw6OT+7m7DbJwebe256mzbDwIcmzKhRLduKXKO1Iu14Tjs8a
pSaRTgbBaBvqrBdqlyZVTnpXjcLk39AWTTglg8eUdWr/iRs0KR2xU3gv9KAzXBfedIYvqY0jTpn3
DeJuFPTqwxY7jf4CJHe7om8FLQ7Y0O4iqOyCJiCr3Y188SHLLPldd4lJq8jshMrHeCYoJzqup5cV
QuYnVJIU9JnRkvDwAWIAEE3NYwY1biivJJvWzGEONkDiz8cMfY4FUEpZmfl0MqQQs4S8C3dbmwGi
7xK1nrrXFfUnjdTTkCv+5IP2indwxRGKkXdoxIWxm7SXsSNQAEBYd8C/r45mabJKgd1DFVrJJ6bl
I9RdhArZ3AADWQD4+aNDX5NbtBqqqjAliZGiwshL5gc8gsRtk1JDxgnmSaVtrylMBe6FwvhG/fW7
fdtkdj8oj1WFo+u+5JtS5e0mMUMlXVlXzHI15dvS2JtYJUXsXF6ebudSI5JGQ9HzNbbYFmdi/kW8
3dHRglRGp9ZvnGRKBOXHscU765YuWyZ1ALVp9WI2S7qnr/4txOgDf0ynrDz491P2i2AbVMzvRgvK
RI3DQk2jqfEk2Ertvb8WMO8Xa7mARQMGWJ4ePXAVl3Rwt6fPWp5299Se0qLZThUjoiDL/0XQBSDc
WPgds8iwb11O4eO1ZGDTDy2ohkrMjSXndNHpzJd0OBHEryf+1qJgzr8mJ66xuJAKKHX65cb1gAi3
rsm72BsRDEDq/O0z+VIRSqVU7uNzNdjEp/AKBq7Ua8cy1Bl/zHFLY+9KVHTkeo9xOKtFa+cvMBPJ
KW2vuXEG0edpFiaj6QSGI/DQ8mpGyV3rQVaYhok9b6HZQzrbJDgfHwzed5lsHCLCEJGc8lvGOVCI
R3G1dbtuSts1y/uT/aGJbSc7YdBqyH1wNrI0LE/O+YKhQif03N4pTYymRVAW7MIPKfGtPBpR4NYp
ya7P+JrfQzGm/ONFQUoo9S6GDaS7B3NwRQps26JGfcq7xaUYtGYM28UTeKuL6su4s0da/N/ZKiuR
Ah4B8OqwjdFp7CTE3Be+nAhjwx4oJZFsisyh096mVOY6hGhQMwBNPnnf7+dGbgigzX+RkJEH91SQ
thjELU2jVgryJWQtiqbAR62vx2DgJwCd7ae4I9Nc++vU2BQDk5tRTz/pDva0I5PXh6ZOXoTeH5JZ
j6MOHxGom2Npaz39IV2h5iscMQkdInp30o8K7mqugjPus4HhLO2cX/+ep8G4GCf7zSGExbBN/+HB
39oV8XzwK5Dv0NAul94/SxrfJ1VK+bM5HYdLFz9nj2dOxoBUIqDOnGoyMQsg2i+wkzwD/YWfPFAW
DUDxrBXI900EkaZIK9Pg7sqDAAqoSpS/bXJw8YMiO4FliUXTg+XUbVh7lfox6rQf6IYizU1tvYaJ
MQWAeFfY1Qtk9mp3TOIrQYoh5iJ4J/AfkA4G2LrkWYXmB7h4JGAfeYxV01+Xb/xPS11us932Jdpr
iwvFFnrjjKPwT3fryg7Symf6M5IL2KK4a8tqCVE9fEqXtvRW/2pIiZlhlFhCtx3tJ7UDpS7WNx9F
tC0vhQ/0Y4++eMsFYr8R1m3K6RkXm7h4IOm6QY6osn2gTqR9UuqcbnBTjw8SQ5FBNKte08efcP7k
ytYpUwJinZnoaRq6TK1L2ETxLkNs5wYTOqPmY2/MUOFPkVwcoPNvNDdkZ90oapwWVMimOCx8dCZB
0URmvbSuDwFYbAxsPzQd4yTPURLUHrBowO2wShKApzkeZ9oZv8XtxV5rJJJM0KgQiuceUCMD9duJ
suZ78qUh1LxJpb9FG8+ukb24y5ViKiqQ7HTfYyiov+cefA9CVFNgzT94Ubs01Ru+RJgpnRs10uiR
QdQH43o5H3QPJ5zfj3ywNzRWeAniaCvxDZ7rcQwEt6dE5am54QnQtp7GwYwnO67qboSD7xQUlbF2
h6BRb1QaNnjBhlT5/hZvmIgqOp/FAuSAzoxxsRcEI9CeZd/YgvTmZjJsyUsjV8vKDttinkkNDm4G
lPzd12gzcfdU7mUOZsRzkxf7aQR//gM14jIJI0UisCpUHhmbwKPYR4LM437pJoewyZdJfggakMz2
T4zJxD7m+ysVsq20hbGSxgyD8bTxz6yi2HD+wmZYaBkXa/15n8foGoXXUmfVYwiScszdy3LEYTNC
3RCU/TgC1rlHkVxeDCpmGhaP+bKrg1UdvnP07i0Dc1oQsrXDCyeJTJCOJR5MT9FQIHsafbrqWVv5
p03Y3XkQrMEH3TVIUyZqIIi4KPLacWZcvDDLcb08GYCnrr2uU2GqMnA1eXBhUz7u0wtG6yvoPaqI
1CBYiHTFAuUsCIwODlW0AbComZn912JObpzxkyXh6MD0IUmrweN4009zbb2Ptiqkuuz6UtBPUZS4
dj4VguxI+marDwZJx//zXNBkcV9J7whDIt4c+kgEVhqrCHYHtIBQH6elDy98swtmsE9ZXLMMnQkt
UqbLE95LADXy+K61QlBQbKiaAWegg5QY3FZNy0pFNfwGQo97eXCiGt62HWKRIds3wMc4R3LZL655
96BKzvKu4JKMVVK4td3UZQLFUpbpLy8KKZIp8JZ6ZG4OTgPgG30nP2Gsi/y95S10U83tMu+9OfOI
pjeWnSypTcemkBiI6YxzGSzo+FjqUS2KTULm5PjmgJxF1QFJ23BtPJ0xrv1l5ecVL4nymVWeqTu5
UVTwigVfNMNyRpE1CDv9wJhCtXkWuekjZMel7OgBv84jFia3pmR9Y0njilb5VNk+XKzYIlaF1BL5
b38b4h2f0dH2iF1bK/Elv/axoJj1HSx+yfZCty6xiCCHJdiTH/BfXsPi0GwkUV44Pg74q5aXvYNZ
qK+1iiohgzNMcMXTUDwM+q+JjYhjrP/drdeajED3OFiujFAaNH8RX0AML7zqfqHlv2MTRSF67uBx
60nbDfbKpkJ/q5KFDoQNHPaHd3oZxVldTJveA4B+Undh2q8yLSpIUeL98v1cAHFKP0l6C4J5xQfv
EKCa6zkDf1nFwlsKB7ajvHSTEK5VyY271f/EAl7v7dcKly74uzYyVb1uwu3qPhPBI6Sm2iSH8r41
33PIwhXJ8YISt6EW3efzQPG4RchJcAwY3WcOd/6pnHgbX7HpyPo2HbyH6pGQ9+nF9/RTYguRuc7q
ZY/wuFy5S/YGYBqvnjXAR9LfdtC4qJwNUxXtWaHrWBZhvfWCjV0A122IPJK369m3e21u4qxgwmEj
iP0ylgebYEB3ib3kwNGUVEFR58sNcKzQU4iWG+UjVO8qf3pK5ViIlrqaImyk2XrB07VaB1h8c2yp
1E7r7jj6JOGQrJ4k0yX2V3NY37LokkT4sj56Nxd/w60fNO+VT23CL+OcrAdkqogjZra2cbFnkMBz
34Xuq14boPVYBvyzVNcl4irzSYU28D/dnXOFc0ug9dmVps5YKIo/4OnDahL+Z9fag4dR/0oI3p+s
t9NLKCbRH9qu50X3gcKwElQcXi3120/C6lrsNmVpluZ4Z3LABdHEMIxc3U5hzdcF6+r6Bd9SdhQl
hLQtzOGVnIcK3R5ELIwVidoTLx9M5+o7/qxgh20N6Ydrli+qxF0nD/gdYm8sq8wBSZC2339+PdjZ
zBalvGjZ4UwrOv0nzxMZIOMGuxNFDVizEJvghoUSAzTTjN9Xx3NXIxlWmRb/daWH5M406exjObzy
Tx8nFKOGhb/dqiYysb6QZdH0FsoS6HmM7QTacDwD9EgMnRWMpminCDjyCjFyhE1nSZoek91xcRPM
GuZGgkHwH73YPnHFsM4im1bzhLjxaLT3tiFp5Kx4zkaYqPWzBguf8DoANpMmxs6dk+SXoqmXrTCl
XYlnUizA6MCgRgALNvHCUiuALUVojf1YZAjwhikgeFSczrgnOOoV8eNz8nGtHcnPG3/H4oW766/G
O2q5u8IV4/J51uRZbhlaxOjbt6F0axu4o7q/E0RmbKZgkERuVIh/KqiQoaezf+EE1xq0lECyV2Ip
DS9PeP/Jzw17oTrJEQ25AzANcr2Ck0AcInCP7ztTpRBBd+WbEJHK395lCjd43BvsEBHVE0aIkbgp
zRxSF0+nlLQKUQoalHo1cMxUdVhDDIlYTQCn1B8xhVhmNS+F7qm45Adb7gissnDWTHm50LMj5G2e
fL/QSQkoN6xBy8x6koqkFXzakek/VHJRwTu26AqX5x2RIwguNMGno+ODthoIZ20LkSNq1I36S+Py
TxXq4z62JGTkoFoFRxvgvJMlU/sJtSNOrrwP9rY6f05YeZcwsM6SRVjwhP/WJXM/R10arAmJcsHs
iYZx1fJMgorIRWY5/hyxM0heW9PfzI2/fjs7gMTX1GLnoN4iB4W4rf4OKXX5xCEzL2dNfh+uOQL5
+Sbf+mqXA0v1WiulKEvtXnO8AONoF/Og6VgKIawQhHZtCc6CK6tB7HBLdoNLaoJCZqAyTqagUsiD
lOzxzcWPZPpfNl3AIafcQGZQ91xULM0h6fe2jb1/H8kS1hWuU0DT7WGfDVJQ2qdZ3xXsM8ip6ciu
5Li+I6oY6j9zoWDvOKkWouUXfarZbwBcorq+xxQ1LAgmpo97v+gKvI/tsaOMAVH4Dw2bz6oyHoK4
+WleDkdelNu0zuYt/+3z/9FAAJ3juUz8gAVwW7H2Dw9JEXsxjWkFpcCAR3IlfsuQ5zizelmLXNPA
D1LY+4AkWAMgX9LwvLobaexCJl/FbDN9ZsurNOdLrlgpBhHujqnstOxDGWgc/sIm3S4zdtNiM/YJ
giU94XgNeJg5r5/ubZjcVFvHPaLXUrrAMw1Wfy7eLwL1paVlh8D7aSzHjVVfJVBV6weuCIRhxwd0
DOt8f3TLox4wxGdUZPOj2ChOVgfUek8l0aZ7D/kqlEQXUcPaCqEjTsdjfFjqo2xHgaeDg00/bmhE
l4aajLVKDXExp0hgk6LahWZYFI0O9g8a8Lfs3+ei5IumVjcjL/1nUIx6bAW7RR9uQWygKrmM2sFC
edVJk66O6cE0QiT6BJghFI/+UakbfFtFt6ISx587ekn4Ws/aVMZY5ofAc7auApyWgeqlMDWTcCEI
6in7mgKEvMfPq/CLzqjt9aqjMFaZtmHaPfixcRavw9tQQfIsGPNF1TjtdPHZyXobHOoMUODaBFA5
lug/L1QkgVrhsfbSmpB08StONSV22lWs41tTLFVsnG93tAOh443Eza4dl1Tu0FXSEwy5zNJ85FRP
tKtOx/Ugf31evY/GUkZ4aS5kxDPN0SriRB2Q7TEJnGNYjz6i1yIsW19QaqY12/Gjuagr8X80yjol
2uO85e1AdfbWjDhcaqg1S8W80EPfgvxqy5QjLBcST+N1jY5rE9vym6qTt75nU9KaPCl8VHu8zIJe
Zd36zsge4e92QprWQ7+zbnpr4hdv36QPYJiRQvL+t5MVGkP4PnTd8GaFbHpQckoyBUUSUpdA54qC
mFxuKncW46K4EwiDNo1m4leKKsu+azev3OiwaWDSJV7LeqrZUTNUm0x7zMn9f7ifCHkVw4kNUeDJ
oJwd5H4wNvMRqN9TtgAW5I9bU/hM9eXIxeIndRfP197wbTM6X0F9EWSi641CTI8Ns9xVVnoa4TBf
6jQT6HE2/YG9FZalOHjw2bq2wtPKr34nh3QLOvWGrDZ55g1Wt2K/NjRzJP2XQUkgM6qDThdn+LFt
NERh59KSbqEU3iRjJZ7KNeybo/4U0Yd3UA9uj73d98co1hCR5Ve7EQCXpm0DrPL3Sy+GGznDBsEo
x+HvkJMQ5BsMPl7BC3CCR7nJahsQ+YJ4A/tOKYCNi8zC4eY+J4Ux56PRKdJDvMeWy6YmhPLZg3vE
TScYQ3/iUPXd+7yHm89axKoEcySAPgMPsKpdlR1VYJesiBelxomaPDK5afO2MYl3lKqiY9ISDJK2
Tc8z58SvmfbAAdbMIJKNwTgBIUsoS3PerYDq43P5ML7MlHXnsENPJWnkwluSKE1aVp1mOUUTbtpq
lnB8ZXz4A0xhsTjqVk//NsvpHx2xeW7h5Y8h3iQ1GtVpmN6FphmnyDIzKViasEUQQ/r9VuqUPJEQ
4hq4FXMkaFQGPwFwMWDj41yl1j3gPQ3VIegfjkTa5UJnPd+Eg68AwCX0yXnrDrXYtBJciRPmqg60
AcowL4x6D0iEq2pBe2xNAuG754OObcq8Nm3mGjUTXnPZs2dn+cTG/E899bHMr1TUtinDmzxzw7Y+
bQSVp1ids6bQTd2YgbW/oGcegzNKpkHL02D9mTP2CLu1LBLykHS3Hm0n/sa1ui2KUXecriqhYoQc
XRk2Dquy7S7iXCOieIJcAw/Z35ZTaEWR5oWMMXM/6DTGbWMO1j1fzZlYsduZuHHflkvlfU9+cM3R
ieCS6Y0ElYBUlalRyk/gLMJCZ6G9tbGiAtfq1IcYf1/EPIelJLGoXbxHCHtYZVml5wpz9Fy16JJJ
F6wVrBwea2E2uZjdh9zrbWnh9Bpqy/COUZ7Oj6LjXsVJoC+88HM+TUHsUTQWWkvLR6xQ8Q3p/AlD
SHk3B3DlSaOhCGH45YK0bYHkkyGcbITCwhMsChyiBeh2bBR0EH0eP4O1n706KnaJTOwfyL8gqqCm
NnOpUlN96Jhq9xe7dwM1QMcKTQUqvEoCXc9oJ6H189Kyps55U5Nsu36KGST89ZrizN8Cm1JBXfKG
OGp7fzy0/a6bRG/M1XmxrexVZH5kmgGmPzZZKgvkaWSbCj6SGxZLOPKrC697EdaD9MuikpB/vmII
DPoDqVW2biTeYQQgIjmn+ytUROkqAVr1BPGSkrfPc+7Zj86ck95qqAFb98KedhNUC7jCssLJvTvY
spZ9a+l90GQdLBRPAvB9Ow1aEwfsJo8jXoP5P7cCx0NCfunTOKN31bwpPMdSqSw62g19aMn0OTaU
eonUmLpaHw5+EcFNRTMy1E9mVxx/C0SvF70a8LAyIRZ0U/lRU+IolJULcnfTShZaMCeCG5UhwYtS
uACVacSrgcUcSH4Qy/ZOQSa3JjSLkrpMWoXfNFlOztuEK2THfPNeN+2OeyMy0vz1xp0HEGzCHvBF
39A8wmklCaZ/Lb7gKpwgpLSJP83oId7FreVsVh8Pm1UFtUNHgGm8hsSRENq66Hugtrlrv67MzKly
vW/PV3ZwpEi0SQMADgUWjgLOO5aiLd27OsJRElNUFStl0omuIhrRoBu+KSx3cuQgyUJhHs/fQLhD
UphFGZlhlVyZ/jwR93Q7FrNl/o8qJFs7RyWWR69ADygtbtC08fN47gyk3AuJ8xlJ3e5INg75B4yW
06Wr525qmN9HuG994OK3W4BAG9LvogWLOVRPdJ1OYU3dLYA6rSBE6D4YQzezoAuCKmkRaJTyyC0t
hb2rH7rCcBex7Dl62Y5cXGkJL6sCc0vDlb1fugpx0AFvIcnNTUJtnySXvNWGg05j5ebCArLl5Vnq
kRZuRyjjPVkYerme1mEM+5cbTIy+crrqKLb7SKNj93d1cg2kZD4ut8ZZuvKL2jysimKOVVeWq5oD
VdDJNgwUGxCnS7sRF3l1E22yYgfY6V8rdxQ0YzeNbcBn30EMHxGxsEjLXOBzT/TnKQO7ITs276fB
WU+F/J9vnPAruuckYZ/0lmbRPYLKyxMX8eLVWWiBN3Xvh+NY3UiQMmcAwNHSmixvDD2d1Vq2bRr3
5jyAyrzBP8/abmZU3JEFMDC+WQeWWVcEI0TBEwQRpi1qFxNlOKARPG+SXPGM0ku9TiQCdITAuioB
Ot7LKTIu3mj7wlr1t23+I9sXKHUEwyHOqEwffIZDHbxS6Lz0n4CwN/cF/aDQyiy8j9pLe9xJIU0M
PQD3iihs2Lt2Ka+yBYbj6a8IZfQUCN4cP3VolRbFLBdPVJ6YbdziBBMyA2w4Fi4v+EzFVrhh/Dz8
/0sno0WjuP7Lb94021MQHhYx0xxf08a0V2xjE9WPsgCOwjBp5SXNhRl5BIhsBx+U+1tS0gndJIr6
3crO+ThYj3VyM4GhhwU3IKBXfSndI2Hsmb/NVQGe2irHzkr8yP0UpbxBzq5sdhGAooQs5GzObqK7
yrIgKFAqA+aEzXf8bIE3rpTNT/lGWReExsX56O+hUvOHewBQSZGsgbbhfKpZPYhJ9SMBLN3HgtWm
U1y0MERZe5SMrocCcsRQ9qMUEG6EzbXTpCzJYxr9IjvB5tZI25JmSEmcHBq2u5eCMmvb8jAYRuiG
tpocTHl+A1vkLwNYZ0A4hxybhgEIKY4QB5W8VXLt+7kYq35eNqkmiyo5GzF5wouOBG6gxQxStTm3
mjb97eSCKsNoW+mQ8fzuovnmIsO54SOLTs+GCCFajsyIGNjZRrV9KqxLp9XMEBoONVvQs/EPeCjt
pb8k6xjzdRtcTRpd+3xQz+a3QKITyw2oACtZHWxYePMXwoheFGwIlavK13MYOAXSMy7j0UJj1NA9
lRliLt22drEauRYgQDo0w8y9IkgB+Skq9MosFanmFy8hErc3O+XrDcu2Y5Jt5m5gIm3tWF57quzf
EgCNdhaovD6zp7LI7fQYLabHVqz6eEwKhQ/m8BHr17csyLeOw2NgPZMLPDYZqsT/YJgUvxSR3c/Z
VhrJD1Pn8jOG7UwvVhvSCugb29yOLQjxvxi2OUUAqHjHngjqR429Pe0ieVfvPh08JqKXrDws36/i
7oh7avWNeVOP2+iKu/0wBVercX5ZoxL6JZnZwP6MhorTOy+ciglkEYO9BM+7i9btr6K7e7Tdf4QJ
BwRLa5O3v3VK6UXuZV2774iTYyh223Rhq2TdSQ8Ytnibi3turI1MRiS3klxelkuFwAbXvtu9eu9G
LlFd25Txm2CzXBTI/Vp5wwLmvW5utK+GimQsOlHLuotiZpvRy5d5oXmO7LU4H//k8nLRsB411Ll0
K7o0x54gEXOT8aojNwlp/bPBSU3O9N8vYRTo3h+TA3MlXO71SzEMrNyE44qxwuJCamVE9CIs28GI
38heu4IB4tW5OQ+6kKvD53C6UzjO39iY0VDfYzvCiOrvondjpFNdhWIcG5zxCWNE1rQxq6mixMXX
KvIaR1VNLxCUVOexIRJkyrypPrF5dZZEcgOE99//UViesMMw0iR30jr2Amqau4UzR3ABNkAkDYKL
Se2NtD3nGmlP51v93yKquwxkUAUGcKriqBx65nITSTjv1csa8kjelKOkQRqQ53DFw+AbcxiJVcnJ
aGZfWMFIkcb/+DQv3ripr6ZrfB4V82+8fSe+i6GCxsKloza7WgNpYL2NodqG99aSSCIF8ZyjCoAb
SW8jQgF4DetBvT2n2sZC01ZwiZ1B9AxcV+YVSEggrfhtg1AI13kJEyzrPyi3S8PhpSbHP+6xZeBm
kSs99gskMa+qnYKKbDDkLLYAQXz+PM/81MP+atIl0VjI5haTsgUSIPWocfA8KA7j6XvcHWjl1Wlq
fDzdnFXbLqXGHfzwoQmwzEi7sfPkusGt6C0N6ZIP0LrlbnKklviXYCLepiCGkKifaQ5H801Ompv1
m3vUoLm1FVCDI8/r/7Sdv1ok0A8jG8RlM1rWb1qVgqvPgaE/NAb6WaluncOxqS8h6h1YlHjCcyLQ
xfTXCF58MH5e3O/K1+zJhUptNEInfHclau0MwrPuym5TOH4Rg5WA87yrREm1bJBjMnQGyDJQeQg5
KCMW+jWLPcFOH/qKwiv+8dbtQvqNPKV0Xm7uF0P9B0f09qCh2lyXuAgHyER1/mMLdAiJC2aHeOII
fq4N7JocxU1WkGL3r7PPeDaPK/XYFx9wHGJ1tvaHamKFAFBRM8yv8A0cr6WHsW6ODKZHGkU7NiTS
VEnKyvNqZgjsDTisbVEO2XdtVQdMaiX0UttLnbQZN5KxJYoVMawUZGt71ljvp0Jj9130lhPMIkjG
IdWfZ6xXeEkE7S8ZoXg3oxjn9UHnhJl9ghToNrOMNe/MvnSf64owPGPP9UeeKC2VER1liFIygu4X
1gxEhAqeoTAWVtTNuKUkvOvOqwuo8m73Z2i/GrMMlR21KqfcWH7PZIYXyPwh9VtrgJFU73pC8ibV
cZ4ySHOy1S+DQFqAnDXd04iFo+9V8G4E8yomGEd/Llccsiv6J4YAdeO2b3XkS8zLIYpasycMJrXy
Ug5mvWn32lbQ8Uy+AkKVe4/d4weVPux3uuMPTYgMH17OcoflzlWj6mJa/wow56FaBO72bHuAJj6V
g/hmorFgV63Y6SlM9of6fdquwpodPDiwNvZ7kSExFT+16WfPzgbrTEv/JIRKbcdYGsqUucTW21Ex
AONy+Na3/yCvz5PxoQws9dvvIWIFeyyY+0IYEepjmlaIuQLjFgthB2qP+wUukZaB+OGPDm/hNHpr
TQJdHCK2TxXKn0N6gwuR5crjhFwHDE6aScN2b0u01pNEPlSd0haTFfRofGwp6P6ZwerCheMiI18O
3erE9x2m5rG12BinTwSFh4LFwxSFbnx2y++YtRZ0EkOJH2cAaRy/ki2BJ43DclkHrYWnEpfbQPKn
1C20ij538bddnG5juDApYxiJdfv0I3eVz9Kj3cME3i7by+rWU7SHJ7Rflutv/djAHEs4JlmmmW/G
b74qJA/+72wYiYhsSzYr1zF0v/OygTjZnaCwplzni0sgp8IkiOs03Ci0pEtszSGiW5lvN9FXDp1M
bzoqX8FeCe/AmQUFWyHdDOLbKaCy88CIcC42oFxSbMJvyX09YHbHP5xNqHn7DdtzMkxqD0eVBf21
OEQdx5Hn2HFBqZqr0wTM27J3tVZJNsO3Ceb5m5vHkr1mlaUUhstflJFc/EN+uwse7KN/6Sg7LdSX
uolRcxm9g/nX1Z4OBOf3PHZt7Ftg2TzUq21s/AB2+vjOOzj2hPB8S+ymp1BEHDyZTsZkSw09kx2c
P67OgmXDNpQLii4WygeOxuEdP+m/bKWh8D5NfikvSk88lGvwhy6lmvPS8M/3CoW96pAw4Lks8/sm
pRMh8gboCyQEXzDvA6ZocARqpZ8Uj4CmFbxYnWS+XOyVYUmWRoibx+N9zBrcS7MwSfDC+M2Bsvit
h9SE9iUA5cOsZAx38F9kS50ackDAcrSsI7RKxKk9z7HN64M7dkEBw/KG+PTorkk4G5irYQdpFTXX
z1U0QSglGmZpu3i+y+sN0g3b/W5mFbAPGdGMnJJUxkHLtX2I+d0LJhIsbte6IdPzy1F4lsBO02Gl
k9bqw6UrsysQEUjagvGcaQITxkcansTB0szjsnD7MrZdyxcfpMt1u+Ep2H7K6tsYqo4u3cStE4Ht
orPln9fSRD29IL1a7fi9OZ+5WdattN44LOZkgzZb/rcSv9m6fU2ggC3GoEdSudnlQonJb0vX6rng
jZBCiBDaEN9sGd59vm54koGqpPYyk9AK0GJDtflnrglNWvOJga3Dbp6A4dvsfSscwkn9jH/gHZfu
7gMFvz/lfZVCyjb03Xo0XvqHxXOjckIA8hSBwHMPEuIio5KPtKsSU7+qyR9a0EVEx9IycAtFZ2tD
bZTraY6jfeowYtPDCFsFGXXupRIz9dO/Q8Tl3nXVk5V/eRCqWlT0ipahwgt5hZpU1OK9ci4G55g8
an6VrJ9+d4nlJxEWyezkqSaKG8/DpCoSsxOPvTO5R4Pr4s8ZAu79XIYRsiXzt8rVuDVBbL/asc6d
gdYNavOdIytnZ0qtXJPBHGsTM6/sAc1atqZSUHmdOZSPj+GMXcio3ZG6bGSYPP/Z16LcwyGpbdot
ev2tNDCbIMWYZyJY1tNjJK8zgb20DXYHf2et7TnUjdQ6ex13I7n2I2C0CxAJC002V/2vbPGZf9cb
4YJslvOjH1I85wDTvnWHeVPP4g/4jsx5wknhxvREw/1WebCnAqJttLAl/JJdfHSpfddsD/bqaqN9
IlxkIZ9cnvMESi16kJ6EQIhvAYa6zJYx9SIDbN3KydRIYADKitiBITV7bYiCX9/rJuRnsCOz0XYt
JrLcyPYlefRc5w+NBQUy1BoVnocjbf6S2JT+YwLfkedKTjbCifKSRWx3c/dhrZGrPHqf0zTDTihX
UczszUy2mb9PPMV8636LUfCz72GnM9Hzy9NkLu79UxcwW6zWcG084l4ErZ5LelDLwWRWjthYv5vR
lVezG/Ro4PrSfvubIYjCnfkc88yPMGTDrapFn3jZdWCZmulCwa4JygbnOzLu/9E8HPWUC4GBx3Jj
TxqxpLWzEca2djfgJ6m8wC8Wu5wFpsxTyB34gtNpXfH0WjVvQ63nfERuMJg4GCV98zwy2kKHOdae
gCAtV+jZX5HHYCP9ZbekG//QmE6H+FgnVomD43u3v6EdwDbF1M+0EWk4l3w4+wpbLcpFXAGPfZKD
6P+awsLWcw87hHlK7cf+fhJHey5uTaUpou+uAMgZ1cYsBtYVXLH7lX/Tc/Fx18QITRKLa6NIm1WP
Ja6eNn8BwHARnoR0hHUofunZp3A4HHcq5UXhxpmgLtCRYBcEleZ5hWPd3k75v8ZN/B2xd8I37Ej1
V60/qwIJ3DjGxl7/C32bkQh83NMSKAZiaylZi2mgUrkA8yxyiIMkpF8CPHxdrH5W9xdVe5/K4iA4
BJMkk5vZS5r+pl2kO9bgqCgl1ocZYX5mG0srqodGYEcNhSxzt1decmKbY2lZ/32tUalQfxmxVw4A
do8pWig1ySFkNJiAAAF+jUn1JHChppFVqn5aAFOqq/H8dQCrfoMwuyHvro5arjO5DxBPymv5tlhq
d/4VDwmly30J91u5LB3XRdHV0bh+6JsCfgXdFtcHOZEsuq1mROG2w7p3ClujWmjXR5Re9JCRZHF8
R121xwW9l0Vmj0F2letej7XuryCg/FLTgajzGa+5mbXvp3PTJsrt3medCqpxac38Tmt3Dvl0RG9j
n0TOHpBk7iEFODFENUfZczQqJDb0B+fIi513GPIv33Pvw6aGn3Rk9FZ2aug/6ru6joxPnHEcmqaq
G/6kImleU8+YTFaPrZGsG91/BrU1Fj3Xb74lzJmDXWFRM3gnIe74D/MbJTVKARIcLAc7mY3yvk9q
BDcOWofttxaqB+LaxsidW882xdXfrdrfQb9iS26QQPQ2gb/cu9t8u6pRXJXJlAE6pWIWipeL3rKZ
aoFXUB+vrE8LaDcwaeWG9iR/5fkYdplViRc+vACClGbVhv22p6GtQNXao2fKW++W+Z1TAn3VpX+Q
iFgZJ1druxZXqXm8D6pEE9jbT5f5lLtvntJbtULomsBFR+3H+g96WP7xCGuIMeeWBQ08Ug8RL5P8
nFpSpBka5L+cd8O2wN0BZj5oA2gFRh63ttUmZoIgrF3s/Xjh1GdwmlcxaBkMmFmkKbnqP42DLY6A
U7BA+dD+j4LyuBHWHTb35XJEm+efz0qPYJbMXBnn6fDq/lzqRdjUwycKRUmUpT+H4l38pxeijevt
7qZgd1gzwjtvMJpd0SbNOvmCA+LFCtsu93U1FL7hBd0oOGR6W0Fu62a4K6OJuzmdWAnZ20XqV/RL
dN5q6K/JdNReHViPWWMXvBW0rrOkz9lWopwN+GJDwErZQIfhXyzwjxXf4Vt+VSfIgeQTSIXjrmSg
4TyqAR6bjelx4vWRQrjFYovizG4nlEsw7q7vh809ydWw8N3gffJiYg6VSt7EQHHP+6OC2dg1cmlg
d/A+YKjwnxzoJ1JBBhq4q1gAhV2EiQGstxR2k0+vCPUwZUIZYodU8C5kivFg4dp+Ji3oyQVEGatA
T11dTPI7eKqogwdGajwKNXqxmmdlInrU5Ix/5p2+fCnkRT8urnlJDuv3D0DDQByRHnPx+0TGARc/
OBJy649OMabIKCcTT/c/M4RHQibe5HiSXA9pMl+rAjHLpFcMDmT+hyyVqrcZZUM/yxxtJv+7vwdI
6tamEcuoHoQplN3lVEwsEVI/Fs4uJgvE1SfXkSIQOPPLQ8NpHQTu2zJD3JidsQAs5jypn2zgPAE2
5mAF1HXHOZcRI3WHtjLtXjTiTmDSuPAiZm/v+XogRyw7YUPkQfN9V14rEsqtyJC32RzmfEhxoKgl
OrYnVWZCaf9yq87zvmMIhB9AtvtdczDtdK1VPjzn/4+/tBm9hzkmpf+6bVkzWhbG0lT3/stXG0WB
QfE3wpS/e999D4512SYZMngP5PFRHpGJ/zHP1ZIDHMQeh4GYPo8mFE6B4lmh1IJEUMlBmxqfReil
jslcIf8byrzyNj6JkNBvLIP2xSQHnBL2ynRcGxWGNrqX8vb5qvXW6Z06RZbZljgSukn/C1eCIwAc
AcxD53us3nqFKrnxUlV2gjD7UwYWp+muzzj8dWaOPOQUfau+h0swIEWA9BEay9zhPuh32P7WwJVJ
q8wxxFZnzG/KcKNF9aVtYpdpfRln1+1zqlC0FaDzk+t/c6u8fPFsh+Pt5+jycRfp5/10sAi7oyVT
Yh3bt1tjdeWOFt2ae3VeGZDCwsajB68kd3PYlsJqHyd/ch08D/JJuBVbyXf7bTTeSyh5dNfowOuW
ID+tqji+cZa3buYq9KEag5OxWC14t6cVyMDR4sYrNdO5eNat92bItMX5o5h0vQwAtl/AhF7o0xrm
UQlKvmFRYDKlQh1VdI0QIzjCmoFCRKUEhjm5n+QjXhsoucypF85cYTXsRmFWIhjrG+sLeoGfRqRu
4T105Kj5bhCK9slGP1VkKPKGRF36BcuVTHAOxtEsSM9RpnxKjNmpeK8340faItZdCuZry5fxYI2f
4w11+NR6GcBMWdMOl37MIg79jon5qocSE10d+0sT40nxugQ/sabiF59DLrtlpbqo2uQu0PuSAXU5
xaUx3fFdONCj/i4jrSVcwZixXtOJxz/utI6IVztZkH07CsEbt1hrtkbKRqJGNU9rs1mAqaLdwmuo
6tEyQDyPUp/4RgVwy4u4c9btnDsMlIDDyoS3AMd1NBEkxZTHnQKgomNAl1AhQM1qbxzxj1JylMW4
WqlIpszpD3lPhpAp8+gFl8LjcAa5inmbxPTzkK25la9pXS78GDzdDUxXU09t2Yjij656FFG3IXS8
UJTaeZzcYQ2zMHNynCA9KukE5gY+b8csn0inPUByo+8qdqjTUcCOUBP1sdafjrMX8envCkFKMkAy
TXKvRJ2pILSEYKPN1PILSsNS0tvuBS6fBo1O9GXmjjAmM+liXz5c0yjnGaQaFUuzveJxi//UESFy
V9+dhR4rMcjzlxpWpGYj07Uc8oj21Z0LmU/Se6TmJjqpiFznor5qUzdgEbYYno/gPGs5Nd3sItMX
CwMgN0O9Ap1LZWiR/BV02sKQUKOYIN7A4bM2Jsw06Am9OWmS6SD7fsHC+g/hB6tGdZEirV+fZz7y
9bqL6pK1bydz0+VUvYyly4J82QRxsCQxtXrji62pSfpgyVgYmaAqCMTnYeO7XctqMe/1I3q9kPEg
/sTpq334mxn/uK598zJM2z5s/asHSqQf5OZX9JHed2sNtvny5eU26BnWW3PjSuuDEVF+QfzdL2WJ
sniEwGXja/OnyKTRrI4StmPMQ4Kq/w+IKUPiUY8Red2bxPE6lZc4mBmUQHElhlqMVYsgOr+5Gza7
X8Ss+X0/fgO21fFNJaMlCnVRnUOvx3nA2ap+dOlF0++n71Wo4czyiIghHyXLi2euL5vRs80x9Kca
B65qnw4n1j9nw6m1hWlVPfaBBIVg0r0S1rbWDLeRyoy52YvnJNvf67bVkPPCzq3IjnvCJwDwWlNm
5UO0bxpbJx2OBINg4Ta8h5GsBcB0CwjCxvMLTHqGILCQ3U8rW29tx9Gf9MSzz76AXKjEGUJgR/dx
EEBDujsc+dDsqQV0GsMC0wuDoy+v5JJZFcyne/IObDFjHI32cRYQIT3KZ0rx3dpXCIRPbRFu9f7W
KILP20JV34yAEjtlzNRIR19fkVc09Fl3ftQCjiDzEDAYONbv16afvvYfrIZeeqSE7d3HHSdKnf/S
a15Nxhqe38uLRiqMrfnsB/AY8G6LmcoFLjwDv84O5hn5GPbK7n2Wu/TFjuOtjg/3rZpRpPxhlh5Q
/NHxZBntf03J+gV4D9VtQbWdMs/hiXNRvlPjCOIsXlQhSiRM/lMYEExx2yePHdLRkeFAyCnrs1MP
r1LbMivKpXTjJghwHbhQrneS8kIz7v8aJrN3QjAAXGAG/KB15SFN+LEHAh0AQg53rOafCwmxsKZz
OymE9J3mNL7qcHFHcNchshAuAle+JWT7RjtXGQmkQaSXPVfbpJqi3X/aPFwEMCyDbfsQvSbuzbOk
J5L5eCb+Ox9D85Tcl5oGS6l4Z5Ls2GZ+BNTEnj5rpncvHuCEjqUXZX3TQD7w5CXEYP7d0NPDlks9
StqJ91oJIlzrkpPUojgSBHY0iuLBd+B7dPEcXfHQKgVZxrxYnTXrXe7GWNuEjaMZ0VrdySw2ujh1
qIjEW3KiYKU4wlVCOljRkXaNqByPyX4yT7cVt1E7UWEUCvYMs4alUyq6ROEvI2C9I9dbjbF6cDWW
D/2UhvUWgfuug5gs0fghyFjvTw4ohXCngR2kg9CvZtfAz7T131zickIxLv2dIZU/whN3kdiXBcC2
B/qvuJlZNdJh3yDmaaEHvouI86UT8gnGxTGPnJAecZYuuWhv3Mh2iF3Emf9a+mrMU1PcyBXgnq75
5iw24A2ff88Hch6LcLihf8/sv0FPQCe/aluZpCXbJ64YMNLghvTkVRIwdG9b4hNx7PlFd23qaTFH
5GB78B5zFuHi6+M4cW7//lKuzqxlvZvgesEYiQex5whKA4s6st65Qe0hU27CEUPfLJgG1yweXUDt
4e9EixYyucU0fmcb3+FOzbAN9Y5caLcJJz2ZS+wdkLG3zY04N4t/fwpyzYq/QTmHN9YQQ8He7JYd
Af8aWNgcfDgGDnb3pluhT87weOuh5QSCxVR01d+CVDJpZwFPjEnJBKwsfvCmVRTssYvEUFneXQc5
/rr5UwXd0UGrsilna0bmrjvFxCu2k22vP1FtkPmLOW1DDJiJkwaEhIP4L27KFj+zQz+cg7Pvr6c/
pNw+tZe/sHYZVLDknX60Q2otXXl0JV1PmjzbSgcfdYmOtWVLrAarkpTVQka9dQCLWGPqzOc9YlZ1
ANQ/ufgCFV6yfqeFAIjB3MlgGUkCJtgmOoc9SAKX1y3EmU0tcb3eAdfn3GmDTRp6Dc2na2GdC0yK
RgZHqfqDTuG86yp5E5R+dHxmyGxG4I3WMEXsgU2e4uy0KpUEEU1Ccm3E0RfxeRqvNhI5WKwVshoY
OHRpgQMsg+PYvk59uuTf+OFtbLzyKghYgM2uGxZMDNeojdyXxaXKx83zopeXo4zKajIm7w+WRlUu
paltPM5djYY+xAFYsHG/si/Z+fiMHazJs88Nulgaai97dpH1s9MfZohquu6+TF00zXrR0VNB/6hM
Tq8okpTIaKjXBr2HbyV/qgLA3zGCQQCzxBL6Cp/lXN97f3LedgK/oCC5R74B38NaumoJh0poWq7W
igZN/Y4pQQj6cdr+clNKyOmnQ8VvE4o4ODrJlRp8MuG6FP2IpTIiG65S+SdYk0jpvgtLy9POijj6
PAMuB5pRmAwaV6Ci/M6xs29kaxuMkuaFN16wRmilwej3aXtvpzgagqvNeGUMDTAjEzybAHzlf0v7
oFrVsL9QOSXIJbwJsmSs+BjOmQukJdLVR8HOky54UT+flhBbOesKRDYre/1fidsfjILUT+pru6rb
jhtIizSgYEfTUh93Vxy+TktyHIjNxFe4RS3enxn+H42kRqcDAI1XCbjDEchpiJwjybFlZNICnWN9
hCKJxoRWPzqcegT03Ua1B30aWHPQIdzVRxYROcssBN5X+yjX1fmFKdibsYyB7de/bZa08AOwxYSM
Z4oONexzLA12lur2z/00S0HMMrLGBc6bTNjBq74fCmJzsDt5clwQ9cLp+NCjvEeJ3ZF6QwjZqm7j
wsqb5ac1/z4wtMbCcX1Nc/KBsggNjSXTFTxGrbk7KcbhWAr/uNdUwBHXoRzUIdtReTnyLq9eCnjj
w54mjGvNXuZb8UAbdE160cK+qX58Zntb3rYtmbCzXMhy2VgnKQHbieCQsYtsxVIa7c+rWYrYtmgb
ddl7AEcieNIf6VfM6sO1DIaB+sJC06GbAVfSFh/DGasErNudeLl5c0+2IXpU4ZZKMlTIo+Gbis+E
OK87Hww0nuNyyzmyAeHJ0EdNwWxG2WTV/eA7PpwDkiSkY7uvZiyHtNlw6r8jw82eDW3H9cLY/78I
B7cpPejj8uzKAY40kpuTBwOXmJ/meulciHyOe/infNLvJRnuDZWu7L8wZmBr/xfUEebitGH7mztr
zMenyKHEvrQ7g/gYxeL1R1cRKCChxrW2aFafOsWCmJSRjfBVWnMVtMyn+69CvjSdJBxMqHqBGAFT
fmPOj1kBvl/OnKsO0g4ir6tvtTAbrULM+o2Dqf4v9ImlgjUsDT2cuQ/b7T/KtzpWaSFyrkUAKiZz
G2H1KAs2vTzmIdUu/j+WUS9JpMC1m+ncINP5DSibICLqobm1wL0fT0HiKjtUznfsGZ0MEmbycpwA
QAPdP/7dTBP555vrCj5nCqmRT3ucOcRxMDKqBBRWLsbmMwJDcjzpdfNGidNjfqrSiwhyhGe1uuTw
hkKhi4/dBf+U/sddTRvYOaWPwjjk+RoNIcyH4dyEDL27NRtAugRcOwz5eup4mvsXxj7i0bJu1bl4
fFW/3XrPVMqOOkiW1WIEK1GaWbwHpvrYyx6zvgxnbv0K15LSqg0FbYQdLucKxJCsgfMITNBNqgjE
X+GR3gqE45vQ3doCeTFlQldui/imX+PUMEz7TU+Ku4RSaYwGO5OlCKHL45EizqbE7GVnmHv97Oub
VkIyVTvBHHlBYQ7HV/MatN0BnVuY73H8os4R4dy3cIFxxjMgdA0bpylC5ae5inAldN79hmGoUbNL
7ZokfPOYnVCyGRnL+H8rYuArc6ngbIDJJNtGqCH/tItSybniDjJL7wjtJoclEXpdoAEmRIqEpsGg
nwuatOnWDQvmxDCyvVbz3s0s1RGlxCMHyzmOMCfnuUtodwDxqPRI6bTXViFPZ6wtWhS+/Y/npwaN
piSk5iTjxGYWMXBMWUHulvHpk8BuKq5m69FI+mTYCcbfMr4yKcWRBV/+RfZSBdBBu6rjQt6ppBFF
0QbqWIMDa8KdGmnsGWTckEbOvX93uzpp+eUGTFHVIqJ9uRrMMTx22XNi7NxaNahRbCmIrIIRRO4q
lEV4SXYLJm4Bc6K6/qaJyN5MnqQdTkreTOK0wDR4M6hMYksk8xIU1rddA+gR+CZe2l1Q9zr3wlbs
/+A9SySKSyjC7FuA4WRn135KG+zc4/Y6UDQ6jyouqsnla8SefLIaiY5hlnBv153zv3Wv7kzoBCmf
JE/covtnGk/64HJ3s0C1e3IHGF9pvEY94aY4b5tr4AMK18xMVNVbFketF94KybrKQhAOOvraAqFb
euPFpJnrRIFgwE0y25xUHaGljOqzvvqc8vjBKiUP/rblX6dw8d3yWw9nl2N3GG+S+5DoL73BDRDm
wDTQXrZGDQYgoCQmvKPklROT1lAivqOjVMcr8radI6Yi1ePhoeyqcuijg0Dpv6EMq9iynhWzQeVe
LV5nnTt6DYKOAHYUgl8CN+78kCvmAsUsakf/q7YX6ZPbCeEM8ul8OrrLMHolK5KpftE3WkZdIFO5
5yKbDfyC8zBqtT13o/3mzP8sW3sOGo11avET9tjhhsfoMj8uzYC05uOisXSjb6di4CPyuGaaUQ56
HsQkIS10onpYC0N7dc1Yk5cT1d90GaVt72JRfeT6afLaLHrqLKv3SqgCB5Gym5uOqabwxN9B8oKG
BJ1xDhzjCOHwIdMTBvgh/uh0y1Uzo0X0lh0/Obi8yfoMoLpURWmqAI5Dx7jVlmR4IeOS6waRWRG7
hF6hmkugQL6iC9LRjtiwNEpxsHDIqwPjGmJzlI7en27NyRmTEo+UDRAPnfqIo9vjIg8cNHSP3Lfb
cA8vmKXEVF9jb6Hv6Og0vc9+RxDMH2b4cZ+HxpKmX2MuX7tbpWwf+lfRLcSZA5PwrgCGiOBS+FI9
QCx6VNJ4kOthbXxc02Y2sx/2/sBpFpfI/HY80tWJJnngpymPLJj2x49L+prVl9aEgpjGasnZSIME
1qo/bg/w/j6sSO97TFJWUVUbourHAaReLecxIE5mjPtjva5Fq29O35gxbt7TQaaeFdxcwkvS1FwP
nxgDr5PX+E7RGZlXoMBYfv7h4HXPhHchFj1V58goDJlmu/IeFb8iKIIhXlWbnW/lwSKAcigJPl00
FMeYbcoE811GDqjq6uSeB/w6pjATyeB/DQOvJhmwThTq3eZOME44KajifIFI2mXZWVqxJBKDnP+y
C82TDv4dC/TPA6/SDc2k003jeQlHow7HTRIVscHT9YolmclHY0dEQRfYQXepBq+27/72OO9JMr2t
Hl3Ohmp7W+gA8aP+uk2W4wgF078c0mc2+anMNaiLocpH5nVieozM8cJrwmZvZJbHb0qX4sPM9N3D
L5djnDoA5dhS/4OAYXrPsoLyAhpCwJgdQMMbUdCfpDejUHxuFu75R45MVkQJ3ZbiAPPSrmetqiu0
RO0mdesOULXcpz16oAKIyYU+FeUKAveSlesCAdiRrQn1JSk33QXsY/Q2sQPMDb+kgtQxY+B8jyFc
C4jcrI/rEenOabx/FvgHmpQENqSByGLcjTTszD3bny0UmlI0KhhHjdkwj5mWb6A7jj0Sp0jQhHGB
QNEfXNqochDLk6TdWaBoIlTAgbMo5OnfUNjcblhhWTtgG0TtcR+7QL7gHtzg0VsiFnVG9yPjOM1c
ygeqhBxsJED02lW84zde0DRO2f9RDc+xslcTaQnjpsuRrEpcRVOns0cXnSyxfXOxFy5fUqpaSEaA
iQVQC5nt7cXtZR8nAQ6o2u+NTqRGRDvbHfMp9/xBBRbZ0AeCg4Stak4YV4671s/ZAU/FjnFJwefm
OLLLizs4k9Qz5nT5PY700opOxuvy1sVakwYYwlCgOK+aWqvnrixZDASRw3WawklKl4MM5P/VUF/8
yW1zeH1/Y9/a8auabu7yDd4bjPV25YL2MaGqGrdwT2atEin8TW2uMg/lrkfZ2q1RUyVP3OX0qeOa
Jp7fbvgADej4J+0jqN7MtA7jmAiSEnYc4Rm91v9e1vYd5RBaqPPCwIwZ8o4YgAWKXSRR4z4yS0P+
2AN4Dku/LGWE4ZDmLTQW6oEkjm2tHV+6anoAXz+FaTOTiN87rwwjpnh51euIpQ+Teer14ttJhmA1
n4n9AtWvVubEyHBWuKtGbJAcx5BCfPfYSdYCFmT5FcMMGEIC4Z7Y35P5rGePd1TH6+38YzicCW/i
JzMZOHwM2FO5RyDKznPS52AKJFGGlU+sG+vnyXXDsncpXAWk10tyWkeIOHNgWB7RePkZYyu/Bayt
gDiFfAJAP4qzzeflAWfGDfM8VB95gDJmP3YBzqsthwbYMI5iJvG3EYkQCPKgac0Gio0nGYGXG/lI
8sjOUGGkwTIX4QXpdsrhARANukyNlhO7iZkJUcWh2r/AasZ+LWZ7fB0OJNZbxy48OKD7WS/fOFSq
E9Xcs/vexoUlx3W+FyawtTwcAFaGrzev5gH/VshFNIvWuOSYDeTXCUzy0CpAwr8EuEtSwuM2FEDE
6T2h8/yHUUSYm8IWa8cNHgFDV53xWes6rL9Zbjqtm/64yVMsNgRge3XcGPeBnnaO2fz8m1X3HmKC
Smja3gxHzZOD047sls3W2E8HO73MVSAzRziEyHAyfRJ1Fss3MAqAKk3OnCHrBB4NfoyU214BWPXe
9lRdmSOanON6TIlka/dGWD+cf/Db51uyLtt+o+O4yAYdV9DEFr4tm5UW2+UaQg7j3ZbVaUmuO3gz
tJQe5sk0SNMhjUvgUlpbOk5r3mZacrCVdZVTWOvoMSfWRJ9AfZm5Wza6KKKZvIjwLpPAQW1ePKoT
pShsnErEFVHDDoFbrSX8ji5SaleVdKFP1jofinB7wOXM/JtCXdR32B91ofFv/pE+VyZiwQbCESu3
0QIyeo3ZnZrxbePtlmfQfS0rHwWhVkSlNA+zg2+LooTcB0VbZSgBj9SJTOiCa67JSFAxSF3kiOhZ
0WHuAoRwk7xvDI7fms555VjNP10MhaDqXZivfR1mLqtyHFfhKqbXnRFkZYcMAOvdSrn2mvvTZ8pz
ped99hXiCiP/52cWgWEeSGrzvX9i0CZeoWl2crceLUNUTMG8bjTKEXFbCp7GFAN6O7f6yhgwtV+c
S0++mhUOSonKPXs3WIcPmyR+QPdyBY0r/hwjQZH/Z3ykWJ4d5AYupKWwyTddxOQaeszjbUP8gNrR
gKb13FG/b+37zpFMo63wy7imakZFBUd35BYkHXaEnRHSCWtvOl6rJCDPbAy//qi3J7n9DSIH2opK
PNhKqzs7UrTpXh/nqWiKtYsb6CLnioL2A06LD62bytMfViQ7ramnn5NA2KDeb4MwBO70ReDlDoGf
ekpPNhYGWL1CCsn53EYkdN7oaHW5y/0COdQCgzN5M9qXhEgQpJH8xaff1nQ2iA6zL0PDXIODz8U+
BlvnMxBtQ4N8G5fKkq2BcD8e5JWLBzgtPm5+I38rpUlv6TOo/uSIKPUlWIRapYnQGwuKobxMEmQ+
kHi+bqeVWPY3/7QJqtxSHZbpdxF2YurYHvCfIVCuTQ6dP3nMtwqdZPB+ddq5IRsxE4pS/HtJD9xd
fXjDUx9WThY0JmkMhXDT68lKPj6GCgglaioOwKFjhxV2GftwaJlI/5tAt7PlxYWeN4aQ+UzqRFcz
D69q3D4lEL1ULBJ+NhSFrbjsH3g4hoFa6tKo0ywVAe1jvmASRLqYcHec1wKCLORlAd6i/heHGx7E
ScGd1/8UYA8iXMD6fgbzqQPNM+1UfuJ22sEFsVzc9fqDHyIut/l8gZPFlHQtA7J1xeDRCBEA0qQn
0Aghp2153dYaEBVjpoxJPOPxs2oJknDORaKFn7ztkOQyULqXFtwaGA7lkHvPWrw1loSY700kQ0M3
P+fPNAT9MxHlLNcSx9FC44q78dV53Pc9n5QWz80gDVQFGORTTbJkESjdlSckiNewgePjWG8YGklV
coNa0QlkQfm1SJDtmkuTt9FrzV96VSJkC1kjsdahTJa/apgtVuWdJIS88KkmNZ7HTYKootB39CEt
l5JmvnI+7PcnI45nh/kZ2esHIk/RTFFQrYy+wfUOgZ0903bJbZv7H5CF/JxEa2jMJLwyVy4QvlCC
QbpwiYYFROD9BCmC194sa5Aaxzdwgkc2v1FLBtFS14YiuIIdrH8hdo8qpRVXrOeX9PsJ5c1mPtcT
4VTnGrFcjqkZXLJa2NOyKVeAsty1f7l6GbPpdP84GwZ6hPcfcNrRcwXdz7Yfz1tzy0sULo4cUCZp
HqutfT5tjXQ3AdegR1vFp3yCGtN3gczj5qJrHfi2JQL4AE42mrMICKuQS/sNPA7Xxz6BA4M6KdFz
9dN5lLVE7UenohqjYkjtC1W+hC8Zq9SfwMk6EdVH8MeI3er9TgHNdpc4Yvi3TMOPVNGiKLIxCB6P
0LSXR6TyqyXMqqj+dqNg+zL5NIcrBWMmzZ6R4VedoEgp2xsAm9WOs0RY7aDCzAVHxxbgi8//JlRV
QJM5L48g/A2PKgHuer4JPeOuRSe2X7MgEjZns7u3p8h6qNb/CS6T+aapJolmCkFLIhdfI25dRsvX
a2v5+NvJcVsarLQZcV1qdOIzAOO4iDBXDBc6VTE/OTPXdqRNkIpBmHkWyjSKdzl6WXKjxMRKPAbS
dEtTbYGR/uE0b/oF+kj7feArt2DccZBuAlRT3FxZ2YdgP5vNudxraSAPZyMA4m79QHs8CDDLwOyZ
ZudA4xol1h2Wruw14LVtESQOgE7BQwAbciqvmnVZXY7WZeN+TA2EpWeGeHre+pVUZ3ngocgCoIQd
9mIqQp6waD39fWVCCPQ5WT9aiHQFJqEL2KuwXKX7mf5kX9bI2ASk+ywvPpTgC50y82tOIzapB2qs
k8nHQzkP8nT0KFGsavxhqje36oxNWKplqczbwnyPz6mKz1rQCxCp5TGJtfZ7yCgCbRcOf0iptoZh
w/mim3TJQQukSieWMupuxUaDBr4R6wHgzBxbiwSoG45NDFCgjcfH24hNKN21wOsVDW5rG+RJJ/ud
e7uM/H47hug1xlxdDZ9rZLtPg6fx5JYeadM2XuPNsi79qqG+TuRhfI4aze2gxoQr2baiQqrDBn6b
tE5I6deBJz3GBC/mqYfRnCI2jkggJrmkguv92KI7J4Tx7VCG1aiKSgoHHeLClOXThsa5Kg2d8BDH
OdQA+w8zcapLCAf7MbHIkgZT/O/XXh6oZ0EbonQM50LfpZKDdDCKFJyipuhrSmYuE0/0Nt7ueZrl
7+l+xmiGD8XJx/Ipw2d55OA0WzVx5xG26EcKRnuEQa7MgzsaqTo1Dt+vij0riG8PiJ6Rn7pIP9z/
GH6Kk/OvttHMVG1qLVlk1YVFmoOlm4Tau4lSvQTU0nFZMrrjyeT2EE+IimnAaLjy7cAOnUS2XaS1
PODM6cjtrKkPh7BcGdWiBkPzp5nSn0MNdVVIEgnpud67wKRaSK/ewf5JtJJ4XhIYNJMx81K3VQe0
JvO1pC5JLwlzWYtKKqtqk1v9q1MK3WaGkma1BZUzGFmdqO13wNurB1p/qgk4o2qdU9dALglGYKqX
Mk5BHcXuUfKmnEoFUKJdNqwKacz1th82Bw3lOKVKlG2JjLPrtBUl9uWY4XISGD+gmuMozYjtM0PV
azTkSS9QHEyoNQDsYQ/CMDBqsw0pUnXKinLZRDXySfA36j10ltv6gYCXTXBtDJovcZZo4DR2nmJ3
0AVUjQzSsfR2uqDm+Vg+X1kA67gegRyoVzZaljMxsnGXSrocm6L2PPvwflTySR+6MjU5xGMHqf2b
BMtbef2ojbv/bMYYp4CLadGfecdaQjwsYZYMCeDboR/dral7mRZpjrREe+eYZvKeDTqfg9Rax4JO
/KJgTPHqG6SBdVNNxcwI4TYKYTZhCM+vpma4Mc1JSqInEZspprEW20hjAW+HwVZIqCxcF29ZIUR2
7E6WPogNyvGI8do0z4tAXiXDLDs0ATZ1Qsm1KLON1b7LhvYFOOrmwp309Nb0YnSHZWNhm/SCdrPw
qlo7NLP5lU+5HSbMHhyk2gQAjp/FyUaWaFdOhmzhsoZGcXJjwxbKvoztxFuh55ixzRkyz0Z7Ps1T
EbRHZGnW4qTQaniOcquvEOtaofJyh9lINuvWEmKoC37rdr/3o3Rw5Jg6jVgJOH06SCRtBvfaIPBn
Pwsbjj0kcK+ElFif5PWlhR/e9XWvtwYnKEPHXUDFxjlXoaQ/hsXxMxwaWTp7x03UfVZDeRfOTV68
gxT2Kgny1IabX5GiA7KqC+tMPTdkxrna4Buiu5xqm6pOG0PG/wHyNSbHG2ouSa6GzRZe/3kwR8bD
lnaisVwYioqO6+eh3j0VV1q1sEwdKfXtSOY97vOhbGx8ayBQJnWKmtso8fFmZPbqnTNnrI+RUpUT
9eH2kChMyUmTufZHtDJR/zxRpHsQgOp89bLuB8ZF78LrsX/tviAUX1fqwwM+XdYyywdgNCoEVkRB
jAxQtFyFoF9jQ5V9ZRYoLz5x+QW88DFHf7rCX5AL89zhQ52KY7lxPTapgIgNGUc3q8z6Yf8GVgIJ
uCZoaANPfZRiqfXPHEVDFIhKh81OOwsnvfJF85fjjUyH9nBaSnnsMlPzM41eMSVnuzFc10rr0C5g
MeTg2vh8VQSOk4fqxDPFXP92Y71Zs+0lKTe49a0g5tTjSdxEdTiRNziFPHlGctAm6suF2GI0YrLY
P9FWG8xqsAkUrSQbh0b3BTRD2iRMQsz2LertSEPs+flDpBjwqrpx7cv4pDb1sTssspeIje6sMXoI
G+ofIwEBcvAGnpu8Xh2HM3SjfaFShc2OLUUnR9gRYqnBCL5xi/R3heh6foOpLJGAV2BPKcMB/n2S
bS8zQY8WXq98zVJRcncTp2EaDYLiDxXSC3JTztdhm1dE+EJtB1qhmoQpiKmHJeHIt8tINRRx6Gjx
nbQeu8ztuwI+GFOXCfGyvS3T2s9skAuG1cflD3Qu8Nlxmat6tJP6k5mvNmuqMGsrugokWsAPVjRm
Irq9r3LB2Dyr1q4GRmkrSHnKH0PulEn1u4ZWtcKRNdugc3JJgNtm+kXYRD2MG64ZiUi5r+oW1DXK
gjuTpNxZ5PEMjhgmoSd6FQeLU7coq4tMkGqUg+HwSwl0iXUj8xn/P2vzL2eyJv0L1XJfCn3ETsus
/yrwaIJwrKT8H06sbD5d2Z3hMlqwvAgcMWRMrZO9yME91HSm1sLNDNeIIhu0tXAFzeqwURCgJ/Te
oc5lEbi9kuJTaASCiqWBdfFULKvmGsmhAVkCw6kXPxcjRPC5bvlnj6dV+2bRFU8FijwMkcO2u/pS
T8C/dQSIT3ghV/ISE0N0rxMmWIPbMAnXZzv5Yn21AF/dcd8vLwMrvMozROKOjNBOjVTuw0i2Dvym
8zArGHSK/9Skkv7OEw+Z5KqdNtGOx4gxaX4UPXRjA8nvQq0f6qsd+oPfzYoBBSwxYbR4sCyB75vR
/WljBRpRSRIGo77vnqMwti//puMglr8NWYL5ExpsWzDj5shAdnVxQE8BEhl1HvexNkQPYUZUGtBY
raM/uxc99kVBgoCV35DkAsZLIa0sGgq5uSFwVr5tANsCHzAdww4v36TVs7u6nLkVtHk9aenXsH/3
TtWUzXDxd8U8nSBbc7XPUZYj3pQ30HK+9xmST2gcJHekbk4Y8SS/BIjiB9w2JL73h1PLy6MXrEJW
DgR2hyzxzQvnPheGKyQiCLnhq0LCHYcWqOFAMGLaWRzoU7k4EJ+RTn4g18WeaHccCidHXn53aa6I
KKo5nuiDP7sfRN9cKtHx1Cu2j9vYtlu2Ixg6mHH6BcYXxLW3FIYnZWF17mqPWABMVEZcZc3irkmB
e4aLZn3ad8BWR7nZ5zLKYXVOm0Ms6qtgwUQ3vLOPAG7aMGoU0/ZnaeMJzbWHqod9EkQHUjLu5XwY
v++G8bambVSgx+FMMOL57fsrAnJhgrPfp5msbeAmUTwIGwv7GNhxW9qi6om2dBxnH/GeMchM+iY3
i9sIlX7O6ezWGYD/hUi8LrzDyII9sWg7fhwF8icuVuX93osOk91jLpZsjj1D20AtQTuQT6r0jYM7
d8zbUHqWDWaXeArbt3Ikx3gMy0/DlbImGdJ0Jha+YQUo7Jkxt5KyAJOqCO+0+xQXiML1bfLST3Pj
kjQ4z41Pgd958hhuvhs5pq+kQkktVLDw5csultFXkCV954si/wnP+JubTVDPlW5eTRG5jevCPxBc
Q2/OwobRAxSMjfyMjLTkVWqap2S38+wcU1a6YTeHslkShJZmFHsXo//hWS+iW9cSuVMJpZFGdgnx
ZKXaXFxaxlU/hBjPLtBouxEiTvPQTkzsrnTZ18SmrUr3sibt6mrZJ1LCJ2inNdoESUoMLKFkdc0Z
CwRgmkCZ5qw/+4TKkduE5/2+SDxC7rSUbLVykQ7BIS42AG0x85xSD1xnV/UIv2QcnzOC7RHLGWtV
TqBk1i5B+kUVJUuPn1hfz/di2BRXOAyXGI1lYhHUOGs6r5ZsGs2ftrJs/eJgDm2EkwcKMW5FTY1g
cpRY17DHajUVX5YM694zuR4pwZzQFty4ePqjSDqba/zChttEUr9jNKd93yCalzd1aKeDYnUnj8oW
prUA3UFu9Sb6d9Sk7GX29FwnErDdMKOVNxjAStcRlkd70jkZdufd8thJJZE4uOx1KzTG3F+9joJL
2eqUSaBRQu4dpVGtUY4rvTolHnDF2IcTb7WrJSvNU3scg6hqXxf3tITIK+xz7aXxLdMhF3eshQ2T
hD2xXqRqzRO6B7eHGmsWdvr5nVQNS7J9AsVeXt3kIL37SOpbd6B/KTvkGONBk8VHBzUMUkW+Ufif
FypV51t4mEd8FTjLrO4BWd7cX4RNUrHF+nKpvjIrGCxTjkS67cA2+V0OwzhdCC+sso7mcBtq2kYf
4Q5uiFEELed0JSa41ESbB3RcianGYqcC+Ism3obqUQHClYUmIJlLcIR0HsXqXYwFyyLwxb4seDx9
AaLML8zDKUcbtXE+K99fx8cvkHumdT5uzdiFjS3b+mamkZdAoFueJiQQeivV1t0oe0yp6ovgaMJh
f+L9oOj+DrUos4yuzbVs6m91vFzXD4cvgC+2wJOwM64AaPsjNVCP62DCYOsEzhjTYyIPd4ntJAEl
XHg/8k7y82MJxxqe2c4q+FH9pMQwlxWpr0+7eYXb0gA6j3/A1uDkEq8QqBjQniUNUST1snUzrqnp
MEWJzLG4le8NxbtRrlvDAimFyz9j6pJ0wlu0er+pjGq8ZpbU94GG/OC3Mbl1+JXumGL7Si261dVR
9aHYzjf7iss04rnORAkdwFyVVDbqpKRSvIuOJDlQ1P3DsPcW1MJPSzZ1GJunaCuxAIfDkMT6J6xU
BPx/AAs6NIyefSP/mCUStwp5byW1OMXC65Y2vDvp4D6XWY0F7UQ+NRc0UZBTWc99Ba2+7z5oZwQ6
3Qq+dTVP+0RQfugxfH7nGYiEQcDU3ajrkN5W4Q6MCYZbFA2BT9yLkwC9LGqql8IFHTj1qagfLjy+
VB33/2m+wMEjiCIhNOs23xKNcpLmae6Madu6YBKTvdbImH9oCzw/RqModpjk3Ybi7dDXOBRcovJW
ii4/dPsRBssepIZ9sJduvnX4LwlHBgkPeuG9tW9zujcX1mGEIV0FCVv0w3BB5aJ57Fjnu1lSpct+
FuAlUhEvqiOcjcBFBxqYx5887muJkBsXAqP/fw6guOWVS2scMYHyVoqXiF09HTHSX19G6yO27ifJ
1MztEZBPwfwLk2xmypRLA5NMeUb6PoU+UQ77s1ITdxQRPat+aFRD3pREqDwXj7dHw8bbEamVIrzH
k5N8Ei4gGjWjwwTlmF9GBNbi14YYyfylBqD4xuyVcsda8Beg2q6qKd2D3blPnU2L5Pnmq8uEq2GF
na8NxK5k47csUc5xZpllIvvDYY958NarMorFPdDUBz/zksBz9OlSQH2av5haJf8bjqCOdu/mjEP4
Vl1tLHJvEdGeXVHUHoC86pXjiWKPCyIa0NpYdgRmJFFzwUSrsZBdjZTj8TYm+GFlVnoxWZpiU5la
7Tlo4cEEOLiPIJzY/6dsl7Jrnk1YxIR5wkoyR6Hhh3ZCxD5k2+CdL2MujR0YNSVMde1NK+P22cXY
Qz7kGmU759DRu797Cd0r6Wae+4d656qx7jOvRkzpX4eGOZ+bArb3yIlHp5maa7dVJh2J7sxBxnz8
xr1RKJOxpIaA7F2G3cR30BU7O95VDCWcFu3ztf8GWs4ZdHgB/Cc4kvg9sXlQtlUxEHCemwWPv8J+
olkF+U2QVAemtjO+qSWIsciHqFZHr5Gu+RXejvR1SAJeeXZb+aXcx199Ohq9OxU04tQK96EA8O4E
SeaRJ/k9kt/JELsP4JljyciALCVNJqJ0P6oUCV48bOC1f7pbUVqMqLL3pp1PFk77Q13E0DJUH6HP
WS8eiasHdN3WiYxuxmPB+gQ4fxBoY4JHMfTR23sG2z80Px608rf50Bqtg5G/2HMOzB99mCGOfQVT
1ftNDCPcfp2WTkM+8cdLRpKXmSH2H71HYw7+hFwFB/twKsPLBiN3g1ZI2EzNh4wn24HXwQZnyOYM
pGoql0G0QorEcXl1wLpIdLs+bC4tV58CgGpzm/f0gjgrEzkRQagARb3fU83P+frYMYQQx0zUviwn
LsiWRUrwZazzQk+hYM2mxRwNA8oFqfw3hAqlHBDewIHKjl7J1GV4MvxZwNTh71g45v0ZYvnoXRH/
QGBWUACOMptDhIVbkcGCJm5lTHrKQ9IIPmx2tcOaN9JJtfBaHUuD6jkzo2Y7q6YYIztdUBAUT9cR
rV4kuCmRfZi24fQ33SDcmB30zfKOi3gcIRtD4wU1j2c+7CW04sTuLMwX25TeW6KNL26zLRQlAm0k
A+9o+AT6Jds+zpWQJ9QeYwRR0OQ8LQcWZKVwcv8ZPx/c7L03fz6JhAWzaRNdf153XiT9q3y72xeM
qEcYZkwwurhwx4SFcur3VD1D+BT2JuG4cWri+ICR8JKaszQpX4ln/5oaRrSe4VMwvbVDvPr3Au6U
oHgHYN1eiyKb/TkgcWL9FKG1AGKE6EGCo9dTbnN5gKU4bRxe0lYHVHT+4IRo2RqGAnrVcNwIn3MD
oOu2gj+GfT+fvSaahIs+TLxwK8cPohuTo8fqgGvC7P21tAleSyrVY0AolqXZoVl9f8lctOw60KTg
baUC1gYyZokMrCyBub/3UJ0++l+P0SUXUsoK1t5ln2Vl1nWU8g8s7giLW/g2BVXLQws4qAgZxJd7
XJMbG9yTNdpiHGuIas2HsVBQIFkMijb9MVDlSEpOWE/N08ICUZjwAF7QLtpG2vFVkSe0hmSrA2sy
5StVaxBsicNZ0oGeAFFb96SwWdvJCQrOf7l6xhKVcZ6K+PPZeATCHUkXglp84ZGDqbnpJZ2mdA2u
ZjgFLyNSZD2Tq1SBv9SRHvhqPkJ3DeMOw//JKBC0I2BsEmsv4nBX0KRgGKEUjPiJpeknZB/sAblx
k1JX+3uuOLQ6udEOWcL20TeSc3agtipPfECLY462lqdqpf92q6rV+SRjBB43agJN/Eeg/1I8sWAU
k6N3tB/cQZxGnuAkmCs8jFpl3aa3R71zXWsph9Dp3YUclgyDNvk029wDIeu/xOE2iLZVvOwiw9ji
BcMYTyBQX+TPMIPvvYigvuAL7+zwrIULHF+S3+MFiqJi3nbMo/iy7mT3kHlOunv2rqTehapt3kQG
8KadVM+aKXtatBbhcp0vYvg9lwM3okazTdb+XoqKRRTyn8iwBSMJKO4MkpgIIKnwTvWXEoNwsMz4
k+THQ483AfLu6krMybuLpdZ6+XhNySBv87GiDDAwWt7deKBWY/MP5YOAOP0lCpxcSEzPGxS+DreN
JDned9J2mcjEmQvi5M6ZlNVvNPxPJhXW5sRQLukfk8svi9E3HXKxqWWWtbQucxOwVmuavoUVI2AR
DMl1zDrARF0bzsJ5gAR3b3+EcNk5e8zT4BBMbmr2V3wtVTdigSbbIPogij4z28gJIFOtjYT5t6k4
dghF8syfK0a8L8fWhxoeaSZgjrmGvy66ntYfNF6DuWtJ/29J8g0ATWYI3kyd5q8G8HT97yZZl8C2
CmVZ/quX8UzB5saDIZKrYC9dyXMG7nh/X40dfoi7lbbyUbmp0Xwk3tfIKW8sPsp00tC65S3doljR
gt4gJVf41YQL/0D8+YlflIcAypY4eeRD+v5O7d5sf2BkNNIZ/o7K0Y+4zFDSHdq1ucvY4DhK9Ktp
wKqk8EXRSUZa855pwR+ndnTQa4dfS84VtNDFbXD5t7zMmo3bOW3scy3/PWdOQH8aL6USGjNzJzze
L38b/EJBDTFvZoOh5IpbIn9Z3tqW0QYrbJPy/+8l/dHJ3YL4FYGd7aFz5ADe9cWhSEy/q6oALFEw
ArHBcnUNJV9h6ryu8aDAr7RQh2z7mlVcjnUaZksebsUFvIdVQJYwFmg4e6UxkzZQOLtyyCoz9eqn
O7nZxwUSHvDA3C9DWFdAT70HTV8L4MZ6IKGIF07cg9vQL8Tmz8RdXerMgvPRV8wGYIl8Q2m06SF6
geN8foS5xCzcJMJLgfoiBrNAkfjKkdVgyolrpebHE9/WUcJjz763pmybmPeu536kSc4UVpLhNIfa
vzV9IKiJF5aM0xdALRknMPdIU4rGKgHXb4754Vgs73f6j8ZORyEep5peCRQtLiwYN6VEnIcP5AmA
LhE1hD8jNh/1mntKHxtdLAKNbm3VYPcFg55r9Y1I2d+UsHhv3gey7OUwrNJeGwCkIwjtRKwqgxXJ
oXQjK/ZnlLETx+0UV4d0jPP50niLl/PotAt70dXhDS8LdLq8s3VjELkWkitP/xZMpwrUstduFIpX
6Bagw9cx/nf9EEKFI4RSgZkx84p7t+puAyDudvgqy/TKPGNC2gObGUIoUuJDN6p+Vb8wmx8c+2Mz
44qDvz36NPtkL9J3wrERu6JW6shWdypQQiHcOAdYacKndSjC2CQk769oEUBPDEYspyghLeJThUqF
IIIrfAr1Txe5q2s8J/YGSjLrv3eXgWABJaJw/2EJIY8TIFqX468/gAmpvXQgwrRRZE5QJoWoLtrq
tMcPmRcNeGsxxngYN08gQc/F12ZFRRP4lIEyWvP7Sxh1W+7MKPrDslUJYRbK55dPRjUvnSAql53r
Wb1hlfcuGXbbdT8qk3ZePagLJWlQe9BsMxJby2BlfOkLvVaJa1C9HsSBLTw8nrwQA+hBeE8AMF9k
DwE4B5gO65+VnBfp62aTvwC9+upemSsSIgFjg5pnsw/lK5lPlDR2K15GS/zP9aLK1qnRaXv0Kb/e
ayw488nX8rVdrxNvVQ+hIIgbd3gsDyBsIYORvoc66P3ZyNPp0AT1UoqfPzSdSbZM6Wx8kq5TsCQ+
ZtAp8zSUh4Mr7k4HOPLsa0GzK2y6MyRCy5fstUEH4jdRuLYR3avLtheBCfXjVtp8YrY5l6TgJyxX
P8Z2xoWXdUW7W1XlLfBSu7r0kUDBDoMAia9uyo0rYZGIv2alMaBndGhgI0VLumqHfgkoL/t7PwvO
NsgSha3xrkFkuQ32b8TURTMYX4oiul00RivXH/ddKz+m6OecrSCHz+sqlEb3b4Fv+izCjDsO40o3
fiWNKyfoPD95eDqv0AsW79sxc+rOvtSVd811BWl0aHR2iN037DVVh5XMPrHLQyImUNfl/eM/8l00
NsBGXTE6AEDGol3gaRnnzPBHfMAQYI1TyU5WbR7jwgpo4xxwWCsDBWwcjl/YKVlKc7qA6WR7j1lI
LF4z2Bz19dPv5+DljPl+sI5C+WM8dsJeiV5+7WcFlgcAQL5kejO6w8k9EtWDDAvNJVLAIZ2dST55
8Q08bFERH05aHIO5gjWWH24F7LAyLzYjYUTEXiM27UkeMZsgEoV+uFi6jrDTALTHaWji3xmAvJzK
Q1ZIKtYz2unVk1mDJ3V+wA/a6C/XTVzRZNvYUbIzUIDMZCkbzrYPaNxhqkezIS35m5qbl7zKlxA9
3NcomB5PQUlFtu92bhcsf9pOSho/JBOHB9V9YtIWyS9ptwExryklC/8Rk9KQp5m9voM++5McteHl
v4VXKkpRdJc5/qGHxmjnxkCjzRtzGEMh2sOVDMgi1tfuBXRwxBUv7hQi2Zt2BEX8dJJma+OxkgcG
qq5yOpfloZl9pJjZuyAKmh81hT5of8U/DtowxlfmRpVuC4lXw5whaijySHOKKcbrUDBtNTDVd/78
RXtkN+mDr/R7F23T7mZlK/eAhP6+F5e71Y/K7VnEduux26BtKveiwMD663d/eSCJHCf20/C3ZAO9
KqXko9DDe3CGIRlTpIHlwSkTrcgn84pzRznfiASUhAsfhPfKVhLC4RLQHeBucDCP7rnrxPlPTC5/
AiGJa1q2pv6vHIvyO5ERfxZqS+eyza5eiLKb2zeR5dNjgchPNZCtC+i1QzQUjBMOSivUug4PlZRr
mUbyS/FJ+l64s1iyf58ENMi9lrcKSqi/pJur5qEG2yohELuD0ocRDgBATct4P2toPiaZRvLIk2sz
BzrrlCyhsIQPrhhK6rLRSMF4RgDwngjX5BiXBrgQqPTclLoy3JpMJhFzkj2IRLhvbaHDOh8S9OdJ
tVUzqvX70hPUS7oJLWOl3HJqq6lHxN2yv8LosfQEWYjUB/fzdxDu88vky7y0eOzOJNQyKwTpe6K8
CeZD7mqmBC91WcJAYltwO+mK2UhdJ4BjLL3du8Iml+4mbQjse4GGgkhLZFhpYeDxlmUeW4dazZjv
6ntocMmFNnYXYV8be3ZjiRGVzfHwILPOVElThOgAtzfYxic+Z6er5lIsghVdMKAm1ITgzpXPPpy3
3UTPaAQYRpcy2LZ3e2zQ6rRq077xFe36adV0cA6RGdFjNSbOWCth+HRhro4RNtWxxrZ6V87FGtZM
bd9cdbzmKH5dPd2oxKHabxFfX79i4Na2tNxIs8ZI3oHE7EZksWaCiGlKQGxGXg6EcBYuzTouLM8x
tGQFwRQg2esYP6fUzESWQp4uo1rZZxCr+wuC+f0KlZRnMF4cCmNswy33pBWGe4j7TLwT0TwAgECT
Pem3rDgsog4ho4d5B0G1QcbiXf55tZ7Cuf831xy5zziMMiePOevNCKrlk+SID0F5LdhWL2Kc4BF1
djbIjkqciljThJiq+aB311FUql3qsDZZ+CWpzxauonbi+yxLSbWHzjIOLAq+gtn6vkTHuBYHSlDo
A+isfQcH6dr78W8AjM5DcRXNWi4gHhOq9cz31T2qGko3i5rf0Un2UM2tJMDAI0cMEmJYg7/38JJc
x8BHD/HM6Bvu5fKjCBuE64Xiw8fLMTdIX4lcGEaUVHxgY4L+NlQK6hrBbuBqVnFYhaD7Cs/0K3ZW
DPyvrdKKyjOjGrERvVThwzmeb+Y6DzQtk/0+BuOrqi7TN+VFVwiA/gvSdFSTtAHtC7f/aaVjGH37
1mA5rB8GaaAzJ+rXpjpqpBeDEzjhWkYHDgsoZ9HyNFBqTaZgVVZzxBZCElTHrMR9z3lLmaVWvLjM
HoTt6F55qJYeCYFfC7gPQ2xGDRsfeK2rPSiRpiMcOsd+phvKcxiTfItcU3kbA0VthdlrXqo1VMEA
5anXeD0lBzo7AZves8QFM1mlzBqK/M2tkN3nIA6ubhipg8yFEdCdcQWRZD+JE7V6Cd03k37DXNVn
I94AibcRxzaXcd8xinf2B5g7EemfzOReIAUih4aveqJsvnKoZNzqxHjUIdM4N9hm27wkKjWk8V8J
xEkch71SmdrFzN5zjb/N91LLuH9MdYhnGmlTZtACILdojPLqztNsqSgEkaltpibxJrfx0Fzw9jLF
i/5QZMbURzLfntymI9zPf+K9SLoNtd3JZSESV1vGSQivo0krdO+1N4SpW6MP/L5V4OxBHOpPQsgF
EaleVD8R/I5PlLk6zKV35uU+o/H8jB3gd2jegRo2tS9xMR8J6BVKyvvOv3/B7kV81LIq94Y8BAXC
eTAUfo3NRvoZKudm4cCLhrPRs0WDJ6McmkiIKJc8M4a8/UBUophKtDWYkZpxRtYQb1B0xDMoJVmm
jqcxKmXb18S1ZPG19pyezfA1zf/zt1aMdxzsgzegltDVj3h571y/+qa7QtFCLw2ERJzEC+d1ne/H
gGWX0bv44e+lvy4gg35/2Rx2zsDPkwEt/CKWsZU+bjNjNxbcSxBTIaoTyVQQX8YIcqUx0KqIjckc
qGP4mh4b6KQYq8sifg7ITjabqv5CPxNoIiQP5DD8dNq7JgyKHvWwNnTsMfDWAdsPtB3dmQdIkDrO
LMcIaW2dDgtIz8xBcUfI5ZdcNbbOTVbFLpzNK7qH2yZAUjQHtRadFbmlMZU93z854HUichzm0wed
yMeSzMpKipJmmap21j87t2ROkmdcbcdonb9g1uGNb7TVS/NRNBB8b7f2ryLwileIBGE+NShwuSsN
zcNZLEBgnU/Hf5/+wqRlIHl0SnGJ3dPnvjT1Lzt5dVb7QXCiz+I4EzvRlAOiA5NlaUWPrDG+KOza
GY5a8GdmMk6yg9m/5GSfknCcGgEgJ+Y67ciotctY82cHzKY3guGwsm35nEg60qv3lGRa7rZ4znxI
lLkrlmVwbzM3uY9FULKguL3zDJQC3hSLiOGeUyJr6X24ZtjraEtc4Tmxf7loWdIujNft9gFbeMpS
32xei9DKX1n9/GDq3daNLxzmx55Fc6IInu0kAsXE01etAUMwC8pXdwIJ50eTpN/tM6u2hNHTUnLc
/2lggv/IGSOKBg6KCRsp9kA/kwwSyxXjgaxu7qESP7vpWzBLcaC0adJyVBmpAl3yZ87ifqNoGWme
cXA8COWSZBmtWZFQ/mOv/cofzrXkfJx+fG/tJCXTg0AP5LpI/xsjCeT0T6S9B/6ZhlxidThuncb2
sTLCEFFQUptFtDFmoixD/QGCrvB/igz9q1VsNBhaUi9HEqwgunIA96p3DFOGbuP4/l7Up17fHdcf
xQAEtElvCkkkdQbvtWzwl3kcVcVVZ0gkegs7QfqDoHcVHHa5+lgr5UmLLLYYTiEHqF1nJV0alAEh
srli/Q12f/4VO1f/0Jiox5lbc031oA615xu0fU74hNzsbX86/ULS9BMjtA1VWRyPsuUhEVZeVpS9
nbVhsHuQSt6hy0OcAyUZM5zk5TCg2mBMIze+oxpaexWPBKTIVcPvJBtA4SqbV05p0Q76PIuPRImQ
uoRKPP9fhRxXoM8Yd8QZSuhSpkflXEBNkiL5u9fOkj63vwOBKsidS7gIaQ8762HS/D9kVr9Pe0zV
GUVPHAil9OEYZQ+kGplynLBsP4WgE7vZ7v+iBOgLiT/qei1pZHP/2Gbu2Q5lOzUQkvvooymQbTD2
BGOMjAOoFsEDn/UuvSD0bMfVuEAQYbxPOIvw06Yelbz8HBW8+Oj37Zg3NIhkVGIiArxN9+3VsZFC
UMY2k6SujUVbmhBoY0pfDibRVU+iyWy+JRcT/5ScVFQRrYsTY5YkZwAnc0kNPOYVVcdjZa5v72IS
hbYtAc7bl/JLnP9ubHvpsehA7th6i9fGq9q4oqGgLNhManEPLkvPuwYmMkBmCDhfSmdE15iQ3IUW
fqWcPqw+X8jXERxzcVx9BsTGhtDxmJ8vR4uihG66wc5I4C7rfc+/rgrzW3r1ueeFTzx6D3CfZ7O0
/he6y4Q2biOc8/gHzZpcZ8P1iZJZiy5Xl742ElJ83tVoOdFB+yCS2ywNxfrVw9SsLbIFKxrkZa9m
96u5SR+CC0OR41bMe9Pp7rLb2xMNIAJ6PxsU/PG5lxdHpG3N7wQtuOHnh8FaNe40xSluNLVer0Pu
asksNA0qEBeUfVWx761AUfX4OYNZxpeQnu+mcey1TD2xnU0pa9Aw5/Uh+cN3OnC2o4qieWcb8r3R
Te9I3FkVws6/aBsf1ZMpOjpvZERExXf7VdeAfOJ4ndzc3sqsgFqiY5CUWntF8ALlRqYPCFuFoMn3
ETh4XXss8oSLofadk25UohMX7SNAXTEYX8rjswmgtH4RY4pf5M9b6Q5CvVe+yE4HdC1xcxi4jWNG
U/rmkmwuY8CB0nY2tofwdzwr/WMW+R5LHzb+hYaGqDcsa2bDHzg3Gn2+oN4DFOJnPl6tVchBfm6/
fUIX4O4ffni0LeaxvcRa2dJCrnGdg6yAnIi2k24/B3jimFUAinVyAQBtvTGYEhRwuFobqbSJPG8s
GejHd2RYcIVH1uHQVk/XLL3RsXFMT1jd9XIZcHseG6VZGNf/1Lw1vDkbigUpcDlsYopxq4HPC3fB
zxoHxyu/sac2MG+gp0BMzkl1KKBdOipyQvq7powIqmaukNxOB7RSp8ImpIlzAhjPk4s69ozAE7hR
CLA9PkMw6UxzGJ7+yHjLUxo/Vk1IB4BXwgeIiUc9BL0RFwwWZjpQZzIBl3V8WtpR0nWEJx54Vgj7
XiPQ5AtJjLMEPu/8/jEjjHntiBDDrEsQcBuiTWjRWNJQErjMhO7D4iIKOjIAUh7U2S29idPOZsql
8BAuCUkmsQTM74Kjkvliepc2yLYlSsP/3eGHrS7Nv2UFO1EK+CHGIXMVTSJK2vC2xrHxyezI0opY
DBF7CMK5ZwKv0MOBWY/qDNYzQlZ8z1rDiRYDqUJbTdGSsGlWMz55oxV+dUd1aJrMbeIXxjXxAtce
/LLVcTM9pK99KXE1XXKXkWn4OYNTIbsc9TSUOPYOf5CHeRgRQwt6FEigDbZeh7gHGFdM/n1cZOpp
tORbchZJzIAVtF8PR1NZXK9KEpTZbq2bGRAY0r+Y0b0i/6cB+MdqiicZv1joT4gaDuXT5kIOG6z8
6PA6F2Y4OxKYI+h/IxhG4nl+iviA2w9VIkNgU5NMy5GkLZU8IPbvhqcao4u3N/KxdCNGgx4hzxjN
T3DiN7pdWzBk6o8sSeMyt9IqQbWyJYDw3eG757ZwBiYdKnWh5jWNdo4RHUkvFb4akBRxxpKV7z3P
TH6pIVr/2wEWLm0CE1vDD8Zvqgs6oeIHOHtunJehVOoxQX5b9QkQnPAnfE7p1uwTtch3pzwe7S9Y
JGszOi/KhcKyhUctAZCkd7gH5vv7ZsuFUln+G2nAKuSpoSDTanvihH84PN8CaYDUaLtksXKCta/G
E/OuJsVVZnDqES9sRW4CxMFoJ9A8vLQCs5yi1pnfAFZIzWyli05Diy/N+Dy6tb0eFXb7vC/g6gXR
WEtFlqYNkUEq1ajX3OIuflkqY5a35gYcNoDxgQFx+4BbNHxeiTW7cpfXyWmQBI3RRwoD2IQ9VWd/
dLnh7w3D02pqOXKVLgW8C1cyCojZXeTw2bInjym3nGjPZXj8ZBZftR444gpcnvJ37xGlq75g3at2
GtG1BWJEZdiTI4bAKe3/LP8lOvfXJ3N+F+OOMhH2HK3XQCOGBX+/PDIPsda2dgFfiTiuA60dffPP
fPrzFQGmIZTh26lgK1aobDDmgu4AX3ZNW6QlLmrjj/ajzhT59lAwW3haj2YCPaYVYIi3bklS3A1/
AzwlgNWYH6ifSwyGk7grnJZW5O+vViMpZmWUqlT7sIu5eRZqAdxmDCfzBxTziWSuovo0h8dJFnHJ
WN+42VL0MF8trPKM9Irj/oloNypOsaB/J2BKjGinVQOkY9tHu4lwQvv6KxgE7rhrxcShFQSYKyPO
IerB5ju/uQZtJCJig5worBhzGphYvXr9Z/RWJYUdAZKRIV9HklvWo5vdAousIAzHOmKOiBgZIXom
c2WzABSx1eQKdD3FUO0MeHNbNWVPEgk/jqV3w1DZ32dwrpew7fEFWumuF/k03vB0wd6k3abpLVl8
4cuYIrWb1J1qmU7ZQd9u3qhLu6xjDo0dbwpjuZMpPd2B/mPjHQLCJX6l9VZyt7Fzn7eth9wQ+i2X
o32o+FqyNMevmz6LSiCickvIptwQf9VSzGE5cQXff6Wr4WwvBUHdenpslLZLNgB4o+MNW8AEQ7kz
joO97x4uxAmpYG1KTz4cA0JXPGV8ylbSyvUZrsm5Hm7v9L0Scm8qh22bt79ujwi/m0Y1/WVAsGuA
ohf7cMapRS5R/5SRZhWwO6jPHTYhtHGqZ4oqLazpiZFBGESAZENnbXWB284skwwp4y/fxuI9Xz9k
CmrhnLIetiXnf4pi1742HlXmljiyM6JB6fyT0F+f9/C4VOXU06zWvqHS0bmgKGIX5vLA82GJTJkV
iVAuj9iv1RV3U4+/YO1ZvB/t+kEV3JI70VR+Z5c6BgxPtWOnDyrnyBgRAAyS5r8CCFzUfwVigOHx
Wzezx9iYYGCuvQgb3i5+CnCw+iluWJq/qlAO5pn22pfa72PDSlUPGCT0J54Z+ekGB/3WV7yyGUTt
8ultNdnJwD8Sy/SLcH2Wam62FzOKOUptlN/LpWWZe9N3FXp/3rIpMopGzg516gyfmVggBbyEhC66
z5Db06Mxd9iIm9PJDKFKqVLYWdsudx81MFJ9vF9Hz37dkxUxt9AG04S8Olh7qlEo+JT7PAvG3U7R
MAHgBifENdj1JxOm7+umEXopx1d/g3SMHKgkm1GVXAmUL89zVsHPqRthPPwdc8xBNsd4Xr/40lv7
w6N3cRawewvw7eMRbvk8YzNWh/+8ziDcNrOY0K7m20JT6iLYALUNFQG86cAwHnqee7wkV9gOU9h8
TOnFbZNYvKVbWqZrgQ92C6Kp5XKfSLkU3geNQXmkek/y1wLvlEBB9y9oy4Vg+41qee+w5tmN2D6H
KAZlXTpJpeWrDB5BQlOtfO9Uf+mRe5V6U+ZhfecC97yT5wqtvCNoA74nOJtliK3MwBiohdJmLG64
oBtfpQRbmSqRn5tkhCv9nPHSXu9MawjYCGX83yPCe5Alco6on1LV93XsEds/4KCfNw5X9UHQsTjP
XzCw50NQPaYcy6LxWl5+5ggtGXI6gs4G8XewkH74z3CjLjXM073GkbglvVOye5y1vh2HrkBgMQ9q
0LDv2yBy2CeiUIE3SRVW3ypiftTP23DB33BusQqUVoRpKMbHZFX5XBB27kAMMzmnnfmydxiLR1VR
z/TRv5tYFG3Go+7cvQ0U5HtTk3AGicOt4ZLM4qny+ZBVspm5WT4G9Nq4E232PyP/EWlDvtl3dyI0
tnijgQnlO2+f0bdHXHj628hTLk+a786B4XMIUIz18brFkb8zjKNxRpuouxy51qLO0N9VutbjVdXm
DaKpe3G7KGdGrihLMIAAiMNZA8l1vhi1hnE0hb/1M3d3RqvkkOknJfUgGfhGUtYj/RxHLuZkV/xM
CVfXSlFNax3X+JC1MsrgHRQPYGU13gvZGdQoOjhTTWH9nEyKGp+i0LlqYdMBSaDTJ82Y6R9pdMoz
g420x0o2kOpoL/0AUTQ6nGdHGxPsWOWqhDS6k2WyhEpkZ1SqsDFt1CVPRsAOOwCjZ82J+eW1dGNo
rsGgVP9+h7lxyxFpdvxWD4GfXgyIQThZFzJig9jGupoSd06cWeu33uKS9vQY6P++vLdgCIj5Ryud
Po/60p8JPI0jZlA4sgIJPvCmUr8d8dBHh1HT4dmTa9HbyDSH//5u+iGJ17KiETY4uXILhs9unMkg
acCfKCZ61vonVFT98ksJFhZcz9a4QzfMIxAdh7VzqShgJKXFj8TUCpHorma3BT0Y935rW1JjP49Y
vIibQquxtEzbGrta31W+plK9RaPGDVwzYb5hlAECU8VzV5NnOyziTJu4u7JiaYLNchVEclHdpEEs
+Y65WTfEg6OsiraBuk6VFhw0z3qnH2ojaXdT/CxWHXqMK/ucE/mADjuuP+vIB0x4sWtA2StfarSv
i1hj08AISqSFlDQryqHnRqz3/UGpPzTzTnBYr/ZSCO5DpxTQ7nAW1VjduuXeEuBALcRyNUpV1xLQ
ie1Xf82+r2p47IL+tvo+skxM65GHL8kQShfJuF2Y6JhxbbrSZnVMk7smxbj75/hU2hN8WINNNcNJ
RvOjJWpFNDnfK9FhTdbkAlWCt5MDFnXdFw9T6N9vFO+iJC70M9t1RjSeb36j1bTKvgS9jvO3TuLF
IRWxeLNsmNBmy+w9eaFTSX+P8XfKBQI8y2IEyVTSGPhCZrULeYq39Xg/MdJ3SXXbxwof/fLMSjEa
I2vYanb69BJzqdI3VFazJ4wpHQ1YPpmTj5orTa4rnSBOUbOpB0W7Vb1b0fWHOzrZKAFqccTW4WGG
3SoL7gDjDEn4irshdXuoHon9RO9JIG/ZXeCjCzpi1gjRSSPMwkzIzPHZkdshl5Ozw+9keLBQpy1s
kXuONDL9/QXUXKPtuvnjDp7JQgWpVzRpPe9rXIJBXxeL7XJ5WoZI3ZkwCuJw4GR2fcvWpv++zDdx
pjaBykeqzCccJbQlGoRsqI28ugnyM4KJohRu07Okm229jtSemYxJ25/go8ZbajAVgq1jeJ/0Ryew
MD18A50sm1OE+8dehGFptQnZw8yi1EohfgnVaYanOxVrKi2pBDLKl20KBpTal65y42GqxV3rdUdA
hYlyPMU/g7ZYlBT1fKKTfFIsOW8yhdpH38aWNGtX/Csa6laG/QE7e4W7of/72MdR72zX1ec0AEUC
is/aDIVsFFshknKvGwjSyde2bGs5tTO2xrGVSne/VALnQCOBJD98K/vLPfx6T9Hpc1EvU5A7KysL
UnfpsM4dmbWuZ8T4mcIwdn+7GjBopYRbywbQnJxe3SIjxDjWlwB7O0WHkVjgIq22jyFllfIYtv+o
XsnspRg59L/H7nUbbjYeACF7556hyL+ZRDHJCPwWG3zgyZHGCjcTnku995VKGZIArFseZo85Po8+
k1Zri8XEmRZG4K3yAbKHtLrU4AMalUGg1PR9oY6i5Wj2k+bGyjIKuAgxr1nh58fjF1tjpTqVnPar
HTU/wDAm3wJkT66A+zIWb7gKoOBzhO1fXlPDynr7fYZHLwEHSkUgRxRBkFQqf3T1hpvds9yXSbTh
6zIiW+IHSNClMKqbJJ8aQI6j/d+W7qi/idDu/7kJFvGJ108Sct9JGvyKmUQ/+zxLXa18NpKh1FEA
K7wT3pXraHGZLvNytCSc+46skJ5+G14pSQAG9z/T0WdGz1J9TNswD4FSCDUTJO3sZmSWPpFZFhvb
xSDzdD7Q3m5yxzFQ8WF827W9uSQ23ehQVEcrcDnAFQYOGjXOVA+wTsFhou6FuL0pWjSQOTAbWqqt
R05CiiRVksKvkkelkexfs+xG/0mQtYhoPQoaqrewf6I619NqUfOTSHhnROakRfVuzSyNgElaNfaH
ifDsOjMpfhXARK7BLUdDvkl+0sF2ZEYX3K0V3fyh/Q7rqzH1sDq/X2csdN5hdGh2BbxXndYahpr7
ocOct2j0pj+IEKG4E+/bnnFvHkfsfc7m2d/x9kcIuVtq2oTGaZxNRlMnJ4NdDp2iUIubBv9FLfwo
0+GmGDZ0p+EmTo9EnqOWLdy/4lJis86prF+b27di5fU95jZ6wye7f3wYy6qj38qCcSHbbjzlV3HF
kVHjUvrVio+Rhniqz6KjQjjkgvphkUr+xJq8qX+66q/xtI7mfPxpf/HQGejZv0XmObf5EgVerzu2
R+uOd34rMZD3niqm6Cbg+nA2t8IrZYNc0AN1f9yZgymChKhkSJB3ChmzoN0wmYNfRe25bv/FcVNP
udzOVjS9tBmFWZTvIDJe87o6RgnOqphUTiC2IaOVnrMji9pPGkIOwYyYWMebFhxGEFVZuYimWda7
ZpjKguNRSt3LCpDKSLSm4tycw2rux55Lp4xVoSSwafq1+ITlWZEAnDz5QWcs93aljzJX2hqwlV9B
Zyw4ehj4fObXlqMy+N6qOsu05MWhSuR89NODwEbotSCjSfTMV/qw4yhtGppzXRBN+BEiN/ZLCLUW
NMHuKiyzrMEtCK/SOrLQHrUGagRPi5WH+v482WAuJ1l+zQKpAfXWw4y3UzqHD7fxSTGaDUgrZlTz
6E1qBY4nd8tsp40fp5ta8iDq+LtxP5/ghqkcePm3++YsmuZKvdjx4QbC9JeMjsgshlWVCuli1B60
ru53LA6giFnQBKjshR3368Xn4AQDAA+VyntuKv/XXNu4nO8sa5eHqFYj+ksUgkc01U2sVaDZUyKQ
4/9c3v9JUM2PMFWTS5VYbduCDKLw87EGuzG3z3uearLavtiar1RTfqye9MOnnmLsy3RjqK25Zf+4
+wzWVKjLXAyg55RpM3zA8xu9Jym+p16IPhQn1PVqJegNKIb3e+tuXfrd5Yf7smC3w7tBGGzzUwVf
BolDnLTdgAYfB4SR76zVxZxwZ2PfBUfdgpYbL33gG6DF98o9vANLJpGDj+Q6/4VA7lvqXEmJCy/Z
VkoVBjXGQjqFNjkYFJfvHp9aYkm2u4xFSipNQRe2i0FHOUxy0cs67B7BXGjFSpfx1jY5dcHmY5UR
JBWo2kLggVtbZAjDV2knRZ5yARYANMRvYs7tXhFiBFrOI4cO5UswgMWlLpyrxi2Hu7cAtVl6fXmo
gK6G1pvvwoTKY+LBb4NfVsag3FcUb9Gzgq98iGlA17+/IkDGeYvTLEpDP7D/MHf/qWNYxtD2Pd3w
TI+/XlzAUw8Dm0R/LVXyjUTjIwlYJp94PkqAzTctekguump9+rRqwtJ9p+Kh0cqFQX6bP/Rd4wF3
jiYwHpXwW8/OeBHWYkmucvPtfBfERZhC36LTaILee4X1GZy9tkrynXCQjBNNmpBYYQ5gDIq0i73b
XTMFw66YL4DmY6gKPwAHIgFGHoK0x46gaRCyUg8W90C7yCUynhFFX6wQER7V+QZhk91dpkbanOXy
Z3SsFQsAlG7OJb3yJG8SMe/rbY7rreEPHRP8UJ4mHPG/OjVI+EnPL14ouMzNwFyOIh52yXPTee5Z
Uko/18/fnEvbbIKzh/oSiaJYUm7MUAIKOkkN0NSWOEdi1Vges9oO1EcBYVdFx4aoQW3hVkMF+c1S
zfOTIROrbFbcflmV7SV/Advb5NugCudMDP3DwMblWv07vH7wBZ6slhaHjGTzqmO2OvYt6nj6I+Go
jH+IenXrfSBgkXn186sMgprozfMkRBqw/6MNYTtfIllzCoe9SgDCaWgDXU8u0q0uYJOeHLCr0tz8
N8uUJ5t6GBfMAAsqhmVGzqy3B3PIy/xTw04LzZSzfuGe4a3l4uv6cv1WJTsWmx3yNhLlxH1dGgNB
WvH5lHR0w2fwgro+h8XtOdpV7T13xXKFNG2NTloMsFpNNfrOVmAinq7pG82f4Zma653XbMyryzrA
edV7YzLib/ZrBEwhf4ZKdFqFC91HXWCEHJmQurYdHqpY/e6rfGm80vT8g2MiIZ5OmTAGuPgbCvWY
l3QJ/HnecrIzKwCZV1l3LENVpLci0EENKBt5/0WFJJaY7Qjbg9yInupaGLnweZaJVXa8LleT2EVR
P85EbJl2XmAhWJkeLhPwyOEArzzpy3RjDbho3/xHQilgmYNInDF+FuW7ujdCoc0ihKuu0yXREh89
hmFUG7wCpgpcKEUyAvMk5CLX9R0596NsCalHOLXR2bR+AFy+ZakZZgW6Rt2JA1z9oGvhXNJjvEh3
RXOdLfUGqWuUfytQTQiefZCoi8BRP3JcsAK/vsMZAv+OOW8/vxgybEOp3mMdSd42EXGSB0af6805
IVbpPMKpmi0KaQkEaEw+r4zY3W9gFnSfItYmDpC2VyQGa7J12irvVNgRtPQIrHldNAMPl3OnkYoC
iLfnUwb1eD9j6WDPmuNflm2S/hDFpwnraVGlGBhqsxZ5DtpipdBrA768ic66Nou6Sxs2d7WrQ2t+
4jOXDmAFabkBosWhE6raI64dER2dEiGbblQ+4U5MkRj69ryPMlIv2J3I9+dKsEY0qfYzSxtOHZin
3TspTQW+FlyO9nOdXrSPrDS5P2Ob5hsVJ6XLYUExlicSxw5S710I342NVZR0fc5IyGGNbuMtxztt
sGLcoOpgepbMXlf6tU8JFpfUjL8ihTVTi2bmSZ9Zn++FUGpr/5SEzMUPS8Cb7RZ8B1A4ObrdtdjG
GztvCejKJMSBWciODUGZZxuIdG7blGCQkaysAbgT5MYAXHhPOAD/3RAXekCVYjj64jOSKUw4CAOm
lL18u0RtQHI3H3j+N7tB5lMxPf77RUzv8SVcSFHM5ALaoi9wAq9N2GElOLvS2R54O69p5tJusMHt
Pp8Su//7CDpPvwa2+Go7nvGdYYK982D8p2GjRx3GXqYdVp2FekUyykNIJTKATaS6VqVKJQKCHK0R
/E4UC6Myaf9F6INY8wRXQpyyLAlKGtl1Hcw+Aos5fYdnSBuK2fALFuyXzMK3qC3yinTxl/9CYSno
DiS0wSobMFugHhwqa0RjQbHBkjsRhDK7QEdedYldfDfcZuVl8PaMO3Mk1/ZhP+ifodPOojmf9aaV
Hs4mZfcDChhxSAIiWz1j4G8m0K2wXY2JLECYeomsPB4EblN8wbXXx180GajoHkU0Z8XWRy7I1VZm
I0m123nsBjo9BWd/OHdvOhDbknsBrhHS95mwg3rGRuQYztzPyR0rFeP533iyIulPZpHjDqBURBJ4
g1kGsLbGdaJ1fCA9XC0rfSiiptnLpJRcKtVERlHyYGY0Z8dAeGc0hWlusS3pmB9GImE0Ek6dwqtp
k6NcIGAD6G2duYHqEumPQo8dyW82lXFBkZIt8X5hYY0+Fq58lXzBCs3obQxV3D3mArXyHxd8Hplo
lNeqoLitT6NZMCeqETqq/3m1Pc0WRFjmUlCBShtrQbWmkyTs7jY3RwgTOzNkNDwHFjyk3wU1zVzR
QpkkvE/mHGQMlkk1YPXfxG3WDKJXR20J5Rxk9n7Zipe8JDQHdQL6zcTWUcvxUyw/qyJhbczBu2AR
pVBN2GbXI+2m+9UhniA2GXmgNeOyeGqeO7hnq75NJq96qZwpSFL8J1lKX7U+65s8Crnl7YLdkL+L
p2zsmuBnn5M3kz8PdCkjuQIHiqaMw7EUPg5M3hqT89p0PGbUYEqzNnQyTgj2i6YHehVwLwmNzOn+
ekhH2keSTRiOneW0sytqpF+T1yOO9Sa6TeJhzoCGRt+YO/mUhb3EhVKHQqb69vozY+zBbFcUi9M1
EHF0JSjex1CJkSMTL2w79jqe1kYp8m4G217ysCw8his+LgKrnP1YEfYx60UaqsdjSWgrmH5zzY8l
gquVtUd1XQ5tc8LAq622YB2XLjZkn7WDqmz3p34S9/gnt9yxXcrQEazjTx2OAwoyMLjMt4/gelwr
WdXkBhC1Jl8yl8DFiiPKtgN/ilB36kq4yhdWIHtdt7CwHVwHi23IvbOsKrG5Zus8JExF8gGHuMMg
nSVsq66IhYs3vqGjF+w0GSOo8mwkMfSQRXp0kqJdfLPydZ4u7ouPVvs4agsJDw+ZHNFBlY3WHpHF
DUgDj4cBpT5H3Zzbc4Cj2pIyf/Bjfxa88OE2zlCq7D9RSMbnlwCsbEE7/kJEYk8H0gEtp2LS6rtn
vH6SZ4YsGLzJ0wFVFkwU7qWxswmN5pExhXVfi1i3j26a5ssLlw5PgVedLj/WyMedTP/7oOIDx8Pv
sD0M5uvOdas8bixiGIv73sinVvd4fPJPOeb6ir6K5KXaCYE771QfBiJT3qSscVKgPIzeQaoZixnD
3Gh2QEZTMvswChj8isGlupjTRwD5ndXmym+/rmJiKfcI2FaJYJHpayIUMma+jIj7d08mRZkFoAgT
zW8GphCsoW5rC8ch8rKqhvoncIlROu25ku3cqVV78LXhzeue4QuHNV+q28wa4gFLpOQMrjGBUnSd
T9HbNHuxOF4AJqRd7yBwiGAIXCI6CgeU4l833BdG+COY4R+ACdDdEyONq5PWu0vTonHd/8yJ/hvv
fDYuln8Wot+0MZdC9IakHg8Vb0cbxDHyhO+er8wtmoZ4b3rs5mn/p8me+J3trS3gNnw6yAihOS6T
7HFBXN3B2iX/tmOg5NONvMIxjI4YUjhc0qyA5hRm1aYbJ/aQz7pGu8NHl7a7pdpVjwvc0QMy7ckj
I5eHlgkgtPQSeAEkdk/Y5vwJ4wvRyuOI1pNwWXixdMUZr8fkOpga2VTW4TgjLTUfSLz/WnRSyzbI
USPM7aIN8q72euzvbJAQiHIJylZkVhv6/Njy91lGuOiEsXLkU0i+DsYr7Ynhej5VyRLRjN+Ek845
sZn7j1nMTNILqHa1dcfLVflETnTkPe0hFlAr3Wnf5JMSEZYARLvpBDMgYpVO8w2IqHUKmzgbwZTM
8H9LkN/79JgSdiVrxzhxCC/UOWBom6UxuTVGwhbMmnedPId5QjUIMQqCCBfKLO9Aftzx0LYN5R4N
6OOmKILdxVpOXn4/dN5E4aR9z/kb+9nq6MsIzsOuHNUQdO9JZ/IoT7IK+G6OKGKLw4Xv5VdRt1oR
NBjOjAEZz8yu3UKa1KvjDB93j6vFy80X0+chUpiCXBXxq5/m0t4LVvS0BqbP6kbVmiwJlJnXRpPb
aw+ZswtGCb93eA0mNVSmN9SCxOs6Mi1D/8GK1voJf0OhMCVaTIc05LD5szMoeoYAccVvVH2hNHKf
OHpSp97KOD9RCELeKajWgK6JnBKpFzVnSbJXmaPeNEqCZWvU02hxUmmyDvC5YvifXD+mmvwnZny6
XMaYuc084HcIEOlnXvNLAS+LJ4dATG9YvTmGK92sah/9yqu10Uglej/u9km4KHqAuqsXYSX2+cfx
GOfAMtoSjvEtHSaFOIrLSCpZ6TnVHCVWJ3pp2i+3iQLvv3mDSyBnyAvtaijO9hwkSHBUhv0hhZvM
csbPxwOGYmz+C+QsnVAnVHweoJO1RAe0z4QdHB7iyn5pSZtbsefaJwda+r1TTkSeY06ztq9PMkoL
0cBkZYS9Zy0apIys4mCWEiIRz7/ZBPOx4k9dfHbVvI23Xbcpdv3YTJfJVgawn6XDLj1/E55Y7+l1
kyp+XqAg7PG6Y/DmjXuILV9Tnq3VF6dyCUl4+8sKizXrh0QfWmIzCPOKIyF+D2yCcz2vskXanYSy
ub4wclcm0CDHu5xK3OGYa9EyTwGoTXDl+rn8q8Vs7nhEUfqDkHDdzEigHEF9jzcxUrd6DPX9KpSO
DRbc8I36oZ1ikzd24qYrrgg2EZylHtN4xtSxA0RvK7/sgtrlNtzAfADkqiGqNvCq1y1qeabYNHY6
50xD9Kqm7+w23+iR/vrCqlQvloOD9DjaIMu7N61dkh4Iu1fHp2c9X1m6mrEFylbAF6U7xRz4J+Hn
VhE9OsX8ri55Aqlu85fBZ5AiH2OaOWa6W2n0U4U0vgnawGkpQ3SN3s8u4o8aGABtCSsc6E+S03k+
Lt+8Kx3NpP4DVpClX28SdgLOld17GZGQpN1LQ01TzTE1vMfabGqIILfOYnJBC0jhd6HR7f773lQE
1QS8+mIfyuV6ME9dwY2aqxT7hPoc2/Z+hw37a6PzMmZLmevfxrn2DgsLkVoRyj2vhVMVVjnNIIMi
ir0I7w0lllUV7pi6N+yH4IkrVMCGUmAer3zTVkbdpEB6DIQNgQg7tJulq3K2osCLb5vhl/l8hoZk
u9mP6pOHj0gti/Zgm+Ce/uFz2vQ2WQBfivsLdqRcATaCRmDf6rDKU05Sm1t1Saje7MHO5oyBdFF2
OvJUf9qAHTQHwqrTuNnq/XprR1tVv19ZIwIwxmVYzdMW+iKR3iTopjfMB7jucqzPgVGBcvM5RwWn
iVivSK60+bb09W+O5wQ6Xd10Ey7BnLHSKrMM96zZc9RYwVt11WNIYhgKBF5BsehSqnWmmfN7JF+T
dJOvIaoe6bMF8sXTDCGjsNu363a1fx99kc5OjZzFAAsVHiQJEA3qL1L8wQrVwYKZN9k4v6XQKGw6
WogLS+g1fm5jbCeLzK10AqNp5ZhNr8I7t1krRivvkYac7coSToQDsRO280ZpdCIoem9uvNAwnuH+
7/MIWwWKtcbvl3G034z0SiM+iEbYa170F8ONrB3x59J13+cQBzRiCLqUvmQpYLfZi8VPzvsmGEKc
UQMYoBuU9eKHc8/E43e3oU49LYr7rvCPC2W9uY6ZoiAubFewAr/lMn5TqQoJuKIbjwzPPymU0Dx4
cLLZdbKovx4leNqpVfPi0nlGHKNOHRptRrhyWAqBA8m1cFVJ5FBIeWvV61uALK4Ih8N8nmqr992o
z3LT41I5kOmDRqGjd8csYf3+Z9pAO9Rkb+al9qWPEJKQ/JnXVNH41MkiQyg/3zXEFX+9gxFZisp0
pTR9UtwPMUwu2PYHxU4rkBgKfYVIm89xmhMIo9poi0e9wifc6lxhJ0t5MByMFH4mmv89JeFhHjU8
NYJ9GYcLBo4+iRvXVk0ipS05GSDmF7ibtph87EqSVn7aWiF+IXpoJRvPQ/8pWlsah67BqbmyWS4H
gqBLaUhDuygP6PyfGkyvyYyZ5NUH8OaJLMogqRHtj31fWn6gdAoB0xjiB+koVTTaC4GnGI8hetLA
r06UAl5QXbdnM0sSziTn4oOGeISdvodm1egNFwbDeLpGVRFoPYTIruAMNQo92wkyhxWkzyiT02yO
D6D9oOlQpvABA5/Fjub6R5K+2zlPsZzkU69j0gQU889Zcs4IXYF2FJXhrQPv5wH4gZLJKJRlGz8R
I8zoBrjj9VdFZuG0d1RossoEU3ynFYy9PWI++zHlvjmc4K4ygrIRq6cI2i8YsYMP2zHz//+bCYCU
3BPJSOidZqs702ahKxFuMxarB1yKE8hwFMKgerDsWbvicWLiCxi4/4RFyXTP1vTr1Pf/kdzLe+fv
rnBMQrWgLtbEFEKfEPUPfD0PuS+J4sX8PW0fB+9raHVuxlxHwY+jTqFA/LfMBsCcpB0EN7doJ2EU
HanmjcXRDzV9C0BcDvPyL1vmeqcIEwkZp3+v82LGpofnGyc90D6neyiLmo4eCM+ir5ljRFJtymRM
X/NmXnaqNxi3auF8gjUrCU9UFShm9RrsihgHYkP9i/DQnoHJUkx3b2uffcELRb+GmKKyMxFDHIO+
UZlesmFoP4XewhwgQ+2ZR99RjfERES9v+NJUhxk99RN/Z6yoXMgxqNusGblfRb8m4URAxi7l29cU
H1f0sDas6BzZ3lQ2+eky39bFBKPyZXtLNPeW5odDbw6y6UPT+ZtjPKp21d/iY7gEgIevv1woFgdw
pHhcKMQcXTGXSkVTCJBtvhrs7iDC3zTYUmrTsxJwMO8VXHY8J10rIT8Ig3RhfTcsJ8QS/cuwSco0
i0Y+lM3/Sy4kg8nJ0/J8BF/f5oYllHdLHJ7dURra7M7AvK4rjfO09t+mlJjhp+xRk40qVRwZ23+H
Rw6ohPM9klYmMa4pehRxdAbCBaq/chjA+6t1sCdHS/OskztyhSf2QKHjBxr2wcwWrt6/H/XWrFZu
GFgfjq9Fp4N5p34Ex4fveE8I7Gnn2vCnvcv05KZql323lmfSX+1tq6M5zKRalz5ey+EIUm4t6ZxY
F0kG3GewsP5GLY1ZpFyiX1wnB4D+9FiFPIpiINS+/d7QE4qGeBDkv4eDtzsSaRFh7Lewn2W4hscn
KYVdIUHduXdnWXfNNDQXFdNksDytNSP+JUX05M4EWW25Ij6xBWUf259BG5Yx/udLRtGv0Jt1skX1
sH5C2nGYneCNt/1Obs/f1QE3IHXF8cpVBlkW92r47A6T7rmAdfmKZD3TqeVEK95snje1Y487fvRe
yzcfZWOBIAk0ji1inb4FrKtH+DJKnh86DJ3aN0ulyWR5BIvBBev7rNnqM5RQUaIbPgJIACgz4X8n
vOG0hAlgFcwZnvzgjJPCzfiVPiCE85aOxsToRvhBjs85ncOZnQvSj0EQpyyIjT6tfmAp3xzQEzWx
7F98xx7SE2wGNVs6KnFngBM/UlMPI/jMHb9S7lr99pTMi4owV1gOB5R9fxP11jl107wXEsH+aXDh
E8IkXAMrAjS1cN9nbmZpMv1eqmhnhWuUjGyVgq+QRkzFOsGX0FFat1pnk3y8IGbSuwdIcvEDfCdR
n1861Ufep/dY2QBqado14NhR59rTnyPhPmsqDwowPS6hZXM1477CwngjA6Fa+D+pZxAv9cuXUwDE
FGdO7rG0wbAlqZwOIAGc2IsMuZOL7Qu09X9e4K7jl01jRMvdAT1MzYDsWzDRCVhL+yty43dJeDur
hqAIXIHYgpRxBiFqseM09g9YGsjS72AFANqSIBvpVMj8A0R+KB0dRYON7zWv+MBW0a8Kq5ti9mvm
FjWD2XF5MLwC2Ufq/4JdXMWoxrfR5M4ZKBcIP9keZzRnnbbQ6iF5oQOIiVXutf15ovWdXL1il3O4
qfr2lbZf4+IyUJawAjIHzYHlestSRzFje3S19lTPGFhTj7LOUCsitaV0MZ4ss2rS27TCzMty+qPe
EIAP+05VHO3CXo0DegeedgaiAbIl5cG4DyxkBcn8uaT7M8mzmw+baOmI3D6QQbSyyu2YWEWAv6ih
Q1S6/2okyam0KHFMYiFHjjh0mMEmnekiUbIfOYlXqzhG4fsKxEYq+mdvFM5QB7nfDB0S12uwaW1q
jPjFr0cNzZJhUhUSVBlcxol1evj3VY1dDdg8217AVHErz1eZrjX9H3JXIzvy96Eh+UHMLnRfuPf0
ANaFFcVMBcVRRpsL32b5bqwp1a03/1i1gtfWhF8YWVW6OrDHmees7krD+h5ly7S07EuphSHpDvzs
1+Qu73rh/vmtpZpaHkTGdxGgGYOqPuXgbed2W84r7tdYQ/WaLcrVNsFtFboLomPtw9ym5/4Lp5HV
/FtjMyZDuMLghWlNdIzVPvUbURSupqXatEXJhGc3HtorjsibuOeaj7nTD9yusTpatq9md9TfwPzL
Z0UPTr72nNShDJ6fQVIc2w2V+xDww8WNe8EvT7Qj9Q2cPPRf1ImVH8azjYTqe71Xecmyz9sC7Uni
H9vWjLj3/uGITy2QiRobYQJLVeJ18JjYKJfuazAoyebYyl4/C/ZbGg1JyQdsU9YgJXgyvGnBywUR
oDOVMp2PLT51CnfDdmQHNk3mMfjc9nGI/CDKN6GcZAOCwqAWbc0zDXNnbbEaHTYH0p2x5gzMm4a7
KKxWpmxKmTZp//y8SajzB1B9s2FtVHn3ngeRt6WMNBmJ+CqG3eubhqkmpFYHjHV/NaUfGArtHXZ6
pQhXOeI0XpfrAJGOmesNzX6VDMlBYtt9f9jCPs0dCfsUCDcfuC1+I3d4vyRH120aD5A6UPIhiJUT
KLEHCI6wBSSMNpQrlPXaZsvCqDmae9jl8t0pN0sLQFLESCvM/3dfUUoBd3LkplBCS1ZByW3ctxfd
7rZJiym7dPn5E0Jfx2H1G+UTvru2YMWVgj9yB6Xv5mqEdFsOndfq8NSeK2ox2+BIJNigiN2yPLH8
17taBroaEDOPAcZ9jGC1RZ3FMxJ/18HKq9GNc5/RAwgwKsEQ+08UAvohYbU7YOQrwwLtl31oSVy6
843F31NO0FHfm1W/odgdj+Ap4G/MVEQAajuxsUN0/DWkcnMGdtozPRCGq1o4+kEV0kYHfC0GATQ2
AhBhCPhloplQHcV+Hf/f4BvthK6VxbLO5+OVIdHa0QNi4EbhPr/YGki4CP4BMOy5w9w1mDhBTRVf
SaLAG6mg4+8+IwG1QPQEoiEpzF4Mc3D+Z3xwNJCVdtyFSGglCBmkepDNyB2zcBy2Yc3sW5QZBUu8
ERsCUKygmIgu208pjFE9Alhu7SChiZCrEvXfUZkbwNV5hzyV6QQzcyyOOaYMVi+XdLlHZ/zg1I7N
1+3yntFOFg9xUYufXl7lP+J2AO7qcWCV4ekPR2SzGtuxABXJiApNE1To+JVEotlKbmkQU2U6eD/f
8QXyPH5E0MhP/N0R0XSlg4csA2zzBFpk3J7zX8yIGiOGCiJI92z526qhyJmV+/Vp2PHVxdAxP4xC
98l2o3Tcg+LlNyiitCJ18/v6nUmM/fmfJaBny+sCZ59NpG6XxJDpxRpv/M0DYpzeeQygseTJuKrQ
Ru8D29s+cb1m9BTicdR3a9KoqhNzM3rRDZ0iWt7XMj52mG7eYyCo2MRBCw9Mx2WFcoKAlBRPs3mh
Ds9z3c8f8ZtSTnV9GUKvYNIbD4ZL37uw3l914cugbDA65EbWMRfB6/GcTjnma1rb1s1BlONtAv0y
wOeV2/BnluTMue5eAJGohtjeu3ApCaDKlhfpp4Ka4jW8j97CWksPzTofMGsBc/8z7Vr+5a2WAL91
AAKVhunSfjJ+O5L7zszYDxcwYh+S0CpSLxCZBLoOB7Baq+/xZejk0NPszy2d/n7iMpKmNjShX+Wh
PNF5kiNwegU2uH4gPhh2nUKAu0t09zy/iZQjBNzb990bRynV+v1DyWq3WPM6jrxpX+47SlIHT2ig
RQOJxlzTWwFRcG9FnwUJioV0PEBotYbB4TDUekB+86+jOzn7omYF1Ic4mTxMxOVAvuGOyfks6u5m
Y1rjUziSvZIcX/C1NFeS5p5aclBxzKfcV8sw5nQg14BuMN/NC3hZOsGxIhtZkHxVsWUIEVcqzFEe
TSzaNVNzfhKhx5V06FoMBd5Y5OhjIbTjbF1z4SLxUdGBYkqTletPN2/TmOMWI6BgCUk+eVV0BcHg
L4U46esaVgBohtddS2S56F6mhlnixtVTttJulwH7aFY0ihOfJZzbB+s2BsY3aYQgKqP0381GPXzZ
/EApmMgbI2BrWMAmM8cYQf9yMkFgDeib8IZqUdqCQDjCFN/sFp7zMnbS4Ok9CoSMQc6uQ6UIe8dt
PbDal2hQbddlR8SLc6yQ5Lz9MqkausYbW98QQrkU+oZgWhGMDLgry8pA5AAyEbYVUCp7cayCEhKl
SoXig31FG81lsDlMVB1KYUhszLQZuSt0QDA8nTm1RKTSCTgYnj2Cq3TNdBzbo+s0w16gQjR4oahe
47P5XRR1hFqll55tua7ryb4gYxJARvSITpceUgtMk6Jhs3ePPpwq7vGygXsnLLG7xVC4D6nhDE1k
akQZP9XzWbrK90F+pq+WANAC2cumwJFEfb+eBTnEn+qVymu+ji90ESawHYUtdUlbJwRF8vTbqt3t
HteX0ngusoP56+mlMidhUV8sXPMJ5MYoYZkhidLZReppX6txVea4NqI/ukbNlf3//GK0addglEwc
ySyJTyjIutUb4LTibme1CmC11YyeHCmrbkIPUd5dYgrLRbvEgGZgJt5ZwN1I45AEhBZgtEfZDnXF
GeNOlOa6zefFVisLUaAhWf7oaRaa0yUeZVvKIVFZ9zt9CcfkW1mZm0fktMHz1cTqgsRRx5zRrM09
idGg/znkuiUtbyaqfs8K2TPOtlh2ve2vMJ90lFohQupF1koJwJqtB4PUcfAbFyEHNKNRtkog5H8h
wCEUit0Cq+kV3fZmaan5mhqzesiBqP8cVpWPVeY4MSxjT9Wzb+DVjhsQyUVFrlAwepq+KhENNWR/
uL2HE3n4vOR/kP2/fqMg7FxEZRWvWLTj9vOf4Hn/+KRQ5Uq7BJRdtgrC8SLgLbpCliku7QQE57S5
e38xYt72+DSbWkIqd0MSpbjVgGtew11RZ00j15wIy2paOZJbMbNOXWWiKNQZFRDq50StcHGttAku
1Ei0Ltpd/8BFfPX346wIXpe5qLhBh//leZxKoqDhlG5CAdMcdD6+J2T0Idoz5Z4yvwOuoaIMEoWw
8kuTFju6D8CVGrkmZS/Zcn3yl7tOhwC0XLho1ngQ4GFRsV6mSgvoUcPUTdHq+5JyheeHUYyUj0eg
SWSEgL4Hv6FfmTdciwPBdAHR1exZ721rnOsL2+PpwglZnrddQNyD/UNlNWCw7/0pSwJAUnQMnCri
ZuTD05/+N+JQnwExBmkPE0QXpJ74PDURGyXdSa56vr90i1ebPGzEzwJby+tLdpCP/PsK3hWJQdsA
+ek+sx8kFhT/5qUQ4l8RQZsI0uSJYp7pfCMco9bREa0GCh3pD20DIHMxXRbh7FGt5mmNL0ju3Pei
9FNDtCiXbIV1R4jGNBBpd4Buzcgymgru7VPND1gixLa98l1r+DK+mGGbKYYpc3Fy6jS7gauazCXH
kgsDV6g19Up0LxOe7dUUGAXzj0Qn6aQvclmgLnOnzMi9GBVnUHCWsrwTdbq4Tot3M2s/0BVsmkdK
UdWeRvKkiXbAPCrCHjJawjWJHTZfBtCrA/n5AFOLgEbyRydUzBzlJXv8Cgiupx70pt6fCSMwAWBM
VEH1ffpNL/UYjtipRBnVebO1/Gtfol9QVOkgDBrVjnkFi7Imy0WA+DiosdzdO57pQGfHVFFyAxxb
OctvEZsr51U4/PlYLY7mAdg4Ho338wbdtM4+hwT9lFNCdEc/xtBcepKma4YvTOTQdtxgHfIjzAN1
w6NWSMl1bV1Psn06dlP0g303uIkgpprOXje9MFkSKocEsi4Yiuz4F/7oF8auE6UqqcZOMLO5e1IP
TZsiKVXx73cTLAMpo0/D6mp12AyZ2CKjqgk8iD6vgV9Mb/7MxO5QIUPd9ezgf4XbtlaYas4Nd/58
4vErbRVD7YSJ4/DxQcIEMybFDnKPt+ZGnG59AmXoTOJfb72vYaxu2LLfeOKL0ObMWo0tI9RJCWmr
tHDgdqwKywPQJKetWzkswhodI5ONjhrivkAuCewFlCXchLI79QdiDSTed0T8tDZLwPpAZer+tnsW
6LyVRTOldHyzMpZyLOPUb95Sz+FnFKJV4H1h0YG+ygXPWhxIQQ+aunWglLQpyU9nWSqOUU3nIvR1
IGBWN0q5bNVR17V6d2vk/Y24Pv7lDtjHSCL/VEv5vjTsd75B4ZuWgg6CHcaixmWlopktUvflE7Fi
glclEzgsrxk3XoKcQoUlxoqnpdk0FPJ4h3e0NpeeYS/1ZV+Ptr7xPv+W2S7lvf9W4kAg42U5mc3X
KPyhTLUP3cwt/shILIv1BiSYSRbUXomc2Jo2XyyDn+6XHaqEN1qCVQrNgqrp1mmXyFRjfY1eZx/i
jBMeMFVd87cxM/4ZbII/2txNTFQ06yNmt7LND0J7ByJ+jxyIVnWUxgdB7q7C77ocyZscTmkhN7QW
FyYafUuqq4c445HLGHvUc+bJdK+C/UZQfnIhsVtwteUPb1xevYGovDWQ88+kJvNpvmgltBFsKlEi
YnO3kZyKiBHeGzVmto7OD71E2o8zhaKWovcze5jRb8lk24xnuz/qftx8/cGTA38F8l3Dsrr3y5Pg
2ykqFc9nMCeSzTpMPp6InYVLHgitp+e/dodz3kMULcrG2niXAsMN2yoshfp+VU1kUzgWySkCGPqQ
O08XlBKtPoEugJoqr9dHfjWo91Hyozub+579ZB1kIYYvoIxjaROgJ9JvdqZ7domEOZELJN16XwiR
5K/8NXXkmW8nK+7E4iacxHtkktp4tTbK8c3up2yiv36vOMAS+LRq7Oj3taX2QDuqDC8rqHJLl+3f
9NHhiBDYZlgc1l5Hr/vaZ9x5NBWn9xbbXPkun5mdfcFbCDZGQudxafTuyKPlSDELkL2boStfT8Jn
SoZQYCi6WkI9oPuOZOOKD8uswT71Ez8pCF6eonoetWHn9Cvkx8STPuJy+VwzUe1jg/Y8hOmp38DT
p0WbWuxBXvPFQ7KiTbWXAJ5LFdj/UPg8QQo8BVbscuC/CRop9zQIaasRvmMi686HO/uCiAsrybA8
/GLKQUR60X81axxMQh8QlHa1Sah5Lc0oP7PgyRsOgXYyaTHkt7f8OLf5gPozdok4bHYNuCsKFLXZ
OMhLfF8iKkqu3rQW1ALq3VPc9bk5NEfSxfISV7PirU3PuWteJ+qsACHlKBn8fxwtHxvdILElXnrJ
gUFu1ieqCDaEOoOxd7jQdHee86AuAxQiNTS/4fIjgOHZUaF/JYJX440PuQmm04FM3xtabkpn7Z+3
dXDP4hm8YgP4TYAu1FXDGPIZy5mLl2GxzEo9AQq2MGMGeSuR1WbIlr27e7NZTlBC/IPhRJvCra5W
ifcYjnq/oeYLOY6mUNbLz+AaZ1HcGgjgkeeQch3VcvrqZnJfCjOoXvqv98tnsMRr6Jv39VNI1cSq
2o14DMN67lxGiX0WZWuFzNgoqCBhJHpFs7hlkLTLHQHovEZuWxIMf+Y70XMWDCgarF+tRVnLBUzS
DpRGxLlipVWbiiXNDhFCQIn+Six2ZmhBU+4Q1YMN11duiHtbkJFZGnJzJ+nli0CqEEE4tUIQdzvK
9d4zuR49+a8Wyk6oe1kfr38F0H8oeBrfGelblsWYFCRmS+ENirBjX+gHrSETyZ+1pTK+76wVtYk/
xr4q3GnFAxp5QPGjyKgjrWlprBrTKew91ggLE8EzqDymQc2fi1bqyuJCFK34ZuAz5OAPDh4xD0gw
56FuzupAnztg4nMbr1LpJZAYGslc9nfoq8BVW7YF+T+IHbgZbVrwDfSXDawuDHtJrcErZCwmU39M
VA96j+R+i41DybvaREQsS7xqoB/zO5YJK3XrQZbdSIKSZ6L9a+gTa6ENcqeKbcxqPH/qcpjZauv1
9r0E5Ac+ZcW7zvoW1XsSEmxD4TfL4hI1ErHWfHCZp24kWrZT6c42TT8/NVtO8GaLnBJZXq/rV+qK
LPSiILUhvitaGuvUFAQ960eGK1b+F/l+cA7T4dwCUvRl2CmMd4xHKbXH6ku7pIpcyC7ua7ssif9s
HLERL8mUpGBIJCTxv8MtYAlmkfdJOSDgCAAnNv/NE/nQwefWMGRWYMqpgYnf5VmE/8q80SJqhlAd
34pykDsgqqSKJsfYGplTp/0hlBXylZ0634uSZ08kXJ8V9TA3nHG2qq6uXU1U8ofQDdwPiQL+bO8n
KLRJxYcLaQ5dr8/qLPQ+d2EdbFIikmKxuNTisyQJTfbkqTI4gH48mKfoTUdl5mYi3UO1yB/CP2Q9
vQlJF6Zt6VOfaIfYLMrr1TZrrhOCrU36SAEiDcAbYSGtT9hB6jjce3pbIRLRab/MDu3FPfyaaenS
qBHvDEkYdKSOgznc3EJqwJSZyFKU4CxJA3YEhEcJi6eSjAgYSLjB0Q7wQ/Fu8sETVqFwJrlPYTZ3
89DCWGz8ym0UuUjkcP9WPjhsIoYGaw+yO2bRR+nCtWR4ebM+R2P3E/G9fMJTyvi9LbbGpeOL3tmR
ozW1MSSj434Sp02uMQjMPG05BwE/e6e2PcnCKCLeDmVZYj/PsczY9dpPxcU43Ylt3nOXzy12vzHW
IIdXldk0TajPXHd/cNUfr739fY8ojaScL9LkgQpWH2qsHaYluZYXfPsCQWnVxSDSBDCAuk2T0GFA
MSJoc2QEOp9mWOf9as5XDoEPSF5ql/DpPJg1ep+deatKuT1sOcprMJC9KHmszhdWi7mqrs3zex4M
MZw6zfwyVfh+OYhyxlRX2ZhXy3Zx2BCqg+cSDwZkiRODiliObqGSqtgJ1i4c1ZniEUe0KEzHSWz3
dRLYVTK30Reb8pmVunbVWl0MoauShUkorAu7m6D/3SH6TwxNuwl2fa0SF1bZqcDT09IonbEtfMWq
uIB1feIwhbg6jfHO0wBow/8A0Dc7VfHZsnZDpuK9PnFWCsoI9yLO9zCQ0P+VhtaqSrhSSlrAKC1Z
2NsciyQS73enN1UhOkJgkIbh+2b/oJo8xhQKWDzakaYmx71EjxVl4VLAcrkNP5lf67+mxmG54yQk
FKsYgHxUL3+1qDKQ2LFp6SB9IIsFagZgFjghOgt+bxYP1xFtJgaAZKmsQcg1DnwEYlQGiia1guvT
1gdBvexN/Fx4VKryBMrnPyWP4ij8XeKPwnJvDqyXM7gv8wmvPXpo6w31hV/RR+Bvcnfbpz4RmcMX
aBAZm12RDRWITzm8TDopwyvxnBIkbXbRnxT8kmDX6Txxa8pgomYEvdtVxdRaZuBOI5/p5Ow5ubrA
AEH0Xkzmd+U4v1cCJhplyPcBuiWHhlJPtfoeU0SsRjr5p68AuojZo3hu0NgGW0mUtyLkpXl5LfiD
mEaIl3mIbsASB/KinnVBwH+Ke+6DZGTcd0Ew1skUp6XUUTVZWKaejW/b02Dv48V0KUW32elCpPEm
rV6VLKhPe0fMl3lZcj1mm3VCXd5xLnHEvx/y9cc3x2tzLXhAag3llPnzhYD67KKR1C2pd3ktoXId
WCSj+w3Yq6goTA6WUv7YO7/DehqTEluo8+BzgWUP8UyWUrRWlBgHtCJYW04Nf/5BpmPUivOOC/95
riHI3A9Fa02IOvOMKpGPmOZCnI59OtlkKnEpfpFA17Ubywaf6YD4c8lNTtI8CxeayqfPMngoFoJj
U9P6xiqsUcXy3/dnY06O/Bssq7FbxO+G0ewzN30UvMJvflppxw0dfvLCe6gFmDBuSXjz/4+mNyNg
KEefVD+/J2vc7qoccEBxNLRBWmbwmr5dGTOJCXZVS8y0qfl4R3tzE0cNjJyYCccEnwb/7BACX1iU
ZayP/a09RkmvSdmBoT0oJrd2wTJHelmB2K2/txlKLDKu51kRwWQaddDC7TixNW+0EzS3li5hTpwz
mkyfu4+rhRb9zKVR18T32sj/WjDpsoXKb/R7cDfnGqEYjmBpZV01UZNydDrrKbxKhkz5WuAHwMMl
+hEwWdBdTxEmc+mWBfkMRZaf83f3gftmJpx5P/HiUdNbNaEzPgUEvCM6cFch4UIkbiVsimOxSxxv
d+90cnZCL/fUqGMYNNwLQBROmIxvGgm6ts6e9CRFWA3UrlZlNFhFyvfme8/y6MBS3Az+X0E343qr
xfICl1sOQ6ldpwelNawGM2uGPPXnfZrrnr/276g7AHVVG9azrLDxiGZC4o6JIN2ceHti38EWvlc9
GJHI9jmXFhOcxEn4rBaxab4qsl1xWXKGkgoik4Qh/i6mN+3hsEoGgJtyhAJA27AqsJE4f4zl9SoA
4j63878yzp7T8S8fUlYHo3vq7pUwVwXC/35+etLiVRcUdS3kNKXQWDZE92aEpzCTJXTDZlpz3Lem
efXRlbKEamrneWdiXrtWCDpedvd4VnEn7ykj3xDP1ijLq2snpOIX48HW1UPJgNu9cgoxNm/kGKJs
e0plWfaXOtKmxyLF//ktw0zTXHElVvK4tR3QAb32/H0NdTs1OrWEsIHwXwJ7T4rAaS+OOswi/4Kd
CgGAk+4UuMDlbUYCB3bGA6V+kpbNJwguhRL0ctY25ORPVroBbMvOW32vb/P1iGkm00e7bI93ZL53
3GSNAJ/M1FXfhnXNQBMRR0JpB5atOAaqyVQBsk0/ik7hZq8kgkoysAvVcPl2YRCUtRpkDcPJbYJP
wPluzTxq2Z1tOWu9pqb2cXYwXpsSxqKBjEWR4COUwN6QbDOR9tUTidCrg+nk+UZ6j5TWKamDATCw
WcmR+PIMTvZPMmFzOtRkPfelH43t2ys6MNX0oW1B7bCRe1sTh6hfuIq79esCbRU4a4Kk7lB8hwUO
L05D8QjaYwqF4/nZcMZG1pys+tkf7mUSRNJgH37UiezpmJILmNkj04J8vSW5+OKCCjxq3e8T0fET
qb4oNorLowUl0C7J+sBtDmZ9+QnZSfvv2JluSYr3OVXnymIZxTHP6Elz8XNMKeUTOknnOpkOQ5Nx
66BydxBpqvX7kWo0+HR/0SWdjm8Nod5UOZvAZghX/NtidrhHbfzDj1ZpgBQWiptA2MI6UqQMy8Wb
KZaDW5YN6r7foIC+M8yddveybvGngAv1O0/OgzM4HqyoJJuWcnMTHKD6FYYKCvPKJUbBFuLEcWEa
Y6zwR5Z2OiDnmDptOE/1WkKA4gwvWn/ytS/OAHK94GEVvjt73bNzIygQ8B7DwEfvmC+s+mZDriEa
Z/O08y939GaAXK006G2xJvRCzv4VaOmGH/ZnFhYz4J9xDKpeOyR4EQqoSxUhfxeKIaq2uz8fPz16
nI4Uv2wmInTtAtKpo90f+ocIEOBERU6385qcVV/c3krRs+ngMjxMuej15tgOI5mAk0kRYWAya93U
rX4mFnMh1dcgnK6wPoPzThWSXEoO8sZOidWbmPfGdCPvuc4S5XIewkq8VjrqYVa4rvafIV58Rwk3
5ZD/hFxfPD4i0Px62euW6ocb0vr5m+HB5Y73MCyzc0WnGgduvQzsOGTGlWMOrXqav9ZN83oscuqn
d9MPQseOXSDdoJxDHbf/7Dxdx3iVbu4ZhKOX/ze2SkBKiJqai257kH+NbtprEXDH44hZunPjKZSP
LWgIblePTqRZ/wdwISRS5+MFQ7H3mrn+5dIWH+YzqOzIoLxUXHoqR+PuZcfpMEuCWjm0rHNoHgZg
OJHdHNwJsI5k2m0PDV2b5YIYECv0pz0a+FrX/BYDty603voEGmV1zOIIN4JvywaSO3l+7i07uH8q
0mZvZJcbV96m3LHy59KwvJsIjn++4nKXjSUicpuMjog2DjmitFuDQz0jxVGYNrDyPvm+UXHtFwlc
4ktuJlpMof7OkXlWzrv0VG6qxcENu49dkW5lddIIcpceCn3uFnfY6DaYwalvwIF64ma78K/LPHOo
7KXpASwGyTd073FQCqVU8On/77VmTOZM080F/j5Nie/N2HVV/2XmwJApdq9BfpiaEXUi1zaTM8/g
udSST/vaPGj47K+BsYkDhM3m4PaN52cpjmv/Hj4SpTpAd3iLqa7rTfIb82Dpo7P+kiy3Gv3uEQ4v
WkTTr6QNEjrYwGfGIX351z3eG2P6h8V616h8KChjnGq7CBEgkfX+7gN01IFL8t0bnUn9gA8pKTT1
rL5PPGxQWwe9UJlKK7Zy43a/aN1nvgZuCU5WnpU7GXRwmakXKG9k6s2YmtedkfPSwtf+LHNE2FAb
jiaeud4yH6fVrImxsa9bF9u/rrUiPan0kA3HnzT08512YNpNz46vJWoat7h/W4W9KQJE/PmcAgc0
dYbsVEe3PK0gZQ0eQonHAiaho+8kFWQIeYwnX9O7ARH7Mu72/ZrbboOPnifHAiBfZ0yGNItzG8uT
5cX+8nsjClWcN4FfxwUB8obqH9Q8B9v/WMO424Kt1qd7R3K/oPeSa2YEU+0RJThbuoOHsVga4jEJ
SbOJaJA+7pm8wuu1vZAgFZSYslnbJwGaQw5JQuFYNfkZn2q8G3Zt77pmKz++a1yEYzymgc3UqT5b
U3EvK7Wt8GlvS42jtcpi7am3QfhMtZcmfOvbDOyWzE4d9DxB4wwmsNykqKGPoiHXiJ1bYs36KeQk
hTJJYZTPXjOWwF7W29J/gu6iZPpp6n0PCvLB1tS/V5WUsipgjX1DjRAlnVWckEek6DpUx9ETU8Pe
iqJ9P5sCbyCk2x0GtO8G55UuKR+PridiwOV6yK/GfciZ1MTCbhWg1yL57wFxdE0DYSF6icIMMqDP
JXAzX7qTGmo5pS0478MOmeCqkPmm63jogn/pn6Y9ltWPuaxONkUWh448WjCjhRlVxSvTCEikHZpp
++WRk0kAQMFWz40qE2G5JNcPCIW9drxn+2K2ZIbtDozJi/DqVG+bwwLQwBurA7Zcb7CfQtfyGadh
g5dONP1UjNdDzJRHl1sEAAULaidaWFczKHbsd3BGxkFKpzko5hBaf02zNFMbZFjZXDsEyXjt9lwP
7WLGnvBS4nIP7vNDcD0KjWb3EdPz4lpbtFvvNhZ6eLg1/re5OBUiz6HHcaBk78jG+wDmM2DBDC2S
iZ/UqhNxelLwnpV5+F8qAQC5vVtsFYiY64rVY/HAV5v0b7LP+NLLrxUPG7OSOLbiwWdn2qj8FL2/
XLP0Y6qhHcCexsY89sg2D82BplEvguPIXs4mMBpEHRvxoIfOtf827XV6+w3ERkIRLP14nqotnW5Y
QWx6pjJPw6tPoXZWrYDHblYxRXd9YOqSk8f+gHfYFLWaV1aVOsVHU/n64b8p8zGifQ0pUHRix2TV
TgTlTxz/d3GQgBDoPU1Mn7/IgX7w3sQE0sWx9yQ2RF2vYEvLNtBSFNIjBm1TDENIWYH9PkOi2L4d
arkeo1vKMSa5W8duKtb+uzgaptpv/Iy+bPXrAeF+MUidqxlxOOLLGa4xBRxQg2E9FSrBTqz8vksX
efQtDoe4erOjNoLUCeYci/xyCdHRhFRJljG4H1+dpuQ4IBwfn9cm3dZDm4uoEpy5tKpETOkapX/7
M/n3UptmWAOccut7vhGqmALpGh/LNh5YLWtu9PY3/Kc9MWZyb+ErTRXPm02DN5Nv9wa9DeNSpM8O
R2XkVovP4kGkob4PHgiA+H8pVmrzjfVtvLWXx9WCVLsbaOJo2Pp05BzhuBcys1xjPwqmBhOxeAj+
LHbTnanJRaG74x3wv2ks01S09e/3VXVrwVFmPgd2xzoRsj5Pow43jG4DFimJs2ZRj2t5BXV+nska
VT2e+IsIZfLj5JJWD2oPnGLO0GhvuvH+2ONDe5UPU+nnY08PxEw+dLYoCWLR1P2U95lXwDk6SKpg
X3+PnZNf3paIHGNYx0N91gOblgyZfulitmVn2+vsZGughvISfE6hyUfEj0CK3/st/ECyGkbStkiN
AwUPx7e6oP7VzcG0PRKJF8/b2fnq8r8XWIOC0OqUvxsIqZGtHxS6RJY/lBtbnptMa63SkKrI+6KY
Es+cQanUN7gEYcbes8v4LXp/y4liHkQ/IAkXrBTL6JmUWWEW7eDpnuskCheUJW4tgxxN3xztL+0q
MfeOHLAD+AcVC3VtcPeulOQSgLoE4L1YV3tHG7DwaRc+HHL6aX8A5v13UH478+9Zwibcw/WZ3QR5
lHixssCfFr6Nj16ZD/rwBYhE67+DlvqGOtiaoMefJ0wTO1+HHXw4SZ//ZXgQ5uvS+xV1qmJ73hOV
A+NtncOM83j7uUs38RFA1knKrrmjOF2lTeVYbPFmuP3ajJ32Mo2QF+FeDCTkWLJsXlnvZ4BbahCV
9bA+vNCt2yngD7p81liDWDSxFKOGavhlyW1OJvzs9PbHddkAx2RyhIBZ48BA4kHAEgbHFTxqRmZH
qEUFRyWf18FbZFRsdN3+3tED5jmsIOrcdRL+oJhKeWJ7vIlTSw08p1TM54p5tY3gZYYFWu+Jwdxe
Bc3/0QC338sDnnWGRn0ccdgPGC/u7Ff2Itrzgpneczb5gcwu6UVdg7/xJIM2wWdzXGOgoJt/jr3+
KCyLqyO71zohm2M2k8g3dvbFkqI4UziaT+/1QRdlChVynK/89K581d8VQklwClqHzRgbCOe3rgkv
tVwxtAQjPRtnqyUlMj4tmXkjJldhoYxcJ7/aYU3dfgklhDgYi8SxreWLttYHBsoLsb0LVt6J1x9d
FOhNq1xayUSD42f/NSfok0H92z7tMXqmUabZwvvoWSc4L4AAJTiiuTOpVNBSuAunZRrkhgj+vlRK
9u0gyZPs3BM9Wcej0oiUf24Ks2wV85egF7H+JCLD3kfZiQQvxCDhdvfRwDi6FurVSiaOiHzxwfXV
/dyRacKqHYyMc3ATH8D1XgTETwtIE19dhNuB+Z0eiH9J6q2CfQaSRsS4PHJnAtAN9+nazVwIrhS9
7pUY3Pna7c7mFiwryZX8/kdvEKxn+FQACs+jeFGLqGtw+jnP2EH21/htEPlhisnBEseMJuHUQ5pJ
UmfAZRMlzp65FUwpCz/x2TTm0tp5Sz9vnN8F72SAF1fnu4pvtT8FUzSmjwcOelDbKZQ/IXbm4b2z
WoiJF/FEOykWoWUa8m2VrG3fDATDHCocS1Z7kgdehW8shQNjvsHtDHsxWrKxOgoGQCu2aUWuLhlS
LX9NyErh8deTWUPAwarC/SJg0uNiGs7cOwSVE6kSWDw4WqkAYznI+D78lBWohQpaMeVGSDMTu4t8
q1SILyeauEdc5DC0AF9BmrcOTqsDdE3b7yryb8/PoW5I442L8TmZCyiYLskfKAwHnCwHHeXq3TfV
Nqdpm4AxxrxVnEkdOdQcxThu2wVV96vGKkN4WoKFiCbo3SSgo0IC4C3pmRq9m0Pz0uwQGVrgO2R/
79GyWYwz/GzPWbopBK8k63EHqMgWKZZT6yzvzTniicRqRPEWVHYu1umxVpoBANoGD8/M0TbvZA+7
7NF1xDHIzqHxnWoEbG7hrHa/3tFzY/olKT+tKk1uJ2m7D6JMpKSqri5HQcrlUQMjus10FAiInfRm
0T9zUdyeecoiZi2jGYiWC170w0/kCPuo8ui1VlXaMmyDA0mi6hTm7xY/1LdKf4ubJ1Qt2IMU8gmm
yJMc2H9K+ujwLqPRdf5OgUvT1LFJw1lberF6GQKXCQx0zDHMOLESHQzstCmw1OXesyJVgiXcYwgm
nNYLtGns+/d+D8Zme9rXJ84PbzJNh3H8Df0Bf8NoAd5Q/ZPIl//n98O76NDu0yLvKJH9Fbf7XK6I
gEoesJN4FHCfHxnOm4X/UNofPvfUpA61jnYzd+4mnvkFAJ/cbuocoz5akFNNIB4V89cSSORigk6k
0k/kGfNOUYMf8qO3Kti28pm5sImw6efTOTln6lZBqna2iGEm/qfW96l575mt5APPxj5PJ70n1tlt
uDi5pBWC6Xzd7K0UhZTml6Bgsr8psDtbO4RwA5Jl4XmWTPdtObf93Kdyw3HYGpbn8V5oT7DbSq+x
K3mJcupmnqQui+ekCJj/IgIHBqm663p7uy0vLR0wEpj4bytKhbYran7ZcojEzBYHNRBDHRRJ+gqJ
HqgSbQGbQ1QiV9cFCI/MkQdPCQNCa1HARlgL5CR5RSo/y5ehowa4ygn5HFBWiEAOg094yYe97jY3
NGWVKYZ6Fc4ZH9u3Jef7fJdHP6c8EZESUWvGiub2vO+3lpVxkd19totqBsdVxDRtyLcbriRYXcsN
4KG/rTbwAm0YuANv76bFlCJJ4JbmNeugGD/HC+JWiTj+dJKYtqsFQBenyeHWeHEk044lCwOleBjt
OcX64XIvaJAdU9qgY2/e1ZgMgp82jVM7bdP0QMqSrZIg38rVywY3BHI+af1QmwfZsQJn+IFYtclT
7hpF6h8MI1KZbG9PQqrUJTnM4IKcg5dF5VQj6jaTd4W9rGZP4UayCVgnt+O3QAmZhaYBo6R2Ao5P
Wh/NvBuPP8zz87Rsj2oIrYteeFUIg7vkj4upXzedFujRIC35AxOJXKn+i2G9sC/jPKvqC/AALF01
6+0WTDPDkY7TTPc9AEk99iwO4tnqCnJ357CBwV69S6JwGAvz/8SHVqdd8c2TvybjQz083+pQgZNE
yJ3jJbhx1u9I6i8zYxX1u/w/4v5C+kZk0u7oOLAjw7vkzV0bfepE9KwrCi84UeNFW9sm4jsCc1tU
QxkFyAduMkFHUPLjpDcPg7qhcQR+qLAdPhU23cXI70rhYri6pK9jhoHOjd0Li07bK5coCQUHBWNB
N9zICaktPFPOvNeHYakhVyHzRDNeYT4oIMsWE6XA1p8o3iHqvLr5P1FnhQOHaGrKVLSQOpc7t/i4
J1f5+NVUeOvHyGWpQrG4pO1qPsVGgza16lGTnm5WaJjnJcTibMTioe7qHZTHbmEH/vg7Gg9vBKcC
QRNZi6P/4bm5Rm+vq4vX524oaOcjMvCgP/6PZJ4R/P9bD2PYWMfwKK4mi09Y8q7zTogjH1ahAlxC
WGtJWS0+KcT6mFBFBw9LrEjpPmYFhHSVrZ+zCWkCgflWj2YnhXRVbTJTpQ3Piv0PFTDXUZ/azo34
7iD9w+NhUkpsly4CRBkrr0BXF5WApt0AShIMwfl6bkRiElurDFbjOPYhmoN0wARzxebqXF7/+f4D
WztMQPKr4SRb2RGevI1+wDxpyOabg3O0yeNQxkzURurV6UU2JBYHaDooku7EJ7Btz2jsZRQdq8LP
xi+YmzGE72wBSLGeB58CdKS42nlsDnbyUHF2Pxk305xHa+VJLvJ3XWJUdv/7/0IWj9sxOAyMfv/H
viDW5WuD/Uv9l9eMirtcCqBgDO+uOfVA+27Qnmk+JGKMIIRiiyQWQ7whugL1NNK1I+GKVRJCMLGP
Y6YnTiNZWqcwyzg4HRO3fErth677wLUcqitMyRSVMA5Akm6/VHrdAbdlN3tkypfM5ON5uDpjY5uf
9kkoGYjGg2d1laYsmubIRXMYuaWgCnBt4S014U6P93JmLlDEZu2VM+PK7SFVRm5AFaCrhg/jhAkA
yCIfz45zp5IDv11/WKW7mNf5JSTzwsX5/ZRIdBFZp2szHTZ/GRGBA2fzyooR+qdiANG4ruBnhxOR
ZSZ3UEXvm3VlzFBB4qvonwwCjCOZITRKzyUs9J+6XZBPrYzuPWbVX9h9b0Yfx6cyCGs1RLgxG3bN
lgyopx79OxSsuqspaCfreHDGjdyNGWYMDAJo+xRz+DH098lMwZZEBdT57+RnSk+82rogke64mtLA
48afWAbJ9xbZhlQSvb3h8Um/eiwl9TmrlcvIdRjHUJDsvh4hQEO9IuQJi8sEbDwdQRWMogqfrU2S
Fyzc9WdiXl3c1pv9S44YfvS1m/HUVzpCUh+LyCPBliD09mAQ6hTFcE3jlGDy4FLDGlrDcdiuUSt6
LHDN9N1wiH6g9gluHRVaEgmsUxwFjoTpUghKu8LgQ1c1bX1G/OgBmoqHShOMD1dI3c3UFugdJhqs
EpotXGYWtPaDvXYxVfcs2YjzEjkhq06QDUZ8aT5n79gtR1TI/u5ZuAKuWzEAjCFE75/lYp5yodT8
DvWwylgCWsxPUfJ9xkVm90o2P5vB1i91PIYIQPh8VrI9IRDHqtJLV1nqisoXBfcnb46EnluCe6yM
FcYT9+u4dTo5JSZLIAogJGTA+4CaTrUOto9Xgv20gnvleYvJ99EyivkP+q6C8gQ7ZsPaGbuzlDXf
p8FvWXQ4BxE+TTkgRRCcMAbn3a5QXdNhoVMrB0CAxPFj92jkNCMsXkYgR9RKXeNRyQvEpB+t9PJl
Ri2gFP1iJPwUmbydaitpJYDqy2CeE6cVeCey7gOuTBtQ6vc6UDF8DIn9LZN6QCoxOBHHrWMfVBdJ
VBRpsmbEXWgKEvR7yg8iFccKOr7BOrcpY9T+wIgYHKuZW9L5tX9q8uWewmCxX8jy3ShqXiKnzR2l
s0iuwHYeL/53TWYDY4fc1GbF/SqS3vdR7rnPYvP7D6TUNGBbtcfJ26bV1Z8cl1jtVjza84LWdSUa
/xiL2wFuPpl4y+yATi3TMZIaQhFL7N6kblBwqg7HHWxhayraZdpHnOPJNcBSzrGBaOCPawtGjEhD
nP7H70Jx84fuf5EVMqPXrosfnD0jR1nppl546tsWbZnLiiYyTt3Tdwk+7IlTIGYkN4MNGYFIxN2O
MouMdNGLZb/z2aKeyrD3AOU7B9KLzAIeqJ3gwl120xr0IJIVYA7PFNDPjnfcz+5G+m2+SSWsFLLy
TOsptXbIE4vYZAJNtq1D+7o7tFEl1++9bdxQzk7q+5zG17NSOUv1EE86koRUJItLP6X0GPeHN01A
vquuOlKMAM8diRhLENrvxlJDWdtuvzSa+xjDsiObKm43aImIdGBxE3JEUfLfAklHkZpYej7Xzj7w
1dhq1EUhNHgLv6Y/SE7aJ0YbFH7JGL71ROikcmdrLYCndhd6KD+zq4uIf4iqkJmykNKA2a7hF865
6czCRBIN1AWe+Ue7Ck1Vwr6EG5/iwOvhfOP43y7FW3/WZWWdoH9bpcjFmmc3hdQO6oWZBLaupJuX
4sSX2vkGzKRRrVhiPGcVzwNXDto8tGWVfTPi8ROg3J9xLpZwXNJH1zwEASBAZYlE8sgd6MW/NoOW
oAx9kTsNRBWfruLj3sR2uIS9VXn+bdQmIs/KRuZMthmuAR5HkTK0446jVNUmEwqIhxCnPyY/owm+
nCHC+PCK/iMNUld8d/tSfBKQjFLUC1fI4raefj9wPGaBJtYt6aKSIN7ucAGzgCTCuvY4A/HbIhHX
UShYYG0k/lvj1IDCtYSUI2qCdDhTAFVSlBjIQ8re2wnuCrC02o0dWmCFQQYzeMfm+bHPpbJj05QW
TjrIC9/3t4guJfyoOg8uzU2JnIOcT5Wpsu9ha4umYgZ6YcUibAUjGW/94yhu+DVjKFPE5FFK0K6f
vPnG7a1BRYyYhdpjXfPUWsPrIxkMvzjZpYikba9DmtU+d6f0wGamkUtneZ/uhE27addNbgOefF0G
OgRzN/klQobZeItm7wQS2SYw32/VhIk8IqFbp4tvu6cUsyTDzvMujcIQSj1p/9ScoKRaZqBC+JJO
W2GcGtVFIlAu/i6YJQ0Xvz7jZ0e28aH2Fm4H14bLmPAmmX7PAK0NXJcLHG18MPG/Z6MS6wNRbxMG
Mkb8PuihG8lRcdwiMUBsNTpfpwTLn/Bwvk4tOs0DyZ2dOTOBORBx0fyWYxK0518l/zkYSRq/E2T+
WW24FaQVCg+MOsnvarr6JW29RCaMogShuei04InarZdyLnovAEXe1mgQfz7Z8whc/gxxFFILrgpd
i1EXV8E1wXrI2unYIRVe7kC4NvZ2z/ATUdZUGgQ6/P0b7izGGwISjriXHsPl6NSHAbBE0+YiAt5Q
Om404QjMv+d/izzcY86ivhdLarWEorM8RmFDSiNfqnqIjfL+kpCqPeNSOEOh850lmHYaW8A8T13T
1VXdAIxGiIF9X5Aire3yqyduYDzqL4s0oG4DvZqEYcu+Sz9M7abiuLNJe8Mk89qBpikJdx7yYEDi
zcWUej2J/9Nhsc2nA4yJ8vKG7yBuBTaVbeEstadXfUjncMh21si/PguUNXYvxfPKL+CWfeFaAn+3
AqT5YVexfo0e/EDQmh6x4EREhnuV9Ty6hm7DFXKDS61k8tOE71nQLihKrqQNLp+K8/S9K48Elbix
K3tH60JuXy5ur+bejWWzZh5zfuXV+YYyWbd/BT9f66iCBUMnPYpTE5J26sRusrdHG36WzD6Em7uf
yB+2UnJyOwHv5CLqzgxqRSYMvrKRak4txPyCujTazGeHbtJTnZSelHGHSQCO3Gpox4rwRNyznzhG
7AccjfT5J4kqPaTLXDYKwB8Dd+D6iDltw5xfMQ/Co+gxvhQ+XMMshfmD4s9LTCnhVIciRZuXh9Sn
1IUfEwDOPYL1dwY7jbfRT1k7iUjIC9i06ALKzqqwwTG6OS4b0MkF+kvxW8A7y8LvlhISapZ1MtaT
M1KwOAJ8JeHqZfV6B/yIbjrq5ORseJ14sVm4ZmBrHjgt+DnrSRbMLdmWqi49VKCHwmLb/EGqZ2Pt
wDUJPLEqy6Nry8oPMvXDjBiZWqpl3U7q5g1rrYmMI+U4exOF3TiAovZueJb3dtADz1xkwvMFu/Jb
swz5csodZ7eeo52UuIbf5gDooiiKv3nN52qpEPdS3ttSIf3yXuFRKSSi9aPHTms2Ir8W5ZerkNDD
geFVUocAryl5mT6kwmoIs2UtCoFVwZLPB88hjRqRelB3dsRjyy4N/rffyTfDpQcjkDbGZ/eSiT0t
DD6bVdoyyFUCIsEfiSxDyzV5A5aRVjeXv3KEPX8DrKzQ1YPCfhgaxztTTSRcdb2B7wrpA4bmok5n
t7Pgi0ajbcE3cleGag3NnPYA62lRhfV1Zc8RQkCSUsUGGAvXJKi1JJRe5pSUaZEfthzTNgkK12EE
Y/ruu8VYPW1nOh4HR1XodwBOajQIdq9+36JaieEdUBzGQpwP+x1heLoDJ/jT5C1BjRAhnxBPOKxN
HwRQpovOq6niIa+dFrdUzld6u7kmU7t6KOXKqr9tdHYBMA8lPfCseRROvHZNesZ5GHx/x7cFbB1B
eLH29S20N2zj6oJPdA8W5E42swe9K3ulbpfy8L8CGHM9wNBEZ3BbgCbf8LLp3L8DAR0iPZSP77HA
aKidX7eY4g97DHdiPCox+a5Rr2ttrN1/BAPUS5Wyh500BzPpSOMyJi8kkximVvJ0CALL1tBR8IBo
i0OsC/S81F1UBG0Dn6air8ZqA9MDGonawisNwV/+XT9p2K6Wvx3axzZkHeACvucwWAXJYBaFlTvO
/8IzDJlg2Gf7G3OBuE6JQnJbdhtyE47LzVUGD3IC3/AqOY9um42OdeJjqs+A9rdP6wXNVyPoncbN
5ol30p61i/KgGrJsZYmh0qcOpp+Koy4CNWRP1vV6s58FylcOxQ6/fjny5V3kTAqvFv6I+RJ48VsZ
wca33zxp80XTIpsxMRHJ4l3SqwMWapImM9aD0QlcRu9EDJEXqpOwuGQC03J/TAFmYx/yijuZCJ9t
ACSjmQxAqJX8t4oPphrJmG8Ck7q37WP/GglkD4r6wclycNrtwl74RB60iYadZ0kAEZIc+1Ovml4F
Fu3UT/0/DLlkx5ayEFASp+O2Rv2xvf6dIiM+XllyvHsJ/sL+xDlFuAK+tz/Zc6jSAZlDEAZ2FfOG
G3sfwSNM8CYBLHsLYKMCw0V8o5dejuF/QyYAk20JQOVgD477wS6FuosE7yyaMVVZQpmX95IOXhYe
i4N4ab+WVARqIbbzrVPw81UEmCGeGrvl1MnWcEslSH3Ti2mt/WiIw4M2yxqmfvwodXxWqTdanbAV
pOOmBTU0MoqG+DOY+YU/4tLzFP6aX584geDeBi0xTrbmSIBxXflsSqJdSST9I0uqufnWqeOmFRvi
REChwDnWYcZ9QEfVwMpOhV/pp4ojb3laM/otAXhxorKJlOdzf7s4pUiw2q2PtGe/2QK8fIA9BOjX
Oa9Ix/aJLsCGwNK0r2yWPLYCjJxUEQJ9g/wXXFFwsoFaFoH3NH8ncsi3PIvVY2MHOXf68CA/nP5s
kpixeeycY1zlfumtHRH/4dgKPjK97tpVep4Glorocx7Z8fKC2yicg0L8WicOPokL13WfKO26UAfC
J2IsmO6LD6yOFnnn7EbaQivkjx3YZMpSxdGeR4seLbo/pXcK7Myb5AZ8BcCM/iJprY5vKoPaPktO
vD4qxqnT2ZdEW2N+5zHvUjgmBcWA7a9ttSesdp/JVSdJ+OYB0FnoP5IQVDOhHSVT8KHS5nYPR+cM
3GTrOnJYXVcEyKdOiFEdqJwM2ogY08HCuz5nk7VKy615Pij2Q7IU91alI7GHleJCIm18SGZ5YCth
tQG54npGoBwLMHOsAvS3xE5yAuPBCtCyxV6k9JdKhSOHzxMBPYYXsm6nZn2T6P4Wj5o3S5vtxHVF
CfBonGdJ3VpL22FnDllxVKfN7/82SxU9ziRUdxJGJUHbr6qfeMhc3Sc6fpSt46VzW6u9FF5Y5lo1
Jq/CjGfCt5ctMAWwWqjkoaiPplvcdaRICksazKmNtq66D5tdRia7dq93sGH/kAImAuiVouNd8V2R
i4RBDESOpzXZmaeaG4Gh94dSpXPRRfqXibq1wfXJkisBjLaRO71M6sjkBHmIX9iYCnvhJjjjRCXL
tE20dBf1vlETvyzRrukQArxvDDi3GkOuie0pR4zmV/5jxf5Vgzc0OeaaSg7n9vj72qRVY+3Ixlto
rJTPfeB33IHIrqvRaOS+SMEucGX6o3x7lpK+Q2p2rPbTZeeORaSIricnpppCAf7f84VhMRMpIAD2
BFqLZlbjRJVkHhuL6fSTVkurz7xfQcG3ivq5unTWXhXGhYiLYeVybcwFAUiqRTDknQ7YvZHPsST0
zKhTbMjyhTRAawsS4IYvwdZrQDUM+iZu6PC3rijgJI4nk2FJnJOVIJOVOR5eX9zBkqCfG/vO8v8e
0/BaqzUZstZhRJJWKRVRxFwfTdkPLzRt/+VhFafu7crDJOhkY9cV7sgZORSvek4W6PnCv6DZg/SG
hYJOjkfgzc8XB7bU+SOMBbiZaoHOfjf2JNqMJ/SQqh9NH5iU0lAEfwB2tTM2ni351eclz1wjurqz
/bC8yDRYS/nJ0shqSjT0CecBXCjI7KPptkgCWJXuspyrZ4YVb3/L5VhculLUkx5DON5IBA7KO8tC
HrtzJm+2JxJhkT4zEvMMYjvqBt9/k6/mlAbRZF0kW3QOnZdb8uFtI+dG3mDHzhvL+nbM7OKgr/U9
MQ8TXH4X4hnLADfyBk5r83AF89cvJMJhzyFypwBiunxYyZRu5jb8TiyF+0q6UoW6N7GBhacXMGqb
NUnwkno3lF8uZLlKJBYfg3IE0dALtFz3Y9wNRwbh61cuyCoisx+q8hmFFhJgzpL78evBDmiR2VrE
UPph682G3PcqNiHuqJa88M/t40jH3+Q3F+T2QQnCcJXJT3XdFZC2S6V+M+pwdktI3xuSjVujs2ZR
sS57mtD2hjKnz6COJ5mvuNszJNEznPTepBOTeREtMx6J2od/AJeNCDiKvEIsheZoVdidIRncxl9V
4IXf1Y2NpPHb+3W0Ytr+hb7elNW2xvl4LdQecnoQaUUALJQQo0VsnjNZuIhZaA4//KryXFJDo6r7
uUvce0FD2O1TEJv3SYtwZbngoFW0uNbZgI5nkie4H9dtIYsjJRxG3jXtMeZFdWffExrUgdsU1CJr
3Y5m2GEgBPwmNbSWdjNaSkkzaCohgLAcohY65w2XWkSr9q9qJBZS9u4MZYiNogc8MgpZaSrMDopL
8r6BH0m+Ib3tqQyhVDKfEZ6eCFI/+wsMynLUvTSp3eyBu8XcDg1Wuh38E23GGCD5ySpVbXAnb4KH
V1MHl56IzJENwmS5KHEo7tyn3TOsyzKe41hBvNjqt12tf76QeIq3iXmM/o5yZCJvJiVjSmh+qhpE
D+YV0eqUthhBs3RSic7Ym0cVosahZTbG9a4XyHHTyZEa//9O455XlPfysaSQrGTnvG6MYtsHryK9
ZBQbWRNwc5Gnb6EY0F3KNk4HB3drCkjPIH3eG22tXA4YD0EPZwpo7aVby+a8Kqou/2m8eDdpgagE
Co2Fe1PwF5JJfXYai+BlmiBi2jY/1gITAnRoahgVXC6o7XmFbYLIeiZfjzBwABDZJn+at45wRMUk
06PhIV3PyXTf/W3HCiMfCbBRjak8G07iao64WmXH3PHfb8r/+RAWdBPD+672irpgIay0Sv4F6dsy
2H/EKhwxsb3+hFuXcwoHs/JAm2QYFz7+xB+sGKa9T5CoFH5fMvygUw1+/DrkmOisOsSfw3+jZBhH
WCDF38HODryGr5zkoy8ceaQCD9GHM8dWynChT8He2D0ElvkT7b0Iuk7iU2QF7RoaRZRm/KUDQwlg
3sDUgjrE2+hNWHDz99NI+Zil68b9EMcXV9YBYLOAmojzrdCnsQtlqiUPNu+c3WsO2E9fYvKAQ0Wm
z8acgxqQnCe8md3SmBUWDSht/YGJDO9l4FLWAoU5+uSVP0dnYSX6agXeMAYQa0y6T9Uh0pf5Y7iV
l5JSIx6DWpUGjC5qxRAJTUFgfE5MxOmjcpCssoh6c23Vuovy/OVF99qnFJOR9LWxcjcSf2BWk0+C
dhQDoEzvnS1IzD37ZuySlhZlGoI3GuG4kVssTNv+mW6oZLVnhE+TTsGiebyWbXfll/ZYQm2VVfPC
Vll8lBL9A4ZrJt+1He7RCQOAmrdDuKzXvUq/hUDEqmlqdSY6HkwUIBk+hiszamwCMX948kZfDKpS
GKhEizXQ/qy0K14lxT6aFp9DIaPIPhUO+1I3JIYOJYmcFq41EG3lPaFcVCMa4RmcR77Pee56kf4w
fD6BIy33+6Sc6XyjT+1XYJh/qKkv0B0El6WoQrzcAOjMEvE7p17rOb0uS5X4NCZHJXsL0NjefU8+
sKokGKzeONL4jmLPnXLImP/P4vgY5cE/BelTUrYHdQhhQfs4LplpICz66nZsHhwnspr7zSX9IWwm
f2+JI+P518HEGOFbsn6Li8sQ1Sye3Ikmp2VHFAH0SSPfzOvF+QrZAvMI0AC0ZFsMlFz2KF+JiFym
rn8lpb3/o93jwAqeCGSrXpciHp+S9g/eenVdn3I08cYTRRvIfs03pivI4vH0eJUiwkfMwwxpbj3S
2ZT3i+9Z34JZaAa4vk66gdLEckw3rlpS7PTb1mPqn3MD8XVNDmRpk1db4YcU12ATvZeSJnrPJcnX
6GDOXzvNmZNMgbFJBNeH5lIdyiQbCz6LccSKpWQH5HruDIluiUh85tgTiBKzWm7OUCWA51QYJ3PY
2haN9kvwKvpxaSwk2Ftzr1+MTLw+SrAJkRC1nzxQuL2rNAy+96Ckpte9ofOmjQVj+6DAsSCs+0nj
6gdy/gfA3Ck159b4diG39VI1dfa2nfUocvdkaTkROZPkE552ZcGeJAJvfIcizQo0axVUYuXjod99
rck09vjUatNJrvRcOmgnpMXTOrsMeNiNvkRvzggGnRMsv/aEk2MVpTzvd0vbtFv+fVY4ctL9T2lq
lTFy4zXVddUWOHkkQv5xq3YTisWTEarcWLsDPcexI5329MDXS5UhEeHQONpB3mRZaG7sAF4Zo33U
IR9PJdTtOXAgSWpaPjvLLmeswYVa9vx46oI66HRaqSu120vcyIsh4al0zcbYyy+rSZhn0Tz3xl33
GbJdPgfW9YuAcgj29drV3G4nBK88/Onj62M/kshrNkOBDRj/YtuTeq41i5tYYvzc1BKuQciFNl+4
bq9UWTzNvhXLDUARcpP1lvPW6jez4kEpmIS6mExgtN5/kga+yV7Rtdmf8Xlf+kpx9qDyrUhfn9J5
1caWRkgFVgs0eOzVZ76QO4WITxLaPF4J1a9MyHiQsNT8skfozN2UFkbqBwPcE+1jmrOOcNFNHFM4
Uqo2nAJMtMFWQV3bPmH/6NiRTisjvg3tvJ3fMBEjZSEwdyxkxhI7jKPNK03OAj5GxtP4E031Tfe8
ho0mGiEtoWSL9Tl/Wop4DNwF0WOG/VDdXciH6Ta35UqTiCBITclTvgfVla85urOzlWFGXMkNn2il
evmhz39cN2TjKHSWQu9b7Dt4MoUEaqEod9ckchxrkyvVob1siu7RP5Qui0Wp/TSv152gtXnZ9OdZ
AhfOLczYQvnuH+UkaVShPYax63DwTaSIS66AcF6VRmhhDwbj5666G24P9XISmouh2r1l5b+i6T0N
UBLLh4ca+EoPOdt+6dHkaAYOUSodgH39hCSxX8uwuN06ShITnzpP2b+tiDww/ewmirNVzvwxEgu0
aMQQ3zd/cM5LhC1Z472p3Ak2ZrsRkxvAS1Dt3H7zI5y+Upi8TteFzORcXE3EBcVKmqkuI/6TuHFn
39rc2bIt0/E81+DSJVboZ8HZLCLB1uKFnqhzDZmKV68Bb9w56QM0OSKItZLxRfuxG+CBBj+Pm0uv
rgwgvVfqQqnXGQFijTI1Szgz4+f0cb51ZdGQhK+bwEuR3p/Wow0pYIUrFi/HTFhY6sBZTlrlaOES
wHUCGj+Gq5F+a12M7ccg/AwBnPRQugiAe9Sw7iKAmBG5Md7Gr+S/5MBfk1t5bfH8Rj9zUHcQh8Ju
eT5LGikWxL15jlqVaMCYw6pQItIHT7JM078k49zCDRtOLcsb1fOnpllV4xtoFlHkE8iz9CmJsPft
l7XSvzETZXJwzcYR0POu0tRKwoekms7NoqZIK6pXx9kPHjYwtIKxyDaR3ZFAqbxyFHAIjK/Uqvbg
Gq8+mHKz7BZY5jjRMBgCZL42tF7YZ2Kpuf4FbGxzWN/nESOXUxsGOxHAA5ArMJ7SC5pNHtcOUBw+
8RYhNdE7H/6SeuaqSVwwRMQ+5dVrM/WfWuUiXNCGa1ZaCPl3NX2KeYHLnkIOLtoe2uFN2FOgQ5jF
jPPAc43Fq7vJyFHZgDuonrIcteG8dwKxEI0mhAZi6N+FwPSLvwqpYViBObkvHYyvz6Fe0zsAXaPh
u/6pXfye1OmA6+MlB3wPvK1U4LDaKKXAR7GmymBNSwtEWcticvAGpsnhCTnsFEsBWPIHYpfqr97C
d0gHs/VxzxDSuaGuQg3xdZbSJdlxxcS97cwAY/Oj8G1I59ZFkv9g/i8Nu9Ql6b2iWYKIqd0hoZxX
Hieb+TF7gfzSGrY8e2f4xH6FcvYV329uYmNRpaqjB5BMxbVGhnhNoZ7xmz9PizgJdUo9MbvlsNY3
Sj28nan67J7uu3dxKAgBbI8DKhWQHVahnjZ5JpYwPjSLkeyYBg43EHXVP+zc/q2WX+SBIAFcLQuz
8IqgPmbv+9TQaceB+9NVITOSgYUF22MIGrScuAojrtNXf5t/UeuuRJd45IurcC+EwuAr4MA8qs1h
rMMkiCHQsCXd7TaRziTFso9NIrJb1AraMQj2pePrHM6t81EHtF99uAWqwR/G0VmLJmb8nQDJ60nZ
DPWcQV+Luo7D9fSVddlWYtATdoTamVuezfofTL4/xYmne9wvD88d8mA9O/EXo69/cM6bPWU2O2Pb
BzecwkqzuXW5MzaaMG+164m/JxKV53MP+LeY8KF0Qjpg4rX2MjW6GwlKSbFIeW6xx3EOCRhPSPGp
LWEI3loP8c3ZH1TXX16R5+HePp1AYeyzh9TXSQPgh6+0tRucY0r14PgCTrCJhx8UAO1cjw+zNzYc
N2WGZbiRJTm3ESYu/j+iMLWgRzD6nEPn23ezNsk0eHcVPA8EvpD34u//oJn2op98F8u6lId7mDu2
Ciio2BuN3cRbalmNzyo9lgztXzr5J5pEY4JSI2xf5Xgh/mbBrohaMymYhi1BNP0EnLTPkdpxGmeh
Up66VHSurhKCdevthhtXZedJfdhfTDJXWc/sxqcHFRLrDcDPNUZzLDjdLGAX/AwUTo4fB8NAMNpS
xV9tqkmI/Ktf85A7+XszgXhPIaoMS5X1zVE8PC49vlPDbAPR8EGHHzDeQAKOn60OXUkz1lwJaMgl
UCAS5c+pDTcwtSe3QpObR+2c+hjWChm/zWxLnzzQ2+cZB+dFz/4jLubWdF8hwF4y2WMR6q7mRMJ0
GEaH9EWijn8ZLKRR4PdOqKBkA1W4JbGW5EJSmDPS1F0+O01KYHSSyBJ6j4TlT3h10L8rS2TlXp+V
g0PJ8YiGIeY8GZ6vPQomr+rq0AJHtiyFxH+EQsWBMei471YcbHRCC0R5opHclma6Iui/S9bAZsJ0
Jrlv5JkdC4dL1QF744ZtZXwPszrm2B7zLgMKZHIkesV4zTRCPC/AtfSjclUpsny1w57kmIbW8ZS7
HhRtLa+92qf/eoHb1JwHgQBoJC8K3cDFj3BnO1kPnY29hPE6sVyzvaurhb9zEBVXbxQuc7y97NR5
YbLnAQfbD/Hb26eeruUQ0VpLcmFHiaYJugFlf2cgFMAlJu/SjYA3PO/QgS/nHzROhP29DHuYK5ID
xXnH9KzZjB4mxH5j/LeNCeK9MYFJmHt/BezMv/12ZzSDsZtZz8yACl8Km0s/Wu6aMXslkamGoV2m
9vByiask5hiRSCUCUEcC6WkkoM3To8Yfv2xyh/B3E5Xq2lCVtDNheTgDn904M3ICX1nVGncQFZAT
dgLUswoyPtSQXeBBaTg5vVlR0nEPwCnifJUUpVzP2ReYlBEKRr2lgLEMZn/0u6BUcQt1sTEKBRHE
g7rLCsLM7KGdwHlJEo9TaTG5Y2pc5Y1/2w1oM87STl6NMJTuTue71KZtHzlVQV752LzGeVz/mjnH
AIubU1IVAPtCEuVWz0cZ6kXXZgd5xQYelgUVh+AZJFhKlNunEhwWQqKACg78snr6V3fa4Sl14R+C
vFR31y7SshJW4hQzDragbQdZGOEHgpzZbpHEvczZBXYHgPTXiaKBMEdiIAmn08Ox59LF9xT4wFJb
TdFETTbzMaiPM9tpt10iApEFpCYN4sawbvJpd2e+yqw8x0iRyriHrTxdFuBg5zzUJmWYNqo+YGxg
YV6TYho7OltbQAW1A7/3d5yr1lbPiB1MHpRchwnjWLligBETBwrS1532jRmH2xf5iARVR46xWvD1
oHZHLULPZ11mEH5OdHsOXIM1RXfRZsgbIKo8QJedRYjjQaQOlGl9RCFreArrEe23tkVDHqJTe5j+
MxUK91wX6goCJcHDQL4D3LuZAkYrZDog+KUkXE9baMtJHYGMjioTWw0p27reCbWkmucGXZ5ToJAt
E5Gx41CqRaq4pgOJ64G/2t6IxqlQzYTf5dXOKoG6JnUsDvPpTiCBDFTQFRmILPVp/kVDcSSXejZM
ymMxIqtWvZjpwEekcdfRIFArJNbDhpSXAxyopY7U+wxtxr1cml7Uwq5JJBHHoeucAUEPKQjWenlG
4NYVKk++4NONJ3MEiNYtpvIrkuRTaEvdy73NizH9+Tm5sSbKUvoFq0vA9WN+MwHZGP1DVgfoKdeg
9a0/mThr6K56CNPULI/BXZ5D2qutEL6tD5cEJZrtrD7VFO5G66yt7eOcDSlLRvTy/dz7XRprwwTD
h4eajrM4nWQWpqlRbZQ4I4VzJ4qfGlEwhw/6LgqrG+Nq3bBwybq4NQzcNO0xxJfQ1Wv0ADM5KeoV
Ji5CloWJCtcwT6RSxMRQQrpmOklysYcnUeanWDp4g2jUDnBc9ClR3VvsAaLZmgVDbw80JRSDCGHr
fDUBy0NdXZ9ieXVKwt/UGuIR1XI3QZlZ/Gf9NhfY8IWKW8PibAmee9n9SCmM/mUwTBCBrKaz0Czt
3E+rFQTxBZdV8Gb0HWu8Uy0PUj5nXPDsYLZl5NRXG6CrjLcPkXpzrgP+4FedasEiIIox//B33qo8
aeW4ZsS+mSSo48t60Rt8toxQWIFAHTqGKMKcCRHa2Uqvyri5mQQWTwf0z6SiNoiLcZPYfVFXccta
oYuGKZV4tU7nICTC6d/CGBVminNpvUxBkVe3CgzuloY5X0V5n3lxgVyqhZSOOA5p4R8eWlCkE49n
xY+ulsjOboACcMxAyQf+O8/az42nU0GBmxsnDT08Lz3CeQfCaOp3wlyrQafOJ6wr/9lFr0/TXeTs
D6ctHkiXa+BpskvA1UBidpJ3w0UAC9A1Lj4tMFB15WMqrNb13P2onKx0utSlNuTXx7oKgqeWHqD6
HCInHoW9WgGlfrN169N7MXgimMk9s3cImfwUzjJ8JY5JdwjMmbc+OjNjgmwtfRfVt3MWdirjbjbE
qNNU/GL/YBy1asdyYVTzSkQdVJcud1oaTdLNRc1RZyjG9E+xS9Pdy5ivRtsfstkH3g/LcYhkXZTW
1cpg5UgPDWbXTymiTyZYrqPbV04W9e8TSLUBJJQ9zlRJMXvWzHqdda2ZzWpJquPvKh+gCVZdzRxH
jP5EidLITrrJFgskrfowQQshc8rmf1APMmiAc6PXxxH6tbwVdpI/VK59cfwerYCHj1YqugHZ+H8y
OVWZwsUweaplYRhRWjwJwgnP0Uah559z7DoBQSXuN18XZrj39hiVfjci0wnnRXzdpRU1pd1TmoID
nXPeGwedByrMFz5uflmKL0nabZ6OOF+pMnSG5KAdel7jjk7Ypg4P2uYstl0SKgFMcOa0MhoqjPzM
p09gtgysbz+AcLJQEPtyRgIjfpz8M0720duTMawqZPcRXC23MDjkcHbHOe71JKMCp/1NiyUjJezq
V1eGu+luwCi8BLLYOVq6o0ThClOUEq9BEH+YINkmgXzIiPo+bT1A7C5vOLgaeriirQw6jXLZ3d1t
Of/ofWdFsRCSH5gVAdJIwW7vfMzN+kbcNuM2MIkJGpXv2LkxcnCf/WHGtYnxlZktHVaE/m0GnwMg
6riBPcenTH8R3feaFsrNZAVEIadx7+J0yCRw/qolrimQOCnHJbg+2mc795ytOf/dPC/9ZPg7Uzgx
D5N0G41ucHe6IAqr1xT1KwuE2UzovNJCiaGoF0d14YNMk6LSwMHnawZA2rhpdhzEjBxb9UqoCl7l
TnLduiWuFSnbx+0P3dkc5zyn4t/elhUy8d1AzMYjLjHlAm8dI1Gm4PdUJuqBW2rMFmYUxMSSnLVF
CKNAdNeS6uhRd1pfmbajoeg+P9BVMsjkSgEpof887OVYT1JxYKz01qMYvn+C10G0g1+kVbqhILIH
yw8/oOz925zJho4QE0EJu0nDRIi3H8CgxC8boyO2SpT3b8VSac3yIeqqCAIHEqT7bXj27LgW+s6S
scCt9CU1MZHRjHZqpjSNbsvZIequgO1kHxl1PlO/It42LUIf8QJ3fbBmSFy0521b5ws0dCmeQ2mK
tL7bBebIGosuXOHRZdApywh4CWSgUhuZ/bJKpqd92A/UkqKtRCGHte1jdltg9KWY5kGvpXwd9VDd
GFujHXbkyPBU5HOnrgHDbqScZ8qURWpQKDq1EDVHTrucXVVN+Sc3zXdbASJIN6I7jfXGZmLR7b+r
HcUrIaRpQBEcU/UfMjb3Lqr80W4fSf5NOjdSLcGi74+7vz+hfFASmuRRzQy7zQwYFT2V2iTWW6Qz
s+3kQDK+5fLtA4rypxtbmz5Sq6Ro6R3A9w3O/2Uuz9PtlBgZSV1Ab14hLJxJIOcslKmNkD6ru/u0
82ZQ2GDsYra0YY+XOELjKDJmvmJ5x2Ey3ZqwwE4fMeh886LBbIhgnjmdtPgU3hB/XgF5+C4YM2wF
M2ftsVIVEsk/zn8qGZ2jjm/zzSdhw8OLPxslDyxLOdxKkYOSayshanJAMlnuOcPpZOLsYEIjbf21
6IUkPoG7P+qVH+mLHSlBDaEjIkVlj9pfaRJH/a20zOCxvZJ36nS7fQQoCFPzkiy5WmtCPrpqMGeM
P0HeSSSF6LWiydQxEUBmJ49Ac0FQj6uCw4oUQs8HehGFRQ/kG7QcFzbPgfH5UJmAbXDCPsFFjAlD
SZyNe8iIGneBiiHOemCti7lXXd06edhtIz7PIEaPor9webpkfWP6nBua21EQC0Uy+mUdjvOgHM5h
v/Hl0JE36WtKps8aQ77XQ1rGnhcOSTLZTpfE0NokyIdCDrAVWHv3nzE/MpxIFj4nNeRTVSUeZJ4o
cuauk3g3DtouxX9LAjk5UCnu0XhkwaX3oBXVVDfTF/imKgnyy8KaDR/z4eFIxaBLkysL5HBggJhN
xYsL9yvnQeN6ysiLsvSW5jQCLEDom6Seg/fZdEDtcSusNcxhJ/9TBZ6kqvPlH72vAroW4923baK3
VqCmTuWQ9FqJ2OiPIeItEVWmu9s+1OF9vBwE8BIfgwsp51kjMlI/ofots+ZeEu9oZpJq7mKAGRSU
WxO7cyjbKDU2HHUMCFgh6X22RxquziKE2sJZYiHC5dy/ABi2zHriXXn3QR9RqEgiGRd3c2PO+O/O
Ts7Lo58z3S3otPKbxgXAxPZDSHFThG+zfT663PP5T/uQJm1aRTWP8h3tOF1Emj9vV3uiL74fQtTv
ooTHLjKcXwh9gFc/wK2PptwyH2Lcz/qFq/R5h+B7jJu2Mh79KzIOTxQ+w0/GTmP8ZyaCDLJZPL1o
QJbON96WGoBi61/bF3DWYYh0WAsAKy1PQuvQ3w20I6lvtab9Yd6eQ+QL3wGWcadM2rKC1FB1sosU
UZ4PgOyQWMWjWC0l5Ls8e3PLQBb/Ti5l4Mv+Lk42EwQyNhtHdfOLjDH+KsYuOAVqpOA2YOaanq5v
MIfUyPuc4BGrU7lPJpbtrFhXeIvDogyaQibaL3WUTF+iKkvEP3jJbczL1cIbBkS921Q2sgC68fKc
vDam5V/a/vFymRXpohdso8ydFfpBRywE/dbrffsb2EEGIEEZMyt+7L/GZB09ZCaTV2JtvpuPD9Kp
tCc9KRaLfbwk9IkKmZs1ycGHbjoj7eEBJ3qDYDyXqujr8QTvEAo1RxNKhTlLD4a3JbBQS0aK1lx1
kxwLBYVY3qmKQF2Nii/oDIWePIRgAxEzxFrFdz0NcioDR+G+LHzUjWleoYKFWp1DtMWkn4QIee1Z
PNOpZAt5q8xhng9FYpATYz1ZwpKmMcmAg6WB8zn8uSLKMqu8E9aB4RiDSMfRPGG2Ti4hvMOXPyb1
rwQE8srPZFX+jZ4eNC5Ww+WldT8nee5fZZPJAMIljh2mUhFiRIyfA8LvSV+bJ/9dtfIj9T9QvdbW
NQPbbfWFMb/8oXnz/79q2TTefkJylmteE3wis345vJ5hAJ78/ZbqJislStH/naP4IAabC7peTQ9k
HopHnEzTUh2/aJKiLB65mW495BINSVksKxEVlu9OLzA5wSbKi+ZZ/H+ODOdXOX7q0grfAuH7GYOv
NdMY/PCbDnSaYya6WiJ9cUiyBuRdvChoQLXXnEp4g9VeaDlGtdNuYHzzXY/0E2q8Fn8fBIyATyOe
jYYcv/SbDGX4tivDW3XWoUyxt3sRo3j0zA8aYzg2ImWhj/lWGRPfIPKHZgooBglgvnI698YFjlbl
08IM0TEodWJJNB8JAJIGOi6yVyqmh0eTwiABOs+kMYU5H4YiJqHB9auyq5NkcMqKLEBozcguTYOX
+reEypb6e61vhH96/h5DJVvf1bwHcTmyqHoIaEUMp4Bm8KDd7lh2cANoM4d86gI4y3XmQGQa9Fnt
BKla84clXnosKYTwcK35vhMDh+o7qQ48TmYLUoTnazqY1YgAOazPU7SQuvMzID66aa1OtlrDVBjg
Q5gJftfD5ZbclyW2E61YLd/TLa/ocmt7k3lKHYir5JeH7Z1AukKnfoKT7Jr77lEqur8YegGGbPxH
0+J2hNSdPcD/dMGShSjlI5d+zSkW/2+TisTRGH1JjKDfBnV0Dj3NNaLevtpeued4j1fZDPUohxXC
91Qt84wlUZomi+OOzHKg1AI8e9bAxpPVCjEaFxreZ8dPTcE1tjpjS7MeYwp/7s2sBXrJxjmGXW01
K69O6b+11LjgSHR1YWJcphxPewNvR0W+UCX2cV82XcQwo4ysG9mVRrNEXtj7UKRuBHWFtfIZUI+Q
u5xgUmM8ny3m/qXAlerWnKunuNlRCzv2fzD9EazHRgoT71mkIdZrllqhktMrgQgevFIgfoTeTNFg
OUc82t0GfX98WCpNnBj8ug7lGQgDGfKEHkQGHm1ViaLJIA3TLQ9H3YtYsWmE+peqRYjmPN6yEGy0
YZz151ixRZGfetfwexkP8C4k6WMEq1Z6HfBdVy6hDVrHkGQQhAkRrMEe2T+BtwDnhTGJz7Xhgdof
J+B5LX6FtMysgK6y11dHB33Byt+5WiL0aX+Ylggj1m0Lw8iWePuoZS7d2UhO+HXrBaKfGR+W5VYn
KGJZaRnCUdE/Xsn5sN2ClwwIy8Mz4Qcm5CsUcVdLOqeO+2IUnSFpILh7bVhXa7ecDPIW95jfrdVS
YiR6OP2t0UKMq7CnqLspYNZEGkMZ7gi9RFRw0u0/zwekU9aoVCGX47LlWVi44UiJ0xp1/C6Kjpmh
k7u8LvnyZv3yIo5jodG0vd021f+bjEOeNTg+Xl/l6pSZiaslebDsEPrgDNnLw6WcV24fABMAiW52
GdZbwjy5OPyuONdl/2d4+CFq5vp4QR6KI1gywqTmxuruKmUCCrRk0UUW1If3zwo9YInem+gxO1Cp
ITB2vS32WxDI1WsCgRLqdD3ALSjWFJLaoflcAQN8ArLsDc7pl7fkzn1vJ36E6l9+HsoJOEjcOEAi
PfUDagGO7wQ1vhbcGbbHntTAWn30auqELnrLCEmVFxG+K+pfTkgROnmEmfar+qIhPtvGVgPX1MOE
TaA4bWmAqjWl0QUrtUurFPITHdE1CUhdIe/OwX81rdU7nEyMFux0NitKlOc9AT/9LfwA5yhSRgNm
pM8/FZG7MutadwAwlJCkNky+FAJAraBgYPk7umPXDji8i5eaPuDBTbFWzICpGTrfzJcv/RDuMCA7
CddS8epxhLeX9AImNwfYwLT6ozfR7DXsy209psfeFQnJVPip5+vbCQQpsfZbKuhfyaSlmhk2Ie5g
xQYZ9hjrxzARx0RmPTXB/cCLjssUUUS6glDZTIWMagfU8ThoQu6garVhXAydoqyJC3eI4r1TnlOm
nUHUsqOALdttG+wrcdxx/jif4jRl6MifmvsXy3yY1a7X6WB6r18J/0h345FpWBP5u1PfVp/7P1Hd
a3pnXqszlT2DZBpfcS23QdPH7ZkCEszaV7XBfsk51pVXPg5+0ZGmFrpsLbm7Xa84k++oDNWAu4aq
Tg94Nt4eRZ50DET+qIoGQpMmBuum9syVDenzcRQes5Yne3pWA6ZVCXDoZC5RYh3ZAS6vSr85tr2p
DjTyWPjHWTVk7bHnNV46TaQeG8liUky7UAtbcYQ/oBiLJARsv5xqBoJ+vtdpv8SReuOvryXkM/uH
nrhr21/osw6OB2inJRv0RYNi68z2jk2m/Ok76US6QsiZRbR9koUKPbRykSH7zpux1K1n/MJXuzlo
fM8AY7VOUvP2zr6i5fBKOY5HDZdQCPmj5U0mqV45jRwgUJAfX841tH4bqQOZme/ATL34bRJx+36a
I/78GkRf0V6wUfuU/XbOjOp23q4VijGIK7vgv3ebJBv+glQ8smtoFhF4o17L9davqYKxC/cXUz9c
RdyyVM458hG8n+gV4xyH+acijZ/JI1bEHqinmZx62PJ3oOrvRVhPpjPJuTS1F0rh7FkGw14Xc2p9
wrqe98cBCJVAmTgrTrcM+6UpcAEHPwrENA1+NGxjA196BPO8IBP72G2vjQA3+LGQLhM+Zw4UtEAU
5HqPsHYgMrdRg1/jTGCY7w+Dx+0TE95e8hsBKzqwNx9FnscumlWvqhpf6aFNJaWjkgIdmaWU7J5O
vDYw7VvLzzQ+on0IWLPbKLoGPU1Rgr6+mnYIXd2fGNvxd68JxNsWUQ7ujtCDOl97N5SohZxXA69K
auXLg5g3Oh5MPx9RuvmftEehJHBnDUYCMEetP9FkZR1g9LebgfO9TY1kqdMMWczo3EQfLxerOafk
mu6ipmFX94viG9gDivw8vmHbNpb2zeIHBWWI6x+BCVfXtMP3iuGH9dzADOgBTeZi9YxoxnoQgjNp
G2ExX3L7GaBQzOlGcb9SsSFvO8owBdA8iW93mf/Dg+jV/f17BSpGsuPt1WXDwA/TBj8type8TSGy
dTH4MQuEodd6UAvMFTCtvJgAVpFKCaDzkSHtuY1oHtBsknfPWmmONqsfRJKyBK12JmzPzmrU5Oyl
chA+Ft5YOy5V3DV1NCCQ5m3fyuNnDEkciaQAJ3bvuNL//efEPAJpvayFVPYYYRci+rxeQxNAZAqY
nESoCQ045wAWNgHTMeWFWOAm7/ejCgvYf66gpK3ms4Vo5mOPrLUlLi/o7kPqFmkQ7j8lF9a8h2Qh
goGt/iEodmgIc+OYOUv0VE6MZ7W7E4AWJKtjOtf/6N05MmUwY8bzk2NafpGttF3JmmoYH3egZ7EW
VKOBJndc6/9W5hGvfL/KA4My0Nqfv56Itl69AWOe1hH2xvV7TdCZrJVQXzEc3Y1Mf09KMQKFHFUH
jPzLQU2MBIDrgsjvMrvqpgZnu9PsvNelIt9nDsPKYrJTSYGipHlqq0GOhYguXFeNj4mdUwRkFeWl
CYIDnrF8MR8jL9XniFHeaza0F8rqN63w+bQodhbT+o7Ek+l9r4dljI3LkT4xZNDLE2z0cwEYtWqG
O5fQmMbLLPSP3HTLIvuLmiDTGCaGySGPsAi0V/oECVgIpQelmKzvYLB/dC9dDrgDVoeZXxZVVEv8
Xzw55u3kJHGB/GxyRQ8FoErSR7iTX6vi7IrxpDDCrakZUYgFIKw+222kVZTMsI5Frgtw5japy6yO
lhRX9DoXIInrjA+gSMeyYv6ahaudAPHSHXydp7dRAFcYAlR2un4Q3TSR6EcGBXA8anyiJSoqIzEr
f+B6DdTtRPFiW+WK1nSPOUfd9pJNC9gEB4SLRmsXRhHfi3aQF1th2lS4xcFiAvxGGfNXQjohAIhs
9Z0cQZGPZx/EXr/ydkeBqRj9NJL7jF2Oa2NmIRgbaaT9GqZDvm+Gqv3KjUsz//LPLpDXrleo0mSQ
R2WG3gfHEYfKfaJ0THdKSVWVXm4dpbdoYLBNW9zHc3vwECpNXYIc9csbOmv75BDfyG3Fg8O35Rln
LyB6XAlg5PlddVwWlHT0KZtR0KrCHivZO19O0dQORTmKcBKhnlnQL9Pm8Z+oPrce8iaY00/59gE/
1y96rv82mFIkTaxEdqk+klMG6KeLqfN1yhK+SRwtgn1N7K2xQvTl47s1EHm0oPuSp1PGw7sT+nR7
v6qZq1nlQFK9GLa+USu2+NINta+40WXy3VqwjNScSjrdT/RxsoQMlg8TC2EdFiMEwuXhCYvYItTT
uX45DDsx4i545NmJET+M71eWN1KS4rpPqcBBl0IPTveEQmAZW/GEQiHud3+WB0On4OYjtL54BYuP
58LfG2Cp2Ini5xEgzwZcgnTD+Vj7iWLtvZwYFHvwOjQ23SpkYB8YtXw00B6cAhTVAYY+YglCSFoW
YyJP99waUEFwvzixJX4Au9m+GPPV167B8wyJ4vshdYjk8vTUCHsGk8QnYhFqjbpAt9Y7JJSSvqF2
Ky+IbaCK7UcKyagShQuayqv2DgbjiHuFiqMs+f25v49aQOZhvepbZnl2siIsCMUEvLvBC+kdPJSu
jgn+3FPlrhktAWbcrqmH6wHy/yVWS+w2j7Jo3J6+UlwLycx3CvoPwDISZwqZBbRlKSdod+ohGbbe
SKS7xIzxDbn7KHbf55ncWaoVJBvgO981/InBDl9uVRsOJVE2kIJ+0JMWkuhRWcyCfErytk9wj+hr
RHzUb1DsWiwYspdyjHQZ+nyeHcfQejnP2AVLeIL+BYqvRJzfZxVIveQr9wCRvq7Z9eE3O43Bl3gt
/SC9rgSYb/39pLAiUVNb2K7C1tS5ZG/KTf4eppavKGPk8o1wo96QGUWr3caJS9bpoFtCvagtW6yY
ww5mkRr1U0PMxiRPqj/8PJZyQQLCpq6yEem3NisGFEy+DIiLkGTeTUcBn4KMEuXhHepf2rkEGMdy
b2Uhe6LgLoOmA1jJ08cuPIe1uqqQWaJg10podWeqxG3QAWU4T89RiuSXTV2MKvnTGLtQOgI//1fU
zt+cNalWtJNDMUbjcp9z88MuG03JrFRNDvoaDL87BGYgNhiFACf0HvlSob35S1Wq6jn4+y20Itlu
SFQCCj8RhELjmyb5e0xXeQ/XNGyVqldRYjN4ksvGMX2VKpv1i0eSRcGmmyhe3pV1f8LGD0W/zknf
UCx9dGDJKls8llRuMBO6pxcYy6TnRJpXKt9wqzE6K7qsyfFqbAPTVemEZE2HyZxB3Peyv3quOLQQ
G6RVP8hYmCbd2vzwKCN3LQRMbGJKvZiTSDOAY7v/fwoJhMqHQJCqK08wRhAILJPG7nLSW2m28Af+
sYmGeuDHNBVsOpPVPVFjrKt09O6726+hTAJCDlZ/8xiv+U8eHcYY/c9gB9Gl7CEzXs69Qhl8Qrwv
ACmjKXxUZBcwwmVdjGd6u7jctewW18fVIpTkRvhTa8ne2pqktbquCH33640RQ5SZopldYoh3f5BS
3FQkCrXwUWhoIT168cs+jO14xX8MtlVRawlILfsE9u7VsqmhHTAhb7dk3BskonhDc1Y8dqFjzXTz
eV/1t4V1EjpND+duyt9pBGmwtQU3eY1qDbKrhG60CtdcQf24dSkqhwXB71ElPOrA02asssAjwB6l
QEa8+osZ56tHPXtYhxy8tGo1LeJ0K91AtRv5CjHq1ZhcVkMNvAsw+3y+gW3OTXn54HMOPeN4ZH7f
IvOrCe7Sy80ubE0kXy7/96voDVEWBuXMv7szWvIUS7VPkvjdwobtOPCKEhCnnABKJRJnQsTv2F1A
kUyaktcRatyPL+kosDF4Gyk6rhPh37pDXwa1/7AatMHCRbKWGNiJ5hIAwdlFdtB02XitRY3xIasZ
bP/X5vzr0x/O2VV6xBPUICodzjwGZ4OscPWN0Kd3ab79hpxHTGjahN0IXtuw8tDkpu4QWzPNN6lZ
Kb0eP+aASxP8NsvHFUNJFm0cWHiRPcOCGrgZ1KLrqHoREuqIK64hUwD4LhTkI0flqMMxWgvsxY2p
2IEAzORCJoEUNeZ1u4Qa5HFad8SE2LZZuwsBbr/nNNfSky9YpdAr/reTXvmIi7KT8vLZwq7N0dTZ
PvtSh0g+O8ED41xHbHKaPWAIevpUee7lScpZ5lm9YrTkgTxeZWIiFMNUC1kHHwrOMEf7RCao/Vkj
Wcq8jCRrAouuUFS6WInuHBxn2DqiHldCnAG9ZOHK4RQGYY3mH+M/Yqleoo+LkyL5CbnL3Dkzx0tG
7qw/jYG7Z3UEkTLXTac56B/VoficYkpPMieJwyFV/RD/jE3BRGN7l7UrlT6lg0De1lLKT2droBGG
e/8OHxLqEYtoItM/nHUZfW1BSGgl7g30ixfYvMCwHxOAy522S3tswIoL6yC0QiwHm2ytz5oWuPbO
6OSDdy/HV5BBbS49mE4n7/rLvAE0ftVW3/cJKvs6korwu6qC6KZ/0saVGFeItx8+fJUJPLylAjLy
pCLtV0IMzAsf+In2d79rYi4DkkTySFOaol1ZajYM8O6oeoQp3Jd+swqWPMO67dnFwWN6eCKI1feu
pxFE/8al9j2c4AfmwXqbNl76uTMhOfUpyxZDAhZxRFQZhtBym5iSq+CZMScajIjQbkYTfhl1dIsd
BLAxbrFeZ2z4cPxbuwXWcZFTLqUVn1UUj8hyqHwMm1Z2a9aYAtHLKe48ESC+6wArCaexKMEPRUnU
FL9KTn65n5oNn2Ut+zW1U8ttN3/7//BlnmaVJUYUXkikPPpcjs4vdw7rBqaNgfxAmel1EsIFvWTd
SwIROR2zl2ERgQNukOdMnJSRghQ4ikbZ/cXlYYSNxOsZQLDUM4Vtvz6niG3RalUSKb1IgB18oS07
VttBFx2Hbmd8WQ2/E9z6s7XBwwOz8TaD+kMxccmYleenzXde9WLBSab9OisK5udl4Zv2ce0TPTMO
8ACLhjAsK5FQ7m9J+k7dJeY6l9SFlI95J/2VTc/NXydndcwljvTyAErrUXrNJnRyDYfyjX+DM9Oo
XpyCxQzgg9c8HNs4edxq52ovUKVa1vgDD9Xjk/U51O6X6b506Oekhedcab50mBnBj/8XvDKAlIR2
WryLwqPzkCOVo5USVzLtH7lE65uf9Q9uDbPFk4L14QMg6sQA63rgsTev20nKhaUIKd3t+lkNpjdd
cQtbzRFxb0wVp7i6Bqtv6H9erI20RhC1s89COz9zFWwZToME+RHGTuV+Hc6YX0ju5Uhw3n1V0dNK
S1yCF0bl06DEdtEiifVOsMCwyHnRrdGKJ7z49UONk+9m7Qa5fud7/rWpkpCHJLB48RZTYJzULr70
QbegXSlqGqMTj+lNwcn19NM6o298wjXHAVpuqiD6Pi2VPGIXM4QkDk/2vCLsXZgsRjx+MUulZadi
O6jAYi7eqSh+ZEfcjrGXb8ALD06BLRFjbNY7T8xUJrI0IjEAekFpcCx/qCqsOEp2uKyTbXV8PAqY
xwucJsoK6q9GJx9kzHEvGztD4VUFkxymrj9+KpDFhRc9j7pMLqpivhoBtuQPqXMLL1KN/tMPhySh
my6i+GoRMNE9e2eO/3GOUeWr3RCkIFv3OtX3NfEec0H7XDADeeNp4+lcCR/EcsMqLRUNdAN1inHa
laiR8XQ1e28YF0yKbTyjNt1XRYGymlifXyy3CFNgL5wDkmCL8+2SLpW+jL0fV8vuF8TbhcM1ZU95
E9ymkwF6G7aGW2jbqa0wJZ3s1ErBCuxKLtMmEXT8ZpzjGjS+GJtVm7kTlb8UcExeaIvUvJqJotvC
xSsLSwtFO5qP+oYVtPe38qn6W59Te0SEz5nSYrBud+Nwr3gHJYzQdaugsFEq69szw6igIowNkaed
AQefafo7m8gaJpM69d7mq6jL4ewSCipGulXrbhoz0bCWYzP+3dJAIGc8xTo9BmaQbRi4nR+7Joq/
es3Y75uCpG4no6h21AU+024O5jIRJDScCO2WNpaNDiNmkoEnSTrWMtuJkIn+rC9G5rH2wjtmXH4v
Z3F12OHPerenDjaE4eF+7tOcg2hXq4vSmZPhK1/56tn41lGA+/MXO/qc2WGe9sXRhVv2vZlly2jC
Jja4q94v7GH1bgPUpAJIKCCmXCdRiWh0ocfkD13WIY70EAXZ4QEkbtsCwX7CtDxQ+CGfKsXg/2X5
pPvT5L6ynmJ1sck73bn8Q5YTeXrg0l5QOQRtuuCL15kD/+2py2++QDLGPNYgDDCKVX8kp5bxo9YH
Sm6NllwmR0FHUUsGk6DKOVK1eyuKx93SvD47o5f/nFHYUNpmEcx+/8tpE1grfdPaZpKzjilf228A
/rxY2HyFdIJFo/b2sJqfbFHLvqwMHTrz48P75Jaodvw0SYOtbKBHj9EJbtRwGrsfHP9XJSDroRdd
ee461JlGDD+9sbxV6T7N7J3h4YSqWd14w3y5QUyuRbvS3j9tLhpKUl4c3aooEJ43Nl7julcFD8EI
a4a5QLQgXPayzLywrDOSYhNx3jbLdnKq+vTc4EVwfGZ105GszEUJ3XuBEpqa3NgNGK1hsapqsWMp
WdbQWylJQ7ghO5S0SXhPy8SkAzf/L6208mVfzgH+eFs9ETxLyrh3ohmADth9GMNUAFaYA79QiCV5
fjDGfqxfW7s/3FJj7adlZsY5eJMFL3IjbepfFq+UYl8rKkhHVwQx7Z0yY9RCZtfulLmxK6A8Ryyc
myYnshBDyRkesuswHPKfWyta5uJphh5nBF+tGTTjVSxadx9HlrjO4hG2IUy0MHDyR/FfafzPPJC5
qz8pbogU8Bc46guIlx/FBxgs0n2N3TozWlzXhdRA7cAGTn2KbRWZx+mFQtjd+fx3l3+yFchJODT8
YwesHcqoTBFLGON4z7M+6x7k2HFCxhW/2zObTy8WN+Zrp+PJHK0tMsCS5UNGCOzti1QB4HQ5KSj9
VI0AW6Fco9uA1LVjZZD7YOI/fTOZAsxUh51VXVwl4c8Erp1p2H33FpLaZVgFjjW8cYusqnma1zyB
jtKoIlXczZYIWQeF5zP8gUO61gxUFgYmNECjbiC+xnNThZAy6vXgM7h71sUbhZfRFCzulWQ8R26S
xxXBIrGv3WdZkNfB+PD/1rYTZPj54GrRptxg8wNHCVDFEgDwkfap4csJ9kW4OFOKi8S7MehsbNYV
WFdGI3UGV7v38U8/W9mYp3BV2qChz3cNLLE5bI4Js0n+0u0SIOzD+8Iuzvv5OYMx8u3z7RnQHpk/
wXJQLiSGS5HknqCMYV/jGrHheu0875APGFPUJAN2/dS0uoYwNujVolMPbSWk4lP5+yYb1cMV4DSE
LJu0Av2lfYQyrDpvkCmw11AeWPRPE8P/ZyRFozAyzAbcd4t0Aj4l7oHYOPwynMtgVMHHZWuy5Okj
U1sG2YL3g8xXbTVIE6MImcHRYG1Fkwb9Uh69r5YbJ2FYzIrdz8kAXoAnnZcA0HyMs3eIO26Q7X4l
IiJ4h67xESkOxGdZsqaB3nL6DwzAKrfLHYqmr/t7GlBBjB49UYJV7s9j7VKwc+dWlRzP/FPn4R4H
abvvtBCN2SPKAz0vTJYD3NmDQSn+mqoKSoLZvid884M2TzUZfffTchmB0GcZXf/95+1ovig+FaoM
2i9HwXtMdniaSkRmX3urv+UPMQvF8B05AQTACmcG4cCqtvtFKkvJNLMnkNJEdMixbqyWQgEsDuhW
DdSrQ9kP8I4WIdLYSw1GBQXGxCJLN5LpzMftb9xK0md3dtTSPczTadecVHyN2aOk2Mx0Iz+mykza
BqRVg0mnkxIQcFnkkpa48KHdWtAQbfip7hO/e/ZvIlahSrGbxZQ0mC2afPhGfRDM8PubJ2XoBOEs
q1dGIIPw0nHAd3Oy3mmqcWrqFUChJZ5hw/hbf0GPDZIEYYA50+PiGXS7h3rR/C4tf79ffm5NO2vA
cSSC+nZHLpcFNbZZuufJ5yZ/ehq2vKJVl4pOSDFbDCirBpLfB1+rf4/hvWPnlrcQ2BnXa7myWDFP
NLsS3qgLTTqFyHvFjZNPYDFuWzxoLSJgTFaMKoKg0SZ/GhvoPUUvLhYFwqM3eeDx8kuSv8IFOvtz
cSZxv7eQCd+5lc7DxECGllpfyU82pTnPZ8LjlxNkvEUeCHESkI1SqOTMCToWGuyVkFLXbGKBUUhw
OExil+YujXtxzsCvV1Sb2+YZ55ILTyOXApYowgXjLaTi1Xa0dN6uI6+1xtq6P1NPSrQwLMjdfgUc
pwbpy1Mi6drOiKBHOGbkqfYE6ShEqbkfUQcQelPZfKBw3C7aSaaKsABkQWTPciSk7Dc4FQZeP7z4
qLeBalrtzyTSiyob26a9K71QXexSiKvCJ9u43SgJMk5Zyau1TX1njNQ9IojiUnPI/am+2Tk7am5v
qbHMSK+tcoZwHgmsRHDROvW8rMhTWte7R2ngMLdQ/klIsi4EwiWR5VLe32AGN/lHwx334JEelb5l
RPkU7JwOznAj64P7k8unAwD4j2OE3QL1ZQL4bz1n0tHTBH3+pO4wJeJoheSdmD3h8+2CunQM75FK
HgW27kZnls4Gd2liXpc+wzso7IuAoQ9BgF7ibXUy0nsCDYWb7UOdbkuzGlSHcxiGjnOQPW/Hzj+N
LmvYo8dazpOlLCn4bDBF6kzggDDAWvZGEF2oDyi/VA/S8wI/DTGz/jsdbeJxomX8pM15M4ncbXqi
gZE2bkoBgI4WlpIyOwYdAEM8JIGkZiDFA4u+pHles0lNHaIh4nRJZfWtPT7D8vEzdf2IZ9xSoyqa
PTQC4TMfQgNRL7bvZrYZWEpKYT9xIRAGXERfyPrd/lvkkH4iK/m+V1fHIeYSPfwpdHAB53bLwQVC
mkCTFWpgLxaKcpOLjRURs202uA/fbDAL1YI93l0qrlo1ioodIiPFFqvsCfqHFUKH2az2wof9AFHr
gjuXArxjTNGm+dMyIAna4ElqyacdnO8HBRyav5esBhk19rqN1SB6DUPMUOOP3fbsUD0Ao4vkSB4n
lHBBdtoe9wzsAAGRMjv3RGRQqfR6a0HQGZ9o3pw/qaC/4qSKMTlpddRWTFepIMFyrxtSyeGYkuxq
Z/dZZxuFKaS37rL9legXVMFRTsW16QRqkk2ZoM+Cf1cMG9wed+gHogsYaL7CCk7fjaHJRn8YcXB0
nuNIsG3y2MtvXAUH1Zm59yWWE4LdqWMS9j6hIieMg6AqWdzeGUVUnIs91t2C5wI50QyhCNpsjzqK
DFiCZNPf/PIxscXZqTSnoZ+JpvNpb0tSQr+jBUgqj1/U6WHWq7mf+rKMBVDoepIUZb89JitMrujs
WhAApCvQEutWSGYp2ZKM119rrW0DZOXG60URxJM9fmXGglj7OHeA9q/KEAy+sCkiG9nNQeAdCn7A
3hKIKL47tHiiF0I1+QjExKzHJokbeBaCr2NWra7Tprlh6p123Q7IIvSzv6Q0kQ1V2BOaI6cJW0+2
cfqgI6WJPij2JBLKKY3iB7pnHKO2uOPfqEnQNd7ET6OnBFMWk6eSDhc63Gq2CX6Pk0j0IedEbr7B
QtdOdD7vX8Luny10Azb1GcG5QoIQAHQgg+2lzIAARFEARw3uycLSk4IPRkDNVhe+dzlVRPTmXOmw
Kz5sY74Fm5x2hZsGfKnWfGVP6wEHHRT0ipidkaXBkEJ6wJJoHWvFOCD38hZ3mjLWQXrMz1rt8PHb
5PInW6b64T/c0lo1mkRHN+A75N/qBph0BNDJWc+Hwsjwl4ydMQYRiPGjFTbu3fzSdm9/n2FxQLzd
iZDISgrI2UKdVrOV1WdSLMM6dSBQGp1KUNaT3riGRP4tvnK/iyE8vXpLQvjYPiGtj72p2kyiyHQU
fr7woZwHKWlMMF5kdA7qIAOUNA86uzy7UtzIalePF/lEw19OgJd+sTucwWAGHcb9rvIUUBqqi1OV
ycq0vOt+JkSwciMaX4aGpa5TaCHFmLnq3UMFoHlxUdrrcIi7DUJHo5c3Jek03LgkRIuLBdoJQzZy
TqEgJQpofspSFvf1r/akwTo4zqWxjntWvdGI/YMg8NQ/WZ+z4FGyl3BF/u5AV8Dsra7QOJtC0YwG
UMZzsG3b8boUXwOlLb2CQ7BoqiNVRG7XkdBAbQXsu48Ri3KYluCu5MmPU9yUVPrt9MCfuZt9Jl1D
azJMKT9XWow0ILi2MEYNa3G5qCC2RDS04jDEcSAxyL9s1KcOHu8KO34N5PQm2sT4kFqkRsUcWlT8
IGrxshmVflo67BJEmEkGy181i1oWwmHmM0Xj1O3tGmbMcvXT1xVaaBNCrfnrjWSPOLIrz2O0ySYy
/yqkF4D+CDpD+2KtvNP8pXF/cj6ZqoqM2yEMeCOpj5bhzhgG92t+aJflfJLOql6dtluPnZUIe1hr
RdDA5LcCmEA1GFMC66FOnfMNvU6U4r9Db4w6nQjtD8XL37PJUIbDn6MzYDb0+oD/ML6aaY2103dM
IWPYPcEa5RfgcizOqgNHLO/fHuCQDxwuy9emBG3WymBq5+QytHBRSnnTm+f31yGqn7VWzap8fO6g
yBCeQKSTV0WkrxALqskC6DZx6FWr3ooMd8pspjFIBjzCMdziPiaZML/GQZFT7gsqY2MnsJry/EBV
FkZgm2Q9UyHLw89rUOgZJteTZVnsMMB14FI6DybAGiPkEcq0XNx2ws/n6x3LmRSM/Y+3XjzIwzPC
pbe/7YGBeiuo0DB+4WQ9j7keYmomLsMlDbWMrUTZ7jYrrx+47NemD0GmFxrtm93xGuExDZFNYYPi
y6cTdOhdK+GNAWZud+Dy/czLE7B5x5pNP073K+flqK5VuU1mFt7Ro3LUuVJkCXwgw+I/1DVPlHqX
nCOOJdby0nFIW1WCWhIwyuA4a7R0MTyvmlJgxtxZgJtk9gKCKzFzJFvphYuWbSoXGDW6kuC9ylz4
b912AYpJb3ukjTeTA/Pb2mwMEB/poSU2IYkIEUBBWeHfU7FtXNbB4TmPGJxyKMKFsKa9wYOJo5Ls
87cQtafNJP+Zs+fZ6diAIFOTREqV6vB995nCFpksX/lqmIlYIDIJP88jtafLQ4VVJt9xCqG5aJaD
9KKetq5CpMYTiNboPjSWVCwxG4eeuxZXyVNGJYF8FBE5EybAQRB4ZYRTLIspNX/puWixPFLtQ+cP
RDYQ5HGiQbdVOft/h8KtOXb+u5b/Vc6guml8HLtoB7Y2QonoWW6RJPUYAfKXNjyW1LZJFK+v4dFi
gqKZRy4l+BdGOlEik41AwHDYJ6J/UXFV4CXyTmYs2X7Eqj8OY7lxDLStgJx/5ePFR8gg4mLEyuys
kdH5J7XsGbcfE8JG1FzJil01YJNLcwe+cfV5KeXW4XzImbKzgJdOaorY8nVwsSWEfxUUuq/wZmgg
+OhF/2jhnPmTJ3EIzuOvWrlznlsqN9GTG4T4ihGk0KhMa3tyEaDZ8db7ihqHDAwQR/i2bE3avOZs
GOH0kTIoA8W+CUJdt2ewi+65As8P/Tt/b3MYPeBAZBv8m8ypz0DQXY3rqrzYDw0Fn9oQ4WixMuHw
fHd6jitIQCs9mkf5WTYG4o6gDsysT7jJORyRv83g5tzJ/hnkbo/GuM5vj1mG5hiX+WdR76TMj5Po
eSgHGC41rDLDULvVZxZlUF3bIXL5zzKdU/VE1ud2uRxuxlgQadQyAcWyC5+nRO4yyZN5fc6P6X4r
My8mynzP5x7QZMfUqEnxrvlr2fCqZPrDuhm4Vco5Ict5uDm/NT6/8BpDPtRp4U1M81kK8zV5YBbI
TeRCCj05IGghpcogfk32IaeLE6XSy6a9bzea8BWZxVjt5kzfA319Lms2b/GF+0GDSWtp7HFUTts8
s/v9dXML7NUqp0hxlX2elsM21TvYMOJ5GGyv8rqWBRlWVO58JA/+kBDzLO63FDJAWU7N/wSA1Cn2
E4mZqu1eGB5Pd0uuygWX9hzs+9NAzFJVm3gpkiHChcMlic0by7+ghP1ocv5ZvCNqta+WvMowXoVU
Lz5kI0ie1PpEGrfMC/yFzvWJQzHChbOx4uCEJZaBZ7+RefZBzmNPFwxF65hMa7Z1OKniFYXyraxN
OgAJhGgcHERjdNJ0MXgBWUvKn8J/AB+dYiGOIo4949K6JsVcH67E3GNQDgYVrJvrhDPaKsZP/PBH
laq5styMrQcCoxIDBMnb6Zs+4eJSgbl7eXWVZSbOHv8+Z1RIZH1+N4u5pIPfxGYNUKaKYVtAPWsX
9gagXr6Xv/vBYs3TZKfv8n6KwqbqOmzowCcnbrkDM7kqCGvAfhVz1xV2jTfmA0Cr63OpFUyZRNRm
bwMYOjbXFtN6TitNuTpuahqgV8O/sn64TtqKTwvMwv3F5fF5O8vwEQF6EgWHxlUE3alXjtQ8YY5p
JqUf3lW2RLMaQjDEQILdaa2jMFVSOuDgziobDRRFoDx2xwlUpLZm+Ux5yETiMllOUcGer+l7Znzs
Kj48exuhyv3SnhSnLIrELpZOX86eofOgSJJZZ/TnjHsJJZ0cWcS7d/hLVvOpJ1gpOVLS8pj9Yhsz
ExOv+umjxg9pidwcqhQ7QvSvuESwc10SliCf6v87+H0ilm2cG2wSHTR0842jlzBfWxCqfuNA1mcF
Lhfl2X2IXPyI2vmRZUL2/2otyw2t+lrzpMBBK8yVYeIIZetBcog92osHvqyJWKUwmJnlajshdJhh
L4FlyMcwhKpEJGkdLRVXqhzJMWFdN+bnkgdI+fvlFz9eMd4OIlkl1LyFhPHvgCg1ehPGC+gKCjMU
FKDrFt7YTNrh/Zz593IzIibdQTQMz6azlnCGdio+t1vo2nCCWL7mb1JfK2VvD24hQ7jf+NNOhUlP
9U/z2Tv/vYIOmBwcbW6hnuuYOndGBZa5m0YNBXMWzyV67MtOaU6GSYXwQjA46it8UnteRUtZtLt4
iEHEBdoGG4k9uWFJKe5ezmIE0PjKuw511ZbKBQr4nG02cVLlgrKJ2tfLFZOVgujgqO9nwn4E0Xt5
CsHVN4eBOE+EgzjMjs83i/YWSTgISTrhfIMCq1mR8YVtQXTO93PiBPkKYGoq2UXrerfbkMCv7XRY
HIKyTBAAvyZ/FqmrDBp8e9yacXUJgf7KwKcPUVkQjt+F9cepdON78CA0Ks/tTCSSRoFBNPpco+gF
cz/2fW2T7+eaCxnYjenmEDSv1WhLHsN7FamqQmkgNxYYyXE99fjAyVaHP5uEDeMP1m4J3rEy9XQ9
/liAx6wsB4yXk5QrmFoCFZRtHozOQzWvHhGGUVBesJSfzgcAwtsf5JmvjfeVJKfBbfm/IV4BFl3J
2lLB5AmEZQWPqeemNECV6p6uiIqXvWjjwfSqwaX6FyBshhaLDplXEkNzuxxwrlN9aPz4piz8QKbk
W3JqWKKoI7a6YiTYkRvru9M5ickXwoD19DhNjIX+rFfiWBlno+rGwD0VIefXR142ov3GXL9Ya670
4MmaN4KsHmukOO4jE+MVOhA9VBmkuvw41VMW+uG5w9KmXh7UwtN7RGcAmDmXTlD4RmgDXBWySQRl
4oq+YvQw9lAmIUnFH3nGG4stqwbXMgG5BaDeeK1wQkVbdQ1IIp9WXHCkspsTFCJc3PflySZULlXK
K9kqz/N/96x5cFqjA0MOfZbl17PyB3kVvPd2S8HOJA8lnT+4C983z/J/6U/OVOUO8/ZFBh8MTzA2
ejm5gFTf685NqwNMe2dXgHZww1FPzTpx6yuF6BGxlMupJjVWMXdTNXUyjcq9B9mFAxWKDkiIZwjb
4PtuU/LRbAj0JA4QDY3bi1Ir8wimsmqOebxZfSuISHvbAgXUR5tqyenzVq6qX/NYeu+KLdfSTTzQ
FyO0tKy5XrWe2+LP9ndno/BaCd9ynN46orZxTSbbHmEa7VkE0d6hZ3wrUpwBgR1j6kyB6RFYTBPk
czY1pXRggY4l1NL91OlTcP1hfQEhf0CgTzMwTnnb6roCOEgJFoISn2ctR7/3pwdUpWLyFThsUz4k
DiB5O0pif0iXAR0tKKV3kTdNBv3CH5t4Tx4h0NX2PUTwZ7EV5Veow1gEj6n5nb+PFqoEA8x61PJ+
4V6UybO/as5kZe4GtMP53XY7X/dDPgwMlNaFloY+v0Bu6FKbB6xZbsvU5iJNnLaKe+BU3c9YjAGn
xvX68y2Y3wCYoYbjWCaBpEVPMMt1YKHnxTEc1YobSIUiVMP/SSn7UCl1BgKkZiFS6dRxUR/9SEoW
4T2woRCOPxFsqXwjYnkuq0U9lgPnsj7/0qxc4lJ73n5Jgo10tecCyoRWg8q2YKUntUIWH2Jmduay
q7A6bmbRIuxaCOGKelBE88D3+C02h4ogbwncZKswFikQHWr1J7BCxX1PqlGfN8yuX1S90S5prhMs
WQOVkHufiA5bKfDNLed+MdGXm2sq3dGSEqrOtLjQuG3b0BP3fGinKKZv4F4F/2XnS0WzohVCvQpQ
ctfi/R85mynclM/aQ6xTUHL1/eNRzl5nfikUfPEADiNvd/Q3LKjibwhMKQU14pevlXD8Zj4OkEyM
hdLkKP1s2qTtS9DUoiMTnegVcVKoZ0lPAP7sj5Yf17vEFjPsIDoFxSFIkQdQKwHsRo1AqUJSVHU2
8KeuPRoD9Wv3lsFlMAXrsoR4rVz1JR3GsUTRs119R39PqcLnWTQgwEVfgbLXWuEie8TNcVTXvrba
R0vyXLo7r4m9ZxVQIiFzkdycRWdzgPvTVo6vKZ9htl5KFP01qwKfj3Q41MVOu28+5jCRolZH7q6H
xqzQwU3XCKAj16qh4pb0bw4ZioL/kfRFkXvg0u7XjHTLjHKN2jO1+8IlrEAbYDpBZndcAq2xPn+4
WoSUt891NT9D9l6HZUj81snUBmRzIxlsv7yi5r7H5duH/fgXPOzIOsDgXUgX+obE6LO61npa0gfO
vbXeloH317HdyD7d11Zvxku/TjbhqC7Orvml2pZSE9MN474a5waX5o9zUTitj7nQykfbvW9vvE37
BSr/Ez76h1Z9BBaMGJG2NXvoIrTZhFp8J3zELQoV7crooQlVl37NrjfxJ/cL58fYg9VWWyEN2p2T
mPOegAoX6sjJPRd4T3pOGPBnauB+LHHKlvJ1ulDhnYPU5S7VvTncLS5cuMwFL9D2MJo923Zkpe43
K/Zkmc2NxVTaOWF7TmfDEJP0uHWaiM1b6emM4Abb0KNfl8qs33d7ZIl13TTMhKVKlcsbqFApABop
4azWhH3l4tmJQKDx8MoMTAwX3vUFbH//4N9YCy26ffL5pSj3o8Xu5+UW7PdtElOEO0tSBJo8Vg/3
NkeJoMo+BT5NKI2s8n5eAWuPQgr+cdx2XPSyFRLEkX+QgHkbICe7he1MJLp1aR6o1GAYc5YwTgM+
kuDzCQgRbNmRWk75afWw4KRxP0ohyutmbMzR/EuIR2hjoASXG51IDV5VXe4adhoFvac0J8OIor5A
iv5KfM+hQ+wifutiA3nbWGFEc4eNR4PUrGDKBgCRR3AG8+F39aV8pMFXdaDzO+uhlJtXPL+JJJNT
ZA8NWKT1rMEpwtMw2Ux3fEGvhJK2xBFtbe0u1erCEYvl08Uk5uMpb0oTDTp24WxhzXcFsu7PHrFW
FWwOUk/nBQ16OKdwUVP9wm4UGFMGtiUIm0JszDEHg9Y18JmSJsEcDl9mBdjmnt1Wuize4FCAlGmJ
CV5+EoWSP6fxjlNTkn5c2Rg0Z4tzPlznBz3Yifll6BedkwhnpSHf7S2Fe7L3LbnbWujbhZp+bgjO
Q33uLyMRaSeDyC+778uwkHLwzokewPdKKppf150Hjl2J7hswP1W9cTX2u3AQ+/+jb3f0ssEOb3yu
dWIrMVeGgMxltPbBXW8Dp7qXfKmIoCwGF/45//IxjVmUzLAW8uyLFOMga9HdAeIqH3W9fSm2ojwN
HxQFRmkdePS35FQTWeTMHhE9iZCVBezkXgZUpaKM0I5nC6aFGDPhtXRCQMEzyMhWX7xRRwb4K2Xs
drLHxy+RzqNuRSwpc8pywX1p35/DPJQdKH104um6l0sjPnB/jBqRTamUH0bssOFopO1WHTBRkwqU
Hg6+JgqOOp7pfYUJVoPN2wkBu38q9NMqPUFG6/8vzNDrw3q/w4KyHXbT3e0RGyX26z+eGlG0/u4p
Phva/2tivhLLlhzT8SxIXzoVbl+LgZaeIihQ8OOa7TaD9SVgyk/v8yHm6VELho5bcZMI4D2ap29B
tqKwg8J3PwuLn7XJCDcr68RU/bCsnH8nJsP1q32MYgoa2ggK/CqrYVJVvwo6Kq/yJh2CA/uqu1wT
org8Y9Pqf2KBlOg4AXZ1yIFj4c6dk1ggSdLFMPsyxRtgkLu0dKvqkDovnNgDFKfQyty4JxqtNmgE
nTj6IZxQJvhyLBUTAuqhBxxTcfkobhiFuasTHcpYARP9P5OfXImkB1oCDo7kLUrVDEGpUvrrXekY
3Qii5qS7hQxDjN4ixaitwVSXnmkydBrifT/WYsyll2Szaurh2rztwq9GTVD4nPBisJvSoVogIkkK
U2YhvN0nDkuvhfa04LaXFKd2RiWnH8rJnVPtEMhzyDfcvH7iemDcUJ8zhWI0/vQbmd6BfbY3w2Rx
p83L2kGlZITzmmAXaW2lfQ8rylewTDgdODOK2jYq4zTFb0CXB55lcU6OudkVV5Z2TPt02ir11rTs
lkvp3CxPt1s/l6Cl8C5ZalxxEqpumnAfT+3i7EhRNUuuqxccaEAaaZRgTezMKctNOxTGzkIIBXf/
yCNHZs0Zhkzu/r6J8SEusu8FZilW23Gg1DbMT0l3kpGrfEyBBzhhquKvwlk/qcirlI1K5sECLDFV
tTcvL0hSpBIP6d0JTmWSGNr/BIzZjChnR17fHUzI/gJHL5UH9HQrbPZqnv9YfrExE+wcSDBKSZM+
Vu39VMWy64COxDmzSdr82jpbW84azI+lyq4TBNguFZFvoSilTX2BEk9Cl9vvyG8fioPiXPiN5VFU
FX0WBO1w+UuYvZjPKsSt0sJ3QRPfSQ7MiiWMkk26ZuA4z+Nqw/e2Dg3oqYdRenQtPPg7MZ+tsGQs
gPeBQ/+p5jrYsZH4aWi1u/kfbq1+0+wJst/KxcJLlpbMibeakT+VzgCLyLZFz6iavVI4eRRHhF4d
o8YyTVg1cpmnwTZiw3vZe1yySrJuHThUv0mI+PdAMrdYTbPuI0Ch+/xbw/bSyGQdrspAeTm1UH2w
HJH7vYkEOTf6cck07v85YDbOwISToNCwte76OyT30lvivqWDbWglh4kbjhP9AZONrgJLKcO5IV9b
IE9UdocTIFhgWWTOhSmwT3LR1LBL8qWZ1ozBW4T/vU/A36ensIiCZkbFVKkDBgfTqveAVyEZ1Qhf
cYZMAc8TTrJ24hwvY+4OAelRJ6TS/h/OQbH7js9exi6iH14kzT0pgMtpowY+EymDGfyD8a9hUsre
ekVHFe7ZlUCz84mdddXEsKwSwhXFi/Vhfa8mvf8HpqoW1LNBiocigoHBLm7fgF3ldVrSu4Jcr/os
7hwf0ttmHYxBAd+8PbmYhEvqMd55E+G+czoLCKy/ag8wz7ElS/wJWo3KAkGuQbaa+JBQ9fQlMJeL
rqWGtkmUv4gcjX/9yLwCJR5Ys/m+7lkJrzCyuaWCQ1MDK+7iAfnAtmt5jtWRkbtxRaXjqiPBVdYU
ib7H9XX+N0WyWpa2U6bKdYCBaA9YwGiZTUIpP0u5i9Cp7a5yKtjI8UnTqWDe1GvBOzVgUAIFUMy6
o3cqvQr78zcj8OBL/fFvLweVeTrlpH64S3NnwRA0ZXfO8DWYDbCzMKdfubdk8C4J07rC1qVt3YNf
xZNIuV17iOgExMCNjRKuhSLq5bDdwwSqrLldN7PWh8cbiK+8H4d4aLeOiXosp7B2C6TyTQZiKlR7
v+QzBm07TxZkwN1+314BMXuiCBdM0UYAUVQU/9GiEqux9wvshWEwm6kjE4ZsJUIqA/9Fce3Hq8bG
/6pk8SnzJrfTnElUSp3SUYVdRkgsnazRa3mXKXEvoLlWNCfVa1KbytNrappu4HSZ0C3PfYoVEntq
ZbGiu7+iH0TjUfLfrubgOFb6XLDUocK9WP5f7m5Pk1ngoW/t18aMbWGFxCiXFkhRUqtXjaInDyZ/
WwvaOBlkWEzJXLR3KsxLSIQHZPQcmM0OXnUbyefiNd5eOXAWphV73IBX3hI53im23tkEF4Cj0HK8
MKnYFAqPxf7zV+BP0HMcCwIVjPIHAiMd5zRh9+vavwkInCO+kclqTn6QkV7xLpqfIvvnQd1nUXEN
uGtwYkMW8tT/N/I9oer12ZixFnZEyYznzJAAPuUsnPsHY7Hphp8VTrijRl8DzIQuxRR8bmWSAALW
N1OEG4ydzBcB+Of/YtZL3GxIh4C95b+KQRVkUqsqRHYr3LZuuyy+iI8QI6QsnLgH3ZO6zpq8k5Cq
w9B+GC5bYcqnKTfnckf5+pZCVt6v9VLMg+f8pWU4qQXRlqgJQIG2bKkbhcmfh5x7F8B5LRht7dwt
JVqeFnD/DWLKwdRsNvLBB0QrJ7kJCWQR9dZh5QNFKzy6hUPEEzhqGC32X7gvcW10YIVTXs0pLyEo
bFY5vZBAJgoPOZ+IJsHm6fY215dBpT8+nQ7DEZ9E1GLJ6Nt59YmdAhN7y4jp+JuTvrUZVmRBnaXQ
2doYgBQH4MgJNIEzJPgkV/3g7VoQVRIcIfvEjVZoy5Vsle8VAjbEYedLRbbCU2ljFXkr45En4eEX
lzneNOPFec/YJ/33uR/p1MNo4r/Nzw8GhKF2ukyzqqK3zQRVUgY5WQP1Vb4qfcmwQdqc7zliHmOk
Z7yEmqdBIfI0BJeiIhtSF6JQw59KojvO/9lcuei2Ur7RTukRVTy2/dfz+MYsQhVyp94pvt5lEspW
b+SDYo64UFw1uzZCsdK+DyjL5WsfwHec8PPDeU1a82XVSxKeTyO4qdtiWuDTj1qJdAM0uBfoBmkX
IZNHkP8OfyakhTos7IlT9od1lHrYEo9dw0IlqyprfTIlf6ZNzxAwDx+m2hWihBuJbeO7bZLi3MhE
+QTrzEc+buZpHzcsKo4sAIj5m7Gr9aUIv0HdAbxoUsCTKIDyoDaiKJG5LHmAj//PyHFcvnr5Vb5r
CR1vZj+UX4E+ispk/TWiASQZKJEyq0lczR03PR5wCOPGRJ7Q7q7mmBnjJhF41h6tYJL65jrnev88
rerbxUN99YQAOdGw5xPbvMAQswhpBhzjIPze5GCbX7RRT710Ug7wGI6dO3/wh2b9eghhZTsgDhef
hQdqHiMwiBG26bVm/Lam1rYG/17F+z6E35c39y+YK8kMuNitykJNjsjWVyg9s01HzsF8QoidFsu6
dhBOER1AFJydak+LSH89hjB+kb6m3fNzibZqxukOJLyNhbR5hwVpXXe9mnPu9J/D0ZpjR8tUCVR9
tAMdTGdPDyeisdEKSv65CP4CNW2N4MSdNm6w/W89kCT2tzcapnKg+j560/cmc+/1NrfFM0zywODc
R0avKxCigBgM507TYMm4PWjOjQvfESnrDUKedn4EHPpo1hIn6uZtl9mDeY7KmLgVis+8EPVzs5uQ
GnQ56c7eM1EPOgdIL6PPlFb2tCbXiy9pHG+d+Sek4IzFRFHg3x0x7jy40it3cucRGIEXOphNe/3v
HAM7VxeaBnFILSuX/mTcCSDukU4jX311VvHCNSaGDxyxCr+pZMWsNzuXtI5YPdAVrcwLrq5wTfyQ
nNuN4NaOYqLG+nXY+KWDY9MaxuPQAZKRQLrlq/UJElmohVDTHRVwigHndGeCckZdsuMfP3UDocL7
DprcWLh0yrYLIwvFH/wNblALUJ+G2/DKxTwvKFcVXH+/vGxRn7cmWvLKu7KutXiyNiaCaFrmNBcA
I6a4mGHV6gmOl0cYIwcUiACkqUqFCUhhsse5RTUHJGFyu+CzpU8EwKqQScbnJK9YI3tg6FD3f5dP
DGFkgiGhTYq1kuM+tT/Ag4BccsYzZvgaF9AE0atW5U+enFS33YX2JzetQGXnfzrBe7ckeTl43Vku
XqdN3HdJ4KL9Z9w2Ulf5wed4aFG7fNIWjfI3OZulBvHYBuQm+SNxKF252OU7SgX7bEqIy2wQM55Q
AJkejMxVp2hrK5B5J53isO3tDskpLM7hMAyMJFczub1Db0N+swk+hYk6o+60V/ctBlhUja4nNV2T
HP/Dg+vcnioROBeDS6IB0Cw+S9l/Yt8aFqG7uf6+cShEFpOj6VukfVC4+5vvFdGcIX5LzvOwvKbz
wueom7+ayXciMg/hgW4wdq1abT5AMLnidATQX/tzrYaOBT3wmUmOHeIZ397l+kOdh8JeGOmCem7P
QAnZU1w1YzuiGowfoq/SFMppZC3w+dXdxM5LAVdt766665vemukQXfMpfizwssOwc/hpATQ+6DKz
qNCJvTB7N3Yu2TutrPpo1mrLJtfCguv+Bg6AhSQsAWGMg0fLyg1jDOyBK6Nv7mFlskwkCNlRRipw
nNL1WwOGlJpOqLZya5C9MzURzq9rHPxAz4I+BOXZ4llbYm96UhXXyjgzIIVuHn4f432szTATimim
bUt7/QQFDqWSkcuC6dNK2WWN/QR6hPA0ONea15sC9Q7tQwiU1ZQh71vZd7AJUEBLkF8Sx3wA5osX
9k2XcVsccMzCzs2BbKVygJ/2e3iG+nUQonVf2sCc94GT0mX9VTEVO6OdfrOOMsyo6jXI3linUuO1
ksjbteZAa796XHp2RhGUpPAtugiuyxROYU8vncJD+pnZ0Xa5ydjYcKZrKYTmwiDfmkenTrznLK9e
HDMC5mG3ZWynIT1n/04jeDyXdiFMytwAH5HoUjunavNGMk80pi71vXZJ1pODL2iqKs7DNMPcaa+r
0dFR3vqFmHVl4yAxS3KoUodvk9lujrv9j7L1TS00WgAOYH0gogAFWBMfsQsCfZUqEb/FcMNkBmfa
VupP03XbuEb5QZB7A9YuQSSZbuHRbwaeLFpumWhB0W02AVBwpttw7mD85VRzOfBwwSlesUa0lh8Z
t3QIkcNIog7B4cG7iol3SVtEDrsIYPRPCH5j4ULkwPnHqambNxFzbNPekedkmWcbIHOhsh7Gt1UT
bRCyLZ+WPu1SKzun0QezXCkBfrR+vFCbIwpwPATdXqUCWe/WYBIngYYgfake8PzAK5cKHZarUrXk
UY24keIaK9YwIaF7FcpRAU08IF4vhVzTbcnpTm3Qm4rOVjytiMxk6Cfolpj/BtXUFyJLhmt7VdRy
/J4q1QaMHgr5dppNX8zx97GkU+QEoPOHArS9bz/Z2CQriAOgVCah0hQweZzRnzZucZWQkyQjMxT6
utXl3JHUlgI/VaWF5PaUIofCUf1TFW4MYWUxt4n0D2q1q5/lujTEGHVk9gBZ0Ut15eI2McP2spE9
KIou9IHARZ+84gWQy7E+LEwbaN/viJIZIcBfPgZD2euCbNqzH2HNHT1FVHCq+RbEezi2+db9ww/2
Z4vX2Te5kLKkZF5jw6BVEo43UCPkom4QoyEqFAGI0rtyl2VmTvPtbIMUXZpBQouVe89okR+WT59T
3Ok7dMUmy5Y76DGWAVsMKz5tdV5i83DxIV7Ulzn9I9hmJghlOVDY4gykJu6aT2d+csBJG2cVaFA5
aOZMCp6Ty7+4MspkOMxo33FcNXrhdAg8VWvlbXTKbhf3tdgkSdH6Y+FUBBoUeLUSTpQ3lNUbK+NJ
HPTJt9MpfpaHsc2FPdviZnEIgN6PI3dfuC4dbtGnPNB1zWiBj8VBZdel0QcjA4A2p5jZn94d19ld
cczWNTCv0yPS7Me8H7DAVkQAGVVVFHwMhuyZMVYT+654Md3I+lJKBIAuaHx5k6CwnsudfsUERw6b
9qy6yZfbmEgvh5HuUz9Y3AuVF29wsf2882rnrMc/IMWKXDjjnNtEGnrox5zmfpSYU2yx5Yst0i78
DN++1NM8WG6CU3VDPUdc2cJvkB1tdihzpOWHnNgbAHcW0OOnnvy8Usp2H4guuspvbKtWTbUY7oNL
gCFSQXEmeL1jL1P3sm+iK627OzW7DDO+hRvZMN1DRJoOZuBYLzzUPiTZ7soDmEAqHmK4H01SSSqT
Q8B2HAE1tMNqLYD1WVfogwnXmjnGOI7SOVGyg3mMMffUU5g7RAvyfYS9d7UVEjrvzJZdB+qlmiY1
Ii4nWHaQW1EQE7HZhrcQnLJGoTrdmYx06VYFZlVm+oiZJSEt77ILSdcX7yWipBPgly57JqvwKEkl
heo6rYie/GCSHgxaa/QPuAB+DDP9MNO1RPvL9rcrJR1fylzly1mfxZNwyvQqxvIMJBT3nkEP6XA5
2jdfZnVMJ53InZmIL4iSyYnvWhQrTjxy5Zk4W1jRrOuwV/lSxRAXPUiydCVmjCFSLQedk7YAlRdu
A3WJWZTGIcHNUKbX103+QPV8Wd8rgH2o6wuOgQ9HaEVhHcDE21rw3dLKZCwvkYaqrEXgJiISFW8M
a4/ZgqBlwUAhyUPTFuXRJxpwVGp60ZeQzAkzxngj+u7m756ICzYkrair2W+r/o1gN3ZhRyxZjUIu
H89KjSpM0iFVT82hFhkUQhpchH7htzUedwY6FGrvqAlVSpoXr2zugrLHNgU/riW00j5uB3JGVwJ3
GbauZSfrkGfoC5ErpMknOUG04ogRl3Xfccr5G8hO00vut5XIR6yzpY8SeEs7TsaS6FxHVucmO1fN
r2Em5JpATKyCnB1z5vMBj3G8Pjc4Ct+Bz4Ba47ihSWm547h92cw/s9xlGXMs6UfWaQm5229ujrA/
mdV1Tqk4NUmvjVbRh1g/13R0ubfIueZxzjZgXpq5bskxwc6DJ8OUxhzXeZCEK3IQ4nhaJmU6Z5id
Vpz6AZ0kcyWTf6fSdZJHgqDgBMinE050cr1X7UMgqxwaqnxUzFrzTI/3I69M0sKrx7tkVGi49n4W
OI/0cDybIuqAEQAb5pF24chfUXf03V1QkioO/cRTYs5rMbgcCz4Dmnze6GwuatvEg7XNCQhtPY4u
LArRaWKdRpuD/Tp/eayM+jgVOkJg3BimwfiXKsY34XoGK/CBwu09MCgfP8Anx+4y5v5R5g92oAKB
gMQRmZsaA1fy6TGsBZhhZmcjFpxWnlXWsCKHgF+vtcAQgXUSxIJZcRhtOGWBXgAJjqrIWmvEER8B
iYoMLzvvHYcqRGboSgN1m+dE5XD5L6F5WHUOg6NC3H5jjfaT7i7ScUzbG/DsTs/ygxdMk5/iMypP
mB25T3v04Nbw/He7N4bx8I/AScJPPkTHjcYu6PtGIrca/mzab+Yd+WwizaZSglXFKPB/who+TwjB
MgWL5yJeO3MKy2b79cfLocLlsxA5OnjbF6itXBPq01RsOpujGi0V/KIDSglQ3VVQ9MeMCE2ZG+Xj
P3hDft54LF4t77j11IvPTmz4zt2nAkrQugyWrjyLT+aMmGs/jBWo9GBPF8ZKw5FbD8+71onZquT4
421huz1zKl+SDYyyJqA8az/L82jPDroTqWK1m6bzwf07m/ddtwgnGbb/02QBQyVpJsNLNuBXdJQo
RNXU78TDJK0CP4v9C56SWYv0/hOcTrVghVfZokde7HKs0E8hfmALT9ZStz/D0sJ2p6Twq0l7Sr8c
hp1qbOn0mKhZbzW0CqIfxPdDMmq09qzTc6/ILEC0rJvPhZxeK9bfmtvWRHIuvvrGP1WV86zN8Qh0
qxdN+PeP4/dwMP6RjXsU0n/buaXqgx8i+5QZPDlsHqE5DLkuwfGxcYaK33uyFqk+4UMUroAKGCLT
9JGyI0DAjiJ4ICpPn4E6wCsXvb88CVB6z4nz7uK85bsJWcDpE/rztcNTkJdW9pguBZrv8Jqik4en
VrQfngNZiqnra6NVTyNcFHVfRQT+t26HXeVYxQFbT8WOS9kmH+rFVduC7VjAsd0OWurszYy5Az2M
BH1PeyCG5jWMRFmBrK6WpIhy5qozg+V05GLf9A89Tr8JtAlKmnlQQOS2R91XLq5tFluZFhqrHQYc
cpdSZnfmG48MSXD602xBi/SKJtiAXLH2McPNKhfae4V1pCnx7wmYniOZ6MuncEw+6PCHMFyVfx8p
+14r3EczYdYqmA6svUMAXMFdampV+N+KP2qtBl9PLZsAn2ST7ZIDg/ReYcyXVqmYLh1XuY9KDrQi
+pBT7Hsm2eSdeY+evhv8dQZ2udB/AI5LOBr3H133FduOX8GzKtHuL8ufvhQmTvVHzFuG74ADhKlX
JbO4tEukbTva5z4QYC5oX5/ikvIO89D6OLNS37F8mNJzg7Po5Iu+c7xHhGV4bd60YlnEuKTurf/i
CvpAPOQP3vNha/HbyxLwrZYb53mQdDkcxMDXUHqA5v4/TGGb8spfHTBO2QCIjRSHXFPGNudYaSsO
HmCKbCaKXMkuDOEV8g4BGANz5oyFjyV2+wMkCf9Ejn5A6O+ew6Ge2FzQzTV2Oj5rM1mM9VxS4lR8
0nKKezz/k+snaNxNlCEUT84NGkrKflObgzTeucUW1JTD3iu5GM9ee2zu+fGeTk2ZioO+yg/RdVa3
dXMPgHxn33QList0hHsc8XUsmP+uwgg0/g/omOox5u22tOVIamvNgctDcee+njM5F1u4E+G56jkD
2IbHxERsq3ZlUHGYVUaDxdH5ee8O19bRoVmRF8aYGNSJp4lF2tO66VjvfVUoaoyfNt4kwXsAOmct
1qlHC97iG8e+BLv/MqzflAmi3p0A+8Qq7kh3vjlwh466yIkTfNwLC3L2fIdtwPM1gJaiEywgwzX7
7A5+8AQRrpzH6owA5D+5gyRP5wlbrbPzVEwtP0nhd9RiMC1LpD/IOe7EtxG5pYIfMNmpP0J6bpZN
TjI4aEnqimMdQqJB93f1BzaSunKSKdLTDR4AHw0bo+WZcHqVJ33lfIzzS34pFlwds0goq5DTPN/T
GJeipL7AMnJ3M1/di5/Adev+/3BqXPhiJUgVM+UHCVtvhtAD0Ojmipc7gKNk+aTIvKB7SfXMNHwu
HQzxX+k6Ouq33XlgvqIBi12sDfSPakntrMLHSrg2txxZbkzNZWsCY/ukskDjrjSeBSQIrnA6+stn
I6pR1Gv/9LX6jDuS4QiSGwR7P28pFdk/TZVvTgBE0TCy7EwnTOVm+WHOhdRgIQwb/GTEyuCWzrDO
5PL/MzV86bVoyIui2HUHXvBDRa1ri9kOdu3NuslFGTguKo8/JIxx6hrW9ynaHmYooqFYOfU4lluD
SMiLFu9onrQbMLr9LvRCSbFaXsuX/iurMDyjUwS0T5YaACgaZhHvX/cchbJpqlHlnOB+HlAucbuC
26B77bspn3U2kISm5mPZRiPAVJYkjlYgRCzI3UAUBJTPYwHA9VF8KmE/yLAzbBhG6dDq5SwRbGqv
EKKMim7682l4BITBRdxomlBOZfWnXc/1vU2lqyc7zVixF7/N4ttwXP7kxVGNCNhREqeACdfX5oWT
hOegYxeAANokxtRvulrubgCfZFtkJCFJSpuvfliS2sMcp6MRY7nYcT8YAWvxW8iLNDBUd6Bxqk0j
2hXYCBWej/+lo047lWTFXiZA8JsmgUMtZ4nCSssIHXqb6po4LYJNIhGEMZ8IMTYGuUKIXWLwD6e3
5/Z/ieSMk5R5a+bGXfXAFFeuXICqoLkG2/PjSBQMoTOR2JT/S8di09oyYRCVWPLgAQI5/hs8fh+t
IyKF+022zIBfFhB0tz2Bib2BKAPPSoxRZgcPHufvIp8HG3mDp1AVO93JuevVZVINTCJSA0FvFY2J
1ZgmO72nd2OfFqTTHGEy7vImPFfzdQKPX229yKqVHDFnAKSiY7mEs8YNoQESfODSiX80WmUb5bii
vpnr654e8dwEp8f/zP74/wPb0c9Xh06qjHfeiGVMxqT0qhtoJNNdEs90SkChiqNz8GGDlTUgVkie
+gAEm5px3u6C4YZLSMjRYjShOGUyzXIN4HQFLG6+4rShjTAv+g6UUFSkUIqkK6dOtMT6Lx8J42jo
DcPmvyZGrU0CMm923Hf26kUDBmiQ25JTLvqvwIQkQAEdWKSO8OQE7Ys+k75lr1AfbCX97NOAsYRq
NAUHmbsXPimDEK+ZDSaL5kWikm99b7KF2CjbVorwD/gRkqZ+H/ip0f8foDN+JyUYRZ4tcy3z0xxT
fMHC3bD5jiSeZ2T4gOqIWBYJ8u0qLLYo8vvJVLYKnuhiXp2+WBIRm9kcnzME0uUiqgZy0d1jEZna
OrzeZ5E94+k1oARNgqgoxZz2xfGtPTM38LeYUUHsKtEkw51kEyO5Tqz1edP1O9RjHAKfrWgUUIbe
9oFhLfBeojXJkfpkZZ5fMjci/AwKkTZERN+0LhFpnIq/8SATdhndjeSeiSA1BfX/qmY6Mcj8dZqm
k+/ROsfbKaEJKNlaBP6B/GQOa/TSxt19vxywgu5qJIh8ZB9GP+ycLWgRfV53u26IKnaa7UVLPTfD
jyjNmjh3E3XCkz1Ow4xxyJKwfHeFRWj5EpVZkx13xuFUO6+e0y7QgtrL1VnSTD7BYJNsZFakZmNR
9Jirg0eZk5UN876KkGVOpMAwi/VOlDx61X57lxfJKFe+kPp8KUgf2++VRuLGd8ryTwxtl3bDyQ1M
H0qJAYf19O83tfNGLi/WZ8OcSercVGqRZy1xDlM1KtFTq+pNA81g63t5jMjoQtS5q7oGwGoZ5N5Q
4Lq4jPn5pXlwGu5YTsZZP5w6O7joHSwrsAuCPo8S/lWaDvrGDbIqzFNaV8FDsvdag55CzZQ6VkO+
hXXJOKNLN412TgDNQ80jJJH6TM7dZJIgbiYVMkxlv2qcqQhDpkCYr50vU7D3GKBvfRGaLlGx0dRX
ICf3PAOxTdnvfFRDa4vql+azx5EtAiU5kllYmNJQgaQtrX1mrjw3IZ8RtMRmCCqfzcFvjzBaetIS
FCTFdIGHQZqXHjFLS9fVVqsexl1pw15kOKg3lyENr2eROFvSdGOkZyBkiOOirArdDWiSWdIH0f1S
5asqS/Htfhkpf+fn7FrId3r5j/K3recrpggZ35UBcZKJbR5vNPffPy8OIw41yUDwRn3UjHpG/div
I9MlBvdJtTeBJsThpnXuptBtnIZVuglTTbHy+RSsDAFeXbXVoIkWUZJJF30gCGy7BBItka6fjOTk
NHXCmqGaMQc1uhQHba+CAOjqmkehxa4jMnOuQ3HTycyRsE4KqVFG6NWvPUGtnc550QR/6kh3Yhtb
C7Vys+XhLARFZZPsgv10O9RbAMfPl0dhSMQntAmZH+oS4DbDLZUaONW9VihWDQ+RdHaOLyN3hK0A
+wtav5yxVWaQhrJbLcuqgggLADteJX3UaOPfieHG21W/Mp/yL7hbl+xWeL+Lvn4JAvqL6zPxLYHP
seKi7CQxIZu4L2fB4dnVBE+w/PsrJ7KNLP/QyUkVVRnb1U5+fXDBbahev1eSiWo3wuQpsTWpIQ72
lWIaU3RewRk93vwX+WCHWxd8DMR/woxk33a5Rf1se9/KhwvDHCDOqH2PsGSNPwYE+gPZchQp9JyL
ctZNb5jJnQoTL5tV6pE2XCT9ERr69DZcNqFGE5PwyOOSC5QDEps3oOkVfFW3tFN36JY4s3MgcyGV
V0cpEEUpN/VuaadxhYMF73UEfG1Vs4cHGdFSNqZG4lRlPE5urvUYZ1bDsJ8xrczqIz7tMhtkOraU
jND27t3BfoFU0aq+1ho28806jDvT6duo+3ldLRoThyf5zox2G384nZr04zy1SKTa0ApzxBK4zYUZ
d665knKat1qbXARxinWcQ9wsmrcXoDNhAfOigngUXJiLZCA6lPScE9+tGfYsksDu73rCq2I+Y3Gq
aoeXK1A9p1/gxA1LA86blii39CS4XC+mBwRSSl7GcN9aZV1qmf2EjHogKuUglayC9ZMiOmxWrZx8
dl5AERAKhrWfY3qTGX+Kmsu4ekTSuB+N5px8kQQAoLDNkNtc63/QOTnXId8gW+dO0uimUFq+MX16
gIfPtlp0aqU6yET8CqRJU5JfF/jnqBnNoFJp7TrqmbBdEFH3bPY6+tKpTiq8L0aykwTWNcW1g+Bv
7MJ8IU81cNJIcOK1lbaKKoLXucStGbAs4454Zl0Yqsq6uBV8jyNl5KcbxOmDyUOip5U4lgKPUWi3
PZ7V9cSiSOMBNMzZosPb+hBMixuJHOnHrcDdjAF7wyga6RV+f41TVBcQ/SLp8X89FSBbzrrFqlve
4nrgzNoqayhMitsOozOMu4kW5tSKcfmZYZF5J8t1C5gENG2lveA84DUQ6xTjDvJBx9ZnxNi6t4UM
Q54hPQLUw3L7wyZHAxKl4oUr6jZ6sNkKuDoUhXTbC5zXSn9JS59EsZ4aTT7bEUDVEoRoQSmH3rcc
hDpEzV8R0LEZZNAc9BpWlCQhP0KJCjHFJdbOfYNegosCfCxxsn+uyOuiAhnQ+IK+xMdeCanWeUOd
44PnKN1+tHHOXFOLJiAJA/ki8RZhwIA5voncjM9Tm/H23HbCpD/nceyRY3VGiZvgMhXm57M84Cx6
Bk2aS5KuKeBgi6gwcDOHJR2XTarnGhZQ1Dm46srG29u8/3oTKb8vbQpuuNFbHwzZpLoOR9kBEll9
EeaqAhmGg7rC1+VPg/H2LcNHupOhaPlyMjcSTD90uL5j+PIHFc0nPXLVKynbf/RjsPyQSFpgl+Sq
485Lep23Jbew2Sk9ktJpUOKV81bgwFI6izPKWtMdig65TSuAZjBEl1xs5lJlDcUdGuQB2ZgfKZZD
n+MNA+PbrgxJX98Etje+VFaYgX/2pjwV98FQq+sFJ9Q/EO4PQjBvN2Rf/Xs58xS2scgQ3xirrtFn
+um93sRnsmEyKVERIvE4E1WCdLvxCgKxnufkxFq8dEzfrXRcDe16u+SC6Ve3aypnPWYjwoW8ZvxF
TfdscdE+TU9GsW6BtUk6J6LuxlE/EOpMDLgHYaf0UOQsUTxuhqkOG2Ww/NT69XrFQLLPS/4OAEKe
2dY08hKRPMMUNU9Z93ANO50pFB6GelZHLwWLzUf3Xc/Rz2B/xS6ZKrFdg61OIHZxfwkVx7ny4E2Y
mFQ7I+eTK6/13QJtmBIvVbWzNbJ3+43gc+86XE6uAK3mMTTzYi4MSOW7TS1bV7omuajmfSZkfjv1
5RNrRMIYvStbCSe72+POvaxOBu2FM01xweYFdZMJJowBm3NpwlJ4v9zQdfo1oe5wjEV4WxhFagfc
CQRD4+4HnfoDgHFNoBhuHG1YiuoN4pgdDuAOeqpTF0rt1YbMRXTMrNzJl9elgqenEz8N5ObbkoKW
FqcJvzwScZbs+T2cMVdfrf1iZ1sv/3tEj7TnzugAGOA8HZn+9qRxVdGM6oyA4FmiFBmB/Y7Q2FsA
Yv/tVH5SbzrgOZwK1kZRM1o2e3pis4tEWA2wsK2BS4LZ/nMqPMnxZN9rmckhHGaa8VVFC9+pOUuK
5EU2umpe6osfrtqJXLifO3Cww+wGiErP4apUpI484vSc4uLZLK9XSRC3FNKDT+KKb4BkIHqZ+j5j
Ib3NFJzZB0n+R8wQWDHr13n6vv5fAL6wkK+0uTPApl/uusLQweAeMmazwMBG375wFqW02zFxhvNW
ZjaepbuM3la3nP4kgpLiX7n5me1h0vlW6KGr94FVAAGraJBR/BLbT56VS9k+7MrQZPIovb2NCNjT
rOOiEfjy7X4CiexjDX+DYqy60wzXv3NwCaAV/t26/WOk4a2ojTB4maWsTULQjZUr0RFGAANaB6Lg
dHXhUQGX9qco2tMDO9NkIPMrgOEiSV0XuPaFAq3gWWoRzAldLfPwY6TY/hKXuz2Y6Liw0A+1u1PX
uSsuQJXS2ROFCxS1iBQ77tFZsiE2JmbEqe2Rc0EXlI6xOojoKaaKnWl0p9PfgxGRgOwcz+ZYSgQU
Bolt1tD/hGaAMMG8y7Oqj55CDIQQObrJyQyMdT6gyg7ZbvAd/7vu9p1SJi0IYn+rljWqopqiUOi8
5VKMiRR9nkATjOsEIsbe4sFuaGImcYE2KMBkCbcYcd97/weJgIFooALMMR28p84uHr5QZ2Cu7YIc
aigZ42UVQifWw70XQ8BEcWZaR9XJPYqDjbNQNN85ywLnbJqGnHBS009jXRlj2fEasvzX1Ns7BFSA
E7BHqnigrVToxDTZcZ68hgyl2ZMvwhqLoue/puSXMS21c0H7efh1nlEFXJ3sdn1FetEbNnQV0H7t
SJVRrqBcctAcMVBDXnXOXBH28q9CCTpl8FWZ+EgMMOo9c7eD2O7VmPYLowRlajAL2ndH4ZdhkRNc
Zj2vvBCd+PGo8YW/WXohUQeWautBvnGKBr/uvOvj/lvgnOh6j72UtdSOeTaMoeFWBeVwMDmkTGn+
JNC+PZk03RNY0+eECFYEuWLWZmuL6XtoUN7shf2sPUeuiWk9h+axbEZmca0+h2ynTd01ncWJrsJ7
o/BcmCUQqUUX99wPjJDt5eRyZZimAN7tq1Ulx1yke7Jb9aaLEOf1xds36p+L1gSHj/yroO6ECUF8
lUNPk+OusHoy4IOpo1Tc3NEHWYgx7viAQOrIPvW3q717WtkFeONG1e9ykJ5jz60xGodOs4EXh1ut
CzXpuzWm1tkrCfzTddf64ua3tcUiB7a217ZlJ2IimlZLnExmoCn56O56eJ8XO2lpOvjOSTVxxT3v
Jus/E41qd3sR6bTOtjYZEqXyQDMqgvl5oBn9VCZmbDoFJMUQ0zgnrKX3E6XOBQt4vYt1WFUWOHXh
REe2BTVSf4qTP1OrDDUF78kVrKiu6ajOydzUJhbkIT70k+jB21oz1T1i7FRTUbXyzeSgp+zdjDAr
6jGUZyS3MJoUPQ/hLd14xOCmmjea/4JrpCVZHG2dSlVzYL1QPD9iC2Vb81ppryq/lmNepO9aLRoy
8Rw+ppxBqP0YI1dOXGLKkNVjYBw6iV6XFV036q1gDOCnyk9K8vYA9CvAipW+JDuUzjfGW7DnjjGr
qnE9fuBxB0vVHhgIlITMiIYZJuKAvFF+430FXMxupYI9zkt0vLOxNqP56VInI0xHpE0akQIMioZT
IJaM5i0/kAIjtfgZD2xg9V5oroxvHDtUdPJOVCVzN9XB77x75RrsGBTz313JgkjiYRhxoKPJGZwr
S7T5hA66082D7mLT10YE+px2p0wCgUJ9g4lBFQSLvLUDpDYhXzS8q/jQ+g/VNCSl2HoQsa5cYJxH
6pSPnlyD1zEWM7IyMe+NqidPb7auCRAjaPa0PYvRL6qnm++7NrEAUsGESJXxQqDwm4eOYG5ebCiU
vHnbmQUHfF7wm21xnPSiJFuJICS5DTWTpjMQUH/nfd3QYIercmpTnzaggDUPeLbSYIfoz/zeBGCa
ykoEa5MeBegLMFhqUs42vLShf6YKSdb6Es29xU+AsSswVFdu7Fv0tSVJOYFpccigGVGZO7KwxhU3
x+cvO+u0SJRMqWShWM6bhUZR19DX7I0d1d+B+m0owKOg73hfQUyqK9/xhL86XrTuZdQTGPp1Tgye
jn3qCXD7BXHdplIEqhhSWsMdFLM9YAj3AoAi95MBLP9gQqCKxtVLpGjTi/x+tFsRl8mlA0ZvfpYq
LM6grCfJKfcqrsho8/L0hPeVT3W0umGUIg0S8KRIY6tQuVd2ZsRhDiH1fK3NLGPQHRhmc6N/dlff
uLGsQwCgt0RJEmYkbfO2R5tPREkEzfKTCgY2Ghj6SLN3ESbMvGpYPn5tqmdgJN4v/e9MGMJu8YgY
6x6sE3X4VJJNEqjB4JBEFVINrRuTWZ/Vz+uknWCZpWjWvLygqhmyhTvTcCaiWiieDcfXavZN+hYd
PXmhOn/8iduAMl1TpumZFqNwDHXlcDWKgAc4HIraZS48PNdKMm79GoZuJLMiZshrYcki0jAleCdK
Y246/zAHN3Cbc+eXu/Xv7k58Uxp/oSx+XZv9TT2neEzbEnl7hhwSpGEymcuyyMVJrXjRWzI/iiDY
961Xf1H4y2BxpC3yeAa2JwhZ6RpEGrvJVp5UfmzAtipQBibELTAvdFoG1S+uwWgSiUAt0a6xumFb
8wmASKS11sxYLkDsGcWdeH8SMhlRL5JOy2Pf+QSaHgAZYtIAY7PfNjAGbasXL4s1WxhNkeddUxKT
TUtz2ZdaXa/1lj4+CwOgHKCa7MmjR65WTUtzs/zuAC8AEn2lDjM/oqRwibLokCxoBStZjpGZsLxs
seHlkbZ4COFhmqN/zJeP0aHzozqv2Vat3QQOIs1XwTDymxzd6eB2hFENXAuXL3ACaV0pqIRIN135
C0ons0RufXtDqmBZC+DIj76jeXwwZ1H4YSbOu+0xvN2Hgv20eQMU9v5hfMuzmuplJyCZNeJGLri0
mlmkm/Aabz1NDzgG3JZvWPHVFUNNrWavpgY7s5W92zFaBMp5iv6dwATDOsW6OHFUBkj50fX7dgj3
Z2hrzeGbtdaOgU7YZA81WIUtVQVN03E0b87eai0vghUrut4n+M3MfGi5dC1WlUzAyl3/MzQPFQA0
9nz8qc0MRzO0l5y3UGQAc6RSFPsXzJULbdkIDEEGASU0t+Fc5jBlABrL+J7RY/IZNEms3fOI8/8k
sEp/ncx/EpiRO72r8mPNXCRjhXnX4jKDfL+mYcRVsaOkrAk1T8VNaB9SBP+ZUtpIs6DrZfLWmo74
6dx/aSdhzwHqe/lOrZV59LHf9RhfDeFaIxUTi774K6ZrmqepW2zZnb2fu7FqsopdMzZAv/WBLNVv
nDF91RcfsyLBeHpEKe2TD/AEpuCVKVYCwxweH4xyiGjoKuVvN6ImW1fW98VRro8XXugV4Em/1/Em
E2vbNhTsCTCmZB0MqzVz6t+B9g1TI8frrXS3nT5A6CxdeiZgB/Jp2HANWwaOUybu+Jy+Mzkbez8+
wwshZELR9hr1peXibVT6zHy9iF3bnRIzBLrAzMT8fPqpscj3iJqeZnVWTUH/QLGxwBRZlu18+gaK
eJkpaX8vR6N2cdXvsPH54kw1dIBi+ppcY7iPo9yVgUNXzUQoaSqltnRzeu6wIh7puKmujtw+4h1b
WO0ubzVrlmJNrroEeauajSVURZqNZjIPxxv/OBzMmd3jE7ccTaGNFFVpS8GPGGZom7jJ2KE5ySzs
jbEboXYJI32/9x0eXAOa+z8x3tfoXuk3xoPInZjhDLc6MaOwFqopGtRY5wQLs686E39Hsz8DAKyF
1cEN4wJgei3Szjbvdg95YSIYg0NGYNPhoybrIkv8CO9XcOeFvonsfcgC8MxHzq4J7RYTzBLl89Cz
QnalYuI1UEQ4SdLdRcSOIQ7IsKhJMW5Slj4bnrkvrVjL3SZH/OjiW3RcZG2dB2Oxk68XTsuDqURX
b23Cn9Oi2xd718/MSc5DS882P+87qI0EbmSTM8mjGVvjurprG2ftxdn/E+7oag/r1hBgLiqJkM2r
5ed4oj1pSzhtnVhKJK71toryZ8xUv3j6ao+RdkPJL9vOkQ5vdm354k327gJYoiRv73Lb9G0G/Ayr
lSfCfSwgnESPqMOgYJaGCDfuhxVsPer1wh0ixdi/kjL8kjL6E/dGRKV9sdPOOZPrYnvD+zheD6+i
sExofy/aMG8TrwYTm70kejniLCRJ5CqCI/QOh9Lyo18uUdrd+3gTAxxaINMFdkgURUcUo8G9D6YC
gwLHp8u1j5icDm3GqNtrdoERVafCyRWz1Jcsfcp2obG8BtffQVuaFKtHmDga0NnKmbMZ52fhxguV
ezhh6l6rbTFhJe6eYe8cteuGTHn/bfKJCJQD+QI8JHRBrTpj4adewSFdYsgMd/f8tYMTv2LJU9LV
S6ovFRB0hrp0mztgjItse+d3QY1rwvEzMF/VINlBSr8oThvXp0Std4LgskUZvm5viqDPZAo15WcZ
zAa3kq7WFvpbgbhNWEWP1d21afHoHxPj75++Nek56gDsEUTu+FQY4B5JaaNlmkHedH2BEUnqxXFO
cKnT1qwBMkaVrUA+Z157meN544CEVWmEzLD+wLFz1aOGeemwFtiDCCbZQ/bEztDyMjNunL2OQahS
K6BgmXtB94mG4jFQs1jD+jDFcNt8+kk6DHSsN/jJIhEEc/hYDbsfcEQgsuoneZseM1LjFqnDbINQ
H5GUVcUmMEku/u/siVF+ZN4J/muI5L35RU64Y4JkKkBIh1wjKGtX0IQNl7U38JOyV+ZjnTi/M/hJ
YBOTXttgyK8/I76rIh2sY41EOAdxI6Y/0VPjdriWNDranaOBCfQNSvztU7zqH81mV1IibZwAVOAX
9Hi1ZKdXsZXjQPCHOJ729XsMlKtXgNIwxgJyy5zir8WOdDebGBBGeSKX1mvJ2fJ/9zgi8EL9CkJ3
829WtDQGgouMkzrB5TqKIORb+S5j3vRNthrB/V0MNRSm0H7tPv1zLVLJ6X4qaW8H4phZ8VxLfQUo
2xoLwzRWUt3vZnRqZB2njtgaEDl/vfloZIvyPBUXlzhzdRx7K1aD4n7zTErdnkH6ZguNJokUwSeh
/5kUZaXRzbytxeQ1Uo3TuQnD5kvavXV+eCf3qXtqy8QVUipCmMP+WZTIOLBZSP6neBpIjXLclY1J
MV4sKfY0RFHIqYNo556/P7R5VXhCM5yB83EUawoelkdH6+kQyUOev6ZY0bYIRobf5ZZIjKkJYtsI
zmHNtHYI2Kwuk7mBx4j/81Hv4zuY12R4szJ+67Qc/DTHS/OS6ceDPQ7nHD6JhCAjKTdpo7tUJNvo
ZjRYeXjXNUgxDaI2x12nraatMeKgPM916jV557/ZpsOgyaM81jqT/UK707Qq3Lto5O2wrK7Vz0hG
8MZANvjN9M+es4XwFZpZSWPZg3mjUyPVCagfAj7M/q9S6JxF0AvNFQuWOtnn/FZ2RIZEulog5hCX
pUxpSLZF70f/VCMAE/f5K2PXMZhjZZTWVpAarE9BL+HnoRhvS+5KzNaAPFomYtHHMU3CQvrTLK/A
n/GIsWvOvhfQcfwOS6L+G9XT8zOidi7rhSwimZ+lAEFX1tEIcAn0RlZk/MCYCMq6PgBSopV6y7s9
vh/nS8/qegfQ1b1VwySYMv6n4TFmKqgjQpsRT96DrfXubcEnwHTrKUs4CnlBKJ853y8GeRzXzctv
NnhxBWxPAldxUiDLY4q75DQvY1pdIe9fpAZURCzncy2XiwGXIUdMYNa9LY6jYKj+aCj7e0mOyZqZ
YG6/FTE4Xc0BE4mBKynkk7LUWiO34+l87MtyoSPlQuXyubN3VfMam2WnwwhED61mQ8O3s+S8Cpr3
45clNJNrxDBEgNa6WdAOCLp2uDbUjFmAwPQ0d6n+1Bj/PDMf0iUjZACG6GglL7pCTkj8elDLzQkb
yomlwzKJYbkyAxAlsVNZ6zCjtFxD9nHeJIekxi3uLzsMXoyHuQGRSWzEjMiUBETgv3tgQ79MHlnt
iDvAPHKQsAjP1Z6uAgDxsR/MWIdz2qY5a6QkuwqQJOggT3t2vmQiobUqAXt3T110ugkVITXJyK6V
mEnhbHK6IjTWPJCa9AdL5vNe9Fx89thyKUr8ScZdgrE3FRoVHedEpOH0kxNdRW0P2vrJqSy+yYZx
FhQpY3zK0ZjTum7FvnVy78Wpqdq0HG5TsxB+kuvFz4hloHRxk5tIb17TTmxOjtZ40glDeU4pTxwJ
1Dd2BeSKu2L2sJ1zXxutzbLWHIqAyxte3B5SFgpjalfBa7JbaWSMuJCT5w+U1phnsnf8mGXMWWTR
aDrKZXRX4C+miL4rVs9yhlULXuKTQSFY46DnHpKyewaGDnBgw/J0v7mpf9dH54lTf34BwI1onvwR
b7jmupouI1PotIYdJoqmgzgRp6+xbJs+v1IPGAl7beQIknI17Zd11w94G+bhXBOqRsOEavRwlUXM
57y0ABx3upefYtH/R33UlOxPr+ypftA9xCZfBTB/+lnNKGg0skwvjSqELIN/fE5JcEjpG48znJTp
1Ema9NJlsISFx5NIH768KfMi1oq2geVzO7YSVhsNeW/1KZJpkgxFjNoLO2Ne7hgJVdrCAFoPDXPQ
I8PBtdbXRkh+7Vh7Akoet8MTJORG2ivMkf3Uq0dfUeUtHE8EY3XjSQU1C30lXdf6T/67HnWUIcjy
fMM/ByQ01PS4UNEDTmOzsaggVyZ95b3D1kiTlxwv/FK1bWo5riWOIS5ixTDd3npL7Mpyyq1MxDXB
UAG4IwQvduBTiKEtNwLr3xAMr9BvZKyAF3B+PiYuAuR8fhh17IrtB7vxGShzoZD9DGm1ZYEsPOtN
XY2agv0Cu+tuLJx1SC66ER2GlNAe0X0h3dQRQ0wxoAQbyHdqS64Bl7L6cnrVYCEFrUrWKlTNQOMl
Zbp13RSzlSUIEfggOEW9irBTbPLJdC98KEFxqhDVwZExkIvr2pczPjT7DcEjxuB3fMBmxovzrPyk
/PnxVZp6Zj4Lzifq2UIpGEFkMtWi7XHF8IVMLoWRjek0DVTryVI+p04lKujxx+KwEcPn8Z0AccOq
CSouah+UJMWkmWU1TzcsDkwShDcejv/58sGBteWXpoUng9y+qPVcVxl29aQeEupLuJ48CdlACXix
L+XZHc/sQlReerm4JizrVdS6fI93Pi89m1MlhTFc2U+nBTlYE7Z+aJ9GkfoZXVbS5FHfTWU0AtaF
Snt7mopw+PAZiGoiuWac4o9N1kChjMRcKJ/lY5TMOp4qGKkmJ6RJM0ksSzTT16ImhWdqdYVd8oiK
t9WF7rnKQ1KE+Sjv3IOgoqiUpElsF03ttJViWN9D46ceOz8WEEqZtT998g+zIIs6w2ILgW270ii2
9sLNKMxIP+tPfW5NGqTRUmknfWjbnrG0k2Kez276lY0OEdsj0I6O8CdIFo+t0JxOMY+Qixj8aEgA
byC9q7q9Qlqio48qiY4NqSBUw4FdBblr49L0ma2LCY6fUkEpZ95XiApxkTJqX2nZSZF2dsRm/Ht5
1uEUaqFJuT62tbOuEpxyoan9dvYlMJgs7hlSf9TwpcTUdoioY+DzRjD1bqT+Ut0W8Ew2qWgtFNKU
EkP7isFtvW7KYRezQy7i3B4M9t3cYYIYho6cy+JVk9SPNuGJREEawRy08iVVWxvWl6Etmw3WmrNI
Fk7Moji3/irk4AT7F4eGP4ZEZRVrcfR+EJA8HU9Azcxkxazp4+Azv5EdLj/kPc9AsfrpWCMz/Dei
xjZnzlYiTMa04C2KPIg12eDqXHeeftkGUo8Mac257di/cxOYUFGJb7wqQ5dUAxTuQQLCZcAQH2kF
DaeKW6fSM2Oc2G5Lwj7lXM0UyUrVRqD1G/2ZPApTNUrevRY/Efh2LzKISX1bwZMqJMOcSmJN7VwY
85165xB3RW6/RfzT1TNHCtsMeksqNTLqW399+jqX+qhdfDC14lc8ZUnj1e1fa/vf1i3iP10r/ty2
4TsO9oORLpq9hwTAf8HS8Sph0lUeXdUtaetQ5wR726j64XmJozUrWk4Brc8KU9v4Ptl7PSopIc2F
N6zjpc4p68xj9BvX9ev0V3BV9zNuukg5kEXnCwnUCBRduX0Ya5Og6H8Hu4ojZKZmNvcUXImgh8tU
VKfZ784pr4INXIpwtF0AW/qohHPLvI2fyCzdZJhFme7LT7ieaJzJqOQyPGZTsZujO7ldZ/Xd4dZA
MQhMZw4ITCdult6ret8bLZvlDR8TA6Gmoh3eSnkBDpMM7HtnBWrhIz589O8StzkbVxt7ADHbCIsh
ke3oGFSjN0yJDHvVtFbqQKmpQVsC7bH6NYNVuoVfdXAVfmozkMv0o0N20U8Q/F/iewpKFAzOte2O
QG6wAhfioMSfcSCrVGGKBiHs0XXpeIbtBQyIuLwdCLxJf/cmYOAKkEG0QVduaUv0coQh3pZVKvqI
LZ2mnUi6n2CEAL5cznh0qROAFjfT/yPUd1pKFRW7GJch54AgCqRYjfB0hyWdxOPu1qmB+thMM2LY
Q+P5WaTRqlPT8fBIqYdQPahbUNf4qsG6LOw1Vk70gKRBl/SROQCoVzhSCDBfCKFcm1LiLRlaMnv7
PDms0bhrYlXkhWwUj8a/WvEpSalrzSxhsS22R6JnGOoLemRXY28STLRPQXn94hHg3taft681tJ3M
sbd6ICrLT+VXM7ec2ZPUaXfKIFUz7nlsqeOvtkowsUZs6zEjTQJI0ULfchsPvTOw3gyN6Gv8VEwf
eaYj2l8M3B1AkgpzohGPKvroJpBU+vI3qxDeELD0RoRyRXMwOVefM+qlQM9v+dbxWKL5MlDKil2o
L94/KEhdIz2TdNRyFC2Ko5ia5LYkVDttwzITev4UClYEDyodmZdPqXMR0LD7DYoNHofiThzfG/wj
Nzeu+2lV0wQcnynnDR+cwUKtRHHse4VhRP6xE6N9J1I3oX6A8JaHU0F5AzTHrP+uveSv+QwwbyHG
MWc+QKrGulcfzCvdy78rGqedynUoeDuY2JeADjA3d0S1dGYM1yhxvI7KkmUmVEbeRfV6tywqeO3o
3gLL9gqlpB8pHClRAvzU3NRPq0VLObeTv0AcVWi60ytybaujWXyfyqDldx8cTGLsfgdAfyusD6Wc
O33Kt3XC4PZcQcwdDqI9OepclnDEOui6KRK/nXCQSOtPn7r2a15tPsGKK8hf4ttI5h0cKWMohoHw
md1j7cw9oe3f1VYhN8epsxcZpRkyzekc8BLKAN42s15coFZkv83yjX5ydecjobdRmL6ebOAFv98U
1D+4uzLqP8CcS5mRmschMdTWEKOyHjAVwkmju8Tz0MzDAaaou5iy0CHNcBY4W42vy/zLLoDba1G7
bLDNjiGac+pDftTAKnDquhXxFc/Qs2R5s3BxgeBZTbQwELj+o6pjkW2IdvJUxQ7SRs7sVn6SCn7V
sjLSkJ/jXHN9DSi5lBnQhJBdMkilRyx9G4jP4gql5dFzcNumDCYCyba56t56euz+u3urp8B4aJJE
iJeGSbutempsWMxGbbUqKkZAwSsy+Vtkt270b0mOD7m4tPA2G7G5KnDA7+0re5uzxoKmRUtTDrWF
Oj2di7sdfJIRo/zzRy1Uw6fpPRHhRCtikx71ftGFVAx1f1hmdXGzhVumgh2o+PB72/bzR7P8Ecnh
7+Yln6SUtNODnOiAhQP7cfnkEcZcrfc2h+KOyMSDYWomFnqWdDERdyKH8QO4NsWT5TxvhP8cgKl6
ENDpryRppTM8Es78SEolyNmLhXZXgJEmdR/lM2eBRiSLcGRUDgm5EQMPjJkuR1Xl5qcALUDVMhHz
+XHnmuBkHLvvIhAmS8GD9gJWboiJzyQzwiwFmxqaGRMcx1o0TrBliWtoP6kl6Ey45uVUvmBJC7Um
F3G8BXBgAEbcyL5vbOgefyN3TfJ5e6rZhvHzefOh7NqFABhb3srMpiyEhc9jsZQthgL3zUrdWEkv
5k0FgxfDwAJ7NiM+EyUKUq+KNWpms945vPhBL3LXy4rBTaYQvA9Lbbhqx3gIE+OWdAyZxWXlsFri
3CFvs87XkFA4bzMHhVEx1YYIho7cBda8GNzMBTN78gWwAvNbisRr6p8l9seg7MUk1FuXN1vPWXbt
VnecAPkZ2uMdy1F9FJTHyW1tJ5mkxhLTYEjhtmWXSCYr7xrMjy3PgyoZRpZnTFpbwPR7utj5S8FY
GKPYwcSEGIn+yA8qWFFjY6q1bOZo7JQuwuXIhPwJEACDw4bn/ZsFepS6ZlprWI2qhyub4sIuo2/K
LpAhobxRXXj1pQ1PhbwbYXpdIozXPklk8WR/QeiEy8Uj1VpL7p6Ojwq5gI1gBImneTteZ2RuK88k
sn/+S1OnHPKyJKYq+ZFdK6pjasgR4X+1+dBmU2H/+YGAkap05cXXVB51WJgkP2kEXHdM9XMq1OGL
iTIOSpnvWdSQFj618CHCEBoTzApfmyc4eBFxAf35fCx/17Xi+kpmx0iOR8ei31GWnQbRIoHx4R6k
mnMTi1hYBpu1FzRupXJE8o8QIVpwiMF1YWRzgsLHjXEFs4ifTWiPER+HYsSz9VJqO317LUSPornY
4yTW4f+2cue+88EKFk1IB5jmH9CrBorxR2o5YPZ+xQbf0B0y2iaIoYQc115xR003xtSTUN6LY6wd
ILYCv2xh4y2NWJDeOJ+0G0e2O5b+BGeBL93ym6nMgrm5yyLFyBsu/FHo1Rye8IniBRkdTl+9+Uf4
7Z8RZ8HyBrqY2vyUeynJkVddFL4nubeJejjoFuV/dC1FdJBiWbQ1cf1q8q/jVbHZvybG0g8mwp9i
6XvAILdwhNJiwvLMtY02NNcxiPA9mfAQvNiGOwl/SRi/vln2eUxMEclesHKFArhPSx/QbrYi426V
0LRLnEY2f+8GY9jCFrz42GNYTISsT3nwoGtOYHrv0TZLdXVZ0XhxyQhIje5I2abNszTL0hNnSRYP
03XVa/4AndcYrjX8hO0ofjxHb+8gDDQUxT1sFopfBuSqgHAmltb18/GbaVKxYinlKwpHyj9f1XLi
gdiQiUj5OrXbVbyh8+E/PrE5BJQikr4vslNPtH7sSi2qtRhTfCT5ge+04tGrXhcpyoIajy58RvZw
Qzlt9dGCBzTKm6glgZdFz/B0S54rVMOf/PtnU1HogkFfkZwxKV0HmOafpvMsSyJ/BmSjeVynurmS
BOMAI7AXInLH15uf/AGb9Pr7rzw1OmBCdC671I0ZiAAOzIlJMkXXsfHF9xZBUUzlFZdxRdFXj7gK
NXQkHu3w5oLqwDoCjnl9/3NiuCd59Se3pvL16a+HN4h1RCWdNkx6kNE1e1LxhVZGJ3y2jypByG1r
URpG/jybyXaErquVkU6xd51kUjuLfW4UuC87UNoflzY4wAB9OGaj6uY4jLVz7eyEXm+Kzvc+9p+h
HVb4FolSNWerkPjUDWAe3g/8iDMoaJd3Wdh1/w8qv9V9uNJBKT5+mrHoKLhoJQLsKiNXOJ3ZsiIh
NYzwuabIwM0EH7GFUzdNmxRN82AVR9ambQ4D38qk/0wi8dEIWdsVsJ111DZE5g4x/CPDffmDRrOD
H4wDK0wOGNymtWzl4UlcvL40dSGtyuyEYo/fR+iXs/4/F7uO638BGEYb0iB3gdg0wOq37J1fBzPV
sOl79VUHAlanu8Up9m2nxfsLHtuCY0XmEP0o+J6j+KZ7FEk7gBegICgTa+0cQc3qBOMR1LkxBovk
eouEuMZAT4bF7Mrt8sC/eEMcBj4zspVSsioN+oRHouSKJL5svZlrfNZ6E9leaEvJ+GtcANo2sGcj
30Rzwh7Ia/SKzI5FE7AjL5Y9PBsaR/hOgXvuW6hA+eUX4JG4IbVq5H49JCyjrsOq6jEyO5gkfR58
dD9gAN5pHvev7U0I3p2WD4l4etb1Ryr+m+oFvRfMYd06K0Tm/K68Dyl/3U+XnYMjpFrCk8dc9zzd
Bu4FrsXjnsfkExhazl1HBsM3l7Yi5oLsxwh2G6SlpKutYZf1Z7vD85V5vjY2quFAd+GLitVjHAE9
rZ43yXQ9psHv68uNhk9LuPzbL08V3df6D6x8RwcIQJqh8DKNJk8fY1+lKgu/cflB7H7pudkBwnCK
IoqFMS1DJub87eYNWdh2PTy91chQOghmcFHrM0x3/UBkl0cg7f+SYjAhWCtxGAVkGcGpcu8SvyEF
oP/MSZQWD5R8W4R8Afc7V8jxghetOaI+X1ho27JevCUf//T2RZEVFRp1liq/NTzL0+0N7v8Hddng
+LpGL4jNxcwMIuPPXMDgwWBafXE4pOSJjUFORPL7MaDau/MznPbwyyNbzkQC9q73XlLEq1dHf6Cg
qROXRWBhJfF/WEQuW9SAivOtEK1B8uPkbJCRh/Tz2YPQaTKFOBz9b+7zuLvO9pkCZoaI+uFjlcPV
Yb7WOFCqOG4DEScDevl5L+HKnNp+b5IZZAQapr1UFMGf7geunDamy7cj4Y59ZpFXcYr6nJhFT0Ab
IkQYBSj3whhQ6ZeH2SQnG8vmRSjkXOvXJ9A5DxLJR6WDQWYjg4QyMozIPbchM5qBpNeHwz4McDUS
lVKjFWKuZ3fDiCCOoLMhJ6vZO43Kb4vgv/6+xNwnGVvJFanO3C52tbxzsZ3XhpiKDFXwMAC8ZUTE
vU8Xy3oiVwCQYO+0oBSjeWOoPCiIjklYzzrse78noI/Q2dl8HjGabREo4VPVB+TpZP2mKCxd6X30
SznuGqMKJmv/kaiDZRvkPWxJfNeKc7AJCW4gWLGySBrkkLU0WoxnMayp5+No261kcTJRIpX/AzpG
5rRjL4oCEQz9hj/iEnOrY2V1YlwBv6flrCnnRi7AvjGRfjxYheU0V7PWe120ctkJno5KeKYYq33U
THU6n3CRez5IfXnsqV7BKgZQiApNwuu52mAGaY08zwffJ2WSg5hn9ZKuru5ZuNlEmOfpiV1/rs5w
4mRLAsIjdqvs1ngEb87Lh++wsygRquBzVakavM9+sDmvpzxXHUJW7NsdSrMIKS9v7VsBZ/iqJrbr
gfJulOI3yiF+i+69m8mB2yGIde5OaS2/73iqix0Vq05Y2a5dKwUglfqW5j27csSFjzwibD3WDM+C
CTyZVWXagCXXhlSzGj9WJeiFdxNB09XF0F7loTWkOcOuZnix1JjAtr+HKAs0hGeuGAiqJQ6XUiXR
mXiF2LJTkSPx2S/7e3EcrDg/C5Hs9zReu/JkyX/Cg0iUtf6JgMQz/0VsZRgQ5EyJCMu4sLOyMqLd
4nnVj9eXQcIYDlS2Al2cF2rZ+bE2285tc5YCf8Fy+Sz/qEMJ/qe31lbLdv0L9LHkc6I6NBbixdy9
kHSIGQ2olr1Spt5CwwLdqbmRAH6iWZLSd3wRNRgdZFs7c8QNR8yMVoIyP09ThDyj+7Uqk35UOnts
t8fQzeexFrDiy2hELwr6gmDhgCRcR+uxgGRxmrHei4HOp2WvZXCFsjIZgMBss8BR4nzSHjcuss5X
3+XChje7aWyK4HhyJyvm1zfGIJRLyD+kc3hT28ApWEuQqi7XziXMk3I1+ZqL0oT/qkP7takiDv+8
w7lWaix7b8vqJWDejM8D+RNjlZrmwzBfpyU4eUUpXydLMWHCSFPj+EznTlltrZ0lppcc2544BKkx
QTSY5csv42JgSuwZwW/qpS4x5d1XOrkCRY71TB+yfz8P0Ci7XsepjyRna1GrsFLOQpyk45y15RuF
v732ZPAyyCT3JGNL3SyQBSAqvZANlWQrz/rhfPUoRdfo7hHrapTDCCF8IeukZvSMdtnZD8j7xH6U
o/WzMqeMlDI9O7yCO1HusDgBGu0E7dEGtwcChRsNdiBT1yNXFusUJvVycbycaer4k8JWI2agDAfE
UmSsDX1DGwCjqS20t6I3YxGddxS7DnMyKTOKBLGK7KeXNPVJzjgdzbwG6tcg036pFhcw0fX08wKI
bNq/RM+1AIyB4XLKngttrte2zxzjMZ93ei/QvjOqVffRaNHCYZiJEawb2+lPDsz4ojSyXB2oY9s/
sEWgGvEPp6AoCwhWg7m5BpgC69FJzbBM1kg7ZFxVljqdGKI3xAq3m+mKN89ivrECUKKsO62pmbZm
GUZw1wOu3+Ti0qeB1Tc3ym2VmwdbFY1zhIa8w5AdGD0sQ3NRwbmMOFZRAluQgkFZKLwiGsByQBSg
ycgSOWtBjG1gr9CccNGcViRaXReSDwIfVOgDpSqx9m8GrYKKqEkL48bW7qiKHVUqDRtKkMvpUZca
6+nGEWijdqeic6sw1cb8o9PppX4tg4RJcfJuEj1FvxfWvNGpgjtIbawHRyzwFsId3UdYK+B5dgjk
bqpav1mTTn4EIMh2bySmP3UVB7j4vFMTaQoUjrpifnnZsEGFF0G259M60PtOGI55MowaO5ywhUM3
7M6HDAB9IqMmIs7cWSdwvOHBTxJHqcR6dNDiwGc9583v+CC/sZY/13IPMxzlIe+RzIm7tiZtnLfg
p4SLkcyrmndo0wZQ0hZUorXbdc3laIPiliU/VfOnAzcF+ZwR61HqSF9qIbEX5PqbD/mWs30G20fS
j1LVYD5mly3ZHYbxLV8Gh4NK26GpmzyLSrF+kyD/JgNym5ktbqLMaTunZR9g80zEBCgJNiBjzpvX
Qs6VswU1kv9MRkabVbbXDuFHGsnnDXz6qhp/geGQd574R7MwxI9OS+WqkDXEwn3iA+Xz8boCa/OQ
xJ47H46DSvbMO/wMJ6HSx6IXyltz1xaQzWSBoeSaJpGxjHDLIsSvvgOEu0/YxPrPjla/sx25FTR9
08x0e3Qe6n11x6I6WyvNpeORq9xroXmyYoBNDYsIkI5EuKcS9h8kyR+WklCZz+xeKH1XtgQxKA7o
fki1SmG6yzP8HyK0GGyFwaq+k84AQyMpLjwieakJJMgkHkiYiUSuZo9YqVOD86IICGdjtvpz39nx
LgKwergGZh24fgzcd/+vPDXfRDSGRkMWdg03WMJOpSRwh5SlRT9sUPZ789IP0sgukqRfGuQM/XcZ
BfJnkhWGlCxCj7P/S1dth5UQ1YyuCUURuim+HfbHfjdju3Hr9BXQR48tiHFB5GwONgGoGjArigrC
hXOauG4Mn9SihgS2hyzGWWmu+Vj7iYxB5qOgMFx4Uuh6rdArxELVRIbrZHsrj8iteQnkEafxB17d
Qn6RaCvZZSatS8uStlR9Q8U14LVNW2r9Min/Tq/sQMZ4Y7k2lAGCroaUx5UuONcfWb8Mc/KZ3+SP
qmly/kzpEiRvTOrFT3QHLevyxKOXa+3vU1p6jaEK3s8ZyMoZIfNMYVDUPJUPwjSqeJcQPNuQAMC7
bWtunplOKanwbafMVFDbZnsu87uuHCyShAkF0QvvFIzWqEaMpll3rMzPiBI6Yhe5QUjMkKh/gGqt
X0nxcvCQJGGhLLCC/FuWW4LH15mBBa3uXtx2JiyB/P+x2cisMEw36Tj2a25exymlUd2jIQzoYHEc
AxSq6CG7To/ht+A8jXcIAoAnUDC9DlK0sgITHeQSvw2Xdh3E43NaIK4ugaIIT9HoXdgeQMV20t/7
SfzpPog0ivyvZ2CUuuwRRq8T/fpKqNM3sAXXI2sqAX1qBvDGsIcbEG5vedWtH1MMunXYTF9lffU9
SzUCJu8CPvOZ5ztd25UQiuWO0lc4P4oYNPy3w7VfWqYRyn2HNY1En4FqBRiZZHMjDeqRyk03sAWv
OKrnosyw1ttSKdxEwEZrPfx7kdD6aApJhx82fhLXtNgSpAKV2fWpXup2m7QUQMlCWWduYNiJDrOB
w4SmxoteKXgpIIiuY94bcfmMYsRVQyZf8RDuBSM0lXflxU+dOYEo1yxXi7zNMmrBRyvm9ZWjnOvj
cqykt7E5UJFoVo4xCLOadkYxT4Xx/mAgxbgLb5HLCf+P8A7TcFL3FyfaL2Zy8C4bIHzkvpL+XIHJ
J4CG/R1/VFDSP5VVtTOnJb7yussAGt5RMv24Exw5kgV/PGwxB5S0r6Fe3rWdaf3FiC9l6YzN6Jtc
ojLwcr0qUPvRz5iGYLkRH25tYbcwKWX9hhPHOSO/KLNjm3Tkm/50Dng4QYdpbvsYy9dUnY7P3wmu
WsTNK9c3Aq7J5DBw3ImfQzbbCZZaABeyv5ZCk5APAwDL0vVYwOl9zdmjmCSHxgZYNK8sHShft2/f
gZDijo9yi7cMfHW4fsQb1olBSGGd8Tcpi3E/zQoibPHA2Rcvc/4Z5ng/4blXI9I5LH0KesJbFyDz
6uWPTcaKOHVMLflAC5vqKmaPD9R9yYnhX5QGliYDqzjIdspJvdCQysI1SuGH2n5veeJjc6+o4hfX
8URKbO1QBtAuEVBun/KRkLrOaqxzuz1AyY6gxbRNI9jurNdNRIQJxKyxzCHfXr2rg3pdQvmJbxac
BD/at0BWO1/bnv8b9epJWTidtdjzsZN3lS6XxjVtTmQW9ZlWGbM6oB3lD4CRWPyif09aSAsvgT7m
URnecCeKa7/OfMsVnwkZDckvrxG7DELGe2OdNICSeTSbUmO/PzQq3OxGMlJuX5X/oOnoCo9bgrDc
D1qKgF4oAcjsHDo26ZOeA8qU59oOuQJ0+OgLdqpj8hvQsYJLWUwMAokK7EFZr6w674KHoQK0VbhO
C6AOfE5+BcaS/Mqz4tdpMLN9BzA6vmf3KpY0wIHKWv1Cp1KV7DynW6XrpIx7z0nkDeJdYGXFIGb3
wp7R3GSsXtLeihtu74AitzhqZtXk8JDiqOqS550Sk4h483QwFMs6SJgL8gov9hQmfPCcKIUNuCFJ
NbiPOhxkwobrWJyoGVXF1SdTpsYZX6kq43CGGtcuhPsnTq5r6PdCAREzGSK+rCaJYJGSBnXe2kQP
h66vEjUJNdt3/cMoq0qJzOgcfFwWgVU/EbAGp1st7+d++1qCdG36g95H1Qfm8Mj6AKSjlDEAthzb
ZeOuB0jWelRzFSv8Ko5jml7Ueju5om3raJJCGeBCxMJOWl9rdm7QE8Z54GdIuygulcxELvwgi75g
et4RqvQ5BqGNFNt+jC4SqnXSlQ2sKSDFs+CaK6cScApxg0NpeUCCxrqcoVTDc2HM9Vc4VEhwdKxh
Dvry40eNq34QGgMv0djlzzevxUuZurxsV7yLyQRT/deVTXt1Y6A5sG7of3lXknMa+edl0UoIPySD
1xfZ+evuffQkRLw0izXLG6a1kDZxdUHGxUul3pu7LlQGanE+CuX3wh0QrvZh2OqK+WbfzanLNeLT
Ud4zkSEY5HXQJh8ZZY9xW6PSa/d2vom5m3MOM7kjU0/o82ksrz5hmD1wHJjMztCKZVvgNBZmniVE
KGfBY+SEBazBeh3sIZnQ2Uq8Ua1F+eHoSsE/mIsSkinT9lllzUjW57etw8lW3/WmxcPtOdQQ0eM5
cnuk3REa3MqNWWp8Z5hmsHaBVq4kB+NeJ6czlUnozAPcmUWQl7tJ2sIPmaQEGufAjd0/9f7+baxU
esWFbBSj46LNiWXHwcl50xlq8hX7fd5BkaIiulYuzV6VWouCI6eRIUQ4K2evsy0FcQZpmwh6g+mD
fPd5+x1EODQF4hBfrkmMHlIgwPe+9Nm/8veixGXmx0OovgqV4/JShird/dBxmwwFLyOO+JPorY4Z
ulEPcmDAlXLbLJZFWkl+s0lQ7HCCb1JKvnpre1Mw0V+Zlc9WKNeXKpMLd/npg/MG4NbmzR48uIyv
RAozFXXaIJ/7h52n3/Mmvm3EIu5UAfU6Gw4io5nQ+A1zhVnK0XzJpP571YoM+8rk3jxyIfwwa/IV
gOIfiIea/Pb2zChmGb2IWX+Hy6TpaOVnj0ZZEJ2mLzPPJVdeJrasblu31vk4/Dk/2an4WsZ/YouZ
RToW8kuJh+0uIkxgJ3sITNiMYu1D1l5Sm8/V0p/g43b+1cjj/4UHqrH7Y/aGlzk4aIQpgf57S9yl
zNr/UG0MAlhmfOZ6z3oADo2oQTh6muRRggyeYCxtGJXkGsSMJyaa5ImjkNzuRftRd2TwKFT70wqf
PyqGE9iqOa0CZrglRoRVca8S8CpQGbVFImKO66xodBB9KDP8Du2xs38Pnfn4qOIhxUZRdIR7YxCD
sIkk5znmYZBDlVxv2DOW40a40q46+/b9S8Ps+I1zmv6eE1+Aq5g1NseK38bdkrzyZKHgg6TgUoLg
o+iRiXtemZY56EiKr8vltv0Et268RKCez9Au0+0HuNMRCvthtWSfnJ6G1acSef2ylYCoFBjw2+8v
tS6MUV5lWpkGxKhLURRcGHUaWieP42Lp6cGQfTtwIXxisHE3St9ebKCk8SMtmjqhevWx1R9ITtMV
zaFlmRU+j9njNRQwHfHYJYHL34OgA8Twe5N/3pg8Psqi2wDIGarLkKPsn2z5rDN89qh7GMH90CG+
Z+R+LGMS2US/FeRp3a143DTONcGiOgKUa791LrISdHe55xvThnfYxCAaCJSQaI/HoLBl4FaAlAwc
UXyrIFXOZdTctLk2POm/KKe8BPWaDHbJnceoEnaeakNq4S/X2XiTvpI4PIdf3cre2pI/P+nX6yVO
38ylFOg2K1Giwdb9O7STs56qHndSbRKTpbdiuHIZn7pHhS3otkBN764hPdH/Lt6Y6OlEAEZQtSyC
ppOR/3lgJNpudwCc5FXP7JkJ1qtrTTHIGHPjZjen8jy80aTPDvus3Z9P9qidN/9hntGLdKY5eI/K
vUrhCc+U/O3dZM0T6QbaI4HBipVkm6MupjbvdNnHQnr4YU0Cf6NnjKxoMNtIZBKHt1rOh4aqfIpc
gH92R3uV5W5Di1Q/5uhCMXC6IO7NqNxsTyt/qr4oMPJk+xdoJj2nX0zLVGALAiyIjPGdqOniSE3U
wk236ntFJsoQ4pWK3zJbX3KbJsCG4o9QDjLTbH20fVZeQ7bH3a71vP6DDj23Kr+HCzUvj2DAO+N9
qHrXEU9v9bAAGrlgBVSNeLtrmwWuXK+T3w2jk+lnCiOsUjg6GGvDG6hoZLKfX7FshF7c31JvGw45
InO0kYpVVlCzN8Cu4RIOcOfSOOwMpt3FE/F9pZGLIvAI2p8zvzFlLX1lOGi6J3EYlN8DWdTDKkx7
wCwxYSWXULmRkkaACJ4aBBN4sqeds6hqapx5ttv8zz3+itkrg09VxtcHI0Rjrw8w7tBHbh0vG6bR
uVPckxwPqRdc7gyxI0rKS5iukamgQ7RyWugeN0qtH+Cu5u+rO8ar6r8pUPkXJdRjk25fe/b/rovH
hF3ZRTUFUq/QJ+JDjek7wQYyTTb7zV6W63YWJKJHC8VGMLtznq5KsOt3dJsZd3tl4AMvSgHUfTSs
6XHG4eqQNKX50LYAVOFlfwza8saKQ13h2dS2vb9EIO/NoBf+ILFAAYxfJaKYhARVYtUUg8yKwWam
22zNQn0Ah3HllB9hYl0Hq8oYQNgL+yNzQQ9Ggn0J46Z94g3Q2umhFR9dLJC2ocqkZnqb8HZIHc3e
e3+le+MDILCzVa/q1S7f7K8aR+b8weM12iOAec2X7rQW3auGBtJKuvUTt4OEhNWNYOjWq1zsXezN
bNed0I6T9A8IeyvbRABFJEr/94tBBBLNP9ixmiFLcLHj4LfdAQcj6BqbboNkjVrc4F6u2MC8KXZv
aKegVUv5WY6c9QwKn4Wb0GGIUjPbFqsXdYBmgNA+00FQ4dBn0nuYoxQJgXcz9cLj8hZ8zWDtJ2i5
Sco+MS9/UQtKAQ0Ie8kF1NSGYJMG/z/Wr43txlfFb/kPlJMjab3ImFiGkxdYBDi7bSiRgKdbRuyk
dLcHJcbrVvlmeNGfpqI8NZ1yCd5y9uaxPvmBQkjHCEMe6uK0CTI0WOaHySvibRxRJRe8Fk71DCJM
R4dFIE5CZltE+ZforO+KQjqdCx7YVa0jb+OzBI6Gd348X+HtD3eyNB75xAxQtDR1kb5s4coWlenu
ajYtKJk8gNfuvnEZjL1Wm/a1TiYmm7vXlu0Z+PfhuNrtftNUp5NpMmf62wRiWczKNcPNhRFu2kTK
zJXnxSgiaxTzgjroqYzUfUre/IjJuwnnhZJjiC9WKDuk4zDJ1l6uj6gpjSt+SPYYjicNdF/ziQFe
8y+zYREt+e80kCiaOhF2DWgOt+dUx7K7H2CGvgCl1HpTvwB46fS4ohMqG2bcvah4BNcomccKCzjn
Kn1y9Atl4nKzIa4ipxcLF0ePbcWgQdBFhv4QgzymuI4JuCVED/Z3ZQnDsiYA2b5KZR6xS6925ykG
LwcacgkUT1DP2tyiadx2L3+re879GBPsqTFh5sjmkaRalKojIHsnLomudOiZrhHznUMva1XDTY8N
+vG0K9p9kFLHk3LgqMzDNTtDJ35XKplbvdXBJwrUsmwUS/hjDoT0XUwWIaL1ovfwfXqQxLcNgoBs
oie8gxD3BoFE3MnqT9tD6TXWmO98BlyJOZs494hOgr38VwCQlgbRPz/geKck9ff45+D6u1cWfGzG
uypVuGK62peUQJA45ezWIDki2J4+4RuvJItN1K9bN1E7o6gqOR+h5TrnRs1/qZKImlLVi6WykNp4
Qxbfoqp3mRVDWX3g8jRsYUuu1DQ38vjgzX+L6gUMC5ONcmF2SI7pApS1pooz0vI+XNbc8FRdM6cL
ExWmFEQGw5gU8n5OBfJawoK7sTVUPEVDccHPDdhe7eJHfuNmenbHOzl0E8O503ygqKXJRG/dtlOG
E+wYHj15tcBgdHbFZgUUoWGNJEGMiptjUpfNAv6uxBgAZ+A2LgoKNzkjRWDo6Vxx5TwlxJvKPcEn
XQmLzNDCGK8AQuo2Gu1eP3QMotsCbKiotIm78WPM43zCpn6C/0nUiLxmamFP0jW5ph0hSoWg4Q6V
2L0M3Wexuv6oS/ATsxFGRhIXaggi/ofQKE7GPPBb5J3FKrWx1QWfH457H4Vfkkl/oRED5+LNKX4Y
oQQioI4YFoi4j4INsGHq/1aqAARtGbhy2AKhT9nUad8RU+vosr/baB6cdbHZZzPBzSTysHYfmw4O
NRwIei944KQ8Be8n/gAr/pIBLXCBs9PiC+Ql4JuiWeJi7JwwO2K6ZBvjyOAvkCyWKl/5O3AjjkY0
VSA4jH6HfxodaW0i+OVaNGVcGeO7fLx5znvgrGnqA3nmmT71HUp1r2dx5he0zVHXvl5E58Apd5Wl
Su580yNw6gcjyCD03URNje0JkO7ZcQtzH7pff92+Cl2FUyya7pgXfOTkYsdX0CUGfOAgEj4ngPKS
HjyTLHM6C+t+HHfKHYEkVbrgz1cA7g9tOUCvguOZ8hJ9RP0dqFcHlJonDtZfPd30kgc5V/2Wpxk2
2kPXgDrgGfHxiyuKzh8YzeDJOzIQuZ3crazhoHAJY4Zwf+nQZCgS2zBE2Eijw7vpdn5OCEJIfkyy
K5jIHxJ4GGtT2O885v+89PrT+3rHPeYud1R5rfFM8yDdGpAktfLTrKN0FkuZAopj9zNqoJ5svy+s
xj6OwLOynmtdpEDEMMRTXZ3F34ur4xIovbZ7sZdz9AE4ND3ifo+PIy42jOuwvBolqP5eolG5vdKY
EyhR+3Yf+/NYPo7ZDlfHFEZmJI/HvjWcdVyh4OMrzyVSg0tfiW7eGoYrlwgy54mF+dyzvZEtgwH5
ltcN9kzlMfmqPuSl2YanLIc2fDum+ixQZHfrAYQrZqTiDXBlfn/uhqVjxMX7cHz7nRQ77St6k9x/
J+4RX/qjsq3tsPNLltu0+M5nvHUK9wJ42KNK8KUaya1QT3mjtmByc7lXQc7p7bR8RHfLMIDlEwWq
cRoEI235Sl3LWyoLOC0rqYNyp7zYf0JCZo1Il9dOizuvEz0dh5FNWDp8zjSkW4YArZaP99qVLDgH
sO9tJoybdWoN57obaIsaPtsSAok5Tzflt45Ofd5ysUJpcTnLaQgvXCgllB1elEDQ76hjtLmqDizo
sDsOliQV1/2PO4OjmiZJ3a1iULhpKyPockDmzKvprlBomk8ffblkC8VFyn9xzv/9c1YsnWowCLwu
MM4Na7RJ6OldDKpW+9OqomO7ZZsSsOGN3Ugzw9FlAkHW/mzkCClWBew9ivw7dgXn6dEMnuxTUnag
WKlcNOzeR7aHloZ303OFEC02Ubsw346w2Y34xR1yWdhcJBsmZ2KgtAB0lA8Q/3/FjqbhadWXikw7
JjT3VcPOUe46KS4g/Aj5oY9/x99j/Iq502UcSeLU9EZU2NzsEGFn7vd2RXjv8OCEZN9GPFgKKfKe
vhE3S/3kd7HUXKB3gOy9XwbwzfZuevCYs+DM1aTx7QI//qsDElFvyebCqFlPnYi4OHK7bJGtKC11
K8+ipps+CRiToMWZXbQyE7IQCXcC+UQLOPk7xIRyY45tLmAJKDiUYqm+TATu3sf88Ib8kiDdSuJY
UqPrhyCv+ZGEabbhGjiUQcvYqa6Kb3OnDJrwjPT1Xt1/gRivNFK/dhtFpT3hLFsnlG4abRNXlayA
YlnF/m0BDgRDUYvrg9cv8U/HaSpw8dw8l9wfoYw8a/51oTLHyoAj5VYnmLmr0P08zeJujj5Q1YVI
HhDMyS2scuJ8UTaHU71denUuIjepu30KWV89mEvjXZwveDqm/BuMEsAjTcRywGzq2DLw+sF0BM8v
1PVR3CL7yBXVbYEpMZeyK+auDYciUjQvX4bCUTLXddfwCK/+YJkXp/Qsw5h+Tv/+3Ed+S9r7CpJO
EY3NVy70YqeO1d6GPfkrNCmTlVUTpLNbSI6evTQzVL2zF2FzRZki9hWxe6ZBuNBEbPYZEtu9Qlyn
89ZRRHOtVbgg49xeWCj3+x6p5MfpZJ8aHe4npCPBuRF8PrYJWPZ29XuMoKKJ+SB1FlLoj8wZM0DG
JSxBT54ar7hMWn2340QycZQd63w0B6aT84Siu/C5m5Rq7OXhvb5udP3PSWyAkbCSj04RaDf7y1wL
z329Ua+J1lYb06Y7uHXoJl8z64Lf07GqTH89LYN21RjW7Bp839CpBZHibvXUVF2jlmEEqtQ27S78
owUZ4DLxzFNvzM7pXK7GS2FCHBN0j9w9tOnfPjlwCCpbhs/OCbvZni8OQKoWL+nxgrVx19Yd6iJg
O8xpmuuUJa1i3ybeUTvA3vHQpHvIQdRjew5+xQpI1aNTeCg3wKQxPzpAMv0hY4f4R+ODxvT4LSSL
Tk5B2M3nOungl02TSvJCADEiWacwbF0VKPM9lmZba27g7WdREdnFPhMya5jShwaO7S7UaPk1j0A6
uKu2zeG5VUPkGvNsJdJdKPrWTIj/UNHNPCAsBCrZInU7a0b0COsb5A5coswe86t4i+NpPz+WCdb5
ybEubPhTStSoUOyOTrh6JS5V2eHKcdHeX5owgqVa8jQ9JyP6l2ksKhb2isPruR65oasUpajZYJiO
0hnpfRc9DnWx4Sit5klsbFuqu+SfXIKg1k/59sBgw+mK1oOj7Cpe+IcWUwqKdWLEGRu0FoZPFwLI
e9Ca20jswIZZQEfx15d6//jhCrnWsW/kK5h8SYCQrgXUzVLzUgdyDjtuS4RzNv3V3JLAvhCJ74MS
t/U0Bl4qDKrxU6K6/ibAFjJkNfFiZoj0YeFR1ZM9na82sBHlJpJCWH0hIZmv7fpyxEitoBFio8Yr
dRDoDf33l4ZAoR7EDKz5BRN7S5QrlqplFfO47gHBfJeZlOsOIRTGbQ8FrZ+fDuIEH0nXuyUU8JJT
y9AO/ow5H7bMpzRYZSbNWmVMPQRGlZVewSOnhmCjhebWd635E70/iFdXriCOjxkERszQHgwmzNx/
1pkOwicWlQIJhLgzMTy0RXKoW635aA/SBY3YOmvHRN1IAWiGZ/8Hnfyo7k4pP3bYjciUcHUPCckf
RvsVBps3yPvk86WsSzY0lG3TgZmvOYBizNkTnwJXOq1SvM8YJKIZEA1vMCk2+MojgmFXwFE/LfaO
CMe2kcx6oCPhiJLf5247JPklFX7KKPzE5RTXK1kM5UNywFNZmsEUQwSqs4dnMJnLkybS7/sms3+G
awKQE/hHqKhwQym/g4G6Z1CZArDT4L+yQ85Q8CBTMu4tHnfWc2mQhn5sUkkHtxrLmM3AJR88nckr
o+Cpc4QZJvr3YBas4kcZFjkxl6ATKRVvvfz8pEqjLx/3odKnV0JwrtWRIZOMPYYS9c4ibATiZhyF
usqo+3MfeGHUmSuqjAHRrLgSWs7McBLRPYBaQG5+vtwQVOvVSIpwUJDakKm0ncG6v9niL7LfdXZO
h5W49aPk/pHMvegCBKlDuf/8Sip7hSFWcwHy+Tpl/Vu3xa9SpGWeiBvyi/Kf3GjELl7JkjiHHBxn
gU+8uHFwaOzyJJrZEM+adllGHN8lmX9gGC7D0Re+pKCvTZTZUNvHvPXrikMaeXwRFstQBZAjgVB1
l1T7bCkQFqhvtjySrMFExg0AJi/m6fFMzlQvhmiAqqcdLasaY2kqTxLo3twr2dtUFoGx7v6bpiJS
7xfuRNX2iJELLgx2zy6zDVLVOYPLfrfMqKqDtTu7e/Ee/3Cy8t+gMhasMqHbSjxt31Qk5g5g+Av4
YU4Nd2sQMuwk8px2drJaBsYK2cRZf0/SvApst5g4m/0G436vWr/kXWVhvoJO9o3UKaSYfwk8r34b
+88ufETfJb+1nvYFGdzz8gYSnAugSjA7yKrL3Qb0t4mUm1PXRW5bFYRQD14L8p+7EzyTcOax0BFy
a9s70GWbCDcnf1jt3NpTwVEFpcH25sGbA8ktP34FdC+rXj1rAMqq/7K0ZPQqa/ttjRH3zFTgTcL5
+/TVMRTA4wfQtcu1gdPAWehpsOOzlt+FWAjW76nc8N8qltWTqiKHnC667N+xwCM+0hnypO/N5JNi
0+dAeahuNMxUoj9lxpngjjHmjHsnn3F47uWnMPUPrh5ODzDIrppBgbfqokWZVlm7nw+ES7CNzu19
EWivrXHO6SxMaTGve+X1l23B7nrfqjD54PUyHKmL4AOOyS1zCUkDkBEIcNrW8DW9q1Y6F4dSBUEs
NV2LTDq4Q/fiQQgEXAo7jhHAY4/PhHKLNttbp2ZCgF0OdBolpTI1unRfxt0BilK/jyewlGDoDS3O
zvXBQInx1OPvyQ42eVU2it9RlUMYf8huvxyHeVSMkTi2VmmMIgGw/vGA5VqYoIRnTXmm3bVD2i07
X+Ffn9rzuwH16gd0KOGYfheGV0rSBOXWbH6dO/EGC0fZ3/RfSOZxoO3GNu+4dmV3CwhkEoUz34wd
5PGFiSbJzdw2razCmD8K75MSn9a4ckftI4k9KL0AjQ5I/UtkWu7cKoXo9vYmzCkCdaLms1mjNoRz
mo8pgnFQ/yjFuxLPcbJmeCUIfjae46YE4JepLlIC5gA1ukyH1mSxJ9bFMcP1XObCHrRM3kqxnljX
djn2wUkw5Zkw38b4guohcc+xz4f7V3DhOoVBcBeSoWKvbsfFZIR1RM0NsMpcqfa0DF8lXDvQ99MX
Ehy/BkhpBbKI41xv/pGMoOTdaddHmywtaaFA5VUnKnYjQKzyIehPbHuUlp/iGwoyM5J8PSwlzdKo
ICRyypOLUbnZulqq8gjWUWhnM3fwPcf7Bg4oBv/XCStJTZmmpfBqRbaQx9dgOxEw7j1aXaPR2/mD
Ofp61nfz/58B7a3HJXbwMavIr7QEDPLyuPAmh/bejPa26TtPYTjI3YxfAXreDbzDwgwFwsXSS4L3
mKgNpXwWoHnespbv+L7cRPNnAsz3HxQzMyQxetBRXbf470SKKiYqTZG/6Rl+t+5/YGm8Y2QOGJOH
MCwy10gkFoyClL7zvXtYz26EZQQCKmLi4goxm6++eWgm4LgZf8NU+fFsSPGG1bnuuTlLDxm966np
33Zk0WOglPSVp7PIjM/GUHCcHwF+pjIPf+bRvxKdYnLQ6M+lvjSkuQSkPLXslCzBC0oXD8rSWMfa
m7ZqTLyodkwcciSnOO0F876nX0jEDuxCTp9c0tpNiwvSsD+SQ6KiT4QwKEElj8rpz+L9MOy3yU5Z
zfNj+H5T2UW36jydljTBSgUR9vSmbqqORvUxIfREL0AdDTNvkJMc3pSfIY3eL9vr23NaJhfO2WMd
hh6Q5QrIo6BdY88Avc2L9BJypc1TH+7qJakyljYIRYKFmtdCgpM8C7K02bKG1md0/3vaQabWtmYS
Wjqx+d23kxQrNWgPjKp6h8mtw62WewTZq28hgh98Y4SbHVvaqOva0OxLITQyM0cD2F2eGbfrpx1e
Gr5RXJTfjg1zGiHe/iMJrqlgAi0QA+eYeVVosq2FJlr5cpj5lm+L1t2Hjc3pAEzi1qOW5/O5jmPw
0X+eHEyw2ruDWWSNUoibBXpv4Pu2/SavK36d9xOmQ6UNrCv3K0BmNI7Bd4ciLMmoPHaZ57ynevkM
ipb+2+WJuBMUT1BZMs1HqO1CFmABOe+G90hvOO51M/jA0JsPl7rSNMvFT45e2VJFbB/GpH/mlb3Z
0iRuxl/ogiRIUJpQkFxmng2iiseX6Bk+IvMyUsB6megeVPtiB4yJs+VXGDIgC73ZrGBhCR6K8IDh
3XkEY7+eT8rR3njE140AwS6r+8wF38gT37Yt7Fvb2BCHZj69KTw+ixkcxeq2K1E1HwOHFGx7j6TV
sDWFloOUqoFdqJ8RKWQP8y4jMcmZSwb/+S4lumJpt87PhkQGe0Kz3Dp/043CTb8aWad7bwJaKZFx
mx6WCG1DyBBB9QJeINC3+MNEyDIweHE1dR0eLog1aFBips+4h/CS5rgFZ9TL/50bpDqF+PyFmpih
LWMaKQ5vsjJY8Pj5VfE2Yz2Gyshh5lYmrN4xYrE7ovvpQha/crLrM0mzqZp1uBEE3X8jAVjxlWyt
XsYguIAoCBFmn2DGJNS78GunmNyAAnAccqb13dmi+XUkFZ+nQoNswHtZvohMnmM4HNTmdhzOH4fv
ZhN/lZwUZ9v0mMsKmZJnBohFGiWoc+r2kEI/1bGnUQR2ZFKFjqjkM/5J+z2Uca95EJR8zsdMpZnN
UsSqPOhWNDVs4Gf5YnMmHrpbrjjI9yXsD5sKlOfBxDE5jRNRpji6s6QkqFMnjrPzwjhM41eQ1JWC
v5gPsijjbRPAk7I+ODRGlAc7lgx4LRVOdfbzlV90vXJl9EmOmWuyEl6+jqcaOkWkxtFWHU1QxXfY
9OfCRAtjaoCjSs2dUw5la4BAHF91v4JYxHqPDeE5rouRaZ/Eh4yFwKMUrm40UbRBfh8y7FIgkCAx
h9JGtT85E/IuwoFHHwPJpeRrohLoYP51C2i8tN9vv6Vm55+tELsKmnc/y8lgYl0y2YE4tTK1boQ6
5zX93pH+xU1Fjq7zPfTrBlmRzHVXL8PxxJXEUuajAPgdcmQEO5rfEV5Xfcr7BOO4oMpbUi2fI+L4
5LlLUBnHCi+Nn9bRIOJLl/LFCnozx4vqF9wXjP0xhBN1GeFg9RljgnwTMwjUg+Dw2tftjHzpkX4f
ShMWNRzZvvFAso4fA0bdJXYztYQZHnNxZ0EyL0nloed3rnSPWA4UeimVO0d0ZpR6oOvbUEl1zOw3
uhhl4H/1BFxgfCS8lqV7FbzZ6g5xNsC5c0SMV5mzDRlO7KbjLfb2zIefO3rX2Yw9eF16JzVnbu2K
/wsP3Nrn1i1kNUP27nkMgQmj/WY+wbutImXyBB1w848Oq9vp/f62oECVopRbJcGXQb1q/IflhOIh
pzk4DJCJzKvC/c3e5TmabaWkuJ9hN3uJDWNegWTTgTQT6mXuiZ3fMvQ/67XsQgl+YYuQ3DX2ibXh
68DUye2RoUm4C3yF6KEa6yWQUul0is1/cHHODAP1XyFCqizQtV0XMoaJsOlqKXx90AiNVP8BS6No
3YII0YpiSzO1V4hpHgTLYi6M7sKRFBnMZjc0APrnK6arATuPEFoeFlI8rGyviZguMScSRdlGlbPf
r2iacr+NrNMZ+GkdDRCQXMepssSK08rTW90vlGAZyXYwDhUUl8QFq/kXcJZxu3DdA07KXt/8kRCP
L1hnb6/+heJNuxWj1HKGARGmbc3TQLHCAymzxxYuH389B04/SVTFbO4e1KoOkgQcNVvvKiaUgxW/
tF/4bSX7V6CC4uHIrQu2CHbMPSqzIbyF5rJLiQ7z02HxJ22zhd7liKYaVCABKMfQM8s0uEbp162r
U6xcNLi6lBs4nYP0o2NNg84Uav38vvIyCrH7TACMfsL5mRcXe0/O5Uk7AjMEIWH5hcfNVrMQPn6s
AcbrilboMGU0rA3SMkc69XYlGTBZ1MvBKg+subbW1arAkamWvs6NDjLK0oDlX6MCZsR7D92eKpD2
cJ0TXUYeS735RyN1VeDJpgqKrnscfwuXfZkLE7Gf3Y6TzbcR2Rb3m6G6JxKfkYYImpCvLDicvsLC
NpGb/FXIQZas9KLHsDvkndjip/oyxv2+vNETYpN7H1jo3LnPm++TAiSviVJ6Q5xUbOc1kto+0r1n
k9xVw9ozyFc2nsUE3QZpEYVlTiduejcJ0UZ+lvtXMJB4ZwbCgZVEer5DFVw09OXKkYpuuV88BuLh
9/IJyqrMidNM6FaewaUpzCArtY7/lup6tl2oq35r8W+y9gxa1xM+DyZ3rNEWRbnENJpP4IVdAh8x
CrayXIAUbbLAcwvUBNvafsCsCq0SyyBFTmH1R+1ED5yU6PJn0GmCEEjo2NSiZ+bUhBKd0iuPKXK4
nysF6iYD02GMF4M/2/g5TKLYMqCvM7ZH9UCnqe2HljJm01ibKXd2TMPlzxZ9mZuPGgznAzlvJeED
lsvIYoZV2+Pp9NCS07482WGNEupeMjeGtYC5oqoF29/BGqoBebCPLpe2Nv9ec7UO3vpiET+8jHPm
rReHEi+mLniZ+mQwJthQqf9TXN1ZkrtrRu0OgF2ii93YL/B2QwGqpb9FfJGT+tjh+HqVTPvCLbiJ
/bpwCrc9b/sC1T2NmZcM+MVedxCZxQ9yMrTOzgp2hQpSpe1+czp+5j2GuoE2cDKlv+otKkUV1q5J
Ns6zY6Ia8jeM2RTsYD/WiHd8Bi+QpQcIC+X1B6f/morb6oy4Ypkejn6kpNf1BdQRXyTNeFa1xQAI
ykS5gRxYu1FajLQ8xiP+Tti+FaRQi/bz8YyF3YwnwGxKM7rIogiYX+jAGSrHKHKcbwhdzqXwQ0BF
hANZWnl1l2PuV+/M7KKefEQKU1AZ18QtM8XaizvBx+cYrmvCewhEuGvWYP0RKOZRb4VkTRSZv+SN
MnZnJEvUXE9g/8XHyD26IIbIx/aU+W13g1YJ0qWGkEtwAzp3Ot2lLDDBknIJizkuGtjcUYYYmpQn
FgvtelFgWE3Tthu64HZlKw+YKw4dZ6fRf05oySnJkr9mqXK7OcQC7kYOahg/aBms8Ob4QoayebQi
VTpTXmr7tyTAiF87m3qcaWXHQ9aYNIEV5nA7nA5I

`protect end_protected
