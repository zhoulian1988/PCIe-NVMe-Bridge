`protect begin_protected
`protect version=1
`protect encrypt_agent="FMSH Encrypt Tool"
`protect encrypt_agent_info="FMSH Encrypt Version 1.0"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2017_05", key_method="rsa"
`protect key_block
uTm1SZ4dKJPAnBnHbASeYedRkLqxxCvIJUmGFkZdFFIPIAAW/qTh9kdS46yxf8Q6yCW5H2/YEZsc
KEViJobEmg3wn6bCKqUg62pPOl4wICwykZ8Q2EPUKEOHDtsEhtQyS0Q6IKl5VR4nvMVonBiTXa2S
6IwInQpwPgPFfuboV0eXcC6OnOKjX/pEyCz7OVi1I6L3/N5nhyOoT2eSsRHR82ebCvG0L2L5NzI6
g3qyb2a9lk1cjjrc1e9dRNHqr9e3pcDYFP+uESgnO0qIvlusWe7XEtU6v0dyNgq+Jn1NPIdYWUpw
HZhsSdEazcOMnJ4q8dnHPC23duqxa5OU/3oCdQ==

`protect data_method="aes256-cbc"
`protect encoding=(enctype="base64", line_length=76, bytes=23056)
`protect data_block
mDWfYlDTBbLzoaf2lC2bKgMD+Tw8EHPw5Sm5NI22mznaJfXh0x+9c3pKghaFg9gYTc70myaO6Uj7
LUHgENRlJoPMgltJGxv+U/96+JxzGAo8/uac0BgTMAk1GS3LV2LJW67pVrElADlKaWRvVCGm/oCQ
ALRRmYspQ0IEc95gxlZN6sRrmBpGWjStVcjPZ5vbreBT5hF26IBHFAb2il3cuZRNG1aBhhSTDpmL
2T38RU60g7XjvluRFIrZ9Ey3r5GSo9dmsuDYv9+RlfiajRhKdXZ+W42Ke6TjBa+pCiU8zJZwk+Im
W5Qogyy3VP9VThIWHIAEqNUAS1wE1hItqVFRzqfcPNwzJ67laZ/+vXW4GglAi6qX540iFUsgEJSp
hnkAId+8CROD11M3CCH7UrBXLE8qxFC3IKyQ+tb19lznGOOWnpbH24kD1/5ulsQmFxi/pDZV4WWP
zzqxHT4vBFjtYiETuPxR44Yrmp3QXd6AC3LCMtrUD5xCIKZ/EgHSAvMnvRVoJyEMIzZSAE1KoNqk
ZYPG1Dt5M3l9Zn4UWX4P06Q5MUPXxPh8HgZ+iHnyyxp7xHXeCjTssuJvn1LnCYTYPx7tcKyDdLOZ
DYhdvT6/g4UAJv3idZ7eSKenGkdYupguPTjHklkMxxuCMqp9DAVkH0rv2CzF+N5IfgIW84fWW4ov
Ry0naZmE80UxCw5aR4zBDetGS/wBMjSO3SV252x1AgGV06pEcJ+AwGhAI7wuInecPf1pygKtKYh+
41qcL9Mpx/hKgWhu7SwS003xpaR6io5vIZoUd3VgAnsre+M8KwqbQPhA2af06FrEh3IusaRP5nxW
Xl+exZOD3mbBK8FlHYcuGlMjLDjUJUuFGcNbqBY9l14AkwF4frVZtIZG3TLZAbtCpAC7T2IlYRd/
7HsCRZy93Qn6j8Jg/Fyz809RDV+jE4+HcTsEewj1ar9JtVHT8mtruLeEKEj2upoDB4OTn3X248Rh
bveYbrcwTNcyyrrlu4iTnGTJukLfxnwPV2srT5uO+HNXqY/BEHOFNlC66MNIky3APGvy83XptaT3
XfsKLFnjU5+E4Af0oiuFyJJW0Opk20h6QhOyOdqDyc63PVI+acymfjd9ffXOMwj/4kDx2USKS8mj
1aDX+PbUQuWEuDwimxFxwM6QypkfYMUacH7hM7TJs8XtroaV7SQ/X/GeSmR200/D8eYS6Vo7X0b1
7mw4K72tYQSb9omhHTaN0YfMHbTDobfE52YOJrPLtsvvPgyY8cjv9PO5cZzfHBZ9rCX5Wvr51Ta8
kcKCL2VQt6QO1Ix0Xr/bxuy7cMoGgIaMBW80AHCJ+yt5246qkrDe/acBda0rWynH4ZDFwA9H+RWc
AnG1fSMBqx86nlg6HEtPZFEJZmehp57Dl3jVIYRJt3Tshg2VRx9K0CInfs/Vhv+G0fTRbVXGjoUl
a7agmyS7ygkt3KLZZCeq2trPjPXdt3ZTNQqIwFTInbE652ZG0oNf5OGvLGlLDEsslAhEMIjc8ypR
PNe0+hhYLXVo4/a3ITqenIJp+a/3R8GEi2vqked7LBcnCDl9nOWNsg3nhLMKsreBFvzsCgPdZ1JW
AhLZueCa+88mHe3cnvY+RQLDYXQVngrLOfpXpd5xfEFIirH6IlUvMEcFI7TA82+cxWPZB/bJNc0B
TAbim9O+O0KrKSfJh423G4P8sU0bcItlJdxndRz3c7UyoDXqbOy7Uac7A7aEIwDbf8KJDB7tQS/K
qLdNPhP0JHNG/pUa4HZUo9vPznhdTgTkSSptmH6frHxF970FcLaQMfYx0U+7QxDZVP8/XvVYzOCd
aGrsRgrPX/r05DHjbdlVRkOKtw5vqONDydC2D9ing99y60Dgxaa80UQWW2oHR/UX5iKbsckNPEcV
ljVD2n+cnW0iRxZ6yHVkp1MFyPNgPlK4u1MaWNz1F9Lvi9/ycWSvU8NoLviH+5bUX99bEz8OX9vp
ObAcd93JVuIcLNXclFDkxn1AaV494iqqSmHZU8Ym70PJe8Wr2aboJKa9TME26IVyYLpz9sAfufQE
MsOtTu9kUSjNuqv9j3afnTVRBS9qFvZfhAEBmBuMH5umTDPmUeetvXRE/w8k4ODdKq6iRMbW+qY4
oLDDeP3h5ZmE/l03npkun7U7bblzzsR5yb8vuAAolf07gUuHhQvcs2v9M+P3Xpg7JHcb3MVjc5PW
/7vQpYkeQEcgPvfIEb4qbJApaScCL2nBvIPBy31QqLY5ZriKKeHVjnTHeHtlXSYnYbxyFomcczYH
0FtERAB6McEFRubSA7ejKYVCp+wIwqdsVRS9GLu2vFJu4Ouu5sf2zfuCiGL0pa2VPE/VnRvoFgf9
fbsUFZkSVQki4FGJCDFsPtkC7G4kOdZKZT8ocjXIzr+gELZRKFc5w2LWkHTeFEYcn5WgYBVQ0lHd
4RjvxhoBPPkzVIXHo07KoAuy+zLZqixMXOju/MsIDj6bUZt4HYRX+xlJ2uei3PbTbvNPl8kyqeXn
AjcLPNarvm0A9Arp5wHpIE622BarSZJrKi8I4pIYMfm5hhXHJz4lZBTCahMP7lK0G0hgKvPbscqV
9Le43tFRBfO0p7RHOcCpGDDQVZMagdxTQPKu2YDS/qsuWc/AjIbAu/jZJBS1p8RHyxX4+sHacpMg
qCYJcuLDvjWXaEh98LBQNXToikjlYrqlkdsehcbxSUwH2wpWr9aLuqdb9ojhcw1fODNYLjTgKgAf
/Stjh2YeOHN8PMCMD4CR2aXAnyD6+XiHQU4FwboyJtOuaBfJrau0VGW85Ehcgq296ZSPb687Ek0b
0YJGhGZ4ZWYlEuhHXtr4AaHTUAlhlFmaQTtYnXcaC+y2KDxvikl+QF9URVQ0vaTd37v+Z4YuxObD
hICGWWMApbU/5Pv09E1B6iUKSDgLPNrFmBEJ/RKwMD8eydST3CSMKIHxAr/PY2ptEg//cE9mJT/S
xDTM1ucjoLBLBsSShW2p18W17gqG1uAMHUiJoYP94vYUfMnxA8uWADbTkxF5rKEW+UxUkR6LfKF4
NnH55hciSG9W3doUyI9oDSYnBC+9O1hW158WALOfow7TD5Al5+zdjq5dv1R5HseFR7A98sRm/jAG
FJjhdR9/IYUppYtg5lHm8+YWrr0lvU5adKi6lOWT32GHRQmTWtu7MIrFKTwNBRjWFPtsuAu7c6K3
sFF2PBq7w+fOMZQO3VxENHW/HNgJQ9J4OfLIk3ogp1E3kODjv3cZOnhiVHX+QS6zGWDfNvrFMHkv
LJYPYAyOOdxTYbnqEvbQUEPe+e4hga7KCnsfxzoHMqlqzL7dbeiR/ALeMVgVOrCx87h7NIENTfsA
N4aplO7czLSoSfcO7Vy+axK2tQ4vWlkMjpZVpY3ZGoq9TyQ1hcFxjPR4zbcVHEuC0jEMWKKKW3J8
Bphu7Dmh0RRZouDPT5ZFhOFAAg05BCEFRBcRhPDLbHnl8WpX/qxmzTBUJLEaWmfkwVw6BlNqnpyV
9FO7HBsGJjV4+EBajL6agh+AF5sS5VxrKxJy7A9Mek9lDJaLYsD76pkIf8dUIUgmRJ/GwA+pPB+U
4/JAA8suSif2uFxHsH3FxKdmJPUiV5VWqUFBjh8kAd/74tS4EXqC3g0msJdEbDZLAvNtBIP3YTtX
76S+5pKtRokHMN7UBcXMAACVsjqYs17EMbiQ800HQV/vOHgeEkbFMXspq9L2i8p3HrUmZtArExrU
Ve7sa//Us0mA7DW/0WR0J07kZdGUoPW+LPbeQjDPS+YRiKau6doncnKqQ+JUJDG1yWwXkJf3J+cs
9By1xVWHU2VLGSu4Snwe/O7k6gVRWoiDe3tRjPZdUhjcXvxVwmC1GaFlGj2+iRpKltKHApO9EBTC
3essHJ3scI7K/YYjxvj0PLrLkR7SK4e+oX7+MJqN/kPMAaWWqAShDW7KVR4cUB8OR7bKMQxw0F93
Py7wWJEO3KvhGbgESWsxeGLOtFeXCy8yIvRGvhsQHCgIRcERJKcDDwMch1N0jA7cT2NGYHO6SBkf
GV9g7gT8bWTlpUdnesm7KsuMIKdOyJnXG5u5GpJXE+sF2duYxz4w4sLDkAoKU00Pfm3suZnHmUMu
8oN65J7uPaYNOGt0eg7VpJnwcE+gKHaMw3IomgvBe57qe4VndBJrV/W6TlWUXws7pEUia4Nf1grj
Lgs+I6EsFIWUyPhkL7x+o7gj9vNRVpPAowhY2w/jep9bn3LQgmrio3bU5ws98XSSQxAUAUhrB+gY
br3E8iRV5ZWSfmIVfqDOBISmZhSn3Hk5wO3B5dO7Fx+xgGK+nrj4AQPUFFE6KBVjZooAmlz3dGpD
RnFUw+8W4MariEbna7NtFVugmcmnC4MJ9Tln+LX6oVsuXpyvx3vnDSdGr9AzE8xuGvFNqEwCW6cL
h+ScIudOht1R9FAEqX8QoX6MUE6igBt3HoAD6U55MCGMJ8N89grvGSyJDTP9CMXvlCbvBPphsh9y
1UxfAF5hO7ZhxC+YPK4vtdtN56mEvC9oj2N8tRjcPFnRWgtF+KQ5KY/QnfBvz+yAcUJeaZOKPnRB
HH+StTW33/tHCK3ibGzdm6agFK6N8BJTA+rSuOgmA3N4W5s3CxGGBglJ541IE5vkO2wZrpOrBbNf
jJyFjGqvckWz+iy5xFb124VMl4Y6JxvHovtwppae3OnnblfZBjfAsiylI4V0K+ZG+RCvkROMUlFx
NLXb+nXlj+9FSLAVwa6rImxbwvVBu5s+5valaW8xy14NY7l5lUrdfb8DNWBZD7Q5cm3MXmeaMsM4
LRufQ3ZhVeT0aXxlHgXk3+ZrZOIXUbl7YNv1aeqkoQxS46ZZT9b1wj08XVa4/61ajJXkMisuM0+5
HAzyki96g8FwQVduk1PYwCgAwnWtqrhhRJd7EQgAE4imgCUrSLqN2o1Yc0SSI3pyMpmBKd+a9dm9
cVQB6/4cuv5QGWFYG3aiAY83GHpwifL+84INhc8mPskNTPAEBpYwtSAR14FwdITnMOZcM5k9e3BK
PhHIOE9kybeXeAVQRUT4Xtydrg2ND8L73GF4ux77bWJKX58IT7YorWb89N28jKTpO2i4f2S+gktS
9JT5IiCtAGKzytv4w4aLqb1zHzISbrPNIOeZakwAesth4puDEHVlJ/TyR13o2wMKFDE1JOCT/QyH
MRSFzpzUvOLWb8PVbYvhpusGbPdELBz7L1qtc6vTRVL1moUoKnTUWHj1bHqoo5Vwe3pUc5WcTUH/
m75mY2CzjeZIa45CZMHJmBIIy8URSK30DIZxpGG+ItpbnwFmRj6ow6oS+VtY24k2QsICMcvTR3Pe
IcSk2/HhSWBPzKJ6HxvZbPv6zZqWnYZoZmRqjeS7V3JsNwuSo5cUgzO/B3JIm8kd62hzjGWDShp+
VlXHF0gbSR/sxB+6/7DQh9Kh7+v1rYVbQk/KM9KKYzuu54knt54kSiZCKIIUjRhzPpEKhI8DuS6Q
t890EoqSg5Pfu4Vs5HMKt2yr8IKVMpZvkNN37vg+33/TDGCH4eAouWJGv8YEi0+ttLz2OLwtqo0y
S7U+8hrzFPrgLdV9Fj8yzpcW6Fxs+6xafmjLTYr2k4GRm8RaDaO+/5r1ZPeEoFla7Y7bDmtHVd2w
XIoJOkbfnEsWLKYiwnjwdjtBbDNXnVPz3S3Hh1rydPhmvlcZyvDP3OwrrYHlqw39gGSYw3NwRv8P
GCpere0hnKK0b6xrGR0Y4UD+a1lnShbH+nz3uXkk9y7plepNHMODVEl2L4u24URNsWKgKx3/wbWb
PqnNmQSIpxysWcX0Sb3oU+iDvWyt3wX+9gh12InhGq7EBpjTAKsCBE0eI1epBbmScSbHsLgLi7q8
4nYL4RaSEVWUDrn6IAJo+tC1R+6HS7GAPXFG+4t3kWg3qmKsIy7T7ZZxtd+x/rkzxOQ5svL11P7N
mtgoAHTJtqf9Gsdo3wjLwSNqu38rDjuHoPU7NxK22SEiEwA1/p2uNQJY7BQMg1c6ymOOQ/bJpOqm
pr3yUqQxINOhrcunD0yGFv+QWNVhxHFuO3qbucMBb5BlwaCROliy7gzx1e1ZPX2nYy38W5kYW9Gf
rapPOv0MPKV5SBz/IcuuMVEmr3tBHflgR3q1w/imCCf3YlFJJAxVSL4k834hWSYyxfKlf05RuXgy
A6CylMod915yg3ypq8VwAuxLekFdC6YGEnO8O/nF4jrA474sIRmqC5hSNY35cN9qipkhSsw6wuJS
cYReOg9NVy7XXl4pKUd8Q2sdimvYjOIm3+Rq5BZinjA8ozY77XZeLFEdXCSi6GJdg+rZ5C2bSdWa
+owhRSTshOWBMWeC/mGMEGkF0a4LdEB/8h6AhdqH4zNJ2JZaWgtTTFHVzzvaTvY1CXb2ee2D1sgc
EOd7ChC21GL21SCy067Z/SPFyC6IPFZmI6jKfaDU9IYmjHiFuM6aA+jZmjC3JZQdFg5ImE7ipGel
m3nqBUq7FBsN0zaF0/OzpN1c+oM5Zbq4Q40JBqVs5KOB6vtuJ7JxCdBNy7s53QJ09YvySz3f1Jwq
p0p4r2yvBF5AAOEh1W0f33i3DV6UEDY0GIK5s/V6S7Sc8YTLPZ5siRl/M7SZS2A4KL2RDtML1O4Q
CLyP+G4aHLRHvNZT8zjPR6RHMjFyI2OrrYoi7we1EL4851dYZ/ra/ziq+Vlk7k6PfMaReDXwyQzV
pMiqSLykWNi2VSy1lrYlY1c3hOqHBt7haYispaAtWHdMJ6DR8Nd3iyfMEZowW7PQXh9fBOIVN5E/
R/E6b8xVC5qOtpYwffU4X84sUyU9GM+2N1Y3iwMtrUHWYGEVHqUKx0koVHH4EDJZEE0nReGnPTsG
qC2B9O+tldFcctcNHA0UAO0DOCcMElrSWrao6eb7UHffTJD3lAfhfyPSP3i092oFUuOqeu8iksnX
bTHqWgOT/SOTg1zzQZuD2Bp0SiNbtOcYqfW2lRXjQzqphf2EtnfQZgk9c3uEX2loVzmjoPYQfuGK
RqpQZMc5Bd5kuX8Ap5TIJBWYa/4vewKq2mF09KehfqAYJB08NXZ44zRslhr+M7RiQw1RkXLxo7ic
GlsAL5zxq4aRukDHei6OdJqFKb9zpcQzYXU0ElifXw1YZfApTsRuV5clJAy5eeNzUjYJZ+XBc5pI
5b/+HAECT2ABHqoQj4DaCzmouLAjD9PXhxvJ0r9T+LtgmTLqFFY5uMCaguOXjuSSL7MNEKlwIRUM
tXamrXkZqbmjruUdQMyhEpx/trsLKQt5He8aBQaZJfmSisb7L/UuneRgwh/xvwbcaTI2/sL8NqiF
L6+SjzGkQRXTmKrW4iBGmJKXuZEWWGLBvRK8v5TZ9FmPbNe3zMtaoXvwMRBDcJsAFVPoClWpJLF5
Dsr6bAeojGykRu3ShVtTta+mUOOkmvBAcWxWhcnkSZs1q+XkB62kUZQmYWXFgpBqjMX9upwER3mJ
znmdpcppBjOO5uerinX6dRF04DVL3J5Ju5o2nUzyial7U3dhaubsvc/z6F1oi4f0ai5f2WwXQyFS
8F2qImvKhHHUzAamrpgHf8m2txRyxfhB4cglP7BvrFZeW4mKaeZI/ZxMNggQ2wCVCQoOsFI06NBl
Gzh2g031MPQwxMWSIXNgApPHR804s0TcZ+Wvry9INCvBE9J2xEUP59etZQWKdldKnzbttVJQHlOI
gOeLLLIiSQzKNAZ05m9InvJSlyE3VEZb0ZNM52uhBG99JIQp2UVEWnwt10n10eSySFIjebrS0s5p
3VJp0hUcyIR+6pdxFUR67pwh9LyFBL4JYRh/fL4LoMhGPVwQ5abxMT2ueu4p83PoSlN0w5l2l4hg
nD+JIVZ49Hq3VHBtJsij8oe6yKignHMcW60rGHqIg+MRE9qdmOoKY0i+FAfPRe9B+gWDfPruUlV1
8Jku8f7OqKCuOAu3bmqqRVyur6C1Mj63vdxrwVlV4BOYeXOvxB+REdZQBcbkhbB2SK8VkbYejqUH
adHX0MoPhG4EpZnYjSyYL6HT+PiGXYLmnisOoacbGmu6vcXlo5TbxgtB/DqD8HsiVKGo+YNg+7gx
oDqFNLRFYy8KsuLjg1l6FvH2ir7CLruqmeIZNNeI0MMh2cnazE6c7oO2uhsgysJ3RxNW+1hPPour
+OuNzDK+3QC8Yqo87XXVMTnjokzLil6bvCJDNikcuI6/MXWlW2Jbpz3DwBQSvlfZykyoaO5WLjjk
YT85iPcQFuU8ykqXtyU/fdB+mqp4T2HA5w2a2dahqqJzXdKiV5EUV76LLa4ZTe8m5bQ7SI7GbpxE
HNxU+7AM65pkZcWSsPSBL8zrP9MS/bxjYuw+9oRvXKfzQ+Wy8K6D6/oWZlkdNukNvci4GXFRpybo
2UxQYzgkYnjezgIOw1DyXPMNI+eaLgQ5muqWehbrOA7fTr6fiD9cjZxqNadR+Vb4nIv+4tEVj2+H
xUrBp/Mp9bASdZr+CKD5PEagH1s/t4lZspz67SAn+sUBn4HrdFiLEMkcRd7ViI75hDiq3MmfyM+J
mUBrbh6u5/IvHcF3LlXWcs20e0TH5WHSEKsvZejSzNYGzd0vOrasQ1+T0SIRQaypgiuCXCtO+X4T
aEGLDC0w0YHEPm9OiMW+1/onvImp3E7iI8H+PIB59OENoHeXmKOIFZ9pujald6u/p1gmXKcB7T4/
suZ4FAZjkF10/LkNcKJv3YUMq6/B01FzebKcb5gP7IDuS2LXCqrahwWLBFD9xHrYMgJCm5aqBvtJ
B+ncEKyWD1FCT3I2gL+vPY65NVifPAYvYwrj34zeZsWGH2BjhQucJ4lGaiD1jj1hw1cd2OXRlnFb
cC8Sv7rHQxyh7MRuHn/Zh/aVUugRdGKcJM3kEygO+vD3KYc4i3Zc9yU4VsZ9IXB8+XiNB5pRFbQ+
i8JrJO8om1iTPAhoWnCnuYk+bEcG8tfCkeSqkZ9wlw8P9wQh7HOL1O2uFHZAdLmjN6skoO45ntb6
1/9B3cAjkdJulKNaCEX+mYpy6/cVsDnEE4SM4ZFtvWAZrBv/wjWE45rVcfdQJELW/LbythLdV+QV
mMN/zFOLCPr3bfylFsZnooGTiXiHYwq6JPd7ldw1hbwxZqad33kbSxseGxafj8EN5yQv14pjM3dY
5Tv/tKk7BJhwy7bm2WUUNXBvCoWR2ug8DuKQ1XzwKj/MYq/F/0YoWb7T9hORrE3fjDoVQjP5gDU2
Acf7Fp+VJ9CsmBAWj2liaM6R7W+NENYAt7bLUF4PADfGpp9Bonzb17cB2K6wz/h+nxqHe2JnPzx4
KoCkY4ckoqs+e/FsttrUixDX4ryaPLjAQqB+6Agf9mmvniZroMA4KA+8iOfSBmyLO9Lm4aXWCvYy
zpQLMHWLn0uLsCPt1F8xM9/HnnggX4jKLjN4QjW65W9Jpuu0AAWSNLIrIY+BwMQos/AVuux1b4Ci
Cv9ltufqlKAgeI86TPUuMiYa5qOQU+HSrOX6PoS8hG5jRXHe6i/M5/khO3G1Xh74qU/Z86dkMtNI
phUby60wxqqjonb6mzNfFj2+daP/C/stJy5TQilnG1AJIM75bu1KtO0pXRDvmwWwhO/neK0xrQun
It3EXTR9UqOC46RuBQwE2y2/EykSuBnpJ16NzE1o5rhkc3Ob5rtw+kWpfbiRC35+kttwv1/WumJv
BCb+eiNEcb5JQbruMnYOkbwJoYmgj8TnZJlDnWvt9/5by1pqrWUVlOAV/Gw9HPxbHeq8Imcr2Vjm
WmVqv/t3bRWsAxA5KBP8PjtoqgmV/TItpypGzkDP3BVgSEeDYXyCKlVMg/C6fiShEbuUoFn4o0/Q
dvCIwjAwX/6PlQlBSmTpUfrSmHRfGn7ppShhFUAGo1lrmfPsa8KffjNDkVPgP2XskUlrFDSL1rD2
Oe0e6mupFrREHu666QT7lVDh3DXFsM3mdRQ6aQ+q3CrH6425V7SI0MfNmQ8x8vnWCWQ6rocM/Ljd
PdXzcdbykqXJMfN7nOwMgX1R5zLxJG5bNS5u03KBcfaGLiSoJh1iFMgSc4bZE6gLKAlw7U7YQmqO
uxWzSwcMM3UATzEHch1vKSx55YZiGMBU1qjrbEFNsN0DUfIzBfB/vMxKAaZAw+MUFxV55MPpklvW
WqJX4ahD2diUrM/AfrhgvrKMbXGGM0ygSK+x7Z029XgIlA51w0ny2ze4Ymap+XKRzv/a0b2VnKnb
LFjvx9Z4Hd+kE3YUVHOHz1nZkYvXZOzqqJncPvQIZ71g+sNEhIuMEM2YTof4uytamxhXa6TlHesw
NpObLwWldmHhvHVqidYwB5dcwjyTmbInWYvGlVr0xmOX58i1UJes8w+5gAFXklM5gsVl+lXtNdzM
L97Fwf/mDVZhsVuhBb+S06TtZM9TcvBd62s46gwHIPzZwtXkIx39azx/bwmHQXplwbMUGch/9cfm
DZYZ1oJfCPFGMKclEO+In2mm3ipNyKwHDktmfYA/wM3a8IF6El4Zt9OZU3OWLXXSmP48bD0f4e8r
NkKinFH3Oaf9+qvkP9KJlR3N4GQFZiIa7CQX8x5D5Pht/w74dzBzBAsSV9KQcd7GnQRzOeaIjtQK
F418Dm4KT2YO2ZiX+2Yt1tz08345Bv8sS/+DyxiObRR116w6qHYusnKLhc44oj7phSa/gwZlL7nk
H3wAab3Ss0X5rvqh3G+MgqW5K3joJNMAUkio7noBamGj3on/PeoqwGr3j2Mw+Y96uQ7Gf5A/MDOh
O7KUCnx0X1TYG90t174EMukOYp4KIyt17KJ8jDcXzP60ygX+Fd+PYvxb8oDvj2b/ZQUbPp0LS368
MVniTBVwjajsHRw+wGt2/3xUa+6IkwTB/sKrVVpBE6jaWyZf3LsgQp09hTx1b92hDPgejHyJdN/+
e3meC7O5krCMzePDGatZNarpEHkHfFaTc1A/7SVxjarDWi/oAhaU2ToPFOVaDPayrbYGTFfNIgjc
NnkCYWcwFL5CWQLJy4M1f+VNSYL249rRC8PkJGWGB8Ww52TmsLhazQDH3EBNMuu7xzyBcGMxYcoj
GnVvzUcusdggZGxa8sXXPVmaEua3qsnOt6y4zXdU7rMFc1tF7zNsBEECspKwFcHJiThQ3hoGiJLM
/3QzJIM3VU64AsFSz4oSS59ZN+C93Hole4mRnBb7fUtsnMpp6FNF9ZxLUGlnQ2X3nV1f1tSRcbpr
hFxh/oDfUzUrG5G+9zzwkqDiXy3RHKtcYj22qSAI8XAyztu+tYBI+hYeekV556x8WcijVCXJAuBQ
0zEkle0KTBfwcsnsqZYzSQpVnlOWsNmrRKln1LvYOazN/ohAid1WaWnyXOXL05/XgA0neqMwSg1Y
V/aY8b+phBR243t/JL6w/YHMMpNouV5EAVlxt3f7PtqgsHRoEeIDOOWA/0wDLSuWINJRhmRu7h1z
q2JNCVMRHS3GzVZkkzkET/zc30/j05YJp8u82lYGBR5DCSZH4MBN/kIakPzmYe2Q3Rqa+8kyO5P7
o1jeNqW+srxcE84/xSx4VQLp05MSH011lnKjS7t1EdymHR0GviDxRAp71k8sRh423Hi6xDMwdlYC
xrmdKqxkPryGpy5YNIbngVpG9akk5ChYP292HR8w0dWcvoqtyp9ohJ0TThScgEHeXxEJN3WBaBAl
78QZYgFjUSJcicweo2p+jXHNzuJlqceHQobR8rF6mKYAeOWzMA/PJrCSGY07tt9V79AVaDrxnMJf
6794Piy4owTlziFN8x3U83UsVZJQQh50r/ItIWJ8mAzEkxI+v84UoVScW6ZME9FdrabjwqMU8Hbl
8r/imu9gg1qnYyD6pDpew0EtaMTF3NiHgd/YdoE1mwhv+9a/NvldZ0IMObyt5byXZz4ghomY4H0g
NXQRMWNPiqu/yW+f3kwo57gQdO6cB35JldIWnskSqTHWTjoe+8gSkR+kaHk57CUnvnS/uBnfEIK+
Z/5y40FaH7Pl+78MeHAYqJYGK5AwT7PSw4Yn4lWJ0JdXdXHAvRVkw9uKFuvMiiLuIJlIoOCvPooC
aBG1l0F7xsEVtDs5iT9dP7pn0QNqsO14zP27JvmiVsp9vRw7fIjeZ++4A3qqvCXcjlF8qjNzlpGb
6cXmVnXuxLPuUNBICbMSWuW7sXKUcWtnYweVv305i9i5o9akWNn/Jxn9/dFp7IyZHDCdc1NlhJBR
Cfik6yhq5pW5XK0o4Ixxu8wTBBdrwktE3/eBuemItyn2ZUEs2Y+2HIyspV9fe6nUmI78INVdrrzc
zzGMnUQpVLHTfqMGb2OcBnpPMv+tkQj3BYjUSCgkov0lolqAf1topV0DFzjtpHm1A72BeXwwiMxM
EMTnkPUwIAIXEzuA3Q0hng9Nhn5F7Hyo54fCwqIdTuPw6go2nYQkMwr1SllNiXgtV/HYDj2ULt9q
wG3ZkNVZbg/hMbQOKNnsq+ZZPvxXEo9uALHMMiPcP8qg2wnWKU4ufv7igAwJvs780fAKPP8FhgWh
dzq0IdGO6kORqC2JePALBHp74eGu68CpLKKYjydw2tnBAnzjlEl6Beqixk0jpmMa6tw5l0+Fkm5j
zJTg3ia6OcXVd+HGOP6YDnr6Y5RmibhQuPjOI1ZXgUCyYIcjRv0AkXtx8blxDlpm/NMUha1mYFHH
39byhq6vOj//wd6YxBR0Hh8jFQusRNUvxE15POWlAWGgJ8tHljd2bMzhd+t1aK4yz3wjiePamnTN
KV4ieReMTYGC4c0NAkz73kLvMyGyAwl7F31azuob3hTgCEEKghsRCM3yNJG85sIhMpflYEH48I7R
8UDbVvYqSQIuvJJjg3wBIVNA/jvIj8KufuPK/UIF0u+tB2lRy5GyUcndhJUEaLGwyRXG2VA7z5/i
oCBMbJvYIGsXHCViSCJaC0crGMtnoDMy5BGAZeiPiTWTiw0DpWU0dvEHJU8QyrI8NhHAA1q3HnXf
T+OW80tblvUzx4iHeRbZgEf8rqRFWmcohpuyxN2zRdl3nZG/CF+lqfCqajl+mkx5hb+3GzDKFI7Y
qyaBAPdHLodCuvcHPif272UA/ljjREnbs14xCBDFz5q30LecF+wSR3wVDt7tiVi3Ybz48Skofhv0
fmz9qKUfHwEiWS/S8qdAVZQ8pRyV3n3MyR5Y0/O2/JLqi+wccDRxs9wTRB9B/uwkYDK1A5VrqOrd
F2Y6IIDGB8POxazRnSQJisjn43xrzK/Y5cpYWTV69WDkYpMMdwVdrpvYMzYsKczPxc6NiYtANp39
nksjwT4qIoRlQACtcNnC/WvH5gwKpq7KrMxfMl9ZYapRNwhLoF9n2FYNzXrdE6GzRg6Lg8CZ6n8e
UC8UVzm7kDth2+R4Iag+VWZ14mbDci/SEAHvFzhEHLBvMxhKRgtDZ4QeQkKfh9wpHEzgtQPGBsSe
N5MnweGzYf4z6Ve8k4c6c/CJWOhgEv5Drhm9Z+lN9E8LVjj3jd3iTcLWx/+T+Mgsz7tvmoVt8Z5K
7RhrV8BFZz1JJ3u0S8YasKIQimkgBO0/nqTDXK7l1wEjfSAYTPGuNpuTc9mZq6DjwfQ7m0Y1WNqP
BkR/GAjLC6802E1fUKDgvquXnTIXfBOieHJsNoDXaaXHRRVjrQCp5bQjeL3iXgEMfnBX7WHNEtNY
Hw3idZ1ENZs4wYsk6dy25UrnuMpfnmKhWKenyGMzX76qI23qmPoUJRZeuOhkv5QPw6KNx8Vs7m8/
Cy9DHG57r/htwBsNmLx0D7O6TE4SilY8KDBU3G5hV58EuWFT2bcsSaw9f3ZDleWlgxaKHsD7vL63
UOYp9s2eb4AL4qkg44Il2vTUhLFEefyHKmjkBtevLo+SfT7lp/WaAJi8xyjUSvjSzBnN6gUE2+bx
Sx20BEDto6e6QcWA36O69qVIRBBOhyBsbPeNFMfYcGy+687CpGvMeX37sP5xKrNtfShmNn5Kjjt9
LNBMH+BfUSKO8r/fZF1RJp6/JqVGLCYoCjYFWxsaxNaMA1mjE/KgSkJ2aJMdEMdcUYJmq2JGUwhj
OGCDg+gRNtZF3e3kKlCm6wpkimuYlRTiaRKJgp3+mSy4XiWjuZsI5uPtkPTzaatylj0xtuTQ7dhd
Zo+z2rmw8FnEQqzM8MGxFKQbKIbi0zGOtszR/SLEa1p7EfQJIDo4enPMZFacbOCWbSjaMnWFAfmj
NByMIF6GBGokzBrYsn6BOqWeOcVCydufSoDb/gdL+uNU0e1tbxDuwMP8HeRNfIHmGwAffPtmhQfm
PzFfNwSvw2brC2FpMYN0ch4BAPKlmGmua88wEkiEoPkQL97SvjgZlo1KNJDEPqfCyCXSlPE1pTcg
koz9T+kjI98mHqqGGcklmCTiQ743UDeTqQD5Kb2S5ho96KAx2NMajzPqGIl+S/ZYodX32TP7VJMm
UnwW94isgHZoZ4MPX9SHMGcgZUbAx9LM2Ke/Re7PXlTSttAbhmYb0h2SAOUkNIQ7tj4rPPOm7QS4
npzUeMr3IZiC1uEJ/mIkZKE0P5o6oRn32PaWOR1QErRKtGHHnAn9b4KJzYiYBvGvEqWcu9TRJwbJ
mro/C5eI5LZ2woZe865Frd+QyYu7/qn5lxdc7VmnugM/N3CWAOOAXNsLazVvVaCanpCcmOOYbjmV
e5RaiJ9BvzzamAhpwECMUAcQsDwVO8bgZgh0utphYlYcLlw0UriLtdA4M+mbs65+2L/guxmuAVAl
LCjihktjDnviOqQOCQylrEFVrNPiAT32Lz18/ZqHPi0Cp7Pg/k21LIsidx0h0MYXcOBsjmdT/w9Q
eaBFV5hAhhN27CDWzkkTLaiCtyy8xZeT/7vgh7SenmyMp8eOJXmLCRg4kc+B5uxpDX9XcMS1zbuy
HynqF8I/Pbr/5oN/s/8JNuCABXtWAKjcBthU+u6HNHN+0hQdrnVkbzsKAMFdllbLYlgbwwqHe6F3
AIAMU7yd9V2qd+7ZtqsoDdvX9zyf2h++pt2uaG7S7s39twM1OPdjRCT0RjHghsVrMquxqYafbayS
hz8EukE6m3NoGMTN4HI5zWnbBeTsPwh75owH1QD25WxEXTp2Hofw9/TNFE0Iqq8arXMHReO09m71
Y6F4d+h/YLHPxFQZtu3MC8EVHo5FU33UewYGfmAD4rx/wmJ+gn+cdCJVAvByApL5i5HpLHrIBLUl
5pTcjNI+3a1kWZHlD9BALHBewFVW+IvxJ8CbMB6sbcPNd1WLL5jlM8tFeucd+vXVoj6RPoqdrbQt
YEuLB5oya/hjkBMNjY8prXbkSJKe5JPfmFGmhcZKokqtHytXMgb/V95lCMW/sEkJWyhwi8MhkuZj
vDuCg5hs5AGeazmYK5YWV7Dskd11gxTL1h62EOU2QerBPZ4Ngh29vR9UVuAy+P6+vqoNI1/7hSSy
La6TLdLlXbVJ3k7zQDUKl8cNDw72yyUAW3rv2JVfMM9K8xvVjWVgTIuOO8CSvpzPF/I8VtxA1CUU
+YhhHwvo5zAygcuwCUJXKfgVEpjzfIowu5BUmDhWtHLRgliTfhk8ybmnBXHc+bfgJkdBGJ9yFou4
+mxhSWy509eMNAlzu/wxxUDJZb0hV+6o7KvlEE2KYslUojtc81pKZFNGdNL6suzubr/IV9xH/Q2H
ILmSbZ+mW9+1TABmNR9ZTw0IabXVIxA6eLaho8mMBbpyXy/dTgvBAsiX/uomsphL1KLKdZs0CmnK
yAr3CMATTZaCkP488bgEcGS2BaQp2WA69Hv9YMBXP55E1djabhAUJ814Tsl4FCppOwt6RnU5sNES
O5bqFlEnJvEpCYySRzv1dKnpd81sTwI8tM+djZv7BmEJ+Zi85EuUqZgcO0iztuzgloANj7kABJO5
10w7MqflcmegggHwSRmNPqH6U5/Uo3qpIwOGnH6z8CxBOPMSsR8Iwli7Tgm9Gu7hUBE+i8ygQDw4
zfBpDvaGe2k1IU/vBqT+98p+3A0IOZ+GjxXIDoUYjfX2tLMeoz6Cl60NxJ8EUThNtH4636rBCUq/
ZrKxd5ZTZDEFddlH17mluvcugVBzfHNr83oSnZ42+RDvC2pRgG8PdQisLuT3o4dSEDeYP9YRQ8rK
JdA87/uNWciYBuwe/CFeS+r3AwqcBpcIoYpAnNoT4f7BWWJb84S0mM/oUv68YRr4rDo71LT5OCHe
JHEgbE6EUcLClOz2TACU0OiwaUOvjYskSPY7v6FPnx99BBFdTU9ukdUmBBcBQTzMm2spP6sD0yjM
ER3ES9wwFH39/oGrA6wLGiv5XqoPF2Brzzb+ORfg0rqkdAnoi9nozLDyojZum03+N1XI/9Wrm8Od
9DRWsReBQOtpHamc3PhDNjZx8rlSXbHi3DRVBd0uZ/uzpmoE7+AYgI3qHzZGzVc4fqR6SjYtvquE
TrFx4UxVZyKIXjq8erC5ZBL/P5r1SCRjReTTrhccmbs4ooi1WibGRSUSrpLfRyCk1T5guaS4olZZ
VPyZj+BJWgdQi+tYsGPrHk/Cibf8qveNhwmwsSJd3+4y0g1NPuPVguRvpfz1gPjhwZ/mbt8Q6UMJ
RBjOK7qv6Q6SwdpFxHGqAz5Y8AguBQUpqg1qn4cxikzAcWz1XtWBIfO4q+omzu6A0nkmx6qsiCbl
rC3fJXr02oyU1XBe2jphJ/kKKAuQDDht4wtkYtUBqMCDD+9TdLMkp3SmImQtfDQZmhlfrAcgTotH
t7xVSTF+NbbhjdVB0Q3OlyNJaimDyqBADvECUI0xEDzgcBfzqo0nVVHrGUHL2Gq58qNjfG4+cKHY
Gt4iMoS6NEt/4FqvUIjhjXYfboT16uheMk/P//ybGzAnwuzS4z/VteqeexNbIqZT1aNFWhtK6tCF
vFl4gBAtz0uAWMH2Vt6HTdbyr5tAL3iJ4RP1Ymy1br0v00m6BaPlLCRj6h0JMYm/l00TOVAkgC/a
1ozbS5hlWhiq90NJ0GCFlj+orRkP/gEGEbEnt3kaU9zcrXKovpIy0X1V2vb6VGi1ioNSdTvGqNBT
t2AdCt5i0d9MKpV0sIAjJiXtA1BHW4Gjm7N75DHQ4Xe39xP+AS5poz1K6O5Sgbltrx6Lth5N+AWu
xFQIrdkkXYl929ntBxKjs90cGu2Cwuvgt/Vt4x8/4NZ+KIzJlA9r0iOpdeU7nMpnZ52WaDdKyq+8
gpkZBqth7UKKx8+F1yJ0wMvoFvIvRdwKQoIyLcXGHxylRnWuhmTZ/HCXhYYnrHSjlsd+0fRz1EIZ
4VuIzI+C4QrLMgCI6THoYikQgikB6sIzFqo+qPiT/S8S+AUdcyJ1YeGEhHn1rxv3SepkyFCNDu7N
XEte7i1NgV8rrswk8oNL8O7xGEl7SsSkbmtRqz+IMQPZKhOjmOLmi10BzifqRI4PDFysN2y8/IRs
6gmbEhARgb6B+2YMKKtcEfd8+emY528z5jAk8flfxkvGJAlfW69x2LMLV+alqt28CTE6OSi0Ubub
u6/JkCQrcKrhrFOgT83PrZL22/EvYWNaWppyWlnxVyMXV1W9rvb7Kxtt3hWwDAFg6v7TZ2eZ4sbo
IeFdK/oyUeEeGpyTQtlaIen9+iB9szAyBW5AmSsRR8QFlYGjQ5nlha/UYhe5C6myyaaeE0JuKBNm
MMQLlGAzNJ0eUFnZe/COwceJM2qCkC9oz0TiAYtmTQUSPeuAs624uklZOGA7kLf52kBiXKPpsQuB
ayjih1Vekqv1xZ/FQUcsNfkJpYvJkpNhPeQhYJmt9hkbrH+8fX4uEvRN6GXwsrJUuFW0u5RpfHh0
Ldyu5TVefTJJGn4zh8XUScCRSk5mMmUcWzNzcIbgjzVr08LeCwBTvtbb0kn3HkujJYK6rZBHUxBp
w0wjHvzL65XYcbSzgupbEmmHu3CDfBoDT89YldDVeH9RBKDjxe+0Kwjamn0CR+bNa7z7a38kazeM
zXXjwDFGrjeZP7oi8dt8cL91XsNdNGoWMM9suztWkqEbsUtZyMyUNX2C/k6Zm0FD71LvzPslqrHd
LbeFTo7viWZnRhUjtt9NBkTppOg8LqlILtb6JZsaFzV/IIEctgAptaFzbYZcKQZH685CxNej+oqo
WjnDB5HzVTVk6giZ23h2//QjlNB+546bwg1Txi9pcI466pVsC6yYy/7TofFzDBq3lI6duSpokx8u
scrAB3/PEwF8jdxMNtQ+okjbNRjqQtMLLSYOILq3+X8hQ/FD3FFz1VzOxSo12Gf82z+k3QRjXqOO
ZE25Io7HDhOsULl0YrL48XB2pd2szIqrDjpmm/UYVEP5fSYBOPnfLGxiDPS5Jo/laqczVWCuwOqm
R794QarXdNm7XIq5xtWbCJkYMykse2E8dnkInNsaycFTpaUpE92OnqcHJBtthsgvoIJKNfEl3nP/
vKJpM9PowOj0xxbhsfprIsfscPOkfBb0vvddlqs+NTnrQLDwmDCa29cgQM2yUE7MqaAVqXQnUTG8
urpihPjaVfUo8vaDKkZ0TvfsUD2njAhilgOWq9ejATDs2o/YE7fO3DRkcfKU33qcxvsiPHxKCRH7
WDHd5pYk4MaLO/6w+s5Sc6FQfcrjOvuQAa08mT9VCn71OI0t9z0ickifvtulXLye/ubM6FuoMZvn
X2aeG5xSKGmFuSzvHQ+L0GdzhTsE6rw/l1CcPce8EQ7yhjdknKPnTVHq8rbdzdvia4jVeya9yjW8
FZW8QiAl9O6k7Z1SrgjEsXOYzafdhTmvQ/lBFE2IHFVnNso4AmKuwO6XkcJiZnJ/jIJvyDrh0JI9
1zZLX9ZAds7Wa1QhR+YrwFjPwVUk/pZi6HagKD/ZpaIBRLJ8DVKJqpwgn5TihTz/okt/+skNQKtL
tI6rovnp+aKxn33TUEqDJPQKLGgJZp8+TK7K81qIGYdc0hlh89HYT1ze8szC7nXn+aR68zWJgkAA
jLMMOCX9Cf71niTj3rM1kK4Bzic/yLmynNxPG0POM94MaGyMYSerf+clFZKh6+3Jc26SnpPSxWsp
4jXmH3P+VyZT6MxCOSjC5FSxzbIhWE9hd4Pf7D6FX6BDoXA5hRKEWjXK174iGDPktt4z2eGBBZNt
Ay1k8UzSB1lngCOQIuxvN2UZul270wDQEtltrW/ktbsFOdHdMbvTrp8eRnkNDw+Z6/Alnw/mv3pH
CPN1SN2Cq2/XtlUQhFA6/HVNZAO9/cqDhKA0K/ldk8FKAAbnnOarfaWYbD4Rw4l1StFLmrM2gPns
dOZ15CxFWe3jlsmnHslnQ5c3T+VkLDkCBNt3e1CWfJe+YXFboVnGDzLedNbsHf9SjtLfUe/NbcXt
0RpYMKwdOAfDDHT2wv75ulQbArw/tMF2YBjT9ao+jJ9QsBTXtu4KHTMhU4Y1XwzD0zr8GEO1zjWh
KgoOCHEx9e8Rd/8EdMa4zrJ05hvwhmvKgE2Me8lVaKDTjm1RtpiRwOZiNlCmuIB37rgqmFHDzzUf
4o0EGzuGpfj3qUKKHgu2o9yhCGvordn9nLH31Gt12Yc2wouptwBsgpre4LpxgM8skW7PcHEnWvHr
pUutM5J/bfKTWAN59PhSaJlulXRO9kHCxosJUOhUS4nb1+nxzq0aYcccIrQQyZ2GsVah4alANrUH
dvhdR5UC/aHFMLYEgwHA92U6ZZDa8jd+TuEYj88svCdNJejusYe70h8cjHMIutlSEMHp6AJRXUEY
VqnVPE5ddapIYIRRYFO6U62l3Gz1+m+1O22ZRWGiTqn5QCWQjfxcZhv0dFVZr3ZLmQQDBLmkRxiJ
OOxnTtZHcD3Ocszj5BNosB5cj0Wfpa+ntpGBYJ6GIOsucOvdmUOmOzvW5dEIMyqLOWt8nFH1+14T
reBdhY3wfrGp1fmC/fb8r40pKLrRpsxQhlSTi+QgDvibvniGprGmJ6APXeZJd3VqPYiPX5Od6trd
2pV19i9vp2w66QZRLENCoL9YAK8g8oZ/B7lmR3s8P1TdphE0KRjmwgd8KoW8oHQSgt9fLr8t94sz
p3fimD465tIwq9xw1poYfILYt5GmV6k6ILHyGy44nA6IQe/IbL6Xgji10Y8UczFhttP8HwCOtt25
bUeaQVYIUU61QTUG4n/1WokgYAW0e8noRzZQF3D8PTIAmIjfpFAwhdYtEYBv9IjsYPnAtwFMKHow
CMKoqIEMsOzfKvHEpVsgGpL0dmr/StQ+NJelutuTjFLkV7fXn32Pk4Bqcxs0Ke0jaGqKdpV5C0lM
KaS2zq3THot5dcBbV/Lu+enfLKbXNpaE3cQ8jMpknigfb+zLbquDym0oGoe8459f9r41jKg1GGf8
LTm3VU65W7Lq9lKKRAzJMpSNv7ppYYdiTgsM6uMkgqTiktzklL7XMBeGca5ytNIABq/0bFatmDSM
UHnuh8FPyOIy9Rukd48CiH60cQMBu9puT1yKkg6e2caotAi0RiTdaxvibnLW+I+Hd/Eg6v6ytLmP
kRQLbu4ROXn+xnO7tttgOWxqHjf8C64RyQOV3GAlEp76XAeM/T0/gtZmU8AZtxNcQefszewJxYfd
EK0c0gXCNV5DVq05+Apd0jZ1a+f0O23QP5B7pOme7rIYxDkq+mVZIDTR9K2exJGobMNWQ1vKdbMI
DwxhmWHMzhc0gpyo5jJiH2CYiMq2fIIvXcYZGjM9eT2Syjtqm44ydkh1cNmvFLzNnlq7apb3/H/l
RAYNS5TLUPq/GhV1m7hWWiEUm0APVrbPX7y2+3lh0GFuxoWz1J4aCCtRwZoAOY+A8PlxgxAKh11o
ae33uHQS93wB7XaYriyiTW+mxi9+8GjpoZHNZtjxqdQgaN12f6u5O2REOhp7GFeUo8QW9HFw3pKV
QzeMDn7Rg2F1NpPYXIsognHEhcceYYNWD9MJ62GHheV1e/vwmvabp7KmTiWpcdRCjvjsL6Fl7jr8
UX/JXpF7MhDeORxByYifwAVVbpcd1ATMlyTo6fq3+PqsmYt2+XuI6B1dYNO9jIVc5GWovSzS2Pye
VbpYm2MAn21BuWG6ug78UQzNfbxO8zuKzjy6EfYDZqNXf/VotqjegiPkhj+2CBBO3TccemqTF8W8
FGrQL/hFoKEFiG035m7b3yMRQzFMS5TzWqVmvNgzeT5Tgp91EaGhknbiaaa8Ll7yJ9aZqP8LWfzd
5T9WmYDgx5R84FUtxI68Jn1vdsTLt+Y0J1/+ZHXdg6hjEVpYRKgDexP/Aqro+MxOJICtYgJJ6Onj
RIAXOtM3yWjy01Hdg9R1+0o1sINaV6tsxCdmZmSD0NL+J9U5iaZu42KHcHU8jIyAqaEBb18KQJCN
n4exFvYwuwBphaLRROL/HncToGIsRd996fVLMH/CpGSqYIgglNa0AKYBFPxAJne0rljnFZTRIhJp
PoojmsbfiJtBqj8VRm+ARpKCl6MnbKCdXlbQKQTO2Ose7OZ2YymPQDnJSRsPbyYjioSk4KCxY83e
AMo/t1szZjgLvCQYNw9o3EEQJr77mj4hmfVaxiaFKayPIf0k6XIymMHrkKUEluHPTYnviGEnwiWp
4NSVyxf24XZ/Aoo49UxXC8rjoDT9+DyxsogsNi+FHPrr35hjn2mwUDFm8cNK4uUIJw/+tDcGKjGb
ZFA5g+ekZkURcuSMY6uorOaW+lM2Iwx0vOsHHq8pHADD3LpFbt8QWWQT8cKunLhjSa1YofBf48nN
IgSW59Vq9w5DkEce5oPyUpWMhVPEXfPAqw+Y0TVgIi5EeGd/TKziq7cOox4Ps+VdQNwQ/dSo9vl+
nko0M8iwP7V/oYYvNkmDePJ1CjW9CPLZLDmkDOuhzAI7O2Yk8O53HTgkUq0vdChMYFpl/WgzKztY
0C0W6LzRffDZal+R/9EBpzZDC0sLdD26WCgjLB26vTfhGIHXhguEu+Ai/FNrAcGnIqunE58JZcy0
bgTpsuvYnPXF155NiObcrcuFAILC9vIzbEGSOVtnzPI+qQu2zDAY2iP35WXA4fg6W64NVvzKNALv
AnKLDZewCOfRMVsV8nYJIDXvxNiLRdJSKihrQaSHnB3QsYKIKaGwb1NDQMLMxvOm9ykD3K3Z7K7G
WcNlENY8cc9aBed/MO+RpV0/jN0LqazHSkECe6qGxBXG6GbdheOiQMTbRFpuak+fp6+QJfOqECCg
/755YF+faNS/v9xdckLIiQ+5fjarNP6Yp6OIyMecGu2h8lDauZDI0+bLmbvT3CeOs11YQVlg80gA
Hkh70gCIcRsINxtsy55Bki9kOo/QTpIUCPZcb66Ws8h8G/qZWAHdc26msjI5wjX/OB3l6PHCzSRh
B4KFDyWJXp9hl/TmhqEgL28ikl981paFCpAJV++qfo6UpTb2s37K/nM1Jat9NhcXtPBTVnJzIZ6Z
DBSfOodszdgciqB/8MSqyx6DGHXcGKTiJYHOKg3pkScOi62j/W1HafpkERDIpRYE9Y/bsuUFL7eF
bXoYTNSDun0idB7Me6ywduznd23m7TcfIAomXnb4ZbIHfPAZt3nv/c8snfZAdvhMH4abbpbjOohl
c+jgHA2avuLGdqP2UYPYIqvPAQcfaS1LGpWZ0RbOncN7cRMbo7tN2yysRmGZEdppIr+v/Yhl24HP
6eZWqUuqfu9iHnaDfbfhCFhEeInR2wI0KAV45MdAMVT65Nzl8MfvXfPWzmYRz1gWl108yxVETgnW
9mExv5ROKx4zLV7rFYe08mZA2UWQ8lojDlVG8UVApgSutn5uDZniRTyOHU3BeUvdo+QepKf4/8eG
H9o+KaYT0vzZuxx487Wq7SAZelpPLm9Z2nGZPA76i436arSNov22EP8oTlIYaHktCXx6RK0Y4yyw
YsTK1WSF3hPN2BCXQH2x07N91puGy7Ya3HNKpxz4KLmPE19AKm4oyAMJA5h6AcTwmxfLh/kN9/x9
z46yyZrfw8kCfJO5Et6KDlDfk9QjyvCTeI80RBNlRpRxmbJ9NTCDJ4vBLZr3/XtT233hIqGpHBPB
kCU2MJRDBO6uPC3DCQVvPlnlbNR+qF0H69AehitI6I++faOAjmKHVfyjCxKAs0zyerVbf/LnXT6H
We20GSZzeJBQEHMiiWyH6msPZRmEQTD9LHqszQHzV4N1VZJEnLf97ohO/jUcQxPJT4rHPwhjFw0C
81lZ+TpV068vKOl2j341HY5fL+YsfNS4KUcVS6uGrejhNdS45HyQAI+0orHCT94+VjyDiMWPIR5i
e/7ZARiwTwEItCdN7yoMlP0HFHLEpu4pM+QzDXfDOS0lflozHGk5ipGV9euauV3B3o0azEUUvc6g
s3v4fUptom1uPeHzQRMDkP24wEQp9wVtPZRRqS3t0DA8stq93CwL04KrWROVTTHEddAHblMKkom9
RYn/gaYzZjZjPMCyFH9g0S2F986ruGAcg3Ig3z492D3qFPnpQvLbLVZyBGLL9MKx/lNOvJ3FIJwO
garBw2rMFVqNSGJmbTufLRBgbC2TTPlEPmAdt/1zOu9NYFT+v10m0Jd5F3b5leNZxSvRTjDGliAh
bUAenna0py91m47noIzrfglqtCz5QX0SGyQd0hLnuPB+fpsVJWufHqnBcUYbG+toLmP1hJDDfR82
PGPD1escOQBjcZjlGZK5afU/1v3gXrrJojCDhr2aYIMpb2HXFvPJnJv/1rs7d+6fhSjSXevuIv7s
O9opCkVXjihkHCOED+OcVoP5+2tcZpv1NjGBXzK3LWx13oc7Z/WRa+TgjAgzr9FnPYTvBnqNZoFQ
FRkyVFcbpN/j1Qj/EfFZ92G2TnVfNlLTBkiHUwCGaP1I+o5hy0p+hlsaVkFOgttzC3q93REFVJBM
TQHEMrMGkEEUEhSooHWcIoeJBT6eXIM5IKe21iiW+7TkN0+3PV8L/xU+T+++heQNbqEXWyHJVKDZ
Dv2e8v9Za9NAiVe6Mdw+OUFOxQoi+IVj88gQiITTy1M/SGQkgcVuyZ/zDY+tt72ww/ND8TjHiPDm
ib1WuAL+Qhfprv4rI22YmlcC4+lRnsOO9tv2DhySt1rYhatc2NgGfm+6SLWcvzdQVDYNm9R9ami8
AcGJPOTcP6WlWRX8MmY88mW+DaJF1/40sAQHYcdhU5BC8Br/A1utq948nubMLYcdn0EIS+ybzdpZ
uSolAYq77IFxZsOk9Xg8Oyj8AmO+yolbhxHA0+hj1gdjeqOy66qABYIae11+hQTG7Pc1f02zJWip
2D08HBjobaY0byYCX6ACjSVkl5kWO5XJzBQYhVdNLrGDY0nJUMEAcEktKavNokPOe0+S6lzaxwZb
LdITqyB1ebWqgw60sxJ7jMMi+c9JmZ4SpJiQ/m078xq8WHXyv+JoMNvQ0dkVXgWOY5x1gVeU9GSw
LQzzCxdBQAlRikjMyLbyuAAso7PCTE2DgVMORqtNqs1Eclefz3r2Nc0ro0r2i9cVKW/b/TRUnVPc
q7Rd4ftF1fdOZHydgd/yN8qOqC1jjhcekUohRyRWvWaG0YZtkOJf/0YVX2pZyp+NFEiKYvqVuodW
zLxJkAGP3vQ7QtAsL/NaW/uKWsAbLMI60rkSFGEREMUAeKqhA0nSdSkR9KIZdgVdSCkqw9caYySV
YxCoIl22NeCvECrtTvV/G2xeELQ4DLq0A0LuMQj5hKq/91+gbD6O7KitEHSrqtdxMwozOzabiOQU
qoJS/1CAzUDNrFNoVFIuxZZuUgagTHwTKcWfrkhKepxY9cFgtwE9mfe/0dmUjJkfh39f1mPZ6Hag
lQ3DkLjXs5TQELat6/d+o4zkxTVmrROQhjvG0dsgi1CFnVhuzgRDWLIL5PVmoBkyamj8ZzoMMYc7
YJTsTsbeQS8NgrOD7ChFKAbt44FFAics4hWrKdKYtD31rRxv3+Ml9OfGsj5WDk/MPotbOflIbRG2
spFiOCzeQVjPjmRsworqZd7cDsBxlKVn3brZlMArkufx8sTenztJ00TXZg6Omyk5wOiauAQyqSME
wGmpSvqD0kGFf/G/4sDl1mZ9Zgf0r0SXfFk2r6aQXWX13FYOBTLWB1VNfvHGqUN1losi2UvZ620i
m32xkwcUN9dklAwevy+1JA5Z6TGtNMkdOZt8RfbydxWYlU6flq5BcznbaoC5u3imXS+LrJJpnkJK
+Fw8BEUDvMeB1Uq4VVUHagQrgSLtdpr8gVFPb9Km0hDc55M/a2kdb4J1JBkdIpfsoI7SHu8+8jt9
t5cTN74B7j8KJ2ndo0weWZcBlq8v1jbtwEhVl3abnIuDoNgjfVBFKMyZ8o+4sprXy1cT4aGHquAr
wE5fn/C8+xDzVuzHOhi65A0+QQHgpmCQrwH0ujurr46xiE8UvXzSrEXhCVSxn0s4uAGvcxpaDxWP
4ev96nbMAHBh4G2/lIFvfjJMa2ZJmbBCYP1Z3aH7+ns82WMAPxobUcF/Oh2r+1sG0JR8/DuNUzOd
YMNiT4E7zSPxLfejRXFcVCmS7olMHvqlZgzSo+v6cvTuQQbSKQ/WoeLrfb1HaTjdd7uJzQIT9Ce3
Mk6GonlR0ENBcTUa7iSLUA7wE+eeXnF6urUuuWEC4leCNMWLJd6xTfO5K5Y1Apm8sudM+EuPbhOn
q2IafcI53au6G7hKnSZAA/WDyzUDy3pPYbZvFm4jaq20uDuu4+VigIQzUkKbKUIEPi2QGf3rW1Pi
4g9VplY0061zcRMbZ8MDN8B1tOGU5JU3/fj2DbAVK7Er5xVfBzVUdIRUeQj+SROahnxqFyDO6C1I
ZFgfVDFHQuKjG4n48vBev6JrEJJzAEXJoBd61Zbybdbzt4vuTnVp6fWQNmkuzGsOGtgGshaAiogY
q0PvJzR0SEtdFzpXPcxJHJERVhRmzL0Z3w6fqjMzGtNzLvle71oY2i7u+5H2wgSVHNcCfn8QTFBg
N/7mKM9wVx+oba+b5GmqiAe0/LJMB2eH7SuqAD0lJyOnlEQFvwKGCjuGFmqAA+SOcfdJRN31B5tq
/h2VBgAlhtl8nnQ2IMHUMnfX3E238WltjvGq5TZJ5CezJRmsVG7leHYLZuNjFovxCsgGd7+c0h3Z
HqD0ngtQYzVMUecskXJ0lR6D5cAIQgIRMbPVOkCvaawuKqmWwPVKj4q+pUf83yhc1mbj3hFgoVVM
mBnO2VwvJ2vFRUhKMNkZI74/FijQ9U6Z+Elh3FS1U/L0eAaqM4iOPPD4K8PBdyA6Pk7AYtL2xpTA
02zBhpqPWywJIfJKSG+PVBRa5FA8jHy93Gwh0G5auFrhFQg8jpwf3bLF0kXgl7js319NP43gKStX
5sjRu2bdnP6/nCGc9ir8pDgpU6zAxdIpePGOedPG/8P0tAvT4Cax08J8nd7SOj6GzwZ6BNCXV4qB
WhwCEjksvGaB5LLaaojbIiiUhkkioAIRRy8f3F+FvmOgbEkh/8DFNV3Ft21SWluMulME1TpJjEBO
6F2XvKdcnAebQzhOFXLz/h2OzmOaZIsgjfgCsv5BGpwUIPPHjfAJnWCemevdnAbo9w80EmCq7Jvd
NG64ZwlEfeY1xjhe+quYZvehWD2Q47lbLwUtnYyuA+3Ob2aUFNuZj470hOGhVWYRjRPFL5D7FzjT
/8Cj4gN7s/ppaU06TKPw3ZcT69O8h5JZOseZaONYdIHC/52ToKXf7XvCfvURuSSyWdckjJRHqARy
cGtgJbKP2eh3/UCAKR2oCOEy6mibNbZ0gKxjq2xiXFWGfvICYnDLZutaE5/US64B1Wq8yBECpepu
wxvkk12sMs8KHgOUaDP/4SmHtJLkQaxMCzvHorr9dQ+4bw/5ufj9dnXvofhDL9frgNMEl4ym6Ime
ezXdyoyGcY3628qVk72Q7XYM1mCdkCw357TS7tbu/Ly4F40EqiGb8HbGwScR2IZi/yJM04Cny1fk
NONJ8231zr2NaelNcddCvj+Qhf7oS9c+6Hbw4KiPbk407vFhkXCHlgGE/bkXA+0H6qSUiJx4SOft
1pR1BonCtMA/mRdsYcAiUDzScaK8F+7WvCZsGrxW8NSdR35H+Pizw3oOLlM1/GG4OXeM2CwS+/Gn
mwAgEBqsAIhHSCgjoclk2wcA2nnX4RvD+qfVzM/vDkHIOF/9CMgGsDxVIPLIfxAkpOVyLwqGGgAJ
es/PO9qVHUCG+7FqS1niepnQyGDXXN2EAoR8VeiPivL37Gm6vXcxD2pEzdQAcCwN7JFK/aFHPsJh
7wiiOrF8ZROIYSn27AMiBMxamrbas5cRNbx+wBJoDbevNYVcAND1vw1X+Gx3kfzMFivF8gVh1pWF
ITy34PKFC84efOtiOtZAo8P4mv/U/9HFTNpRYabkLNl4zzhfhyPC1tWmgdq+KhumdZ5PIadO8gZZ
t95dxuEKwB2v7e05iZUCi1t2u2+T7BaGpSb2upcW850mcyRkKc7PfxAhqurW83XCk/7ILqGD1iEI
pIFRtSpPprlAxzCw9TS4vaGzkKHivuEAvjBFHpuKsJIDBQMbV7xeF5j3J5ZvycCeST8BS+RVk7ES
uVW/EUtgW/WJqm9LG75m9sBcyjyTxDNb0WOY+mBqiND4jxmTr8nM7pRK3/SMiY71OVgc7D/p+4UH
dNC9K09ecyCAv2HzNwyOkDHsGLlR19t460pMCM1iLbbqJyAs2A/gXJqlDgwtXxOc9Tt81polPCXI
8ylpRKiFQ5g7y4HZzjqXoBd3sjNuG62AzQWx1pJXbtdmakEvXVXdHyGWkr7ZpwMFR9QkDAFMjdKW
25Iv0n2xPbUctDlMXRPeoVVXzo+mr0TvEulvKhOCPkE0jCEXNCF61ZiAOooJUVI71zH2KLk5MMVD
7FBr/BLgd+UiOr80Kt/qroxZ83NX5jHjo88kD4XZ0tWaN9p2e6CvqrTcQ21ebjevbZgidKAbbCXs
Yf32U2JAhnmVQ/7MHZ/GuQzgt6kd6AjWmaskn7DBaY8jidA89f6jYWG3+uC1vQ52OAXCERmZFw1B
4OwgFG6BMqBdn1B9BbKQnhpAaSUR/Ady9H9vvy/WZizDLB/koyQn9yiQ5yQJ50svAhRkqnBMqxDo
Yh1gr+aJgcvMREdz6XjVdb1VxSQAvxxJKwxk2m7WyZbm5OcpgbkItmoGuGdXUDX94MJLU074OvOT
4Plkto6T4hLsGPU+FDhRWatriUBX2h7IOe9Ut2KLBkuBTYnuvGVy/NryWI5WBLcjsLIx95ZYeexk
Y9NSq3P4SDKEs3iQzlPwm2guOOQ++3qsPF2mcvLhHh+g74sfGFXDaGGFojFvMKwkD7+riTS04URA
mAXgFAzGXfsC33v8cVEA0b6K/3/nWO1W3eae2Ie6sbJG0yEZEP93ZJZoHOXCuEUyrUVudniHKLEc
No7irU+FJAqA9VWNCVUg7I/oPvYetEfikZB29tvXsXbJZYS1W7IYRNYKFkvTlAqU6Bk94QqR9fiU
//Cvj5LGrdQ52ud97NxTBx/xfogahYRmf0gyGj/BABNUtOwYdpRBd3kzmHz7ntesnAUvKQYceXdi
1Xs0ydyBa80+/Sr35jWr6l7CXGsNeki6Yw55aEtjLE3FQbPHcGshfuA7UtjU1kPH7jOHU7O5eYlq
OU+W+F+8nZs9XYJmZHBDSiDprSDUoUS5H618xs9d8TqYgCSUb2jgDVF0Sly0NcLUiXb9GNn9xDgq
mOodClKLLhHO3y1SG+3J930TngkDDG5+BIbmemfXATHfa69Z1X0+zAm0aCjqckb9fcqGv/bzNFSd
Ds45HnLplAPmtsJRv0h6X7myFtItEaoaldzqfSsux1zrtplzOO14ok1IwXsYtP5wfa442iUqqCqh
t7VZhLX0M3cOtuAB0Z9eWBibph056/9/Ag37e57KmJJdZQRgFEjrSl17mF4ikw3NDbl41DiWMsdI
F/zDlp60NroooNSpOPqkWxtPtnei8P+FAW7F2Y8fvJpg3NWqX+/kPyZpbPe76yEynBZu504Jgb+3
4ZG1dFhcRWcMj/5II3R5yuO2yX4nwHk7nUUTHRS9unczT0ZdAst+7wUQJjnp7/9QwOTymqordHs/
BZc9mxhDJDDOdn5k/QIaMKCBJLZHDrkx+j82PskT8LlClet2VMqkKb1nLge0FL3aOmMMaJE7jKRT
vTCtTdb8sj4k1EV5+aqnzP3cjRKMlYR2WB62ntEWvRS0H6BCoTi/YGVKzNfjIYIY/uNKYWuYYtTl
bfG5ra4TGVqm+/NeFM3kxOfsUldUdvLI4NArUfdlDRjPA0xNfil/wcHLfuzxQ6R/tnYc5060c8YD
gN4HWR4P+GertTTtBFuhwCRCqq72yIfZA8btjQBDllmaeAFSco0/qq3F567Olr1lUveWgtGOVfq8
cSDeb0UWP740w3aSTVrlsfpdVgBfuvivCTdvuILTFoxvUkFwFbICsIzN+/5pkuAtmqWMuS+qMG/l
FrUyeb6ClinEVjQfEZhmG5iViThv9I7x/WukYMdKTyurfvpuD/muyvUt1Y8WoZp4zMI8Ppulneca
rcFfsd4qJ/9KONcLyCNqfZSjGEKZMvPTWcUCL4CRvs87NE1gAtG/pUXmjuPRyF4ENLl1HEzK3FFR
Fwa8GZJrXEyEy5IrrduhGvlqS1el17JW3yj5BYcY56r8AJJeFGpZ5RX3xh6CbINop64SSf69Catr
ogjDZE7wrF8Zt7sabjwyiKpMtGVltxGvr/7HjARN38OvZV7z9vYPuD3YjuVqTHV/WA+Gms0LJbSN
tsOpwJT5pxYXnFUXGPJKtPTVBGXsxRqlFvY2/ax/DFxMFQunRRMHUXvYyVkCU1dArP2nNGeydLQ2
LEj5XOsc1ihHcVARjjnfLkDRfdr6vMpZ+mNlpAN1xYSgBvyJwQfzlpBfxLpamufijnhVfuo9bOjM
vp8tw8LUU9elACGod8q0inYxU8neS3U0KH0X2B7T8CCTItgvzC+yq9wt9wp86WmfLqCioVAs4GmJ
7U/bqT2FMvJYLvK5DRRLvvNA7g3K/fxIGpgnN+k23He67JjmxpDZt/V3aZ0c/WMMihbPRfLPDIhN
9YXU72LVnm5ot+WpiAiNia4m9q9uBY1XHzgoQUTKdyrt+Y7TnM/UEVzNdCorv1/8jK1JQk8iAey8
f/MBInm676dMshx7U0vOJO+uFVRs6mJerp3I8Uoi9EorfpqJmlClruza0+MlxcYYaH+eD/AAD5Ua
OCi9yaQlNK1rrJagQQVgBhiMDsFaCX5YpOUnDhem3A1Y+S+ndlVv2VSYZDSeh43vDF4plbTk3U1b
1OHQMiZn6HCgqgPVDkWnP/riqoB3YWJ/WXzG8lfvkQP5ULKUrJpellx8iBKA7HqOgah8kr4yrGfp
KBIeY+nIhFxUUtgQ4o1w+qdy2owKb6IdoxsSII0uBJvWs8FKoeeJ5mPBo7yD/gzzyE4Sr4cB+i0B
YPHiJDWzOnAchrPUjglPDCmHm/xFHNfLybjAEvts6e+GHxYauiQ3cwPY0i9/tyRQD3wSeFF4MlaD
5I2iMnoN9Iha70nyRaLnRJDIT35c+r3oj39lZIODMBQEDCViLi6VC9ZNbC/E8+Rgg/IJVmC5UqMa
xjqB/9soskpuauWfB5tOa9feC/kX6cB5bAazyme5i0ZlxFp4kZGCWopElFKxFRL3PyZQ5YhjWLOL
kiNWlzOBjdlmHtefeh2Q4XA/mWgWtc1LmG5andVQrqL+rDVuEZ3TJtmEJ0NjCXsrtivUuoXidbF4
bYOw6cJrnkf672H58jtEFjTUPqHrPxNxVcMoo0FjnbbS3DwAcHxAjwovIy/ORC+yy2+fliKzpx62
iNlmzNmuYr7rCrkLDSr0hz5WTDb1qHP35hzFyVfkFaVrKZdSFmtoCgc0So/jkooR+i8E7qh5M3Ly
/Ka0M55HmAWpN+R1CMOPw6OTEj30YowsrSVWlA==

`protect end_protected
