`protect begin_protected
`protect version=1
`protect encrypt_agent="FMSH Encrypt Tool"
`protect encrypt_agent_info="FMSH Encrypt Version 1.0"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2017_05", key_method="rsa"
`protect key_block
mj+hj31m4NdSScSlQQEjIPHn7tsmjRkA41yKviQszlqo1PsOFCtLYDn4Q20a0UxySm2vx4SicP2A
d4evmR+O3fCNLUFRss7ZYlvmVCqw26p0yCuu9AJVsmGw7xO6GENXmQEeLGIyaMHLgp3Ojszrajan
nAX2Kwe9kuAFEffCtlvYtgommRv1M13IlPDgYVUcHk0FMjIzCRhtXGnEMSK9yvOttwJyJLA/sZbt
N3YqCPGuRzKidZsxjOYoC8L1LOJc+Dy/yq9u/bwHfwWEWzKC3RI1dWSUF70ECBtWVZMamAF/1BU+
rS3y8NjIq6Vm8TuBGQgJnj9xPbg7TqW+1+O8GA==

`protect data_method="aes256-cbc"
`protect encoding=(enctype="base64", line_length=76, bytes=175280)
`protect data_block
RIOraTNkZNU6VysMP07GHU1szUVvYZbU6XcfhQgF9t1mC/4OhTpmgrIVDwd/Q7pdTQhr+SJoLLUq
R0LO5AQFEvPU/Igugs6go6Fem4HtgEWlAIhw7FDr7WDBPrDUV9P+6pu99tTOtutZvylUEwif1t3L
uJYIoZ0i3DuOWY5clGAt+n5hMx+kQpvClPM/owiPEva353mJAXA+XnPrQdN/NdwM467y6ZDVWEwu
lctm9bi/AJkt82LoA6hAnmHncvU2PdpSgfW9kkmWYHKzjQlkSSIxjUhuYPe0ErgUMrET3v2puGWG
sT5END+SJClWKoZduwQ8yVdUn4jGSC7Dg4lybq9s4G3iCRVtrJJO7rcp6sDjrJNGf9ACFaIbtsvf
5/uSisDSKjExcnCWZYWdv4pGsqSsmazYVCAMEBh+oIwgk7pC8st6C/UyVOnIkXcoYfbT0WRKlI5s
+YwgfWN0Ixftnq4jTwvh6ePmUkpU53S2OnQArNVaP4JM4ruaq/94v4S5y6enHDrWi/YUT/N8+HvG
KVkO82qQkhdG0A+xllPuBPgnRF5NfC6LwhULJyhok2nYl+tE6J4aq7SyEzDa/UV4dM4AOInlP43N
t5ZwC495K98hW5oyPmeft3p/LLCufTwb67OYSSGOd5z/eV46216s+x/L3l5qbDblKeA6htr1uR/n
imQAySEfK5IAmLnBedGpOShcNi3X8a6CZGUPWulmK0Za+OhLtiyUFGySzqwJVUiKqyGQ8k7SfFAB
rHeSWD8wH2G0bFY60AKVcoZ+jHRht+QkH7HhsFII3+pBHBM8uIjTnXZxbDmNYzQg5tzfNuoiGvF8
uEdWdSZ/D76pvY2cP2VeBXB6aklUVOh70/AzVkAK9odvamW4sfMLXs19YZsSBorZUQhJKlCguoXR
+xDg2BrwoH9XLicAZlVPBWnHGVtw+HuKgnYybBfwsQQanEN/8fshGDbu/Vjaec8YUTe0zGmN+N5h
plSNs4syPhF3gXB8ferKtSrFxFIUIb3CUvi36jWmAUrYGotuebhp1rptHQDqSp1Vwfq07ehYskKi
eKa7vl9OyWanjSQMi57wr3QGYPJtKbjCnicS+6eBjaqzCvQ7Ctuog88sQdfZ+JAU5MwZR2QREw/P
t+aYcT3PeQh4pzPQZPQYx28dhNzQv5PNXh3THrj2RyhAi7Cs3Z0xUevgw5cb0jjQJFje0s1UADfW
0ckkZnhtKEbye3mmPTzMsYXf1OphIF28O/KabKYHGcTuD0zJvAAMFQo6rEixylkXfQZqIYID8MJY
YRHk6jqEvKPcXg7xiQsyFipTpwVD2NRkw8nmLx/xW7IqJg1nvdcw7Gv31tUXiKLQfjjFkm3QgP1+
j1aPv9b4pWhh/tRDIvpjNT/Ecq7weyhMCP0Nwi8lVw+pCmcZtSS61GXSYUs7SZ7lm0SYyQpzSyXs
xMLc9rolGLBITh4AAFtIJ+aQ/o1G7LoUWOdbEHzM8wBgJhPod1VNHgive6AOvMDrR/ZGu22tJKxt
4GmDXoJfF1g9Ce9yblrNVrhdbXwyZyrEq+kjLkWaf35ZSAQyo9d8h8WZKmzunnsKz+geX0s6RJ3F
ofM6jtuI6RLEsnyHHA6oRsqn9hU6TskcLBNcELVHJFsJFmWiklX85AWE17cqw3hI8dC+D1MJOCge
e+oyeDdWvqfnfJzdCe3jyeXVXvqVMMTi82Z7dBJwc/z5wyScF9O+uC7XYhN5LJWV+fnBiA0AOtUY
nCNn6yXnlqMB19YAr5Wi7X977XnH0y40UGRKqywj/oAHDf/Jl0otPn4Jm7Zq7nIRO9wEd1nWZDXR
tDmV5MR4icHaFPLVfz97F8apOubDWHEazxo2jhVEI7IfuW7xm+sCatzIqSQmdvpgt6KMg2U19yQk
rbJfq6tXyU33G99d0YvDJ+ai3cPaGlSa3QXy4mGXn2TmgV5W4nfnpKnRGd5a/cVI4pWWwRCkr0Zg
wvk05rWu8fFkvXH8x8BCK7z0vLpMBnf8PfE4ihOsr15Z3N016oFSd9oLbKukMX6bCjwNIsJfBM4n
ghJqOfefNojZwK7VBB4EfnUuxbWVZ6FKZok5FxdO/2Bst4rFMIaRe06s8KOG+x9gqKUmmhzxE7F4
9SXlbiEdAF9cuTGC063kzs8I7BmR3wfENNkStOYTConBAPX5bRMXDYm2AAECc0D+y9T4s0s7IjVF
c1xRIKb84BAjZoTjh0My8nhBpoYc67b20h2dLcWl6JPzoH5/UW+tKgjlUzPbx5LUl0PjYnWWtmUC
vK18K2QVOQkYlNbv1R8akUiAdI9pTgf4EyLdLWhHdKDZdrIsyv2Y4bLrq5/9SsY/DLqvvyaYzr/5
WCZ2QWEz9XLMQKJR81FJv/trAjPOYVWKjP0wx8lLrR/eN8Fiy4ov0bkNefhn+MtwNdGvFBcBhkbz
fHtQdORGUu+v94JqguxL91+Egkgj8FhczVNEa+ysAaA62Lo6j42SL5Pjr23WLtnSphTwkJAI4b08
TIK8EGaeFBwhm061s9RQy2qtFGxj0rUbs7QDgvpdT4U5mHVUQQIOFTIGqfjR8+oTpKwsw4z4IxWb
fOL+nuo0TFkdzFlsJavrsIyvxuLzbXsqls5rbS3e/0HWh6YAGRCHcDU9sTDeSEkBAUrupQIaCf6i
McEvGKk7FJcozl9yn6ggWxmm8c2IpmJtTAzRjgSG/MzX7tVk88OLeeyqszlFGsYjt8nPU3krnccW
NqPyuGw1kiQqtyCAM+UGNGP/oImRF53dCIA5M69S9GwznjveYfLnc6aN8H8aw1AuiXRCddFwLYM0
ftK94SuCUYG0H5MAGS/WghyFxO4v0WPpLwXyG08dtHq0nDhImx2WOrszcbRdl4QJgh3fWdaxevyA
PKYc03Jl8yy2Sox+ajKGUXV4Zwm04Asdd3C7F83VVLtlewSFWPCH3dYFBjdbySc9MaS2unVCwpqV
tuV7HSN3K7E4o9zZGXRuBrrSU4a5r+AcRQ8RKTyLA8F5PyfDxmC1E32Ah+lEUwc+bQicS2cdHe9W
7onHsUwYIJIjrS+9DT2c26ips2sB8HxGLunfLhv9AB8/Om30kNorCoNoUA7Kjk0BcyqmHGQvluVO
bK0TLD2H1kYiPgv7M9mBGq++6IjdMb4qBIXlcEaAak5y3acCP9RngOl6GdJ9IT26tG0xXy3qL4Ao
04CzRnDsGUggOXOwesxw9+eTCOfy5vkf4xLu2UAF2+sNvQCvLmnvs9StP2BULQ9RUj3eFFpqmqlE
gLjeRUjpZgSyvAFp4rKLJHl50zr8wJX6/cRN1yrt5rE1xCO1mQ5JHO2qZSA9glfoMpViXtG4zwSe
jKuhm5+RmEdBbI1bfIj35yuXC4T1sly+D6eqTR74qbVRYHBkRELzqSd5GS/xPRNzSvjjYY3oMHGf
NfkchbFBz2jepxELIV+/cHBao5LdUCtz/Ei8u4jgoGLvIJZ6iYp/tFhOmfBNq6DpEmgF9etTEhoH
vDEELFg39YrBkDqgz8sPW9tSBnSToh7lgg1OPJAn0pkGDbvvrsQPLoHgWzFbFlxM753TGIBQob4W
Pem+A5XWYYQOScUAB6XHtKhEIfCz7D2Hgt1st1noV/oJheg8PojnUqsx7dFTW1n3AcQuBUstplAq
4/MIktcMex+5Q/u4t6oe08Qn7+h//vHbl2u8ToHZXCWRvbRWshA+JF4DY20WJz8O4vCgbBi0Eu81
fu0DEizhcBu/PJFMXSCUfIfEMonmgetAdXLKheQIbavoqv4xwBAv/JYFkBcveFIz0hA2mMMRH2Nd
Yp76V+s0zrFAivp1KwBkatHhp0HuZssLWqSTIqdzJ3zFAdCDq5u96tcubhLm0emXaqXMvQG3wa/D
NMfWqm93PN+4miVzRGfMfV5W5jVsf642vEezThUfl9EsnA1WHIgi7DVoBzU1gDaMXh3AWgzNDYK3
wVXv0CgBHFI+DFQ8O9F4aENkApCZVX1QLWsBE1zhGH2uYhKfISl/2tZr/bnv+w6TWrVA9tkXgmcV
+88LeyfI9WeDBteI1httBF/vFyIewQp1AnNLWktOJABa4VkYzzeCnSNz9or0bh44//X+AWGqYaO/
srZ0rZ0URTP4lkDmNW9ZTcBLHaUiihBHv/zJlFflm2/fgahlJWi8FuPWBWJJGTkhSWldVkBqrKB7
kC28SIjgdDpxdCFycVjs5QnBcvo/UvVwhfZ0QaOJAhsf1Dbw/Q5iEY8gw5X5fJ9Ppnp4yTc7hlcs
VrX9NmoRok9HT5xC9jV83NIg9R5xsyaCSihaHUu3JIkdIYBtDoHuWKsFCfbRyiZ3qJoc7KmYVc/K
pDu6mWOfqTATk9IQhYB/sT9p/shIWYam9OvPA0n1smLLkOsweUO7gvmdURRvOjEDz5EyYZDZGnMr
FwsZp+vul2wTAku2V4b2DiZpoOQ//oR93xcYqbLx0mQhMrrdMfV8FOY4DoKFn5XBkYm88dyLFeg6
oIONIr5n3uipKgx+cdKVroSQ+TCecuEyii4a6p6DFGgynf06UIy1AGeEaXtc+3wSc1FxX5T6ehi+
chQKiXEAzzCh7rtRWff5QUzFValqgNhMwYn9pFUQF4L+uCTQhXFb3BcCrgpT8FOjJouGQnmIIUq1
Q33G/nhjxDp8vOax4/sjYaSC4LKxtvZfgfLW6pT6T5OgLgKNO2/yQzV5IDGxs2dDxK7ONGqJU/5+
Dp2yXFZY7C57mqSAREJ9XzeZBAJBstGXv2L3ArQC116xJ/K8k3n5d2vkVaME1mEt280afK/6LQFW
hGzh6IxOIsZWBZ65e0O62uX/zl7FjIQGJkSUoh/esEnZO83IZrrp9BJAWsMiv+m329dLkaE2JUkj
5nMnUwSIpFMcGSWmfjrYpCRHWx06dIavND0StjUuXz1ydQc3FWE14fTPT7zel7zIJuZqQqK4ugkM
Yloc7zJAWydEChs/UNxyIjDdCzqF1HWiJCcejUrcL8Xk+h22ylZzQKxRoaLet80bIxL35NAngSID
Ec+0ddV7A9nKlK6iIRnW9tvNI1+SGdj5aR3ViRP0MgBm7QzdhOFjEJg5njIUHlU4IFKiks+z4xzZ
N60O63Kml8p7e4dVGgmSwyg8wpqUI9LCbdHO8ygdk5aNk/lNVzXI2RD/f7ADZIL/T4jOtfPkcO/A
0G2CfLulC6BkjSmOYiXeBkf7vLFJUPT1WOgsZqLM64zN0lmqcxuVlc3AKIdDzYntTlMJlNnzMmpx
mKcu2AuQUbGMhHy69g5kQy6BVddnNEO6qDCBnT8h3ETDayurpijmCQ2xHv3bDy7dBru89m+3jmXD
m1+/aTEYDkPsjeUWmin386NYRyIM9MwHNOWW/pWYL4Gkop+LCrwZ2mh8IJtlE6NqDksUkhR7m+jK
iCEgrfEYYGV9SBnj30MrJzy9m6ssTPezQ9Dhj3xOfXD9xFhD8XsJTtBTHqCzJtn3ypAWw/nrPHEW
Sk3y0v4llHbz/RAfa4XUiSW7BNz01Z7onj4FEsTo6ywYj9z1lMLPdoJtcwVEP6bubHgDuHxlAIl0
qzdyCj2NOeleBlFGTXyd899dVF5XT77Amycw2ZVAs3FBeQkep4vAWArUpNjAHDtJy2qVDDr6FhfO
37q6TlAMr8j3k1PEQ3B4m0V7ft4aXQFvNOIUwUi8wBK+6s33UEZ9u78tqmoDlbLZIh7AI1J+3mQb
0nLnoH1B85G/uOMZQGzQE0Y6RWKXQ+B0Gt0iQQ+1ru4cOhJis6FyL914O2G9nC0ikCnyLWui5DxG
y9Nq0yQp/tYNt9IdOTcdwT+VDiPq2QZjpUSwpbzrqsYUEcT8VDEcuaNpWXv5zQMWMM9zu5qllwtb
qlLAmKTz8xgSpusiWoT/x6xdwlTEBc910YmkQgM+4PrVt+cUIFy0BbTwpAnO8FuyfqhRAyhW3M0t
LC1locVdnqKUOmwL4yI6lISJJGaVeY6YTO7iixMjS6qxsLiyOWymr4QfVuAGQzEbuAKOkQZ5Guv3
EzlNGWhn4VfaBRPPCn8k3e2KHVmSjtKgj0Zdc46ytPwJnB+BRsC82fAwLgJ0AetYMSal4A4wolxj
TKt0LiOihRz3VUrWEuMsH+55C2nE0IejOQOQQZevTFiHS1KA+OHvjOrMMwc7d2yI+uVsfR2L+6Tx
dsTMy/WU5OS6oiPNQnMnqmafKXjzoYiAXmIt/lETsbzRhts1VwxSA8rnuXJOZa0yZ396mdSDIrsY
u8RT3N30xnBxRfEaKFmywKMRdcwdNbo+4ZiEXk+i9wQTDx60zLat8th0gomb19GV9ntLmdzPU7Yg
I920tCwKSlRZc7Yf9Onif1bC/Zxpj2/fcpRvJ/WLLbH7fQ7KmqHYIIBBfbLiR3kphQHqUo26jFyV
ja70v/XwlwsnFMAF5kyZu0iALinqmF4EiLLUfjaK6KLxTMvZUCGuWWKefq2gskCpaZIBHvFfiSLy
SGxggT9Fcq392/wzFF8fZ5dkAFHFf8BVdqdo4A+dsrWgSc9HhcyOwhKvF0cPkq5yLlFio6SVrom/
BXnbznXAILrtj2WaKyo6mMHkNcnKBYJJqbHjmkVnRq5648elHCuQo7xUha48nszG+ZVvglR44JQQ
dncb0NCRHj1lx7eZ0CocqOjL5C30oEbI7gPAEHdFQfTVrhcMrzqZ7ONBNVYEV9yCNq/MUxOu3y+8
WesUqg5m6B8axt74pDFdWU3cQ2mwT95n088HjHNL3m+KwP5efdOp7GG7UQS53ycP2SbxVP2o7DfE
UWHZzV+aV0r/wskiyXEIDtWTEbh5MkAx6Dx+E0xw9oRnwztfWWa82u+Id1ykD0Gxxftg19DLvQLe
EZSHPScIpGI7qz/KKUmcsOTza7UKk5baVxchMWoOx7G7KW+ebFgQL1KP2/8VAvvRv5lHycfuFXRo
1jaKjmshS6PgIOFpJXx5bdFDhYzaM5OuaaCm3KZ066/Be6LtCRbEizTlEgQDC+AY5CoRDYDrSlfN
pRBWZ3VRlrRtZ4Gm1B/6UGMw/0F9U79VmaubMLDweexxnQl4vJvqvSXOQCUGlHEh59TE1SKPU6tD
Dzl+mV7flI1QwFoXYvJAwbLnbstj0d4y/lBL6l1rlRmgl+ypMM/DlcAqr8SAYhZ4iIt3yLpnl5TR
BzsVmnMSKHPgY5iqF4CETLPcAAMEBJScjuhs2Js1VvCFLjWzKzlEphxO3JOZScPY85B9K4IPC8Th
WhUwup/PcZbhR4hrrnSSdzuD8wpLy5yKRkKK4Wm+UwIephONjHWIVlamTS6XTgFJxdcKWjJsTJx2
uPI7KoLwOZPSvrPyawNRsS6W+PLY+vpUim3QuNYVWHi3rFmfMbwDHizgmmp9GZdXj4kj2v3JrtIP
dK4d+l0PUeocYh8xWv/wmNxFWZrS511z88gtHQ2HHw9yC4REHkVR4pmJ+zuQteNZOXkfQ/JZMjWI
rp4UJU+6Q4ZTYqmcjPtb0rQzQPxPFOfgZeEEPn/+c+dqJcAbLNNTtXxXAUOtNHw38wQX+KjoupmH
T/Rexk8x8bcYcClTgmCind8shqs2+Zs3t3XlDR8ZSYRqK37YsMC3gxRkaMmK+dPk4jBiR6bfIhmv
kS2Yk/akc9Hfr6DlvS8S+ePr3HNCmWyhhse0v9nllLlGQp4vzx0bNhXMehKjrHd5rYSycV0dB4r6
6hC37VGk/6R3nRzi35H0mJJWwliBk1gRd+fk6a1FUM3NQjz+EgQNDf1EHcmqjwpbGe/a5HMA9bs5
wE5RNH8T4kItdjaYvddgu8lmiGhLjc8LSgV83uVi33ykE+TRAdkMIRhglyYiDSj6TKWcjGLgLKtE
Vn9SOi7PbVVapsb0O2PtJGvBUUW2ZYhIUwgxkuxNUoMv7GCuOw0ppz3sZzNhyXjSoFqzr5v30/VW
QBCipBjXKnTM+oe6Bi90B/FLaVRBlHZB0x8m/ffcdlpcoRbGDyzibKeyGuvBU0rHW5jYln0INVj0
nD79c0YUIhpPU0UsYij92mDqAOGKExSK7XudtXDZ1vgvuKHgB5KnpLCKDnNYhur+lfPKra5TOYvQ
Qjpm9U+phLp1o3f1aq2pHQWrSM/AYh1znB3/nVrbbjpAPMIsmvIcK0gpuRJoT8EjlVmGq97JApmV
1khjKoaQmhqWAnom8LXJnaGRHXAI6VJrFsXM8BKivyS2Wb5rNI8kxS3L1ditPvVGAYEwjFkmXt46
voU2v+f58ZM0kyx3+1M9jfIu0Vy8p7trs4q/B6yY/mFGJtKsdeKTUovLRh7uPnb815cawJELXjTy
tDpRNmiDIC/Nh0oZrAfPUR6lyY31nevbQ0cmydqSjkWFDfWgePjmeUAPguww4XBhrDlB7GYSi954
WUxdLEsJLKOsNHefUXv5C88IwwtM3F9Px5Uu/0vRORFJCHAsOiybmoaYmjNqWHcaNFw4NmScQyA5
0O8ZZMQ+yGsYUgGO8ynSdw5NBvwcYjN+cxTMmz4iRiefpAKVZRaU8mQ9l0hJURDpXMRZLz+nYw3q
RdOUL+9pbyUnbyXxcheLL+nQWjVTBJcJtS4T2yjQ53n2izS+9NDwV9nwy/SGZmc68BiR9Wl1eeoq
MDkVnAPwKe4ls7kRfxNejLOvb9VLCPw/oP5tQcXrKpV3RbvbzTat6jIt2TlrHeo0xuWY1ykN5wQ6
ahTmm8k+0Vi+XgNIcs4GwkB97UAk87Sc2DydBNeSVrtLWPR4plUF4Ki3kxXb1El/NpkHdBtF9bqD
vNo/XVdFLOW+BOc9NCETyNoOOcN5ZfQi+/WRVL950INfqHSai5Uye56/sHwjhYh8bT2kzyiHWKhW
IeGAlR8k3rpaay9LBD3qLoo9j37aOu2qdh6a+h9uY9RM7Qq/t659W46Y3snvqcMLcdjBVKQxIled
FbZeXyuz6r/WxTZZxoqTNVGHyyf6dlA6ksE/3q5JWml59K5aPMOB5PLZDtSQcb4J8V7dvXN33xsB
o/utm7w8yQ9HgFxqn2zukZOnBcQfd/dhAcgyp4iQ8opXXU8dqO0Hjx+E3x+vO79kW77FQVEyFveH
Ke04TQY2OMyAtU9DQxdN0GpdK/esjlnBQVgsNqlzWNEgoliR2gqYYc+K9tjfDh44RrT83E6xngTL
SLzKxi4x8jmqUbexGgEZNLlfT/zeu+PQH4xlO6BAtpxMK3TtznXGwsQr9STDPgDjK/CPpZIDkSCO
3GcB2yc4+oHVXY+9wk6sOxXvhpS6Lp+aKzwqpATcR18qLdmLG7ktpHCp8IEnOjTcm1g8zjnYWqRd
xqNE83DmGyP9nJArEwsV62UjmUNOH5PIEfl7f8fEcPg7z0S9/a4grIf3RcY9z4NBXY0dckYenSvI
beKPdN/0v7WlVWlNnQbyXFNn7N1I4WGX74KwIttFiMMEKNoCgeMV25R612/GFIchdaDXRazSq+PF
kFVdb57E+eRcPqYzsG+gwq1OuvSOvXH9gUjl4B+TvGhZqbfTvL27jODgHdH9Jx0U3mPVscm3os4R
XYoJLZWA7qsvzZAaANDw4uwKffQ8ujjoWd9FYFRx+X+Z/424DECK/3n0HChidyRO19LA7G5mn9X1
PZU9E1cwhksQkkfbLNDQAyPy96vWExrQ0pFxIM2GOelxQFFkQmbz2kZv8xjE/7ylIjW7Phlr0vb1
y4T3wGwwXkdXJxkFnrPXlYCe9sG0/BBVQUv1pfvS+hFaAQH8URzIcnu2ZGYiCsdayD1kSBD7flL/
iy9CmMI5gSgawsf38/JGF8YdUGgJVWKW6YzekgnhYMKzi3tHPdKovhSMT3yocr4vedioD+AHGSqz
KBgwonSYTQsQlpFgtaq9xd9hGin+qU8S2zFnOD2lNWxnso5/9Nx7xmj2cIGNd6ilAx523vvooPr4
lG9VHUR13wsvPG2kKRuA13FhiYGrrqiYfdHWgRdwqqXkUNh8sdwVemvOvz2NXvyeXqL1crACljly
aL9sk9J8pmOiBywhPkyfMJbDHqIQ7XjWhkgojZ/+U/Nzsb4kih6tfhH5XOENmClW8emkQ2wvyBjc
VAFkFFq5MrSNiNlcvxE04SXQFbdT4MZcOUjJ6ODRq7YU0UbvW1lRYDSsi9HXfGPzjc12++9CFltf
A0VnDRPQ4ATCIJhlg4Kgw1IBkhqqcaRIKFU1Zy1EkvCwtp54hPdlUCEvVBz7fK2PZg06svn2jkNe
IgyySsepqzwDlgyD1PEYMx9a3ZfycuvqHUTv37n7+oBJIk3muq8yy87gp+40nLpN3yXx9OFjrMry
aSy/fm0OKoLY/5eZSAw6mvnfJksrlI1JgRF8Xlm7/d2uKpv2oKQrTw+A1qGx6BMsuG+ldKCmbGa/
P6LB9gKB+UdFaxvP7azbZzWLcktStnB0EfXpKVzBwksMITkR/3pHkcGfQx/Q2IhiRt2UqzlGD7DI
PS8+4SVaZs1l2NgcooV5cpvsvsKzb0DFrlGVWq1AmaTT888cRLr85iv26X/8KcQ17RMdlqKNfFYi
AKXokfFJjr9UgQYsCyVBbtiAvHw6FaIsMLerzNxK8YGXkAuRCt2nrF7ndv4mvo0G/tnSfTpEHDOH
X9ev1ntYYI/9ws5waszoTxBtbgn7vHvpsXAJxR9EiX5gbJLZv+DLf+bbV3GkUhXQ6S9/fXufFfZ9
hYqL35JppJUNTwKbqxoM/gN9AgsdlG002j2ENoQ8+zMp5Nxu28QSGJyDKloHT0zUNY4mgsrVp8ZQ
+mEI/IDBKwxoiCfYOVbTFBNDLDkg34oscmuXaiDG7AY6rHsjqZldk8wXAykpu3MIa2UNliGjykJF
dM4x8OZXTMqlnaJrkH41DK/MAcC/JiNdeSzicavdcuOm6YJDbl75VudXIqiTMZYptP5nLviDHkNj
QOmpRgmERAHwK8dCr9Pcbo7comB+CukhDHluKtsLON6AkR7EeMIYrt/y66eogoF8KSybGRLstWx0
kl8eAE5DJGHyqE/pKu8hQyTmIMr3JGgTUPIToImjVor4QHmBLGKRbG29nQDnfQawW5HH5BvbkjCq
yiO3dHj4pj1MrV5NNQK5oMkcHPBlsfp0+ohzDaqiCTbNaA4/lRDnzY+UIjGVae9OC//NQAYr1QWJ
+PNu7ieU7HyO5fR2pONS0GfKEpiMq7uvcEKNYrADyKGk1y1phKKN4EsD6qYZn0ofxParsMmytTpF
ryN/BJM8fYDkjDytycK71e6Eo1h7nHl3BgWXWxWWkKOujtaVX0+HAC7ZEag2R7CGcGyyNlc6JiOE
aEgwYkvSBuxMwdjkslLv9iXiwb/c4g3GRHHNNf6AGQVL+xabgq+D/PkO+jDSK0t4joMnybTCHLqY
BFfQd9YzDwa2HG2QPXQG70NKA5eFr7yFTG+q4mposoAJ9tmt1aVxW+rx5zmYHeGydFVbERP1CXx6
2he7prDIn21WRdPjLFACh3OhCXAQyUFUAbzK6TF5mj/F6vmLyW8STEf9aVPmUTgbuvZoba2K275j
sCL9EFVhvZQBVTQH3L/npIQgAgHIKfhdXdDnc4AuZ4MjJlxL9jIcBn+V/YwMyrrarCZu6kE2O7z9
sBw2ARunTf6RvDNVeDh0hECKLZ3saaMpVcGdjGGEZpLjsA5NeBmrvaIMlpxDxmpcNLsyV2/LQMI7
/LUeAyxvV9+S8VGS8OjchPYc6Em9btB+awU7E1wutPbhAaFkvyV3ZPtSnPOrsBfmIg8SqaHSvoFG
l4pykIEn1D2oSF3vKRRMwI5r3PYPn6ba0VuEMpPmeMKRw4kF1wrbOT+K/JImFTfltH2eiBmQBeuO
Ws7zGSPhiS2/DqhyoIJW3+E6Gth1vE33MxTQmIBLZCda/Ih0Q4NJA1K3Jzct1cC1pEaGzuRacvp9
AlesFmZytCwh2HiwniwcTl1D32v2NP9/Ogz5xEOSLyYq0+GfHvZ3Y9dzpXiLsXOLmfyM8F9840fe
vLRTt49bQMADuP1pEHvm7Llhv1y8uBvFrrkgl+ZvGb0mMmfbgz3O0kJihCe/lSHT+0w+g4FxP178
MWfSzwoz2GbqC6GnwQBX76pZSQdA3cTtfV60/7Wc9qnTPCSxwy/3qRZT5W9WIzu9APk4P1Qx/SzN
0j/RzVCszuazJxDN8yNtzccgzPT7sQnD4gWovytfNJa1ysnelQS8W1Led4R49rGLeYL/5sRd1PVA
lF1M8NqjJU9x6x/eOkTiccyiPwHZYpBzwYeASqGalecD+ulAJPXmN8SN590EVfMJ93d0CVJ+QO7P
4scqeAfWF68zXxfNLvR30INCUxd/ZFgM8JaoxMvQ6ul7iLqoNHX06AzO8fw2D7iAWytExGcNvSZk
8DrxLmkqMoc1mMajBHkpwqJ/4rviz+c2eoA96GiLZzed1vDMSF8CBp/QZpZaFXQpa9GtP5ccvvwO
PBg4WE7PQcrxttCsz44NELr5CWxIXUzTWg7YiuHRoMMZx5TqfEGRL290zfN9TxhUssJ1FR7qXj7B
dJgRTVqFdKP9EzEULA13FWClvE5WBmnd/tgPB1fQzqoY8ru/TYtyop6+zSH+WRz4RlQPCURxLopd
3RpYujTENf6o6SQYxnmIWewIOQoyuJOUM45ghHB6mt33EC17Hp+JzA2rDz+ifKifob5yR9WSyI16
mpQQ5ldg4bepDEtIrxxDm2KrTEkWNriRmEnSjqPsThcr0OVTVZ4N9Mc7+hzGMpYcaLYeQL7G3IIz
39T4woE4woBlj8ktZ+3Qkkq8lFEvted1/CS2rgraQEzHUBU9xDslh8M6sJQ9ZldXUHbgXWPoIsp4
3DlrklVa9nxGZMcczBRxGBPVcLMp+dMBTyb/GmJ9+zYcXK1+p59yTGSjGxptQbjfo1noA7WVEEwQ
QW0GRUqDn4JrH1zdOdhIEj0OGib67xpg/aW06Vta9fSsFIdTFYHQekr+/K7fGU7J0ERHCjpf7+NU
/kHVc9CSnwOzpL6mNbONEm5YU/0Rdl2nGBUuniAmXqYQIFYAW/jzDCiWcrtgqmcu1HNCBfccCHRA
zNP1IN5Q9jH8p+Li5rrKDay3J7LZZjPR4uoELjwhyZQQJAWIxQc6B3H0Pb0tB/H3Rw1oEIbeF7nK
JCWwqdx0HMnQTHATO9H2XWvdDO7l/o4BThrTNXD24xjMzFmfJPZjbtw5J90nwxXizjOrOF/SxkjS
45U9qN4FpzfyO/ybWakSjF4P9b3Ae9OsO1o7pm9C/weCwF8JyaenlJTZvZZD6RERldMpq2jThzF0
XIik3HSN6nXw4jegW34KbzrY6i4Ur2fSYe7rz7kaIAN/FUBQft2uw7lfdI4e+9RcS5VYWHLslKRO
CjFwvjlkVdX3bu7Hxnh7lplBLjS+7fkzEOPJXWTh2n6D7JH1iXg50KzB3fhnKdxC09ocf5jZfgfa
R4m7A/lQ9OAE2w8R4fqLFtwXeM587Li53O0/XsDUcxvEzTrhhmaD+acdwabzGxGbyL+h8BA5oxBi
udz4fAzzZ0g0HNYDukoYJzqJwUqPiXIMUKnBx11uf0c73OjArHNtOXD2cDt6l+aDWKUy6TmK7GsJ
BYL1/1f49igEEr+A/aDp9jKFkK8iP6BZaRuAIcu7+1hJj3FZLl++otuzwhTQiE4PwO1ktyA0zv7W
/Wx9FZcRl8yS4p0vSaid3mPbnlpggrKpoOQ44Tz8O8HmD1K0eL79Jy96/IlNCDTeqCmwPVi5LagU
ys+E0ifm3Sz2UwsBZH9A3idA13Gce8JrkzFfJREuEsASZSolXs+X7JbDiUZ55kzl8aHOniMKFitF
1OyYzU9M0Gz1ffz2LqWrsHy7zVphO1oVMseCD5IBBT8ZI5B9IRMi6Lp5h099QaHs+GxhQpqKAowB
+yVZHIADIw/tJsIC2ll1spBTA84/jzkTScd1p8cwTyMboNmRjzoEKnCiXFhG+akMzJBlptUN3XY3
1Gn447PSAJM1GajdZ9RSWF5SddRQWELtCC4nyKoTBYw5nUJ8AIRhyMKuP0Jzo3XopZyJSULXuCcz
XySExwput/3rEfhfQ/mAiBz11OeJhmNx9pFKSZsJurzD9t11eP7narfRRxVMDvtYMBBM302d9fij
kTbwiiCTtBYWPo6TTOUQpoQyhCKlcFu8SfjWJGazN9Ve4NxGNTpuYaZ92ru7BuqtfhwtfYDu0qJS
MH/L4Jmuc2r4QgzRK6QSf0NMiqvDgxZxgtENMl19UkzQMaxYn1kkA/Nuu5rtI0c5T4vaYcr2lbsb
z18zNjCqiy5DjeYqS/uqWBG6hb25E1hvCWgYwsKxICOvpt1bsDd+J6juCp62fBt8Bsia14bmuoY5
S2jWNKpFoMB8ASH4nsPwt9bSyLkr+cBSTIZPM1IbuZTkKgDPNoJ0dPGD6zagi8ogHwLMEgaGSzwb
PnNU+31Rdlgk0T1XsuxaTiMIcQzFbfDOnCBt5uJ0xPEzSgPW6R/1AxubNoAxMdkT00l9Jddx9qeW
eXqyvDpBxLKzOTGE/yGf5IjaBRCeyI60KrKyiqXvi2P0PC43F36BcVgOtQwb/kkNUCi5LmMXXLEk
zoqT/hiniqofQpX5/cZ3nuLhI4HbhU2jXAQ4FImKs2ScX0FKeKIi5I68KdzchCrBqTLqRtmzMiTG
p/RHiF/Xz1Ro28n4ZWoFteT2YeYEHNE1kb2cD10wxxrQpzQlIn+5v3RpVvGvGiYkycxi/h7YT5Bo
nsclvoWfZzRrhE/zKIW9QftLAuKFX+nNdWAZVOb5jZRoU4RLMllC5kjfBX74ruttwMNu20zcRS+n
INpKvuZpEHvQoUlQEup9fVWhkHl/vLInvf7D+z9wmoY4uV9GH/7h8wqGy7ay5de0s3JRrenXpHPm
5eAE5g2tsSflVsUJjX2ijacO7oMGBz4UinyO7ouZhAHpSzHgOJirTpx/q6QHmjJeT9ga7Ge8Alt6
1fZuGfEj9pWrOh5wh8twzti0/GSNkffDdzsWAb1hOJznKcEh0LP/Ezqz3GUgSKyRfZchEBeBuFMi
5MRE3nIty66JPaD228jS/DmtThummvIkhy7Lb8aELgnQ9Vi/SfDDMvsOjKujqaBc5qV+aSol4okP
nK2R/cYV7gmUHaV4UzdqciaZHQG+MrblbRVrPulgYfUXnYeB5UU0ipnusQz4uKxisymGFcxa1zbN
j6iBP9oIA63RvLX1+Vg4Hs9zsjXmEt/kwQ32fkMomxDRqodXavSpygz3VyJhdbIqvC6Gjz2UAFVj
SCRJpnoyOGxIViMusWm9ckNdbLaQSmBjQbeBLlAc2Gi3ldCxJz9KF9tSTnwZrGZurSU2eYeKXtQl
cEWZzLHgCrCV9/xPc9Eem0+vl6oKTpylTDLUTy9YwE6nZ4x9sJsgRS6t9/pmheLbLPd8RAThaFvc
QgeLt+ultsXnNycwupumQ8LBmt9fG7m6tXlVTJc/uViE6JL4olqJLXEK4Xm/5WukEBr/ycZUuZYD
RY4zX1bTAfaeuaUosJQdF9Nf1uO4pq8bUMcz5Xvqo7wCra8Zh+hRc6ZwdBREt4MnkzNEELx2KJgY
a6yymzVAQw5hYCvXebFOlC+kv3J+jNlyPEBnM1TWFQrKsYM/n2rbkgNHJXL+Y1h9zLZjK/PY62im
W/jcG9yFb654hRlS/blw0wClxme6JDP5yVtdIuP6PHyzmORrQ5ytIqAvrzKdqfE3oc3UGDBGdVc1
sxEX0r83D0OqWycwtPBBPrSXKLyCMyEXZ4aCxRPS4L0/fOR+vOUWzoVg4uv1IXTqJlokDPu+jbEs
ecJoE4Hikh2HzCCDtQSzsIb3wBYEnFGiqKzhpFwSZyD1NxHoG/GfB813k7VbeOAAPuVIiyZj6k02
uv9UHJIgFXHogOJCX5Hjb+ragqnb/2eU7ZRRh2rlMhHY6bclpZploT625f4i/pqvYhmaybAfBcYq
YDnOJQ9VB/lBwF1WWq6BphuNvLYnZ5urasiM5GS/KPUPrSUGPWzPe2ns/CHJrSiGoGYWrUgFc02+
P4MfK3mJgrzfIz8+4hh5iu7DBCzH4NJmQhiWUJB6UmpoSenISfsE+j7dwupejfzqAlqFfpbrZF57
FkbqdHI5fjmetwnlFw/9NAKDwwGUIIxkWUZhhCIXg3jjrnoEf1gMYxEvJXAf49gizP20onR6S4FP
MY8faHz8RhHh7TznN4l84WVHXD/5EXA9VRXSIJkzMx8e/3jpvEIUIDGJx0ejvGaAf77Tz/um2c0+
TmVxdWszl5m+1SbSkHwV0OI+mI5QM1LhymhQ+vv0DJyX85+9lpVQWSSYyXTjtsbVHDRbfSpeHi2j
5+Fsp5G0l39ZCmvGlxQe3nQ1FNur0Mc4SJz+H3xwT/AQ3AEQtJg1R91L1PGlPQ0eJuB6CZov/50P
yoaXiuupWmuWq1FPa8BO0ZRMjMgadfuLOx/XGZuuBBLS9rU/FcGo+4iB5Vuip1CKj3KsXpjN6ktc
K+qI4iKTcUBWcON0NxEUUi41lkycHwPlnHA/TqmUXL11aT6iL55IQnlSRBmdVN8qlmk0gZPza2E1
HjSKGNmc2Iu6h0NcpuwRGz9SnNgnZ2nNBEHEeSDkdlieZiDjCYArS1tBPCWJOUFm++pMvAu1s7ze
NSQ4BMMqH5MwK6qv7ltI9MJORlb/QneUtipNyTkLYtzWhMNWF5QsIpmxPKAR+c0kBj/nECSd8txg
PlNipeuo9lXF/e1s91FgRPFYIzLNwGmS0lSHSPqIgVEqZV2YO/UIMBsTmM/3azUAKmdqyGgoVbkJ
m1ju1AurVkIMEfoomjYPE9kALzQ6tGfmp/Mvw6sbWjdojCAdyz3b3GF/IMKg92asRoi/HGsF1o2F
UftSsJNgjX7quRKOVAZ10VDR+AqoU/ChH2xS3vEmo3U2teiYrE/BsX4ctC1I2+h9yd+M7bO1JJV4
aKUlFJQQOlVaL7ZAVYVwAf7ZsH85CFbERVR4da1i8wxCq0LK/6ARBhjYRVNfvImy46MkDahc4hUB
QhnuvJiGm2jQvvHv3amW8ZsGwvfwPl/tYLYdLSNV5zQoswN49Jls5YfufHpw3uuSaC9b/Swu4Oed
r4cjVCZnBKh+x+c7K8tx4FTevA5uDdsQ2w/lr+EvPzACNxMp/3cn583S4w4Pjj/AWj9hkSnHtcBu
SLd+rjFbO3tJEiMhD6Q14/TqgY5VxtrXChgnCcn8tTt51LYLTkknpeR3PGabICD7bzHn12JMTuLp
73bl/Xkpo3Bx0zAOpR1kwVtbnyyYEklwAVnYe3y7TJ+ZBazRfk5z8VoO0q1e5Uj7F5MxwEz8T1/I
uDY6DEfYK9wWIy8oCWFfrSiFpkutWt3CSN3rjIUszNfNPQTV1mSJyhwWKfVPqAvIjeKgooIMUed/
qZjD/Dd01JD0TqkmYGMBd7DxyPEeMAIogR9qLKL/qzw6T8VAVdmyYW5Pbcg8YKxyiBr9LjYe8EXj
+n2xkqq6kqxTAVgjkLTMyEvR0IKeKZ8+Kmg8I0XEHcyrAK6axoNaI7wnoSEG4IUjJIAtGhatcLtP
+TAkNYLGvoIESchtvHI9M6fOi7VnPp6PXqRJVCh7mXSX/URRh7DkwK750L8X/MXius8YiUkX0dtn
FgfzAD8PqRtAysAgya+aP8sRn+8waljEs6Cirj/lYIizIEdoXLDeFqQ1fx+hXph/X8+BQOjFFLX+
JsHnsg6aSXYsi9zNwyuPWvelR5afimxNy3xabmDiq5MBsjnWRKFYt5jXxc/oXw2jvdgGuTEc6Ex6
eueCUC2n8Gl8z680Ol0Ctptlb0ZYCyouKQ5upmos3dzBxAkWCdamZVVjS8Ff+U7/CKFFZYdeOWlG
b08PWGY9zzxf0snN7XmcAB9DLLEvfvCeP97Q9vF+Q2ZHu0xyExh7ohMeJyfKCEht3JN7B6l5MUbN
KA20ohKePqs1W3rWC5HRoTsX3lv+fgWMEQhMvQwpK70o8SSaBkfkGG9fmoSiWEN3TUGSD609DpFL
mVJ136ZDBvGHjnTfHJvWlVofaulZguWxMwdAgEo2Ob1gdVWKyMNj6j6TuN76+4JyJiABli4RIxBZ
sAT1h1+ZtfeGP6fx4bHU4h7vkAXjHcFkLxfXjm4zokn4dx77Qk5j/Ubwdt0EvAh3daHHCfNU7xWS
ST4mja9/c+MvNdLe36lDyg/XfdSe42i1DYbxbIu+CtlxLVvU32BJgE6szl5rP0PICZbizrTVyP5x
/cxk1f35TnkW0XH4xJaLDEtxnBn0wev8XNecO0tB7x4cDcP1kHOrLN9U2WPbBV2FxT0626mxDdBl
iTqXa3ZDbW3jm+XiKntkojrxUyfdDSiLHNquURhoDW7MHrUDIUYdNMXRDpbWfQk+BP220iUoKEDJ
aVH8wKA63oCOEHA0MXqkF6Fa9HiyRuKaHqQtAF6Dsq1HklAucKDEXNKD7D2pmayXDURvBLe8sAJ6
imDpyc8X7sEI0q0uyz/UQ2QaDTqiebwNZbIF2ziVs9psViETXFKaaOssl3aQCLnHrUuEbarN7fGk
x2otU69hXjieFfNN0JWcvDRGnKCHWAryoqqitu8CqbsDgLGEMEormtCGqLQ873RhMOT2j15dzxkv
zKLjtB7CRovnsDasEdwoBUzFTewNYoCtwmQ8GMUVuIgzea6NTOexQFSIFFtedBOe7hDGvdTqJt06
PU4zFE975v4/oX783T0ml6fWkjwozWtyLW/l1iLlLcr3Z63Au6cDOJU22/NbQx1FC/TEmTMLfi4B
4r+kuOt7J7YS1SGm7qkRU+A4IkTEW0tLXlMGkzhTy5o/rft1NUXVMeFSgipg0QlIYFK0CSQytAWE
Vqw6L5Ow5J6XHEjh3mGmR0tNJDCSgqZnveuC+M1j35kR7E0kKoIenUpSkKnVYrpVW13fbcoZXIpA
8f1CBcaw5MZ1PMc/pXpaMs/hniUW5YopT7IKAgii4RGX1LVxmD2jKi5t/w4H/j4nITPki12wgZJi
TXgsZbrWT6LvNbeVSx32vMHwhMYhL+0xrEtdZaTsu3QtHA/r7GiXl7eleZaYtrDX2s/xiwGg39Im
T0C/RhUlVrOmCK1KntLz0ZMy1+GUgiT6aYhl1Rk4Ry5jkADQxBL52VUZAmNF6ULHmUKzv+bhWpnm
ATWIkWHstGgCU1mJgL1Hm2IYvlI7gZC+Zu2cb517WAxyGYTRrXXWoYMomonJlsPweAaHCAGBuZQQ
LKxnC9YD99mUrP4YtEWt8ZMvz94msFOtLMNyYEU5kCByVKAxuhFaGuFYK3/Wxt2gZmhjXP7u6tcc
yv9YY4L23Q+LKkhXy5n1cvPjH8KWQGlqOxX/qBeCUbvw5iLZPDEKYkDS1MnvolgV2/KpggfyudYm
ustx/XNMRUf1vb2r6mlzJWf/siA3x246P8PRQb83c77Px0H9XF1FKT1mjpkPRNyea9VO5K8GyWbQ
c68TDZnK2ylq5PNAWDebUn0C+hUqPsfgFHetKmOUy83jfy/ZFOrG58xDpLmM09gdhBxiqqSGd9uu
PjEDlVjM2Enl3xJPgEnrpoxjkYcvQr98iBhQByAsBsq63r4/lv10n56nCOZnkn2J6zNHQDRdnXsV
6YLTZFCWBRjzjX/CrVeiQyIXemea8iaRTxriEEou3UxaXNLs8eGbNcsifxmOH7tkQ0BMq8aMbp+j
4Rzk1SCirMw9C6pFsa9nb1gORD/iBS7x2kxaDfpBPwH1xGKmY4R6xD2w6x6RuFPEkZhlmaN3aiLT
pK9gScOxZUXWMNGlFx90U/pxNNhnGkTYe3b2KWhY0HMwLLXsrph/GRTWq/Fng8JkmgzxArPP/eMQ
7O3sTtE0caWIQ/xgDaJT5c5sNLVLQexMnJ0RA1Z1EhVCnhBIY5up4X1TnKwFmDwFJkj8VVayGX21
CIshBeRto4bi3Tq7BRvrWwoqMsc8IF0kSezYXGbXFX0H1ubFrCqMxaApSQbtproonVcq1L/kgVes
UBN8jLjbSDUn9DcbomdVUvGkQtNkDqBm8IfcVW6quOrFwwaL/64B7uvQTP2oNl3yuRS04GoDRk0I
vX9v6EzRevdt+dhVKORfW5mSWhuUT7OZjPl46IDJf79EW7SKfi4hiafl1M/ILTE9UqFqM0MWbf/I
SH1BkXGCo7LslcXXjME5ppIYt4NgSXc9pBINgOwBhkSv9EWC7mR5ioA0KkznC/Cq9sI51Tndyn7T
GtO2yj5DcioBfUnxDCg7KpSZheqhi4/crkspa3cHlc7iZ1MBckRm+YlqzXXnR5HhfsDWR3Ym8D5b
/ll/8FrssEVyReFLe4Twsymso7dT7q6E4BgWkxrKifu+BWDGPAKxCaUO3wc7Tsr2G4F+rHG6tHst
At1Zj35krBZZdK4ArtOEELJZc78n9JUXlwjEwLaH2t0gOAwkLprtkYERTk0oLXL0as0LpPxpk2JG
XSQ1Pkb2M/51aXeLVFC6JtHHtHdWKk/X2Ng5c9ypqXFHDR4eikULl926JgwG98aQ2GcOaekS+0aP
4H9LuatSQCtL+XKrCeu2iVN+WLhy1Np58FUdj+oIWO4+05mdHJP7+WyLz1coOJ+e3SFcPlCByzby
kWwrL1509BMEe9efic+Bp4KQATVsz0TKbTJBu54DZK/X9Cy5arycN7lCHA0/2qaSMOjoDra27t+k
eDOMySJiF6iT3VI4J27TB1gA5Fb8kC9gDB5wYMCVIpvyb6vhZU/XGe8lMPkqY2N9/fnzNCCSOOcP
i6oXJjxUU8zxd1mX8Kvz2eppvZeFWZix9/eFFkFMYLHNyguiKXRjLxCMYZfRtCGY1QlU6EnxsbgD
tiuwYhbRNvwe2A0t2XaG+ATvHzBMzzPXRL1mpc30wldGfsYEPCm2Qr1r7FT69SvkLGDL6mg2ld8i
bfLlzhzLXF8LRrOqeGfJOyc/IpxwachBsPy0ViDaqJSwzmeofp02W4T1gDf5kfpP3cz8QEoorpSz
17chcusgpFqofTK2J66Oj1z062Rhqe3NBRB3h0S/SUOxrbiXJ0mcPojwTJoemSDXGedXgJXLCUzp
AZQpDGd8T1qbdY14PB8f71ikkwjdkWAnju1+Lx3PdWapDz6J8L3lmoJa5925FR8xwWh456YHgwXt
AAdfbxmY5rXE8zfkeXa4CxVlp5a+EHWrkzlBCd3B6Y48CYyeC5QUC5F0utUA9zLd4I0O3T2G/GHM
oMxylIkVgIYGQZ+sSfELK76Sp4f5qtUvCxQ/IWTZUIAi/wIWXJOSdCoxsyHAelwufnn4N2k23CBY
MMRPY9ELj+9FOPRcJAyzq0zi7lrI80U3Xg7RrBqiEnWh/NNYCr+2tCwK1dgy6vfsreUtJ4w+jiIv
K135qur0ZIVDDPvJkUMnZcUWVQI2ViZTU7bd9JZiKls1pIXYsv3wB1227DvRcvpPe9TMWIle5mUe
OzxtIzilc0gTF4bfxS7evKzYyOMVMIy1eenm4xx5GxK1HyYzsTbPwOk64d0H6kZzbid0odjjk2b2
3jd5ztqmzwkdMA/tuAIswz8PfZMSG1YGPje1X0I5khqKu82vc3ghZytkydGDH2W3Gr6RxBeoEzhY
1vcPyaAhMoZY3ae1X2k9eaeVCf0xSOqH6jVSBSxjrcTGJLPgdGXb5+HQxpT8h/cYTvbn3n/dW8bl
HQZDTZxSReWwZFdGPZEYAqxyo7zuwYd/VawCEVSVTAFJKLAZnFWFIIA8p4vb36MA61fDW7YJP80U
M8foWydmaIVnchTL6am5dBBaZoRFtAkRju189RUH8erjZnun/bTnAHhsiudlW6w+OObM/WkvgZYm
IWH336N8s4Zu8SCUA2zd8Y+O4XArlLilwRyQsecsT337T6IfIfK0NkZCELAbAI+VStOVIR3LfspT
k3nySOhj1QicCUu9OWQmPWWgYmQzD9giv+Vre3Jdy6Iu4F1OJQKEb9X4JC7WxizOOPVRYIJCSO/v
XTJLzHnob8tp2SCFenTbRJUKjIBHS5FqcNi1SAMzi9zkgxMjv2jwCIepBYyZhMpNkVelm1ANoWa/
bQfVe/J5jrZBUgzGUQezLPLHhhZPgIBOwDhjJ/0vztcAhY30/eJkhFsYCXMg1xYD8pWHywhhMOco
7fvzVrDsucyVeKzdwnEUgbKFFLG8z43Lhk4GxL7y/BBxrcpm9CvgCtJyKCOtTn6Ev3JngM/7H8eD
QWDswRztzXtF+g3i8dLQ/GkZ/LOxBRDguqLHMPn2hk8Sq/OOR9gSpZ1YX2YnAMqXK5RT6bm0U60I
ZXJoqbBcrPCYPh3AjEq398GTcFRTi2Xy37y4OoV4TMRL/3w/kaw52Dj6kMxF/1NZs0QwNsdxTiC1
KOvFeY/g6MGSqNW0Ky2rCAEFysy0fQFU4qlLM5qq+3TOw7ZWdV5OVSfCoWe1ZQIR/IPAUsaIQMN2
AvZm5Ts6E8SopP7DqIcGvI+sbijkraJ57bVuHlJhum7Fdqu2Wf34lJ2yOONoTNGV67Xvs5kUaRmJ
dsbLLI6XyMj/2eP4h2ZqVaN5825G3/QhpFjdTIpUdmowm0Ji++9KC0MR9XWlpZwr8aRuAsmGVWsy
/7iKhAHTjf4gRK+GiLvfwW0Ik9y7SdcuC0kCry8BotqjgsU2MEvHEZTrII6k1MIgyh335zjQo11l
wgG1WIyE3nrRI1riqNfLmWQAv8+c/SGgtg2GOJ4Z//Alk6KIAzPB2ZcP2uTJVJ94ZQ8jZJTCtLwP
VfW9PiBiVXmfLHOYnmtYaWAOPv9L7p0z94Ic2Lg2bNJdN5DtbExrVLDUJzhg3mnEtyM1CDjzurR/
L1GeCNiFl9Ej8kp1m0rj7m9Ubpdql2AKlEKXJc8gbVBPIvpo8fgJWYud8C//xDHu/3y4d6ViX9aC
oTX5x6TMVPgUKqyR4SrIGxVyjzikMzwxTQ+N6VRsNz8dfKWc4X3/+Z3Qxl9mU8tZNgCHGpaVzGgq
znSWd/B+UAG1xYrTuxExqcLfTLz/gBrGvPAFsIB1Pe6SKp2FuBUT2ZxqonRZ1xDn6vbOpYu2xb6J
FE1kPBFMCyvNzgu64ErV6gR1/lH4I0Vx1td8irXd00dY8QNHX+E1Ye25f5oEu39WC96fzY4AJVtH
G6eUZkhDPkeqDFhqWzmkOWFosxhsJPuoBy9dekMg/XG9vJOZ0uvoLlByCWDrUWR1W4FqeTJx887N
9h3itNWbZgQY73aIJ6zDn/8PxQWMFpYfd7v6QQ2NUfgk3bsYR7u7jHuujECSwAb22iSdqZOm6sFQ
ulxZCuVclCNGWUQO7lTsN0nOaIIsqrvowIELLj2FbsnAVG+35yk00p4VvnLUFc7n4KBuGpcqpMT/
f1UNFO93yrXNKYUNh3sBNRCQI8iIM+b78HYyM0W2RTWhl9ojzWGMwVmnHvqjxJ9VUMqEh2Kpw/O7
pCc2GX5D621nGCzwtTXH33o37nmAzB0vYDV410p5D/2I/Gkcu06Jx/NuSzGfiLduY43KUXG5B7ec
boNiJienZ7mmFTvsgK74yLlMRVvvQULqZoUI9Zy4MveItjybZEvqtL/drTfrS8FK/I68xIARxkKM
4E4v1SvxUyp4/kdQvjjUjFiqfwzwGG4FYVHRaJrWdn7petk81d+1qC4shk/n8DZKv0KiQzbGR+9S
El3df49uYI++VG3hJaYDZ+D+Dh+BuOIVpXVa+8dIvvM0Oq12H04dEKuKiAEih5CX9sI+ENPS2N+L
CMTN1ldtz7PEuWpTysQubJDUWK5+xkyCVvSpjR9B3d9jD5hDGs9kIJtubfLCQDVfFX9no5nX9gQs
lrwMwRNvW9DHagCH1Htra3Zvp0Pei7RDdUz9lfHAU2IgqtQ4m1w4T5qGLCb78PARgVyVIvExIGyL
IvgEEjYgUEWWKZiwT6hDwFs43qg6PHJLpMlyLrqekTTUYvhpLVClPNuROMcFMCdjUKZFP8O0WOe6
KfLOxy8NN3E5wKZnvp4CLdLPEgUr14OcE7pXbFJzBmNR8gw+AcxtNdMaFhw5CGL5oC+fxHNnWSja
anBTs+twMa/pTSb8GQfjIa71ObNNFYINCtRz/Rf4XnhjgaHl1ecUTj5hyI7BNstwalCQgp/G8nLi
3nRhQNdyN/+zdpCBrUVKJozaeCQWflm04vKzaivtx6aclKnwsumPJs5CgQKFZGsGVdWMHpJ9PC2e
7QYOiX/n1ds56pMjTOo8nXt3+StGX2e60Xxe4Tyw81E6tOgMr3/NTjxqBJBBgKPGaG3zT9cg3XKn
LuRwkI1SGFeBN6jQsmUWmYNfvMM+v6dAbQyUYhoWo5BjUfLlyhdZV0qRigJE+w2xyM1vp97YZ7Iw
uOCs+4jCEKdlYKkqYh19c4tKulgu/dXG2zB+XAJrMspQXzzdM6oBKLg+F2PD67Px9+g3gk1oT6J0
iVs3p0WsFDN6nrA5U3FetycWiOXk/f5TDWGSteV71vTfpOCA70aFtpnk73DeJfls6qkSkj62XmCC
1mOcLfUIPNwSmH2GdWPkWQkmMMdjuLWH9wTS2htwH8LiitVZ+JBeF935ND6ns464K/NrmvXiAmaA
J6M2IvpZOa/lWzswS286dSwaLb1//H/XF/TJ7/CG+cKzPXJvLXtD59IEIR69QtkDOVT0EHzuRjb9
lcwCAmRP0S94JqokLKCGyfpyi5D3h2txifw4e/8Cwzo4E+DmsW6I+bDZe6P/5KlYKbZ/e4VDirFM
eOQZelFMJ5j8G+wQ4OoKkmI4MWDZqFMDDsfLS3dck5CVpZ9LlFeTi2qzJi8TVm3P7sQbAXNMzl4h
AVpd5UcJqT9LEmi+R4PVkrk1JtfYg6rHhCU0TIFPP+YiU/fKazeNYAyv7jOQizpm9iUPDkyBNgIy
V/PYlRZBJJYAl0oxLYSMs09FIIeERFJW43HyadyRCc9MkWxIrs+Y4AR7UDXh8P0duaEcpsmqaJ2X
+knkCSdD9v2QxqxlDJKZlf1mxGjN36C/gjifMhKCCbQoOzyCdf4hU4nJ5JJlWH+AdNnPuGTFJVPW
0wn7IiI8/kev4w8SJkzBTMyux6R5nSPX+HsNiFlAI9drFJTwCOFr8GXfr1OQbNtGQDg+RWTSVxLt
SlAfRD66mvNO6GHMQQffQm6U7KwvxV3rMpn0nO1wqLOUGbSA5QDPn68FOclKW7wayIHWHYQHhcON
x3zbdF1Rzq7gNRMEVMuav/AVfP5rtyJgTe14dqFrQBQ89YYm5Rg5i7I1fcs5XGTBRT3rfetra1ws
IYaD3I5AivqsQujWGHK5RGG/aB9mAshOVBhz6ImsDF7Ps1xsKwnku4ohQjMcTDeVRXgKWcBkUeOm
RN+crMQoYOu7kAvYOeOdb3uahljRfeRBV+KqmRibNWOghvHN9oI1I8Sc/rKxE6ndV+PwJ73Byf/N
CovvLnAVeQtQWjXSFUItQTdueJAKr8JiMdZG2gswD/A79LWdQFosV1ob1k7hDz2Y7g+drDfWNGhw
4bsR1DYSplt6XihA5I16qLlA+6j6t7cv3a+scbciFrlU5/JKedwqRwx4Wq4+jXRuzwRi/BRiPTEI
ws4XtAtTd/HBIN7/CHQHCKZ2YkhjfkpaH5a1mSET4co+ze/3jfwrr8CQ9TZLOhAiI99A3IKsHKTK
WePLUgbqa3FTxawWk1CdjdW2ZyNy3IkIimJ6f0bigxfOHr/f8jGBp7ix2PyaV8GPvZ1JgJ2vj1bN
6+8yXifxWTFIJCDMfkecT8XcKLdSP7n5cbhRqy5lJEf1qFztPy5b8SOxkcvsDYj0E6zZvMKv4dY7
MvnKaC1Dg60zp1Wrzy/QfzJhfrxgL9bBipQt14E7CT4M77pcJ54cMczam1Kn+kPQHg9HtDp+QYet
raapOuubogi3snt9r0h7eqEHsPMHzdIKbK4Ed+kKT0z9cgASsLkzPvvmhDH4ydzb5v4l8AipVasJ
FLekKaSxDyEMzUf+TYPl4et8YvOUVSWUS+8foU0lvNdtAo5B5Mhc173pXkkkHLpJREAarL/OKAos
ow7wsQf4/s26Mxe9OPY853GBDHhy3QZtRKyNsh3a1Bywrb5PtkOGCyDpEI7JQ6wG2TeHpZzTyb0g
78K+nodZe5c81l/ETKMIh+GhjFbghhgXN2tl98FzTSMFiSQ0lDqiVflJQu7FKgN7+uMeIIes6Hk3
q6aB1QNLZOZpQLdldmeQnMBov22Lemc1sP/wVBMF2fOMXKbTGmNoApEJW8XF8ZVtWeZos0hb1uIs
vPWQ57B8M98XRbs6EH20gfbauMeouwA/IJbIGBrXRc/lP44FoMObpSAIGzf2X2aEBF0JP+ceZ80b
i4wD5MEcAtvwcEiB6GQfoCbt11hRFUwGDGpnhKXxanXIXcXd0nq6J2FvIzXhfLH/TXWpvIjqUcdB
84fvmG0Gav4IzGPtQUzwmwvcKS2ixj5U1sVPZdSTZuZjtYXRPAvD+qvFfyFzbJ9sPBFI1Id72v5E
A2D3e7+2D23e9HphU5ybPS1gWNOlCJVdl5eiyvFd6PqLgssesYoKuYXc4TSsdbGAiVwpTiQgXBhJ
tqFwEhikmEtgYRGEzysSQ9n3/gFRZfR1bA5mAMD/W4jp3LyXIJfYFf8IdWfm0eqdwg2fHbyPxYVI
lsIG/CVaKTCC84zBdUVJ7BIRS9He83i6+927VbKkRenljEkvr3YleCVTNvGNJsbtO6sDYJSQFwS9
HUOfcECigE7TXUHlHJanoplVRQG8ThdvvsSNtZeNudgwxKrsf58tXdahd72o+vaEwIvWJorCdC+T
YKo1FzbV1gmsAjEiMT07x2vN4gbaweHnrJA1Y2lv02xtrxJ551ei5WvRrLrcIXv86+6Rq4LuNPEI
vEqgMkNEb8nwYF40qh17e03yEfcsW4twc52WdBjOjEu2si33UpEt6scnbEaunUMpApWbJjW6ycwp
9mUxplnVROXMA9FE9dEYHl+hPwsxEc/PW9Ct/uzHn/2V/MzZUs1G61G1kY4TVh4PLhY5oV9bviWm
xc3WD7veRfKhYRTENQOZT6DioFwA4BERjeOBLosSA7xseQk/zGjv76fJl8tN5zL6WR4wCSXRtZfX
taNvyrz+/kk+f+Ui93ZyVELc8kaPYOcaopEdqwOWoGZz09DWXDIEUyE+ZiKNJtIIVlgCeN6kiC3r
uTW9sUkCn2OV33DO4Kvmuz9fOzE1Ji0Cdbaacxs49rQd1eWJDEQ7GnbkJK0BtS0QcESgzaEnzN1t
GLMEHzXz5g9wiIfbtnq9u47ZsbpSOHJT7wyJSoroS6/hE/uaQ7LBtrgtonKa1glreScEKuIXHgJt
iGtcIhTYosWsI3sHbl1hQkB/klyahmlgcMBBOmDuT+5ZPagCJ0UKiUxqaBQ1aSDGpK4JubxNhZn6
lVM1sz+kD9NuHuRUcFhcve6+zjkEb0+ggORe711MCZJZ+kRBYUFFIBLcpkzKzWmjQOpEtsBG/M8J
oaKLLF0e5QaUR5MLQ1Hc6kmmIoJ6hYpPDpcXAeB/115rhES/APeOUUeALxmVqbYqRq7fQQiqDw1C
19Z+KQy26M2SyKUyMOmJl7QXOXcHyrKTvr4kzBWBjMz52JkuC7xQRdDNcNBa7DUG+we016VJCWkC
VCOzTYuy+0K1unvVWyZkMvnLZ2iC4gzK3RjAqfREAkPhRzJmJi6ud+7fmMAvZiVWCJVU57LwiTty
QkXuUsV+iShYlj/FfTxXDzISv9KpKqbDUt3lZrw+meKKIt16Ier4zAzwZyYGfsZv0mlQF8x9lPVq
wLPXdcrIfXJO93DJSrWA78Ssw5wp+T+SnpmJSNTO32m3Q0eJ4mGN5sfPnCU1P9BjT0uRL91Bb/Ho
zgZaCPcwQAaL4xlfxBwwTG5MYM0OrS2lximCX6DfKfITShPvx/b/98ZLOHZ3H2OrFNt9on3YhSeo
72oIcmG7fu+OEd2i+BINgZAX2Eu+QVbveT/EirNCm2iFq6Y+iQw3DKMvv/CpS5tVZ99EXYKzXkrL
9VPzOCiAMOhMiIg1cA/0zzIZ/T0OgYLz6qMR7iqhH9epJ32MqnpSJICy/W+Pt30gxRZ7RY8+OzER
E89/sQjaOr4hByHjQnwSVn5okHb6MNk/0e9k34o8fKcyzB/y7UWTkRMFElFIBqnlm6zeMRuvdCuM
ZgctF+VX3BzjNg1F7WMDAWtREqotI2ngORAnIPB1JvJ0QEdEHvz8+WMhBMZtvTjZNi4GY50P94FM
jl6UBEUwsNojZ3i5M9vVSF0nrRN/OENoCvEQ6X1xqQosXLAV/ZHpqf88wb4D2jgMcwoZP0uO7wsq
VRr9nrLedvjnd37bI8aseU/dNLnBAH6q36jd/8SSF8D4bzb2YC9R6byokg1EryDjoP2lc83o74MT
e6FuGHQPQRX/olbA0tXf4lKNXACAUwnvBxilPqxC4KeCZ65u4CCHDPc586OnXMmxolTGre9+VTZT
hBPRoNGThYVZnpGoIoqLn166hIqIHMu2s0M4XMNJIK60L+8EdweAfgXkt+KdD3u4mblZD//bFN4+
qoyl55QvzAEtrZy7nJLl8xGa4pUkze8432I4QVuYx+JgiDaFpRPMx1dWRriI/sCCZ+71l7gmwfrf
IYY6wl9bKTBB7cw2O+Hi5NJ5Eoq+s7TI8eLyf5bWZ2KB4CyzWdqk29DIyOlpNn2yLN/8s7XASL2o
icy7y8E6WipdgO3GERMs//kR80AtO0qZGgEvWY6Qo7AGBB6IyT/m9Nq4zIawQtv6pDtDHAMVxidh
95uTcY/nq32qecXZimz2qSK+NMT7nHGpAwRfAsjHx8mePWMtJiXqCiIu/8DCixAlC8RIqcEUzlYy
B6uOrm/HKoOm2N1TtKm6OX6gwBXxzflbYW+wBt+gHwVt2FcxZW/xmSgsgANKa3Y5yS8bqMyNwoxd
QiXCy+yE/uYMngrcxF0H6KTbdrJ/+YtjyLkm9gkxta/Qv22oj98hzutRVgotccGNAX79QbKA/zH0
CpL2mkTqY6skrnDdX8OznEUxDzxNvUW+Gm8WrsNhzcY15Gx6bqyM45yi+bM81hSw0MgpL1bTrc2d
iJo6CcXerkVncYcqkkUG318C7WLEaJ0Zvacs7+Vm4f11U9XcBROHO8uSsVBO3oQS6kLTUEF96xdM
De+plsE8S5Ob4U1qzEId0DSKiDoTkzZWpE8fgH/IZhaW4AqMS4viYp6qI6Zktvxn9fxz60bhAbV8
W5Wcl+cTAqFH2ngu1MwDLxgRRkazFH40tHJnqNhnSQWhwQY+yakb/wl4gcktHxUilRn9647++Kx2
/JLq6ZG1yXFgXj9zdQaaq8omdBrO+3GkDlJedpE70PIiC5VhRMa+XPM+9XeC6qV2qlRE+KbLiiSn
QKPo+Ly/77lu4OlQ3BR+lgtgcek/RtSzOYqQgxvg7lS/0hDeVKMx3AN4LeYzWqM2czoxF75Howq4
rSU4eTXlAMiKHde7ksM3Q3qgiSmeF6Lb9RJtE41mKUt+b4qArGd7ecWvzmHUxNg6Qh4txwR0Tp0A
YU1qjIYgGfuj5OTCITHNOBpOaUcLAB9aNh/6a6iWGQEPle3C6Oz1g/NYPIteRS+LnI59VBgAVGXO
3EnP0f0J8E3irgdMoZDdWyK1Tosg1JXx1UIis2V87DTA85jFhluiU0j0WoISc+ax7WdU01S9ARYq
IKG/zVV3frGZxUvwK0mLwRAAgiEtiTJLsb0tUxmL91TIbaFSp8BkmJ/qL8EODCmjecnt59hiPjTf
rEH6Y8A+fEi3kRTv42NnXRTxe4to2AePamUFPHs9iDtyEVhMgdsDL7PppLC9ixTWQ0S4SSC7sWjc
P0xgho1CXCzhlmnOjFaXnOER4Rba+MRUOAXyCN9GnH8w7yOSmH6RbfmXDa1+FVY6LMTleg0lEnSM
fRMIt9qzDbQ6xdnH10730psHH9/jwjprHHlvFEnPUbD1uyrYoUMg3P0v3B3blLMV0YmIRZXZi/k2
0Aa3MAHHOLV/uwW+om/8mHzIZFPe2z4Y/LCkCtzAs+ulHRoBSc5tHzyN8Cq9kJ5a7Lav+7IAqYaI
YdW5l8gdfYwCid0dkMzib8+Ve9O7qflKM0yCE/+lIOwnZJqEXdXhlJFFoQiJaN+MWRSpXpTyJLK3
CwBymAaRHw4cJn1B2r4haUINQ1tA0NvPYQLKEbuP5LlE+8Vq1KQ/Ca5xuOgur4m/PCCHCNLsVo0x
4seQ/DGgtN8ieQOv7O0VVXaiH9ETv4vw3a3j3wa2JOoyYbzxA6ArZQJDnk69OIqpy2YRkX5BK11L
VY2CCbahnKzw74HX9rg0bajaKnFRHcD6YItAp7Tlz8GYQaJ7H3wkd2Ls7TNcGGgh1jUjzr62yD64
dp6ITKa3mByzV2i5VlCh9yZVXR9b6EnIEblVBI+T4ailAIb1QHB1QnSkTYsqqvTKbiDM19anMVXj
sOP9gWAtQOhF22EeyUSmQVXKYIMiyJm7zav18CrDp6IAS/15hIE7wsY1ThSvTkuu5VgnQosQ4RZC
19mCJODtyqIGQM3xQFwNVl4SiYC6xrugKEhpoxh8lSf1mMoQBkSMgtmaDqXcF0Vw/8wfmHBVJZgk
I3NxEQQT1cVmHY+ofCcBcdSc6XmHddBGOdTBi95EUaVkBaNkrCociN126SVGdKaYeilosdfUSNes
YKccp5O+QHXzYam9BxwyvddOCgl+Dj1kuHR8qxmMaNPDX2ntC3CkkrF+rOipLrswCvOvrmUp6jSH
Z9fqKNQvfed/yGGQTudlcOB01PEfwB3AJX98/46neGEHTnZKyhQcLa13l2UZin8CIQ1t7KgSpjR7
t38+JzA7LuJL+JXDsHAvKxEQbaq68bPIAlbG3FgU0Jh3lPKMNn5kcACMkmlHXe0cjcUG4CHR7O87
/Fg8dQpB5ibPxxmcNR9ZLb1zlfMxZbS7KdB3TFK0ZC3XeCwPKo3zZXssuYOUxa4WITaN7lp5SGLs
NssJQsekrpoEsoYceMDr/oXewpYnvCXU+RjArbIC33CxHDpdYwNdoSP2oVi55OP+zrvMo9EhmnSn
4by3bR1rGrKQWWl8Vr8RZPNUdkWuFwb2YAwyIvLH4zhTzFCvTN/7qftDCIfpJwwS0+7QMM0QlBQo
FUDQ/0NGHUHNylo0pJkllTR6q35gsKtdd1vov6mp16XOTwq5GXPPTjubI3cqCXup0N3C680jbrxv
U2yC9AJo0P/wqX7QMYa2sU5ypKCF7J7HwxZ+6C9MEVnisOW7DgHU4u5/zNbTVz4kCr6ULxcrzxrc
J1gNfwP8rdPMMiA/6rJpuLvKn5e2v3LgwQYQg8Og2IFjQ1i/cXeBjNtQljW+YQX9NnGz+D32trbC
bbqO0BhCNZgouq2Ly17d8FKCAhgu4OpiK/ZEb8JVtS2wvFNOFpAPmLySCkhJyeCHRuECOwZTZ3Yx
CfYrME6WMNg/ubTiJYPvm7mw1Zx8ztfBryCWDU47iCGddpqHe5Ap5CBVzi+Co0SsoD1wQnFXWhlt
U4F+YBZ6rgNYbfEkQltNKfbkKt+9dNRgNbigk3s/5pDCvGuPy28jz4kDhRmCjtWddlXK3rVHFSyS
lGAPRtJAX5PJCB1Mm3piYp0JhH8+si4fLxB+0o1bRelUezYXzRyDN8ltc0GHDELFCjkr+vN6x/YJ
FT2ESMYgKXetZy8ucs6JoziIXVHeTtc3LOxWSfBmIvCHcy8Kgs6PfCO+movHwkPqGtjW8U2WIl/o
Qx9PFVjhy2ExVOZkqUTXRgHzmox7HQ0q1301tnELHDqMl9O9nDK1H2qUEvksbot3iWUC3tTLrSX7
koTlkpTpu9aMfvOOcGoHF7PXsjBEKxlTUsgG7Gc0bI82tOaHePRU085+YA2SlSSPiIeRpJk9d4PU
NJUCp4ISOMygS1XhyHsvoho/gLvBPXOS3lLIkdYJ+9/I5oDcqSFeecv3U6tOsVCPp9PLG5gXUJBZ
L8qry5/WC7cj35Hth6naCVctZNOYKtU93nf4wZZFyX06aXq5rP82POSPw8D9MunrFgWPyOIY+Wbe
4vJszIQIqZyGCdjlUKfTPNDuOp4eOXYmTQox6SXnHgx5Iv9zVQhZiB4Qj1iUN6nJL+0AEMWzgCxO
ElqM1Tu0+sMES0rRiOeqYosMHvIl50KEFG28W8+sHs9R8/4A/pLbGInMnWCFWnlOaguKvnvo6dvP
m0ZExut+LNgfegA9F38FTCmi5m/Obch8qSipLboRVGxXF8Aj4N8oQNm68h+omyhtUbQwq3yaU9lD
BGq2JTeVhk6VAeBsfQU4CnUFXaccpRvtcfBZFcvT1WV8UoGyTdhMb4pQx4q2j5gPbKnL8txB3Qmi
zCTX1PaJVGVQwDTqF4Q1GrL+lMvA+FDwkxhwuop7p8hqpeZfqXlFUfUDvovFZTFPHJRtm7HH9RQS
by4DMcdAflrn55DheVy3+JNpfP7rxkJBydzN0PKP3RlPCSNsKuAnELA1f0EhrhS712Om32m3S5mP
adK8J2+a5t85stE4t5i3UZkgMu3/bo9akWUgkn29DV0KR8ubxR2yjccjelVfgo+Q69j3jiPkayQL
7lqAVDs9DbsCz9qRDnm5ujGaUXNZ40dC96IPKbVUqTU+pa22GXy4OVZf6HmonLkrApEBxcXJoTZ4
j/BrUJA3L0ZXzNMXMYXorcAWqTGzb8X9B6VQRrRDOTaGhQ/4IZ+cvG86UJPjjq7NOr+yBWqo6BeJ
aFkO44kWyhTNnQYn4jsZ3C1gRrUUwQHrqCQwucf5yt3/S3IxH+sqlsZjK7ukfdkXzgm35bntmsh4
qGvcCrbbaA+QPULWh9dqOyFNywRyQRErzraYBFiWT68N0ZcFDYoks4mCL3Kg5sL7wUQI7RlFD9Ap
Auc9fdEDgGl6oAN0MY1Kv31MdkR44o1Y3l4iWOAf9xL5IAtPyGmL/8n8eI1h1wvv1gLMlwisDAxN
w36X08sW0P8/KItVtyEW9yjVhwuGdW2w75Myee6bAC0A38uElA/+CTBrfthvwgDA3ADsNaGuOHvD
IQBIj7s/QuI87DBqM4THs54+xtOC0pLa7HUrc6vI2y0DHw4EUCqnVUS3Kluf3kdMXQlc/c0DgQo1
7TZ2lIjmU4tbRdMRNeebJaDOv4gR5w6gprHL6cxMyUd7vrJ3MZ8QLm9gLBC+BM51cjEALXF9bVaA
nPy/esMGiMw0/DPxl3rXLz9wt4v1cW5kSYQymEr3NpNAWWrOCTHfQjljIPbfcXuuiTrMy+tnQhD5
UcNCYPg7CrJ/Ok1lt/gstT8Wr4dPU9x7SfzoeWSa2g56RBNth2/JGKe8qtkwjg+fUfjEg9pBFVTb
BbE4qJsk/dc4wHLmZYObiSVN9IaRfcCGgY3qPTgj2FKCUhcDju5M/oABcQGSKGFNA6ERGxkViUpV
wsD0sGa/Ak7lFe3iZAT+QganesQTYVfSJ+upayAOkRpnVGck1Ebgu/6c4Uikvc6UJycriNAf9Mhn
dCBz4V6i2QQ0YVh7JYi+lfszkjWT+HRx5rJ16T1HFNNq0thJNhqPA24MYmeDELY8bqlg+uxm2lqi
k9V1/Jz1hFOIFXFidbAZ8FnoZ/QjFlmxcv8eZ4kPcYsF8EAUeFExhYwRQA4st9VP2UKM+rbZECE+
WcdqaHsLdjDJA/w1A+mJskECJSwZhvXwv2Qx2aBpMIASo1uTPOIArV0Wnc8iHYdfJYE9F+QxdLLN
ViVZq5ngIYOgBmMw62AGs/c4Wqy6+c2t3uGb8rczrkRSpSvIbAOrqejFwzDK3RGw0AVJqYNJbr8C
MsYO20gB1D6uqXs4DEe1OpxF5YJCvIH6Jc27AfuQClpSq30Id79hgBHFmfRUkpBwASXUPhcMnfHU
We+fIqrRVwrHVvy0rt4T3NMF/tQRFx3URH+FwagsG0b7/QUYPFOxsTo9vzIswS2N611l12OTc/l2
5RU2NCfNWjuXDSYB3aYn6uI3TDruU7pxKXs0yUi0fdsP8l04wUlE+tgkDlEzfCilBa6pK0St3wFZ
/jw/p77qdXR1nX2GL5P6c4CR0pV+vo8B9OzAxr0EXy0JZrgqgKsjepq7aKZ+Q9xaUFFLElo1x05X
RKzgYUv1JiFYd/AhRd0WuLbyFXRvi5vG3+geI4mYluIhx3LM/QSxSbfAfFgV5j1FaTdZ5rcJX47H
UHiJz83r895woX9Yf2Z8pEtBiUEX4jq5nIk/6ba+NZySIZH76gDTRGYlXeIudhzcJNMHecGdXuhz
yqmSfHaND6IeuP+HOVNjOb6UzRxScHIFsi3zzKACm2C/Zw2FiZO46mGSqXhnGQIrvbXiaK6l33II
iMar1PhVMnjdvWw5ZWYx28+9n7hHAQxXl2uuZ9eLMFwmSeJYwJ4Cl/Hto5W4puRXSf4bhd/Avjm8
QX2Q30Ta36YyNhK7ETYn19JjkYX7C2UQSwf6sLaS/pIaPicYJ7+8fn6/iKmWRuvFd2HsjFUMngfY
EvFz1QQGrsoXw/d+V+1y9TZ7PE1yhpwfcT3AdGYbVUtpd3RDypOH0YlDoGOWN19RqSAmn5iQerQ+
2/XA1uRl+lLuahmUJQp6z3BjfwooUzUuVQ/l9IF7hHb2Z74wJEwwGWAk3QpPYXKkN9N1e4PaZghw
9TE2u3v8Wndjvq6mWZGI07852/OtOIHU9wBm2T2L3U00SOamAv8Na+9483e92tUC2+rI+1vq250r
1ZD6JG2VQIroLOOICNOE+hjRcpmZMng7kkEKWNLB7FTcsfzRa4jp3YwoWFYfBICH4rlgtv7KpKjt
+y1xzrNyR/ZkhFdUDxclsvIWbK7rPcuPfYVnH2K3YoF+xsfvs3MHg+DI5mNjgUqqisM99fkoP2oy
+1ul7w6nObBBT2chggHcgx7dcCHvRB6AhBUoL7PCp5fK/GK7HxyAEsCDyb7EopbJXSU8xJgE9mpW
QodQqnKFqT89D8bhiC/xr6OJ5pcWcVqbdpSt0of3QHq628WRbUkAv74XECir7HUoORVE8RPMVFyo
Hx3nRoH22l/w4qpdP+oo+B7SEpfw7cQ2HrY0iQMzYP6OGcXackPVWhwgWZtXu3/SGNAoi40OMvFJ
Ij2rFWUO+Zo1Pp5NnKg6PXRH7JaJa7bZsFJWd+hJI7QGCXJk5WLvXzxzY+0MdYxGZWVGdnGZR5jI
ayRX0P14C1TJdzWeaMKS23sG0f/Cf+5gN732nnaOYgUx6Ukl8asgM21XMPTckjHkMN3W7cz48ntn
+iDwd/P/9LYSqTvQMPEFqgqKMd0Lo+UBFmGgYJB3n6FPFKbFLavT7qY5zhgvclWelWBsNwN4Zlc1
PWFBl/5s2BD0IfprfF8gz/X6+GrPnXmoSUSPBRfhOZj9TWB3PDBuvPEPXBOYjOV1xP8tzP+RW2Cn
q21801k88gNJVi5E/kW/8HGcpKlB+1My6Ny5VPPpXhXSr4Gbh7Kl0X7PDeIo3nY2Rp3Z89W9PsSE
dm33NkqDqzK6JQBxgbcSqyV2b+NTKCL1q1Z3Mlqb+InsrrfgU72nnDFRlQCqHvuCkJHCU+n+2Rwu
/g4iMkJ2C5hpvV8G0RxNgiybt7wqMDCpsoO9zfJwHjBCDbqJWIl+uawPiAExdrJ61TN9JcmKf0ET
j5AplsYe1VtSQxly3E1gbS+RiEwIdHmX1BjQVcfOEtOHAFq8T+GNqlbfVLy5uXPAHC0Z7s3ztM3R
IVXRZj8DalWoxdxFiah5PyZbTVMu+Zt/gEi7ARYiLG9f06Z9hv3LZZ+J6XnWx84fWdk6nv4vrpeg
hQ0wFEjB1boqCg3sr0G/EREtatLXAeT1Dap4QxYHzFj0Wcz/Ls/CNlJqnJaVNpG0717heQd0gdR5
ULSa5HtGL/C/gP6ExRYycXbuR1TDI8hDRdb2oT9cn++//kwi1y5ehuIe9mXUShyMTBz8XVyQqeVi
OPet67HrG3dvoRDY2KNA94ar7UTdeKY6ZilIpjzaqDSUN6LVKdA4vBL5TkUX7cmxxfu42+bec9X2
zQcB6IJ63Yb1F4roo9bK6g37vKBQboicB4FlTVQRacNCOpWSn2t4JnoqHsK4v9yym4g4EjK1b9aO
6vWAY57TnVHOxC7N00LeWxop4WeWQkbhwx5wKbMPHwNOpC/5F20FBoyjiPB5lLNwt2nbVSTgQU0b
TbHUwJABBmNN06SrMJGgz7WvbsFDzJc9Mf6zhgOwypz6ix63acMVlxylnlBqtmWwZkOtwDNBjX+4
XS88FmuUOzweejwWtivorVv6dbwvvRT7SWyVGZQMMtXybvODPWccHEqWtBh9dwtVqgM2XgbNIn9E
1aFG7/rqHsbzl7tUH2d6PJNqMjb7X/MnGzr+/x19edqcr55EO2MY0QU+dlhBkQ+sjDo6XpWb+/1l
YACliDoyAdsxh8+MZCbE94NVaSPHJvue3B5dsOEn6ixiIol9V5kewzuVxrOMrSALSxdW0YMM++wP
cOMuYKpITNJe5i3Q2zEZqcb83qXWggA/jtR9iTq7/o6hGY4A090Uf/wJiNjitM8nxQVVaIMyeaCh
ZEcubxGzZwesQ8EOz6ixURgMP45bewTbmEIY/zbFS3IWHk/w8e553fLupHumBPqPvWIl8WSutHqK
/ep0ZCziJptaNmWLkf1w6MpXwJMRivCQ33UPg++prr6t1/fOzGQMHpapm/e14ITyQq8/ccBBmW0x
wzFZdNbQPxTlaxvDo2SKQHfSpT+242CZcmMya+2MwiVPci0dCMXOQTSujUk5RDyWX+wggNXLJqxs
xm3lbw0ox97eTFmwm3He9+XijT2iy7adtI6Fjou78ACM4XD3CI2OEihDMyGKTxOuvnRfMcPJSgW7
frMf+VKin5Mqr1aXQoxLFMxz+V34uZ9T2Bhzzgxh/PpryfjEN6RCFaRiUqxg7GVyPH3Ha1+sxT0k
vbOurJ4q1dgiftlmZKU+Pkj/3/BSWJ5ouQkfFaCxnL5n228Hmfx9L9Wxa8Ejn9CerOntJDCYsqVF
RM8SSkFmF0sRgdhgcimBcY+yVfvdCFrU65U/RBgFljc6xU1xaPZSvD2kJpUuO+dxCWvyZG1eVfOw
gBWlUR3KrHkpx3hLimySbmFKlWj7bLYQCDGehMNdXW5Bw9bCrxclAI3OEsK6O+yZzlINJcA3zd5Y
5eve+ihCayMlRBao0ntiQA0R2FElABrBFM/Sls7UfVBj1TxDBweveieSEBHhRH9aWAFf0PMrDHH1
ucu1VHvj8LFIz4Qjg61XZyJ+hunW8vHgSLPWKs+cATzR9snf1kqRKQQM8Kv4Kl1V5dJdGehi5IbA
w3v+kPJbX9q8i2fkZAwkASo5aBmB4Q3rdUqV802gIUghIhhBzTOHulH/Ug/y9kIHTWky9xT/vjO7
yYC0dTKXGg8iwTcjLR84Lbww1keWYwQICTjfuYZbUCYtzLYm/7YW3emLk7Cq1LypfJFKI3A5Zvxe
PQQYHPhVStgt0mP++oaGsPQXCXYrcEMzGs+wyxIgRYkE6PXEnVdnI/YyMJHGH/4OqjoVqdjhGJRX
G6uL1Wv7PdUJj4jp7QC7+ijy4tzKfI+TJcl9BHnhXml4XM7RDlQfCIp9Y8SrGR2035JI8Oj1vudE
vPVEN/cwpKmmHIdXmPfPBW1dJdyEfaSrIlDnc/cL3wTL9eKqpbZtZXv/AqqTu8nzx4dLiI6Iufor
LBPzmZTW3i8aMpAPielfi9VEEQzDxbGcV6uFYAya44PnY+Juzx0T6kWYUnTPZv+LQmDW9EdfEjBC
LdZdYxjmjCLsCGMK3WjRXdVCeP/qNXtTNrUvNmEQF/8UYfOKZ+SbGn4RjtNCdUgkFWOWbfqPQCWe
4wZIANT1Gy7y0Q9xUeuSqrxo4gC3CEJkwgBy3T7Sv3b5TD3JYm2VYwSkORTATRsaYJtKJnNVMXJp
wO/yr8QGK5Fd9YiuXy3tE+UwXcrQByJCDCw8wTUah+PkzS6cBUuLqsamf9lJDS/gNWn5BwYsmsQ+
Akt2D2RtpNbjeUezhRsH6HRQDfWpnhTVLXlXmkHD35ioXz/JCEw65gP5RSe+wdLSU9orx3Nm08aY
bn6KlHn/VvdZgPTGDE5Z0ZqQzJU15DZhQ+eky/WH7bS4WpCwknQF64TGmzo8wdikw9+V2gFkW25G
E2mF3XEEjFxhLtVaZUammlrwtPRxAdxVPTG5vSgkZYy3Jl5Y4/yjsOZSvHfLQsiGl3N6GznckhWs
iG2Jm655hCfMKq8R1T9LXcpsfgFPjCAqQp6YK9af3vCzCvJZh+67bMORuCPQ7Qkf5/YzBcRCBK9B
8JH6QG/SBoqF25gHzNYJhjRKl+dQzUssStPc0OP1/1feZ8Sn47N9bx31Q/mXBI0+y6wmSNUmpgI/
EhEFutJpwOGIQHAIk5QVzCOKRvfvJCn1HFIseuIUNZ6LUVzDZfzgprOEef3ApaJ2tqjS9ewfXxqn
BDM7P5+J4SVHAfbwoIwx+9gx+XAjor7bXhKbNq2Jovb9VNkMMKX/RgHzeMVTlldWUfCR7YaHNKS3
8somhQmV4p1R2zCvW+hETl3LvT2Q/+kp3LqWa1auJkCchDcZhHWF62z7n9lVTKtkQHQGggR1Mn/s
UIYV66VSdzYoSa1e7Ffg4/79hBiRQIWcCxNgJFKjXV2HN71I13UfG0jQEWJ71Zt7DWHWKoQRYopG
/3o4kZ5nx8GqX4JhgCeXxhuthaHHr9neRxYOrLGTcvWxCMuXHTrw81+miWVQGNtbK/4xet1W8u4v
ENvy9alJ/V6tj1IvP9TgUyjGxs1ZoI7ELba9nf0rChtQRfz0vg9uO038v3KF4JI5Cg6cfLsMVlDb
uTIu/g6rll0zkn8oCiQFBSkvKfYLw35jbwQcUWj21RNrt2r/IyX3roRg9L2De+o4kiFXJYUI7fhL
PjGA+KTVIbxz+84e9pQeIyDpuzTJTJLozYMbibXxAE11e9eKWMtZSor2C7W7D5ASac4sFDSBcmn0
sqKU3l5wKbRFIk7w5PmFBZDT4bxys3UalEeFepVAq9heWS6IflvP2iGskryZrCwDmWYGuxWeDljm
rYrWiVboWLVVmO0g1XCQaJ/1uLEyRIiO01ISzUTeqs/Z/fBS0/BS1e5ApnkDBJt4e2HxMXvyJq7V
HwvK5Hhh+3/xzrbueLPDG16uPvz+b7LM7JeJm7qqBR9ASJ+46yXeNhFrRJbeZ8v0KHcZERBhNeJy
auzJDlME9Q/HbM0lp4meRp2Ena1tQofFKaYpoIkHHp0YSVvMTW/jLKXBKjxXC/rox7GJJvAm7eIX
pCqwUFEniYWE5fbKh0GGszd3EQXr/ghQo+hKQ7btnVbdYCf1nJrlysLvIY1r1eJtljS9aNEQburj
rX8eh9OKCZ2j/xc2ZPvLQz199Kk3fg/lGVe2H3YolVedp2HUU+M/HAdDysA1/I6MkremtiXuiFtH
v82CByyvo+dwwEIj6VPxZeEfz4AcHbIjweBwzHzOffA4zqPn+9tOyX6qvrOUjNAt422fbUEvWd59
4Tdb3VJxoGnGpElkLpD1tOCV7akDykrrxgt+aW0d8TbyZvvckPivboZthmpHlNGUto1sPb0ie0iO
3lZ+wHYHeqdcjpNXlsk5VdrObH0S7BQjwjuM6ajuXXzk3bdubZK5kODHqNnzIb4MuXiCEIRSvbwh
7PcxFnuPO0gTZALx0YXFW0EQT0OSiS8GJL+Tnc414B47/mHJNL4vPAPvxLjliOCaeABOi06SvMwb
pwtg5gCF1pvZbj/UNH2+Py2bIhOWNtghjJoOd2Dv3BOgeSaQU9KOnMLFgVdEuie1v5RnSgeGCTGC
yJ0Rln/EXYVzvSWXo4mllD7QTu7zoJ3ptqBQ7S6HrRVi0ar2QOW3fGzDPVMLDGMKli4XYBihL6yv
RXBgq3KjIWJljGHo4okLMdOsJnh1zqCVmfpn0vUxnjqVJS7UW0UEQNetU5ocVSyeHSwRLENrgjAP
wBLpAQRCf0kNAEGr7cXjvezFg9sHa9H5t/Dog4gYM/EOdGvvAt2mcBWvDX0+zQJCDC9E4aoOyVs9
mEC/xhaqo4raDdyry3IGrqcliZCGk3sxH1kv51Bhc6bhKj6r5sDtAPqqfgfRcd2/S/GExn47Nvp3
44AO1eUj+Y8daArICU1SqMRR/lBWOtVIalW3vzgzEFWigPoBALLE8ypt1whsCMVBpLRsP417HO5s
oeQt9+HM3gRwfose2iNjvoRTA0z7iDWzoCRyn4TdnBzKq5W2CgSUCgEDhXbXQH9gJMlo++CQZaGa
yuMGmqKg92ox0k3kzXrigDG/hve8COIq7J74UP5Iejc2yDkSNt8YjYrvEt3jxZZ6YnTlx9ZAeQ5+
dKBZMwucU2Yd8MqoMbcxq35y2SIEmay1CImhKOiI/HPKf1C/HAWkmqV55vf1SEXEccxv5J6uwxcE
uBMS5eahM6yu2X1kRhp+l5+r4jG96Mi2cWZqq2X+12s+Q8cLdWw6MkrLOCt2SwTCTrVBj5T5v+RO
vHPUZUhXuRdkcG/Rg83bgm9nBVrw5p4W23DT63MXWgS1RboKNJaa3iiBQzjhshgpgZlDVY7xmC50
CZR/2s/PbSAIhAoncuhUQ4kJx2mlVLIkMYWhtnQbXHBtr8MUS5REsHcbPxDiWIUwZROs+6SW1oCt
9fZnF9lJLBgG0yllbPHVm2kwwRkrJFmNMMFsrWSN6S3+PktZ4eNYQbE4lW1L9qMZV0fl7E44tTlc
2uRpKvpj4qc2JTML1G9qZaoD2NWo9fw9mEo3918/tEZPgj2QeuyEpINIsnF/y9eR3YEPttjytjWG
8VnhUlAmPZocjwXsD+aGsXm7Du19VZn8BYwNGuAtWf/SLvGaWcuthEu1hpbS5B02KpLUOPPlO3tJ
cnY2ChhyWIjp9qlzHxO0FQJ3n/1CjtUhmmz1JXPeqg2DyhlWDL+st0+5juAECmFae6Ck+eUyGEdY
9JucB0Ka9yJ65xnM7FeBCiMhUqraj+zRmKa8yywyrK4TftPiT8YlXlEryrpD81nl8SeW8tnSnocZ
CT7sg1osHtAdHH432zSwbBAwUaPt3SoPkMVGOJD3WPH6IGGDJ8UWKk0ZvtG3r4nmowfYp7z1ntsU
bYKOVA2jTUei94QDqdNgY9CqGsCF0X5YvzCHM65zzNUoStl3L0f3cyW78/3BEtDfSI2u/hbWdHho
TpXMlso3zSTUX/wuBLZbq2ur+Rkst4ughefxky2uHzkiRwbL6EoqUbh/koEW4wTiXejmsIjdFdA3
i3B5TO0ksL99FYf8GvP0X/O3sNZiM8mzG+RFhILC9wQKPKNOb8Uc5dqFKBMoEhWEy0LwSCfLeOjL
LN0ni/AXE5AsU4PLQkqaGUNUV0LBs3AarLlekMLUd4mFgvCTso7kVaJV+Dsz7tykdwd3hCPzxnuD
vBI53swCNRjS/HlPwSCdDi7a/xWIIJWzSWkdgHveNWVR11CQ/ABqFK3GAJTfzU8RBX6AohaDc6a0
h55o/KakZQWjJf3Ni2bYFA1sQHxfeF9xBbUhMmWwOWNiyc75+TpOqh7Dyp9iPtUjizvvloEEe6d4
KGM5ZsfppBquQX53Yl7TiXQu1UOIpZv1OLtzbjqXncUC9qYbu8PlcF2MI6yKs57ewUSgHrbOqUvB
+bM4O1z4H0y3ZmMwYFVIt0lOj83U0otjsle5FrUbaMQD5erm4aBzg6BhwMHrUMmqMGGCg0uPnq0r
sbbtHaAaAEbKj7GOScAQcQt7NLa/NQW3I5K403z0Fse2NvHctFtjxTI+4G4x3U0UBtwTv1ojTnYO
ZNTaAmBPnOHW0qCE7FkrNW/btJyofPpYpY2JSPad/9MZeRT8hqIwyMoM40rtv8bf9OSVP5/vcxzz
JVMlVQi+JajqwR+JuFLtMB/qnVz4SH4xAme5jR7tBzlocPEEvGmBfnvXP7KsQzjeaNhhEJrRHnHx
oVH+6ruvmN0+X7mCgK2lJQneaXcAFVSeh3jnYwkuX+ARcLtTfHUkARKwuIOVqfp373T9zwNeAKdm
ZyovIqp9UTyfNPiA0EJ6VYk/mKOFbMDHqo3ZhPgSH8NiKYs7yAPtcyKOfD7MkLmf3wLbpVQcS9Bu
YPt1nIi+318tH/bRl88Q4WK9fJEAsIihBnytculeXrf9PlZinxsaw7NWbfDaiqdsQUcOUMurojfV
T2FCqmT4ph+Lq8wrqjE1BPmSNvG0y9CpkeGWjcI+ttFf+sw5WusgBHs8gPN//UJ5+4P+bFxS0LO0
x8mggIJnWKKxP1qiIJWeZQZ6+68IZecZ/DHzpsba+grVHtWSP8/fNKTXR6D0++Q+StwdhZVw10JB
gRqnG/NtZO14fi5ctIrqBbsf8KYFpbwEfKhCiJTY30zH/sGXWFxNBTmznZcDD0lgd4vDqE9rMoCZ
vV5eA2GOB+qkMOyx9IQ6P33yLtSHT0yjMojNfr0EKY31NWhZwskEx7eP0dhm5KW2fszj/XJ8LoqP
ezFLUH6rLt7lBzAErgLOzTVZvOQkJVcvnmOQlYSH82PG1/5hvM9EYODi5CjMuamW0vdt+03/P70v
T8DfmVCBtZpzNvg6WKyGFE29BFjO9t6SYbHLxhQGpspZk8c1Xrs7k/Xv6pXNZ4hwlwmaSydYYYC/
nvA5vgJ5xOM/T9q3TWqKci6o4iJ02DP5JYLaOFUpW5vqZQkbULTBvskuV9K5ntcuprvzbNyXvd+n
pUWM2wBQm+mbMjh99ebPj/jSE8Ke1s57rKS686uPa06nVI3r+ZNBVoHM1jDa98/BTDdsq6KZnpZV
R9yoolgJv0f0eHUJzaYNzDlJ8j0z+udar7UFqbT2JaxEIW4V9HB1sfqMuaP5L4kTYvsLFCtduLkX
sfQocTC2jnlUF4b90kD07zKj1H8HZ4U4k3GQWWaXDsTTZ5dI7kC/r6q5/3pjqcjXS6ogzs4iO6re
3eyceRCUGPoFC5QtGaiaaGKWulkD5Ksx4UDHjKZ52jJ9vQi8KXo4ei9mWGGofZPpfGjohInOBge4
LHAHik/smzTWozgSRZ8gFOP8XN8hw+LzBUKpQIbCHNo/k0nctaHBdaoF+kYpvsp2Fn2eNoEfSWtb
Bn684jnSbCpHkxumyKMc8kc409JuXyhITyoVEEeqjFp9H9ZdjstHkiqo3AvTvBXgms2SVuO55oJ+
qFaceeFSiXdeCJmHCGIctaTFlRLYZfGY2tTaQtOjq/c9OSxoGRN5UjR+eRNP2F7pcUbWaAI6sAvh
kW80Z25I8zCr50iJ7V8la3T9UPtpRuQopgmKZSc09d/wpynvTbo0DoDg3/mKA1GtlB7xP/OrkWwR
qA8g5fSbTNRD51E53qEVtRUtS8rZGWmNKHkBnlk1hA/sbyok6GbWnN+aoTvyknPPFeIQsV9a25VO
w+n2Fik+G6iqNUA+gGQRPR1Uv1jJGydFHPWL7OlXEtOLUyuIXccqNqZRmdSzfbeWcaQeCSh3Dbp8
EMVyFzaJJEDCd0OiacFZkdL2H0+Ubaas0GAUvCry4mf1rJv86ooqpci1SF6T4MpdB1PgX/F/dqqz
Rg452Htqp5RwXP5H5XBerns6UeQv/nQgcjwhmcZ3sZy6xDUKMeGy82Ft2i172QJytkhTYmFCK+fc
7r04dD8NhfRlgBPSHIFsTUVDRCgkp+mF+WH/CHdSmXaWdREoOLuUVNKvgkddlZifVlr0NiUkgMN1
3BsQTR67kxqCy4Isab9uVKr4uigCcfnrHqobORKHWJw0Ssk4VtKVpQZj8kL2GPXgnwTo1jJLYMU9
3xXCyq2R8NFSdPT1Rlve2s3tge9X6sHdh44n8ZhEe9xXOfUWgU+RSCjSQj70vHDP1Vt9W+MxpeKe
akRQjp/87NhlkGgmzFHCkBR8COFinZVRP1Kr1G9KJ/t/+GjRob3gXE4bPYNeHoTLBZbJ+0EvE/Hb
ueIiqZCligsFPNvhxfZVxhSddj39Y9trbdTgOsqfooaNO7iXm3tvxAYJxXY6IdqSrvSeBVvmxujc
Z9SyD8XKR67LgZ3pyrIeM0nuawztcqwTlj8nQdWxwqyg1naSN6Kd5icFyx6iPhOzaygDzmOdAhWF
Fo+6nM73Y0lUlrcN546Q0ZapApreu4VlQZ+PJWwsl5kxQSMurU67IKj89WZejDsGXW7Wx1Kgty1m
8ZvvIVeZX8pJHGe/Kg17VhoM4C5VHkg+2dsfbz3F+0orlg930wCgcdTn8DxmxV3gXNnTp4RQBQC0
QGxF7PRrVcYL4LI6H41DjFWNceCsnQwx1lrSactGG5wrjknaRGA2bxHO83VxgHwb/x5G2Pf/Ql5Z
QgZURmRIq55ojbdy7fxeoek00Vx64JU5Y4ywgAoSeQ1LUH8uG72N+bKrYO+20KkcJ6aIpqlentvj
8DcSkUgrIUwHOjFVCa3hEXHwohDcfCGiDl4XhfQ+sMQIlnGjWO2gPYIghBaEAFQLmsjnY9GwrZZn
YKxvvh4X7GGTqe3T9dnUyuBrxhvTcrw+pbtQDFavZTRUnwJ2yFeRHH65EZRjsRNGSstFydEYOgEt
EslYiKZ7/N3QuWaRzfKic/oARogsG3CnZiTTKxRv2H7ZYSC1UO795h3bbYQKF6cb2xbtHLTS88AK
mH/SFmU0Be8YlckqGnnjno6b+VB5Ud71/yCXKdPUrq5t3YOT045bWMf/2T5SIE6zkIAV0HXoHmRr
NGkFGMzPXpBenek8C37q1Hw0VFz/ZJjoOYGrBYsi2D5DVJ4OxK6WMs5BcnsJL4pPNNqYY8mokPCz
G1Euu0AQic+p+K4GoNdpS6aLUO0sffhakgtGJDULAFafs4wo82bDdUWy9qyjDBxc637L4x5OSYIT
+p94Uz2uST0NXhi5S5UWIo1qF+L/enE49WwAOantbWXUgDsjPzlo+8N+oRRD9Whki4mzJEMkcUM4
Sya7Zn2pel+N6x3lTdzxPYRu4CiuIbbfO1W81R3yfMpVv690xugTWpBes8flfXshw7VAnSjVjG6w
/2NY2W4QOExWJrknmPmF9RiRRsuv3pxQuievWGieu3iLfoR+J1AUKYX1u2SsfuufMWh+ML3J2IT7
SorCgPbiLPrPEnZDsxJQMt0fL8XMnu+nQQzpWzSk4ImwtuZeLHGY3zyFKU3A17LrDP3hS9Q63eEi
arviw3cnPamZ74BrR4gk0f5UkoREEMuFqeCuAMdRci/7+R8ISxAUS+LhOwcUyB899skv53E7pLLV
zxz1JzkmsImozoDhHeVhtZ3rReXMDZIbI+1aVK8v6/+xG4H7vfIQJ6Tgr6kg3A7vccqM/j7X1Y57
nTUnyB0QtgBgszfHQZZQAtErOTJkt1Dibv2tVACoFpEUD/o37MKoyLq2Z2sxkaPm8c2Q0iDelJoQ
EONGnJoKR9CuJDgjM5bzWh8o1Ew9owEKoP2dq2jCg0JGypyQRTDR4tHkMu+7+sg9t7txV8tib+k5
Volp7KjYizPaxQjNrmEgOhcji668SQQ+WLslAcUgpum4Xxr1+QetMPbhS1l/ILx/iXrzrBYRVLPh
b1Y60ZqPUmzt8kxGnbTTZFdRiSEdQlYszFM0YC1Yy8njllgeiukmAN7l6rxqt4QEPvGenZ8nBLic
sBI3tSRCrP6gGX/J8DmJu8nh/bgntL/xH9a58iDrzyZ0/NGMATSx9uA3HD4W3BGoDXlN5Q/EAvFg
kBrr1Z2b5YzWaB33f+oSwpZBaKp2mvzx5ArlIDG0xQyz8kqhahhR49Pyn7EHz8W9gDPa1mlXcBi3
C6LrzF1ZXSN7b9eR3fbfVNhKbYfCFxlqqiZaWNyMzzi74A+X+jch9VJcLffucbzJRW9SVga02TI5
s1duCP1MbeRtSBBZKlXHVqAsUjMs/D09BTNeRN8ihE4QxIM1JV06H97WewSZah9uBpHZ0Bzd4mM+
qibi83hL87dvjXjZayF+FCUW5txV5PTKVIH8YPDe27nGdDVUeST04N1x9lVHBkIoJXVZzm0UQbWp
wCNwHsEaZUJqaU0L5jXGAXEPaFHhixy5H4vhm3WFHg004Qvy8q3+roavsBeRobWC5zZlXE0piVVu
4SZFufBjmwf3423EdexSEBoh2/7Phu2zzn6zVjYlVJBKJzGea1KoX4/gBtq3pC+bUfGFUH4wk3KE
XjQkIToXF1oJwDkX9jvmNY7lNvmTAotgo1VfZwc3+JGY078F7urM4z62ILaO4CoogddWfBs46Azg
rTm9qRbdrzyN7BxROVRVObUQ4oYBaCsn74YFUO5jFbDX6zH4bZN7/UAMcgJ08sbAYCBwHzwUEKWm
GwnrsnlPqKKrorIVHI0k5ll6YbFYsPlsqLRuaexA4vQqPdD+bJN2Ld3aFi+aMnHKZwsnXGuOqO9C
JpTPMiwE0SNiZPK3alhpq/HhH+7QWuAOtUO6x5BkeewnauSmcOx3eVUnxmqdCHSa7WxIo3hDV5BT
sc9EWB/Ugfnyl2I78HAeocMCjTACZafHOEduKYZUj6ec3cV90bst+qvcuxOMR6kQ+6kzEDK20Vzn
IGthh6jRjhrAICKMUl9fi49ukvxsPCpSOwkZJgwSfbKjAOjpHhLaIaald3d6IkP+KS7tvvM/vmRZ
cvGEWiBH5O37ohlgxKknXW7y4pmrKBEUPCChKl7+qGqpPf4RjyxCu/+eJpAGB2+pp1rI/mmAqzks
gTlvoGYKD1L7gd0zYbiREaNnNHIxKyWXdVGScqD1CvSlUC9/3SLX0wSHSqXYTL7dE0pbk7OGEUJf
cdE/ziLIQaF04KQrxDl00kd73Na9vl40zCR7FoG23Ni/9WMNbWqlEFABgckoau6iFwQWFiNGNa80
trmqh6R/gVxP2+tVyTxCpGjldDDx6H2M0UqD9/AshUIJlwvr9E6VOvBSpW+RvCuhAQW8rYiXsgwx
ADUbW2yjgP5pmyvOmHcAtyYU4s3j0KvnMkisE7BkLBaGxmjPFzXjGJpwI3aJHKtH+22zb4IHPwuB
FyVV5mL6yEWOE8rb2FBlA8Eqtr1Px00N9JIcXaPXLOx3sziENco4Jq/0Ps0Kb2h8H6qHePHrdADF
/u8zRlLEMt/wllXeIx+NY4x526e6BTWOeE09EP6h44ge4cqzMbN5cojTWXyPx+E5yecGpMZAN9eU
j80imIoWO7t3xu3noME0D8J8QOeqtFK4XwEbO+O1aucGIf1zBu+3QZp4UTfv97njFUy0vFxYQGT/
/CXptVgqqCBWXsYeSrblXqZR1ixWbWsNehiYTVAjwdWv/kXHGHSd6hjrjBIYHWOYgxxd/69dKlYY
kfoCmsilb4ZB4bjksZn9eA7UT9Lg9cfuo9kx2tfBfTKiqHaCc4RdL5GQYPaISkVTDQicaVKYjKf5
fmxSTLN8WJPaCvTPfU/Q6XVWJeCuFocHc3r/yvFPsycM9vICX4VAJ+fl70xkxq50EzjR/0s6QJqK
nSJrWglwXKJaUrPkqux0tlf2Lwid81T/WCcDonJorEoqjKHeIjkawXs5cpd712XOiVMW/TSXhqGL
BoyofVvNHdqZwpHxLsd20A7Z6HukSRF0GZVRdqc3NLoJUajypTEIiHplZogC5Gu/pg4LYNJtx7Px
lfHV+nAfhYKCLFl7nTyiBJp79rZ4/5B2rfWs4I1s//hXz5HlmlBAf7tT/Pwv3/sRWo3cZzAVAS/2
MeOAZRxUXHL8caFAJbyfnqHgCO0OPFY4rzoF2DCwVxp6++o2C01OIuBShR+uYLz3VWVh7Ydlnr8A
TpHlR5q6Xa91NEzn0nBQqX7T+1OGBnT40RnxtwOuku2jDzj59Gph/RQo2DPwpaDGshgPf5YYJ9YU
0pdgbNIpBkB8UW5c+hTsNAPyyac5ejKJ/b2/kIiqHC7C589wmEqtydNEFGVpmBPQYljR08S5Rg45
fI3RiTC4RneXsp61LS+YKh3elKF7RN4/+6j5duz4rysFRFZsXCTJnndDEkmatMZbjyJeOrOtSIez
vxZB4cQwAn9Ln99RRY0TmSq5dvLzEg+nP6nleUVJKzo+4U94ppK1L2f4ZZ3n4lGmtZBlOYKmdfC4
I1f87erxNv3Mj5vxKQ32NYGC+c+FNJ4bz34pK+qWq5lPX4MpN0HmbycymHiBQgxMQFx1GmYUg4da
JGlxSy0Ai8I1er58QHvEb7qUwsJEdb335DhMJ69JHF79esrTuKFNHldAipm4axo2TH6MSM9D4oTa
OPY7Y4Ww8Kksq58NHlNg9PbHhJexRjNuzqHH+oYEswMZEF4JnwjspXLhqX/3tOwaJ4pN9ErZfAlO
kRO1EZk8/1BcOwxm9NG/VNxNKWERFMEAew2la20QlrbJujILm9dcXfdefky7kY0Xz6Y8uIm9V/iK
OEI90xJEgzr5gBB/X4NVkIiccLPlaHnjNa0hKKKOERZdsc8igL+uAdQm8tFR5BCjGoZJvuJHTNWm
Q4bVOxG21TuTBJqFnQ+M8+l5T92lBilunHvQa1aka2s/ln2pcTvDW9B3/rqucUIjvWUVsE/Fs40e
3329zywFP4onjjOtmpkznPl1F5fmtn06qqjXXlsphl5iFKVYt+7sLO6etwdnaY7h9CT2NlTg+x29
dcZi81afv3Qa/GFQZVG0VixSYqRARZnSDIhMIJ0bsH3cCMAmNt3y6WWJ0OBwbqWKpHwoHvBwVhIF
dJ+6WQz4kb1rilq4rK9ooXjQleoSvqTXwNn/9j28PVDWoA5Hb4/7CiNXTmaahk0pzGtx4tlP3Ap4
ksCGsjq4KhjSapehuNMbqd2MX1nRSgWuu0kvsZKufQ9ARZuqMoR6zbZp0tNB8meiqhRjjU4Mkw+C
F9MOHn9kShq+H+1Ah7VAdKpGQsioXFbZCpfQrGpjxbkl+1++fcHbmkRa5u3l3ajyjvFrNxG42I02
miSttvdRDtEg83lCKm73Tr/GZAD//saHnAuqR8FH0I0VbSW9msKg2syykcoKlTzAdSKR5Qu1biFS
bO9HqZZQC18BPLiIRxinOL5FgGcV73EzGqYSvYTG0ZA+a0GJi925FbMP5kFV3h5v0hkRQg1sEqSa
Bxx1yGP+5R07oTbY1y73+bj6tbmIEzC7m2nkGooNthxxQOVQ5lBLYoaVqf1/x6acxwCcySmc35vl
yOXRdjSZyJYkd528ZdQqNIGJ0SOyVaQNzAytEq1K2e6VH/aDa8xsm2x0DKBGkMB1+lOdQLe557Yt
UQeeXQIaaAWDILDVvv/0p+0NKQ5w7JC2W/vwvWhHTcNIoefQAqu4RB7ufLgoCrNfV9e3greYSSs7
tqTXLpG1Qc4D0cPCc2lfwcbcv8qN3508YIun/27gdIletOWWeATyqGWsljbkcCBZVvlbfUofQulj
OLQtGVtMvmlbpJ8zMB56w+RE3aWOep/l1/dindno5mhb2u7jogARD1xr2VOpjL1pd5ClAiC75kOI
qNX8H4pFNqOD+JJCMHnEBoJJ4rYUEOcjWVoy2GHfjg1fzFekeVXailBHwfkVW0Ou4fP/vEz7OLzH
xzFxWIZQFzTpAI39eMb6KeI99Ss6SWPTiFzCwzNMbvuZAgTRZvYvZDaphy2MeOVHdpxSpkAAcJWI
6ytfCeqeq17sG8KyGKdKBrSxQh3ntH1jf9kvFMlWUEkV96eWGZvkEdu+cb81qvqG6JtefBU9/kQN
gscKH1PpaHmo2E+4FofAYmw2okvLKNQwQZmK6EjzTR7o65TJWkdGVIer1mkNu11pCCWZwucf7cg2
lHOjA10D9l20XZoWkRDick7r7iAO1WHdSAm6BjWIF+6SNPiB6AcDaWN0ApM/w/tFH+D0xPJXn6Xa
/MmW1nRFyEK53F/ldqUUYNVAYCN7iaInpUXIpDvmub10GO50Sx8EBCwrQltKjZ99nmd5YL6kuxk/
05ApEAGFhI+ZnlFjgEdhPsW/Qg0jKL2liOfODIOtCcKGw1BfoLkVhrzJxzlMEIW1Coo7vloqlfBd
llwdKy3rFfkayymJZoHk479B0ZOj6vvIAPxGSazQkQba+6YB1OJge9QKIPpFyWYkSCK/c3jMs6/c
pQai67LYAr4Azcpgl+mTfaD/qo36m+4ZOFtky6EYpeX+OQCcNPpPKpAc8egh/1/FItoZ8h1MO0am
C+MGV23+mGaL2lbbNm/NZkk9D0Dz+/WFx6aMxx5LF9Nji+W20x2FwwQHX+TKksWcxEKW/Bsh0p0s
mcg0HKnr4LzWPSh/Fq1HbtyW9xb1oSQoh98AIwP7X6G4BJ20ToGY2feqWRDGPQs8Cm9xKJMTu/45
n0gutCcMXPXSXzYPNaOA7p+ICuxPR7b6sybzTR2ePGHFI1yUknbqmBsF+Y9iDYfEZkZrrGGfpAZH
gkyV7R/X5GobxeHwgL8ymwErt5en2gqx5NiBcp3heZegQQ7BDsPwJBmqIPvQhDWKOk/jZu1lroO5
JXg8IzgUJmLbfmiXqfnuHej0KEzBu16KWGaNJny2StyNBCSDamR1d5iIF+p7jMsiTscKfLDYYuxB
uKdxBtGSgJrU06lTy6Cla36RA9eDRP+7uRC7yq2cwyws+owD8SEQf9QJvKfz3Qftnaaz1FQff5p+
44UAoS9IjYBB1/LqMKtO9nR7HUxb753Vn0JrzrvAOQ8zgfLKqqBUaknQu0h/5wKbotMN6+YJdkKH
enfpCQaALzodcBv/Ndb7hW3jp4s9wp8C718VrDC9YLpyped7ri4xIX6CqLlr5a24EXHB8DnH/aQp
aTUdnv7ljTTYQuM+pKGRsVOwFFIOfdzZwuyHTHQszMiNMcjVgmgVB/NufmTKSguWE6gDMA5k3qMQ
NUcBIk59BazpASZa1CuRsiKkxs8Y6Ng0be5mju/uSq+J5mJ53ME3vXkzXS8Mmxf/Nbt9hWq3InUx
lehW7ezDrcn/aLSCGv2dFOh0d/Wj5WChQEbiJr8/YQCv5rdp5aPMSF/IpQoersEt6cZIwS+1W7ty
rG/Fpnt+T9CZnG4FRoC6MyIbxwcpKp73kcoRErs2fwE9GTpIkNVobbh9LXQSWLYBghnujJ2B54uY
BJh8aVDzw268u6Ir2dKVGNbK3A7HXesGWKdCKjZghE47yavCSDepxyEQXX3uLhUa2IDA08VIcPcj
KWkfl52AgKgiI5/CSWcUEsJFAe56K0yDHu2580JvjJqktopHUn7hNEhpCQ5O5mGjMAmNAXUYW0d4
2mMJ0HBkhVn9oJZFqyBWJgCettRt/GAe9ZQ69G3t/cxWu1tNBHIBRKjELHkEVQ2fxBDZsX+KH3WZ
98SD99ofa0XWFPlUwCnrUd/Q2vYi/nPjofVeSs7Sa/z5WbIWLNXN3XxOCHeeifTY8D7iVRVdBrPa
Yad/iK4WgzbeCzpcgFkAxtM9Ktx+qOf+VYVIIlKjhJFSL5tR2r8rOYPLXVg1H6M4CaOx1h97Mndn
pyPlfBB2b6SPSI1rY91cfTrQ+poSVKffh1udgf+xXLMnolT+s+Tw3eC9ljvBR+3bbJ/98j5cSZH+
b24lEud95xn2HInhhzTK+cJyepwu93Xx2Pe29LNmLJjGu7LKzKj7pcmvKoYWe2+tJTNoXv21r5Ye
mnOqNRzosULJEMB+MgDlCuEeMQHE6j/8+Rykx2q02V/hPbYoaTUjhIAOf1cz8eJ6jJ8slS12xh6R
kQGuRsTljxqLDWP2Lnuq+debMuqXlXR4kL0nT7J2RWc4atI6ngHC/i0isrkUgL+3Yzf1cFdgXSob
nMT7iyV/CyNSQQENy2nBtPTfXaiohBFuXNmQqjlV42kJKJbfM9uqCVYwPouiWcmxBp/pQSe69YTc
6fWHx36hKBieOhvzaLH4PM/TFZ9SnZp76PZRcO4J+XbX6iEtA90BQ4NcEntro1n8NNt9VKYa2IVt
lOzDf+XKh02WUmQc13Pc4Ydv0dpWoH2uI3dXDqXNg3Xj0mDIQJuefl9Ve0ZRuj6oP7xgBqH/FRw3
1v9ZI1Uf5w2QZaJtzfABmwq2mJQOYopSVEsu7kl2LmBJC/5q9oIy2GJ7zrYWBkaUqS4Dbk+danyM
RDnuieb0NzRFDrU0XWJInebqOB2tnziDnBLKNACogKrRZ15N6krdTnhTwOsEtbOh6NbStnaecvwG
v7raFkBROHJ+iiyrMGb5EVI5GXO5guxKiKRF1OAfIvq8P/vfMN76XjDZvMkcuckBGnV4oUsTYtQi
+OxfBbWsmaOOcD8mvRW9qLqB43bnYWVedchvblL6J9N5iVMnaRUS6vRXgyEKn9+qWViSPgKKDn5z
hY01F6cu+o2/ghw9tquqKp0KdlNF+mBEtGIfEeGLIUhJKjeTzi2sP9RAfSFmiu7YE12hhuXyisH6
Bh1NwWd6G8TzZ5qr9SKIxxTAuTglMcS1VSIJNc3AIvi7Yb1XaSK8nvIsadSL81tg9nj3s0f1kGBM
mlaNuO+4fkNZV4ZvDokG6qAFq5/eTVtduhgT71FjXoOD1WyZZaEzStsDBxkaAE9yoIQG1LByl+qi
i/UhDj2qUTyd0YX4OtTwOTMe+nutKWtAa7TdXRXpiCKsvhJk14rl4GrQoAPaDtYGWS5byWtUgkU4
83rxRrc2+growoBAVvVBFRBXRzUj5GXxWoWesHd7rPpNnwh2Htu6ZMXlDzGkykgCM8ymY+tYmY95
e410o5k6yeZek/6KQj4CCorPdiusLoM8xyFcdfS1/M/gcB2KFw5wXcXeVSOIS+HnpYRG6EXcg3n1
WlvETHMJSf+1KF6dxpQgXmtPmlRKSZgJUtAQolZE4B+skCsol5vbqSlLIwAf9W6I/qOGczmWir8B
3IbkfiGZZCpgXHcsaVSw2SmR49TAxsdKc0hzna4KpuP3EpvEos/4hcv3r2QwOM3jNP/ldfXE5uyT
MBtZEBc26W6t7hnR5siMmc7t5XWWMWTbS+NO6LWbr/6Kk2c4o/vBukaIA1nlE6VkZEjOfLr6ysL9
s1My8bYe5n9OAacZopOquCFq9D0yGAOzOKLLfO8p7utAc0FQMr6ltdolV3mMoFhiz8ymkJ8YD1Kt
jWBj/80C/9enw1FqP1wLTZijsvBH6cjCdmN0W2hzZ2emg3e22+xlUPreIJ1hsSN/F1DwfPteaOmr
fypZVtR5YJkOBkupCd1vxRwaSj21beAvQ+Csw37z+QSUmWjX99Dc0QEdnyRsmvTPnSR0QwuS1621
14gkS2XXYPGLKvXOwHpracVmSZevY8tc6qHp1+Yc0altkoJOjM8PNOyOxTWgSsaW3KiwxKrFuBMh
TptqwqXGgIWncPUvsFv8UYq2yO+xTEI3ScbK2KwcOYd5QdnR63xlOWokn0rVR45VMgMsYMCT3QLa
3TafRqG9HeZpF6ZSs4eBXgG+olYugkkecyjE+dNjL/hr9EUlEEJoHbETYjrzetVy09QPPbMiYzLr
KhwsTovJ3VYS1aTuB2zjJEKGS5vcN2k8NAQqPdP+ui0EqAs9FnFnpt7fseN8nu+rxTmgmmx0H9Jf
IN2HLVKlOUy+BMDQdrz7ykPgg73MAoG/u/nQkVEMCkPJQoWkEtlBfil5fd429YB0tU64sLbwq8Ld
mQKxl7O1RK1F1GQREVHXuAP/XFO+2M+m8Uo/fT+dh2oY/q0YkraAy8aXirZSehfxzKFm4cL1oA14
qHIgqileK9ulT3l04lJ9JzvgpaNqVGkmvJ8UBdMuuKmDokyz7vA0yFEiUOmy/OLyGneSVmpEiixV
DQMHtr6G1qAJ1UdMBX+gNP5bn0kRUAbRtg2JvvX+k5LoqS5lS1TZ0mYM89e9V/2P7pnxHa6EeR6t
aK+V+7CUOrFBJLrtWE+SeeguBPhCBW4XvwAk7rjuLlzwko663uKP4o0cU9CWAtS4l7zU8CeK+B4H
wrV0jd4YDVcGIekDHtAllnImAM+F/RYZfHJwX3laOj1jhrKlseUVS02tYEeXkbT5bLJOHo2Fp1+X
KmNbW8mAVR0oitvmfDy+giOutxmXVE1b1X5CBc97N44txT8DOHCtHaL4RsNadxtf6vT6h76ynNX0
ywsV4cqNyrrUhrb99bRbtJd6W7tCuCh89VwdhMz+12NQsp6Wc62danGGpS+MB2yzY9QS0beD+/8u
71yntCUlvAu1vp3X3Z/Bm1QtFVauIh30uS8eu9czkqaVJQ60MxD+PtD5oWYPWoZVXaxO2SlLD9mj
o0ds4sZKb+s9RbgmnzM8JZsl14dUv/VfTxH8rGMt7cULCCMe3iEUe9JK8b2gZcCLNdLyeG2D7bOJ
/JgQuOwPtZ3uff0205/Tib3VslPOtK62PKlLlcf02kNqfbnPoKX8lv36Krz2LS6zEqnN+bjIxcif
BYBkyX9ODrqF/KSxXIhxYVMN+rKfhR0SjJWDAqs9n33utB+sY0OPmt7CbBw8qHCv5iQmZERHM0wp
nqnjIU3iQQ7RXcmiuAOZEjCNAK4vmRMjaKHqnRWwJO5DKGYTNaqVtf3jlanoRoy1WFoJZKB3G6CZ
bATa9TFsoDP2SIX0ucccbZzflv2U1BfwtsxqFsZ/xUkw7RdGSTnjT8mcVmRntkshSZ1bpT7JO04N
fyp7oUrX5QzkwflBIZiezWwqDUTDEkjw2SiHE32idRjtw4cLwM8OcDgQ9eDvJHD7+i3KpILL+T3h
70tKW65MnYi1LRTGIT7wc5B8miBHAOyOHbPfzLChcRBItSn9vTr3uIfLo5X8Enfur45vi3uNHd7V
QnNxLBLWxju5blWnADxbRihk2gL5cNT2LkpBrBUIgfg49vb3XQrlqSnwO/5lS/kyvREfHeoZ9dKJ
Vpk6fbqpCEGQ6LpJCbfcZWTVDfbHg8j58NGq+qvGUS3EJ2+u5JQFBS5yU4jrCkFfxQj6L/95LdNL
XbnXJmn4eK/khrlLRldmxgE/mJ4SLjREa0NliN41XVpqkk0UPb4IazFQXmYZGS4Ut1tIim/wiU5X
0e04UlU9dSu8u1lvRembmbYjMSMAxILJJyGDaQD93iDaU0S/IHkV7tExl+ykwjhVqzp5uJZ6Y9oj
klKafoJAJOjnlnEC9AhnvJJgOURdqS0VBPb1zIvOcuUkUEpY1WtGj5Efu+fUfPqLW5OJ0sxPba3V
zNQDmL8/vJaSDhJybCoZ3kTF6b+7EmlW3wlQysyNZ5pxmB4jm57csBYzmAGKy2Ca3a5DiNQVhg9U
o5VAhPCNDuKbm9IvvvXQ5Ae94iKqs+2XB9j8EcGUxY4+IAzNWIMlEi1zNdawN6LYr2lnQ9T/JYPx
OVqbjxheQcL2ynVnN95ORgBHYlZd6LZEv+/Myp8112+NQMZjxByP9RNZiYluGZNLgj7GDMLz9YPm
4srwOLkcPo0UUA30T4yXsEFNCbNQU+l0bTu8VWop5LANE2wRSiUbmZ7KKQ2odrryZktFendNx8yr
RjwJYMMR/H2QMfEqKi6lKwfqKs2r7GfzSD9tQ1R5MEuRYkZuBmu0OVsjl4Dd357nCQnIeNxKFp0W
4f0xNwT7DW8tLnWE/mTrIVvZ1kOafncbnO73JbO9AxrUVJk7FCFPe5y4H9qG9F1LgIOmEBeVEqts
/YUSRBbNYUVLcQvZ+TO8G45F6/Dt74QKpilkBde4m/NnpomoozxjRJsnX7jMGA8McfDrrSuZCaCc
6LymMz124AUoR8qbYthbwWT8P7Dhhfp7uSp0Kn6c6EnnwzU5iAsPWvltS2tJzvMd65Tz7Li8opYA
vcWn3Q6SXTxdVxww4oL4zQyqtiPB03blkal21wsBW3Ayk3KAvM5LLdfa8ZUHyv05HUk+Wd/Z2+Qa
Jt8ls8zUHSdzuflNZbee30We5ZE0zOIrZ3YcAPE27sBR7HQ0HhmvuvOoT9lteO/p0eoVb+F1CKti
M1Bm42bEQmMNIGzWi26Uty2KU/d3yAwAcEXmsflr4TbBhzdJReERirQdGp9SkX5uh6tQ/nX4m1Xf
ylQ8Rdq3ZzWGnA8tHxBaHGIg5R8uvUZg1XpscbThcDkXQdDDucUheuTuTi9IUrj5tY3wAsho5rQq
jKwV+2XhV8WxMSIKrQ6G1F2K4uVf2f42kKD73Xmig0ySTBXTy/nK2wJwbzzoehRIvRCciNg/Hn9Q
kO/9SbJrd3vU8DkANBvd1rzNnN/y0wqmBwpsbRBOjmksUWgzKZVfSzg1kSV8s0E5iCT+a7DwYl3v
mUxXJ4WBrczflaAM/4QEAXQ0haP39g1gC/bNHmD+5OpSZCYLJckBs7e17Bh7EYMfBfjju+L7MNQ2
eEUu/BTVkcrgo+QnL2xeZHFTZu/aKw+1WLoftISHEczyH6MrbUMoTNDwo5uLJwRtDZoIZ/3R54oB
KjhFzp1XOprKDB27FPTXMID4PdSCVr+E95eu92aufIfOa2XVNH71Yw6T4MqRuN651BRYkms+39q9
re34Mm8CUlPBqQwaZ0SKzs60HY5iXcHXaMej6iRohEqn9uKXCb1uGUPl38n0lmbe5MbMbWm29oI7
rOxBXdhaYdQ/P7/lxfghBvcOHGY2rlWglfo8dSlKMgboXT0klNY6Ss+/v41MjGo1XnRyMxlUxmor
LUVuLPaY4gxBocUfJyTX9CkP7by155Z4VIjatQrUJ0gMbHCDpZz4C/r+ybY/ywJgAZlnOmh/ObIn
LeMJHDM6niiwNM3WDBKYo2rBIH2yCe9TOTbWt3/ob6/VFmsBQYscCJBRIt7z84Uy8Jv0clrDK6bY
lP2Idc9sq0ktJlZwt3+PPFxBFkZSK9IfmYI9je/M5Z4nddhyBnEYZDzNs1RBxZf9YsFeKIceKydC
rOLdXps7oPOjQ9snqqeSQm30WvuNKbessGpvCtNiNR2JOh+xL4dg/rpqwkC3bMLzj4dJ7kiwEHOc
zOxilyYEuaoXbw/w9pPMAnxZXeTtffPrFT1UtzB/mKk37vJ9EDPdqTMa0vDYmCbVtAgyronmryeG
AkPfOTNjbrCKnLhILGv/0unG7muv2V/6QK6pw8BJWdtfnladrmx9Ti5c08h9cY6f+vLJZF0HCprt
nsHTYWC63d8EtZejeV3nSNBPkdA6vwOpkExNAmxj/jYwQQNHVNuWOMdYTT6TRNthnXOPS9aITDby
pVpjaPXbtu3jm4M3KqEfNC5Z3P2uc8XXRgCl83crSH9n5t0kzObGnGrUosLgSfAqcffxCM83Rk6H
Z4fTRsKL8z1S8EQwbEJBkl8nLknWmD+C+aSpxYRQ3RGov6fH35pOVFo+hbuFFcfa282br41syMyf
+ClYGSto9zMQ/F6ptu0eBcLcF5vN093QONrmzNy2zib5Ert6LFsb+n9L/Thuv7i3tjvJdfg4xB2T
cP9nhNbl0t67PNYX85wlFJtI3oeW/Zl24LpZY3aKXkTBMCngykzdOJfAWIt8qPRHmDFXtIbha0E+
i9oFDYvn6jM0b+lRpfAL8/XzJTaTmpL+fuMEIKX/+WjjnEc/2Ri+OybCxPXC/BJyPrKvYC5GdTB1
EjdAi1buQxcCimYMvOlsdBJzPJkOdVWQI0ho15mq9O6s5eZqymKCAHHSHEUWt4uzSnN9i32TB030
ni4brh4Kj4G9gp04cqS2SxDyIP1tpw39wCatlBbamU9/7CsNDVIhnu0lhDVj5Y9Hs4dwfvYUgPPu
9pOu0J+QDcMedYoik4CGl81UeyZHloehhABfMYgSzLcqpbPKvG1hUGkdkO6GaXolSYBhoFP3cZx5
nHGqA6QBYCwVn0/XMmOhAGB8CZX652XVucMgl9BsxWDCftY/ld1+BDPruc2wMPVMpFh5JrWufFlJ
Kxz77PvVlYXFQx3ZvVDc4y5HLeZ79zgYUyfZcWj93d536Mhbjw3MPgTQl6G2IIyKo8t8gA3xA876
wwLILxf/0Scmg62jrAnGLsnFb89yIlR0FZm0Q+4clkeqTTFpBzz75lU4bGf7XNSrtzE0C1EEwWVY
xwOptNB2M21OgaWXCZM2LXE0otd62OTu5eBlSp9YY1HcTJXfw12zd1UA0RYGPWb+9P04y+vVj3J5
0WAMr5HEHwfx81jenhPy9R8gVfborOQNcWfYDI9wTdPrtQKtfGyEZP2b0cifusZv9FpL1vct6jAk
9ZFmSObWXdVOgnKtKwb4IBwLjSh9JUtyAioWN361TgcLX5U0N4adK0SVbuOhoxA+kbv1yXzGsbVw
rKsGpJdk6Y92XbkzVEJw5kWMcrkcp4vW2GuwPXUaQeNVL8ewYhihSNpCemXkOL/Gek431JSUm8kR
8nmQyDIpJvpDCq8WyLcrDJnnJNsIKgrR6mt9yL/tJpGhWpeQMp4hyxjQSZHPvTSs7kW22zh+//Sf
UYd6pw9eqq5EylxXZXRelEv/4oGR1K8zTEu6JjTOBb7SGJILUVWKybuT+krH1pcRR3uT6xKqf8jm
46/eL14+NVpTnGFX25lEflp8wnXDX7+PoqAZzjIW8wn63lgd1ctm7AyOCdhBUgRByn+gpNlw5LOH
DubslH8YCMKFDcgrbKuF5IyPKlp4T3JP8PqpAzGwPyK+S+EXpMzjKtCO2FIUo4eqQ+cbTz6byPVj
fSqIP6Js4LAWCzO7Vs2CGbaYqcHKKbiazMMAIGUxZRe3f9ypdvy/9vH8KHTbhjFVtTeynh9UIuW1
aIfJOGz1KuRDq9B4OToUxzZsNDeEDOGwRpSv0FDRdOuTlST7HDZJz9Aa4oumOSHk3O452JvFQrLt
k59rtGzwH2jvGkrNzxYcxKGQ8GPMy84F7jlz5/GQ5UBTYSPRRU5UXPx1i5hC6AkCbz7eSV8RYljn
FSUDc0/GPFCZrQ3gk6J1I9R9N1kAgFbS7mHvc2flZdq0qWohS24bndCdSiJEkIvDhbbVuuvBl9QC
vdHhvuNi16c7MQpqLbqVD2M211MVsdCA9G2ME3gPcTaDG/fHKi+QvAbsY67JEtYoA4Ba6osaAOJ6
LkfqG/BkSzvw2ii53y5mwlP3CrJlnDguKAy17I7ewBL0bAFwzmc94jcbtHG8soMRsjP36srqis+R
wrPvP0kE7lbTkhJ/RV/lapbvuvuB/4NkhRomxmEYSsD1UbE8BzQ8GkmjuCIhClwnpykrjjDgibtJ
HlZ80SPfchjbjKTVjRZ0bGzqHh3PEPpIEXjKBPj3MQKEDbyxwOHqKUXzj4sqxGSw7/CpTIjocUhd
+qhKHgbW/n41O4gyjfYfZYRQGXs0RmIAwZniO/OpQUrKWIhNP42w4Viu2UqSLu9SZXO9Ob3ZyGod
vv33JwKIi3WIpymFl9a1JfXSa5KSDfwifCR5DmXJvWr3DraZKnANive2Grix4hG1qPM/xPWzYXGX
t2EtkEX44EuLSK8brA4CUL9HQHCsh8Lodknbg6pZc5kcfOmM9dTE7Oqrjq8YKZo6sRBKAkFJMELj
BF8y+BAGbNgjP9D8yE4OgLpXoe6o/oQrfbB+9djTxEyD1kq3lZmaICSExRupTkQexHo4TiASbgAC
XlT3XVD8FTKgj4qcYzzjhhckYmkabc9lrqkqEqW6Jn1LcoKoNmAej5zp3OWMhsOgaB4O23rK/b3J
R/k65V+6ONPvAMyBQO/0kjF7zNMTZvvgGBwaEhHc2ioACuJOuAG+8Xlk4fix7rIDNjS0i5kSUZ1E
PhwtVR/oYF9xH0dSb8jRCS8p+zQpt9p6Cpt/vnG6WpvCYMNFXJKY664huSPbfhwHaNam90O6W2su
cQLG6/9a+5kLEKbQws/DlOVTL3AKQeYR21sD6OBf9ysWh0CtsZgENrRF1UT4298wDjXWOxmMn5bl
4d1Vu9p2U406dz1uTqXL+ztGFOLYXTHXMZlduSy7ejBFg6jwYXk0yV7jWIJdIsnVuHF6lzq9IhWX
oHauMttVEz8vZ/iEd/t04i36U/LhbegiyLrePyZYi+pwnIEQfMVsZoB8vVrIeca3zYjQIUZSzlxh
4w+6E1biNb0C2bp4veHBJJjRdDHBGUc5gQPPJt+UoELHOoLV90ZEfffuYNY84XrFEc82CdIEKeME
gaXNPYStOADx/emUGd7viqB0CK4hVGuBYrDTHLizv6MiYS9Y6JSSfY4SvOJsykBX9aNNpEA/SVDz
lB104nIeiuN6TpzKGPEqTXIidYfagLTT/4h99NnwRn5u1TrG8VgKSHIMDYItq/LU057gX40ld+3n
dc2eF+nCdjN1vRaNREZR27zkDRLGoOfVRY+ScQYX9tcjI2t08H4njTD89aXb50DbjO8DhH1n2KP9
9pthraEDg2sONcwEUhAmFKjccUlbaIDjZlbcItTYhT6e9ylQQtDQj7ItOGF1m856s7Rq0rxUvprw
h7NmbozL+QPkVYMkQUts6ILaO64t0rnuYLPbuGVfB86JrVcBRSOc9hnpmi2ZEE1v4RFVkYwH+eTW
RojFqBR+TEMzOBTACKQZqUx7C79EvaReAHOZlUnARItgkel4CvwMvHXz4ocxnn1vkr2Is278uH5q
thtQrg9x2AYif64uHaCUQRg/Y+bvYkq3Ovo9651G+1NNvMO2ViNYZ+shbHxBJ1rWdqIwKD+J4Go+
X1ZKIy0vIOOb2lVqEFCvCebeigJTly+8lYeDuK8sVJNUU0VqaPvcPZE3NNlRVZPd+XRfNWfOvYM4
QOKe6d0nPacUtoCoeJ2Z5rvYXPdXFtjU8PqDIFIE5J8r/FBqMqN/9E7SExhs7XIh/Cxv1R6NF0Tp
80JDs0NXckCXs0+agAN54R7nHZQkp5uagqRiVBzi5CCKoMymYt/ZdsBqDc47cD6NgsRueXVnwnzS
6ebjhJ0fxUfFYe6Il2yAU1FgLEVS61x0H1k7TCLlIib0tZamsUoCetTXFxE54yoCVxQ/1QQ4OMER
2nJiBkqoBoH7eXT3aEq1np3KQN/aJN7lzNBLr4q9FZpKvqAKXsu7/i8eLaH9XgokGiKdUMaQ2j+w
oY2x/W81EJMltQtaZzl4lyvVenYHJ5wxIBcqZatjOUtVnD8H+KvZbL7ivlZ9FxkegAsogkPAI1Kk
R6Blzu2nGWKwHz418+e6gXO8Bw+wFGOKxbHvH8sO7YwbX0Oa8sKfOavkeVw3Ih4a5GItDSbiBOoP
9XpMG4O5lXnXMSk12SlCnS4zOVuZib40dpwdFIYD+OwgbTl2GabmoihN/xg6hdzW2DYWDov/gM4B
6A/j1sAGaca4vDY6tztoPfwGbxaLF9Bhcrj9kPgx3Zfx2SjQCqV9ZxEUU4pSJYNnP4lmWl0VQiyT
7warZtuQ11svqSE+OU6R9qUHhrZky6BI+F32ZOtJTmlGE/HTfewPebkl3FHkjHFP8iC4hS//9TzN
Cwlz6dT5Ip+4PrJWVBQU4/JEvT6+J4PqQ66A/Wi2dwz4iGuxYv4CJ7QUOJ7KWJtO0rGM8Q6R7qgL
H1IOEefRWO63MVPT9OtbHH3dt1mWb2OTWpF6KqMkclqTnY+k+0y2n/LzAkOTiEh5qnmQbcjGiWA3
/x2Mm2K6GOXtbbLUJ4aNNZMBs0VEhwA4Pm/3pZiY1ruQXIW3MJFKj40xgnYzG3djbKkTQu437gaZ
qtE4AeNRhpiUh0niYOB9oD1SDDtnCjAG2Ek4I4c2UIG5eBb4rqE7n0jJYXeJYsJNllShQ2PO7yT1
ZG2w+Uj/lXtVdFOFZpGRTO3i+nRfXGy4GUDivW1qLQNQkqV1K43X00P4RMxPDyXafWQ7SjK8tGJm
ywmG32mA7syhQOuGjiSpBiy2SWHk6HjSbGlyS/cvSiBCIAr18oBTapsrfn/d1diJi/uH5F8xTgRZ
YbBzo4xAoPsPX6vDDvVHwNrqQlO+pibhD8qGlKbgT6SIRF+PTPFh3fFZIfQ6n/GUIvCqqBK/4OH8
/aMxs3Nj6ASOaEIcdr96np6ng/3I9A3YNVEavi35AEkFn3EZItYj9XpgEpJ7EnDGIB+D72aLboMc
7kkyB6l3PnvDZetb7ioOOLO9691MbT84ToWXeXK9h0tjSxVWkj9SLrBd8DVTMADfYnFh+AI/LZQI
ngfwZJpThhTpuUSR/k409zrJ3F6EiolYbVtlzFSN/IBkCJtPw/fwYJIxsogia+iyzjNm1Qwk2N7G
I/OOmxdE6h15ye+poDzEsCftixg2s6e2xS91Q8ejfKfRGJJEpdzK8I/4OtyQckPH9h1BZJTFr97R
tKY723++ojt+LwQod1rYxSx6G04D7U8KeXCYwEUCAIPSionO/j7SkJIxF2sScrBskvAqIi30NKZI
WaQ93Lv8m20kGj1zHLC9Ok9lad8YbNXfAupdqiPR2/X89tM/vmt7NLR8Xj+tJODUoeFUbW1ICxf0
UBcmA9hej+JKrOSbCr6lMAbgSyjhm+PB2FhTzNbNVznIp8qRYqWHmO3sN7neKxfIqE9gpLBwon5r
sEou9E6l1uR9eeh1HEAqwA/vG3GcxizMSMqX1kGOPt6gqurl/dWZB9s9aCSEtPYRM7wIzBQCGAPG
pvaOxTaxDYTw9PWo9Uw6jAO3q6qEZ4hTyBXkMC7SD1HtCaMtwZVWEnNBbktj/IAzTZ15VLay5e21
DoLMfc0EfiG3rA5xt30T+PpGTk8Jvx7552O74kNgjwLF+m4xRQSx+8LHJlBkEURIFQbGbAToChBW
tIzVE5PTsZfi5RTwd7A+9v8HDIHor6dDn7gM649A78N9zcrJccwNvAn0+YnEIs8OgLZNModKX4Cn
UTocmWuChtrKd0bvZUmKB3F0lULouAL0UPWbNQBdxxtUdxjdeHTXga0zX5xHHyms+WvKc93aTp4O
tNZEEi6dJ1BV4sHIEN+53fVvZvkZPFsbL/3P5UHAOd5JnxrDj6MTZIm/YOtvgIAzNhd39ZatqEcE
xJ87hJIgKfc9cd+h/oMeetm+ilCpQgOjt/w9kI+wEU3Aj28/L+HLfK19ajpxwlPlWaJhbdhgrUO6
oAlugJh3z7OwbpKnlgwaHDMecHe6uI5/AiC/9Qt/rCBGfemPECEEi9ZMijFQx+Y+sF+mf74n+k2K
vZIiF8zXigHaGQ/JV1/WG63iGCs48RCf+qVLEtVB1bouB0YDaZK4MPq/JHSj/JguZSdrmzmc9eDl
hhmz6tdw6dzm8VT1vuPYF/BgTOGUAZJZ8S2bmg8dLF05A01+KXAV3FIy8x8UYxhMpzz2D/oyl+Po
mMxb6L4PZkNwV3oIC6jutr5d9DNxuXgjg5vzqFhf/xngcBSRLw9/8rHWxcB+W/Xt7KN2V5CypaJS
4BM0bH9JV3DCzEusIYRhhUEqrl3Gpc54dhwx/vdQgzuxSD/GsDZU63Nfc++duvrbXfQjtE6ZWlHa
a0stX3N/P/s7oFa0wI+lqvcOqWtlwjLQ1aZDSB+g1ZnlPUI0ta6YlH0I49fi0BizBZ41l1N2ua3z
pBQfCTId6gAvMKXuFUS6DeoYHcmlB1Elc2Qa2o+5o/yp1x3LsSJlA9OuLLaa8zItHKeUTYwUXMZa
+fwocr6nxPrhfBkCq0ERRftcHNeZEuMIlxqfB4NlUuGheXBW/+G+JY5qOLR3jA7mBqr4h77x3EaA
aB2HmDP3NrLGqoF8lsQV1SAGiutdqrGqZKE+DAyD+v5P+xitwco9gBBei46jOMhWROTUlQ+Gt1Wc
OcDW8FsBoM0wRznRsM3cfC6K24OmzKeNXnkgXkN9MV+2I2Uws54IaNMmhZ5cACflisyYNpZ98M57
QxhNp25HvyYvkyp98fMSBMSo+pf9RJvyMwie/ft22Hlq8Hw6mOrrvzrmsPUG8ACc8xGkkFJdSvj1
nGF4VN/m9JbWcCROp+rtif2Gizk6P47Gu/FwGT+eKLQlU+O7aUja7LxZP45t+W7NOChlMRDkJHNW
zN6qAl9s5/+b9twuwE4H7nH6sJNQ1oprRj/yy50kUq56WiFTCWvkhlPXg2uM1JLCqOXMZQiDBSz/
P76lRI7aLbnD+64uVBs7POKWGpQHrYE8jdejOvmZ98s3PT1yTlRDndqQGJ1y9AkLpw5xQgSp8gbi
FSuhjw/6RCS00BRfcUZ02VPCXimmbzji6jxajKsKGCn2SLAgyd1eG2JTfDzVe3G/Hluj9dFie/c/
grlV5Dho9WGvNWbw/naxKPwy3JQrUWWFjdb/72rmq5bTuQxFuFiYgVxE6MVKSJBQWMy5jvkUzQqJ
y3Fdp8dbvT7i17JCBOR7Zn2rAWvbTQ19CMizxgpTnEdiHzQba+3wdtam7Rx9JQbx5YImOLsOj8It
IP5wOyiWtHd2khW/bIw/+vAXG/2XUOEX4quSwvSdH2sT7LZQ4Be22w4Ax6Mx9TQ0WLdIuO4MYpmr
rbsMiSeDzjWmeQfbh09F8yMq0E6W0UD1nbShUrXKzM58xlU1idfjECeXxRPXiU4wfQgoiaAe+wrm
RcJsZPupkvlxQdLjqRf24JbsQUs7YNZDKEIr757LqOC9Pa6acGtubIPbgAWnRIn9ylguQsDWRSUO
kqkwiaCad+MC2/SCDcMpjNHoFJAPBBE8mK/R3fbl+V2ml4R97ND12kSGuSKcD0a4r/cLwNKCvP8V
QrpbOYo20ZtIWIlAza1Z4piR8PEeJ6xTM6rfFUMNjAFEdk8j/cYG6v5zwMC4bZ2wXU9RJw6q+ikt
IGSFXzWBGUVO+K1mB4jStJyISBapbWcY6Nuhj0RPWrjK0/jE9iVoAs52lGzMyM/91+dde37RI3Gg
jJM2tnkbmdAD2xJoA5WqzqIVkfzGtISALeiW3gWCplHmqJIsSaLQP1LAaboHi2GkUz9BuOVQMuhO
NUSEK1gSE/yDD23hCSrx7PBTUerNk+VQJVBUUSHVf2qb1zH3hlmDOS+rkXI72OtMVAeSKyX6YfiT
IjltYZ/uDBdRnHCUXOOERVdAuK7EpOBXx7zWsjx+0y+CtWY3n8R6FALqvgW9Cu8YVLSYVamJLH1Z
kLIz+rmB8tAhpntftvh9wu+mAkMcAxymtB6KINZepd+PxM8jelVrmlY8spnV2oxqJFzgznWNv82Z
r20GDx42tPjZnR2W8gLooFc7KzFIPBxh/4+IBbn9il/3pleletITDZ+ZpoGWS1VvcFI/lsj8fr5H
jnx9uv35AyWV7Er3bUrnLRKXUJW8zYJY06jwLDZxg1x4kuL4LNfHRkxVbferO5HDONBXRxO2xkiL
THlL7IHUf8/a4OnF56qwPOWg5RGvrTheq6CFV2mr1YElGq0lShMmQnGgjL0S4dow8Ewl4TMU7q3B
w57bwnEAONm9maHHp+JmzoVywYQ3AtDIbi6/AkdbBZgIU4mmJvgF+2Tt+C6JeDZy6dLLEftAXgsX
RZiBLZIrg4onO9DXPizH9vPLleRoxc5B28FOrlhb74jfJXl7FNNN+USoJol0cIVk74WLmXxhAPF5
L9gnzg/ded6r3ladHxKXHZCopqWa32oIgBxjgdByXFpOdmLrDkvdi+YaSRGX4UIScCL+KQyeOAW/
+xXYohG96d6SOGaJkPbWJRL8Ud/jZuFIGiBKDQUNy8Fxq847NuFTFksJQraxu1WGOz0DJWwoYKgx
zGm/ieh3vC2/MhfwjRZyk0m6zZiPcmV4FSPb+Utw0Rj/GGOZffWuCF2za4dQWfSncJLmcQgp+8td
DXAB+mJbE049GSJWyPIGSjte+U1qJ97cEsHgT1HMuLh9sawrr39nCyIxL/0qP/1qOnv7aiTkcLfF
37dcqz2aNTrJqWYzvzKA1N7B0EQpvCfSMyXcY3+zJFlAPgQnNDOlZCuRsjcynPFf0tDUBMVo3SGR
RtrlNZu/utKF35SGN7GLl6LZTKjNL8LCO88atPs853Uw6ewLfRxXURlfdBJwgEGvxO6Q7YNFqHBk
frCViumAQCJ6LAuYdoBSH9wMhqNmmo2e+gAt5mu83PZ8EHXJ1jf1GWi6pG8FV5r065EPdnL6LXBO
zjTN48dEcWomE7bvJlDRMpERm61UwVe0F8C1zLX7ilUFVdfYRGDvzgDT0nCiAYAZzlwKvesmNY9L
IZRfG9zxTb0az1vdh1eNpCqmtSIGbvM/x1wzEiqCebliP6fRZDjY1hwiUsG+vt9ioI2GmLb2gFGw
PLdr2QjBbQqV2QxWjPG7UpLPkuvBSbv2d3hh8DQea/Qy+/oYbDtvgRMbJym+25GYLY/rNyZpKj3l
isCsA3+xzawqmlcPbXVi+QJNm4A4lr+87BxAwYrlVuK/gTsV+D538qRn4L6+2BG645Zon5hOtuzH
lX9rtl+K3jehykWW87sl0+c3k9D7ipMf5cTqL7zfmr/1APwrtADOb6SEr1PNjnKJGo2Z5QnbKKUJ
aTKaDqOGd0SqvnUiN8ssC90g8gYIDs31aGK1K7vMYx2WoswEXVrAdfULhW/2Jo5/O4ulLfhKPymI
pgVqblhh4lmEkZLM349f5NCoR96udFT+F/c8DzZAjXaSqLWc5sjiNLMJAclwTTBSv7xxmtEDUqSM
uph+NqRDt0NdDJ+ezyxPDsau2+D9/QYEjO+ZiDJzPSPvmx8R4EocjHqnjW52opG0dbDk5eEjHp23
tgnKmtrxHqjiCQhXD5j+tOp2ulfFIAx+fzXN+no6TypxcQ3LPg+0OUJOe8pVyDYnBCzoPky19LLZ
BvDlDoupoFqyhZTbqycpUEcb9m7hI1Itjl1yATqcyHSv0l54yKycTxKpFHLLcaW2v2OVxnWQBmLM
ZBiw/AcT+mNSF0xbTpMnMDMaSBRs5oiK6oNSIHdN8Jse0ggtKYCk9AhRIrcuBXlr6iV3Xx8Wmxpl
l3fYUOhqI6K3OkyKnTbHx3dKgCo5enoIeO5wMA1QctGhCWlByW3yd6BSCdLrE8rVbrB2ZKi4nxrP
FPeJWydGO/jz2nZsZRRRbMSWhlmoM4XCFC1gB8aXysC6A4izHUKoR3gR0b1cqKeu8aVo65ik2kZQ
0Wv4igqcMMraLwwAfFKNeDaPQmAwr2rftYR71Pj3QOGCVb2ujvW4nhFE+gjV0D3PRyd7bcQXJLAt
iaESHDNm+qaJKIDwxhgigzUAGkTO2lHAc/Qsrw86Y8LPJqgQ+uDFx7XP+y9nqaNDo+qcdCRLBz6/
7crnxY/UdCjgtBnp3sNeM5182zmTb0TwSFmZesQlkgKcUwFNJISXzFSOEh8bPeK8vn6xZh4qOOon
lpDI0CtdQDFqFxaWr44gdzzaBUmzDMN2jqGmmbQ90tvv+NcrHE/b3yKzTDMNhrYWozeLTOBqnKLo
SZisHnekkw6ffQTfT8vF3tyWJ5zBtfceOwMRTyRgOVefny6PYVN1RmNLMn/SV7+eH/zHUnLUqnjS
cp03pEIwXWCNN46a9mgESC5zYnaqFonfFHlVHleC5esj67nyHQReiXriZK0KWJJIXtZAcdpgKGmt
j1TivLUCqTlR/jzy477x+32h6t37yRyHINZtKX60Lz4DmKPYs018wx3DDtOwKDBfMKIX97+PLJTw
QOVS346GIDJX9LpLmHbJBc4+c45W+idAso5RkLFpqhHqYaqlQ/eC562WcjzZIBK/R/hZSj5SU5/U
a4MI129HfP8Vb/0kSTQEkOlpTg5uVa9KVS9NtOhT6RYThgXy/pAdvUBROOQh6uaszW2PSIbGJFq+
GSl7j0L4MIfHBP8p6qaQgdPlvjlfQuOIoxUlsPzhkDhei7dp1l3kr2sWXxfcqqoGcZhPsF5w0u8l
beAP+WFsNV4fhzSyu+cbfKfTa03saoKcEZ4Fw6pZSWOW4y2oNyu5hb3aZwOx4BUorxqf5lfKrErb
EzxFIASdpr0c9XOJWFFFJIHxbYYA2EHSFFqoAoG6TdQEtYkO4v2YE70b2PLToMj1OkXez47eOsSf
fdwNp7DRUwkCisnSVKcLNi7OOCPy6C/SypWvroGVp1O5/xwhchMDMFkUNWnK5soFNV4PXu+n+meY
eIeY61hfOYKgVcFMFCV1SDZdUa14GhEud4xs7kRPohPaVFHsXP+QBaFYcHQfFgU9G+yzCI5pHc5L
HgbtSvJDo9avE6Mise2vfTxBGGgOOPR0A2AVtfDkICoWtZpe5i45aPHzKCiP4a/jmoz9RJPraAjc
Puyyi8Bqm8xvohEA2+wtY6WE8brtmV3SB7EQy4wQ8FYHGdyfnU155F5+ttvyhKmeXsWHYmuK67sn
mmgettK5AsLp33/KiUTflNxhFL/7q/txq8noDedKW6fV3ZkfDoJUkZnNHUiRQ7xadSeeIKboflas
KzSDMiFtXcFIIcowIdvYV9k9m/5R/qK7+H/tVcGFB1MJjlZncjm7/PfoB4crukc6zKqsm0sZ7X8W
GgKUdYPSjNsUA3wt9kToUCPeAOaVqckrBj/xbyH09r/g7JY+9ng39nlgMXb5z8qxX8OAk9XeAshy
VosBnHrM5/b6MikbSc1pHXsvLZ5QsqQvjcQOcM9CJ28rRUeTi7ozJTRsQXaBC/PmpkEVW/j9G7B2
H7yKQzh1XsMvAwgXPO2cFKaN07O1cpEZ2HhRSP2fpBprzUAsQIU38VvoiYzpH0/7EsX+DUXWRlAN
PlHGSvhnMsm98maibUFx0shOHLLQxkTT/hXXRrIYBnxKCFJ+MfIXhRfscgzs3PKBCi4M2Y3g7A7X
G2EMMoFP+MaND6NGjCZniXgLCEKLjp/tfbAKqqpkt9w57SXJJJkWbPyBWDAYWGE3dsubLLOGl1Wg
dsiR4T4UreuPSSg5/mEsbm4PUmior68/lWpqnO+JfsQWmtFhlaAE+OmONzDAVLbzeyHlQdLZHJAk
w7jug79BSpVzz0zEkp/uubca4Tw4KbLwIaYq/ElvH9EWh+jSXqrAPUmY5sFrCrJxjq7j9nyvL1WA
XtDQ42f5oLRzuuame/wspkPlHY5Co0y0RJIQCC9Bi2FZqcb2mfduo7lkJynM9ESP6u926XWWk5Fa
U7In8LiVSwZylaaCiTg8QH78dvS1HMl554fjyd06Fz9CHBiAyK2fqZibQol/B1lNN4mk02T0RYrf
ASeDYvQjJjnn9tRBqVmQap1fsRDLxDvS/qYfrRRCyUYPt4UwfPc8LDKUuHzaKnc4YAOSNm3VcuZ8
dlX9HQRPfg9EoDImevELND4oTkIU4guwZM78cp+X1OYjELzaN9aEpNOBS1Mk4SjKEMzJmWSCreX9
2fuuGmizU18/IIN2lwr9M+LQ1QZpDZE1cVgq3TtD0FBDxiraTMzWw/zshmNzNWf2MkKrTTLME2b3
U8yoGpZyC3UT/hVBcNHNXaMetF9YL4HY20Sr+FtIgeLNSCn7oIz2gMdW5mxzguhhD7tmBucLHnZx
14R/YpbDhzpvbgzVBW1Oa+fyaibOgCx4SO2ma9dfICg23gmw3AMnPLVlW/QB07Rfa45vbXvuSR2l
1WR7J4gBQJfjfRHAfc2U8XZJZMgUSyxq9ZAf6/4FwYvhpX07wlQkR/hqt0gg2r5i2CwvVLkBMCUx
Iuri37RHN+aNah8JpD1XvmP4dNWk28JOR9w3trg2V7/yBwIkbspvOdsgC9RQiPtfmRNa1ebaYpo3
IhdoaXw7NR4B2CiM4b2K91vdIX60LW7+2BL+lTecWh2H7kfaFJBdjRjZkqaiu95EjgZ2U+VYf27k
enMZ965Q0GykSkygLNkFOwl0oB/+P/pjvsqNd1TgtVP5MpMwaMmAjwucbMQOGt4SduLo83PTR5qO
8zuKevogLrnfO0g9e9bq+2aazp7biwy6BEh+GAAcifxekev7gnj2prmJu75FqFX0BqL9bCvvRzvF
/z0OS7sAHCKCuchRERt1wgn3w2GIs1taFA+ZmUmBFQcGtBdnhaNNogpNnBWO0NoiWBZfrq4Q91c1
TrnxcWEReByVVb8iQddfSQHcaqKsg5zpbzUpjRVEird2eJjbR/8Tc0Y/2NxKX/Ot4BPJjDehyxSP
5Gtm5iPC9lCWFMO2vHhPPpRhvaRYF6XTWEUqLAvKs/tq2yZo1puvLOq8s1zg0OTgoXy6pNd7LZiv
gQbtWjPc3nFIhkQWMHGNUepSOlmVANRxaBIc6w+t4Y56mpjPptRoNi0JVtVx4XZW/MdyOdGT4df1
ENhMlqTS54FysiYSIPqfiavoL929/Obue6DTsJqUMKxHdQbJdKMdgMY10O0xF4qjP7AEiT53KH0J
N+4Fr131IAGu2JOp08vJaK46H8zPshXvYa4VU78jP9DtU5jCORHuXVxeyp7khqO+wgGrPaATmhYR
Ze9aZCK7Bn0d08Y1hZHAfYtsbsUAGyjnrrCzI+58UfUbGhL2d7HUUQ+sebgkZXVPLLrRs/brBVz1
TnCET/LxZmjqcefdJCwvUROcjIROpcIVq3BKXHWhYNnNcoM60py3ilCNxaRZxnD93jOoVgkJImxC
oBdfrzf+6ymQQYgxWC29JmUHMUtDwEZUFBTF4hJGyt4BpyRzAVzgTQ8VPtXvpZFJTXtBn6OC3nlm
YLDI3jjgr7srhD2E/OhGXR+wqJ05+MKBNB0UDZfVLxW/4/7M2/dwoJZZ8MZRknhXwh46ZGw1Ntwe
rO1uvW8Swys/7mFiIDw2m6uOgwR2ZK4wLafZEoN7oDUPPevbWs+VW2nlMJhoiZBCDW3zvGtpJZQ7
A1zBFJwSwSExF95mmmhjfCe0pUS5uFbrLljJccJV3hCeKdWz3faDVnj9X0ez00P9thd8FXEoAT8+
D4gX+1GbUz4zv5uU/AQJDnpShSSiG0LhKg/DE8DzQy6hzYDerN3C5/yf3M5iuBCFjoE567qYwHlF
jmPOyHmJ5+woSUwQOCgHCsevG0pneBQQzZuWgxJcNG5ZLvKM30XHjdz0XAV+C4jdZWy2+QDQ7p2V
5s//ICFAZeVUhffCXrmMEt0bqxd50zn/Vw7tNc3hvOdarPOu8OUHKUNWihCjl3pb3VVX/P59hFtA
QYp99qQOIl9LXb/41n4AclNSROOlmKlUY+BtT0lzYgPjHomjF015XodUyt3IUOPLlNbhT9cCv79Z
DY3oR3yyKn+cBzi2j9jQZ5qBy63nVmxIGr+0asuuYMU7zWX2p0UdhTjE0MGwYderPYHhmgLTXCZH
uUKJSONKmm7/+KeqCRwPhdT8X/BRM1OQFMceUITFXDv60IuqTbTluO6GBbBbIHPKOCyJCe5I8sZU
fXiXV18bCjZNOYdVSnrrwJq1n5t7yB7HaMrm3cE7oPKf3MUqKJu52vC+csDTUgedGsSI3XWuhWkL
SpsdvFtFDgbLW0WA+3uBNXkbQeW4HFJvCh71svSoJDScyQMaq/uP6aaAJmQ8VicxIo9ZBstOx3KU
E6OYdlJv/Ff99zd88SdD5dtNIhDE72qWBfZAMYUh6kymauKH2PrjoRytJttYaW1OI1ZB3O4tK7fe
Z1t3X0ljOILn7NC7EhMmy07bpPQ+cqFSRrqceDWcsnUdm0CHbUjDQ4RJr4qBlxAsHzIf0xFCFCUi
thMJ8gsueaIDBJZ8Gv75ywehNKBlumV2XxS6jFURVPo36UxhzoQkXSJ7WheHJpMcXg+cZENAcKVw
DGhbO+XfCERpYeVdGYK4dGNdlyErUkuRDkDWmHBrNb/5E37yUk2luA806EfgbQIqZ0gvkKRDVKcG
6tDQy18z02KkR2GoDMZBo++pwIBxCt2mjTyJlH0zv/2wHsaOmxBNMdxv7AVc1EU7OSZi8dsy4vVb
Cm6lXntEaQzmX7mh0sHV+ehOukJKCVFtJnf7CzCUqYvqJNy8VcNAWJUedrGbLDnBs3BfhHJm5FPU
SvhlPmCHldqPi69/1+7wdJjHSdc58bCWlFr+SkHnRhRFZw+WC0pUPW8Ayxj9bJxscICGqxF2pmbV
usYGJjAa09dnGu6q2ExupxH2Qi+4nTCxCdUCqt9ejsOTVuEVCTBM1rdDDhNEJexO8P0KtSdV3G7h
u3Xhm7Rknr+hi+3/kZNVwJf66rRy5ea4UK1SgG4SwVFmVu1SLpGJSpQ34SdnKqSkXGBAZP+mQOik
mdgaQdkbw2b0aB+WEt68PRaSj34LK9IKxTAos6Unt3iNVJuvve9sZNO/Eh/kZlF8rlZsqgTonovm
eXcuxV2HFdPss04+L75C0mOnmfqqtzvcg5mJiwz4tyFgWYBb9X9X9mGYlUzzCrMQDlJMzd0aQreP
wdljlrRg7fWHGGX/iPQKkXpwmBZ5yKtIZVHl4dxftP0B5J6HvUhRzBhS4oCuh1ARuYpUv1jcO70o
RljvhExU3WmcMkHm9fDS11u+CSZbR0G6yoAClbB+9xrDqRTl34bFkw5C+B7yKZ/Ga4yOvORVWxRy
jH75lIcxy730nSZL+C/rPohvvJHW9tqHG+u+/bTeeEIYtRjs09gJUZfmYLWFrc35bICm404wsneD
MHZ/TiS0YD0q9Je+yLcy66K65lEZulm0TIXrBeNVZq2/EnkR5yKVeSgRgogn6ugH9Uam1dJ3ptc1
mBNTKcmpwwbb6dbsvWnwdJT0gY5NPcay2QE7QQAL4jo7oY8qhSX/vkLX2Rp4CJDu8ZxJJxD18KCw
sULDxkXucQxhMYGUeTS9vpTB2LvlRk6G+mgs9HsBNhUa985AAL4vzWdQqN69nEvx4k3fjsQJxmWi
liIHJsI3JWnQMQ5B6T7EDghv3fUqPDE7thRIHN0B7Q60kx/TnsyxviSCiYh1uwhjYD5HqHPjUttR
ZgJlGlh5UR1rPdI9zgKiK5FcT74zV28rzyp8Bk3RVDhvd8AhqS3s9hvYXMhljuaBI4pGLPkwh4+x
b1suMXidYk0tsh9TYrRU9grvsXetERsjxk4pXkCB0/NdJOLO0n/CiRrLcIZwmU5tDz0Xfl6ZVWAy
AjsqC5/8+4Ye1iE33Be4wv+uDhDscvpBV86mvmF8v0O6gEmf173TbB2hOMdzgvcPv2DD5wZmLdQs
6FLM5V5sCU9MGHHURzFv7T2cWmfioozhYLcOgjjl5kCO6zMEVWnh2JSKXi6tt6rPtlGqeAZaokiY
v8jMkqcqC2o28UZVPz0dRSRHfTjSga+0B4vqssi6UKafIG7WB9A+Au3WiVIxQNrVoVMm3877w7Jq
4vruObNsQEX26NUCUOI/GYyyxt/xbkoHsbkjr+yIKuBejBwcosJ8QNIIbuJ8m7qOTs9p5aUNGwPH
lKWdAAqpwtEyPd3x5S7qTgGAmU8JHPcijFDdzrBKO3D5dSYy0JlrWA6J0cX6pUuTCaxwt3WEk6iS
bEyQW5V0Dx9LggJmbplYCKhBdr74taeYqliw3JVNMyn7pIjLH6gG/M+TA2B565CoKTEI9lbMipiB
FH0DmhN1ieyAYTtgxJzU8AffpKs3E/Iub/8BrRyNYVQ6BaM13ubr8Keg7bM8vCPg0Iqz8nb+MnL6
QLPVr/QIc2+Ov6+a4ZnvmmIDmg0XMhSyvcrvsJ/znzbOLkClTtwZau0ohFV6kJhbi87kWHtyV2oo
vqZ/Hc4GHGLn7FcZYrxyDqffmugWU8qJEVzi4rVcwcOWtxq+sToINQTYfX35yg2kzcikRTle/GgV
dJTmzTCwdfDSHEk0hKk44exH/Ei8Jds74ZPqt+WuJIG9P9S5csTq7xVDOGJMI8AdleuiHcEQJ6JE
quy7wRiWhWLylfk3yeXoM4Yiw1dBB7gzsTe7H+bUKl8zPbAB7rovZ1r9cwXXfjaoOsfX2v1An7Nz
kCTozKFr5hj7NlhuvitiqO1vxN0LjuIV02/Kp22Exsmxn1DEHHZ0pgTLo82T3RRgC18NwbvsmJ43
IYoC+KMM2TZqeEaVsrQ9v5ZjMJFcnbsyK88rv47P388UXKBbfIg+aYlQ34QW8pKVqSsRIeL5V2uU
PJJ1U1ITVlwzjOHTU8Ju33kDJ4Cj74B+GtERrnS6iiuwSmWWlSIuWrnNVGp5aEJ0Qrp4xCqFDFP1
mQoSut04eMS/Svls9KPSexzRUvigq3Xf3O6z5MvBPfVC/uJ1dDb1IA54aIe7IAsiBGKykrIf1Nyc
0g9Xt/7XvE3keCrxlhkzM0WasYfVfqaKBa9+xaYAgZRAr5JqWUTSYQDshhWyzidyLXY7A76FIl/P
d0d/w4iwetroGo5K5/cGOR1WkXgmzCYY3xg4yxHlyGrbXbs/yamdNmtr2QQsWfOFRrVyF5baKMS9
8B3mrXHwUYCKPSUnbYJEaIIyOIlLJPPIxUr3CMuk6ef7pwJLVV7Fv42JGkL2U4CF+077ZbIK+wUt
PpnhOY2O0E7hIHwcG9pNF/LcnhFHtpU+YQwuHTkfOA1nkSPtcIj1d4V/mfEMGrd0PXSd6MBqRINb
eVTVeyarwOG69s/KZ4cGTRaCqOTrYwY36ItlgO/utxL3W57o3OSHeOOBBOAO05PdDYS6Aww4c8JD
YCoARuh26EpM+6cpiL46bnoqIY696IoG/K/0r2+7szVRif6VUwEqvSdXybZiQOVSXiAzv5jAmg07
v0SNOs0NWYZjBppS5iE9mQKM5As4qFkMCJXa56gpbixrYY0bQqibin9v0OfBW9L6RktcQt9u2kfW
DMTWcIsS848YdFtzW3QsyZMikhjM+p3918QSPx+UEZkzrDPQ8BviA/9ZcH30ACjp5YFLioYzuYry
u3n6+uJIgCbX5/WFDSlFsXdOxsXlv/oy054SJgN+WOJrIRvsG34vDHKuCGc0upRuVIsR40qDIBox
ksiFOwfJ1tLI5mC3yfpjUqfys1SGkEfs89MER6XMpyXP80UuDddsvC4sndBp8LXwgwssLE+uAcFY
/PpgIVEiDA5q/ZqsawZMNSD4Pzg25N2Cj7wUM4sWkGG2uGTWNiE/mg2/KGOH/K9NUXGY3so+c2EL
Qzenhuow3I3ek2SaCksnejNXhgIh9X3t6+baVBBhxawMsGYiI63j0E669AKP1+lgNZ8EPN02qPuu
sfoq1eyqYS3rT/hk2EvOnHO2DepNYVcLrALmSyQgdLPIoZ4ozu4qHNIinSoQDXL4scrE6R/BDabJ
ZOHDa+JZ7rGlEy46P3tfTk35HniS9/ppaqixD3FxZzFURV5u0w8Qk5gushe1MVDGxIfGSOpk0hvF
VwCliufYT6OMhHa48KtZ/5TGy1DlNfHS+PkubNLlvC/1QHXJKT531n6J/pzf1e0QgQopT/WcrhZx
jlF70ChQcNjKMfEtyMSLMoUgbdWuSFmaHYhxy5cpm7dx8EOG2Sj3pytDDCFvqpjswwH/SGV7vqQB
c9uWtTZPQfiOXv6U/jbeFlo8fiVOO0e/8Q9YwwW+BVQ5EdxJLM0obvXO8fkD1bldF2kzVBrbXHB1
w1vJMAc/+nWMCCER2IQDm4q/z9VXs0PIa7EniI/h89pHVPr8yLPDB2LT90MELRDz3MobDDdlJzeY
Ryk6vujqCPiF/x66zVQ4a1gkc8fOOqi4/7q4Tw50VWu8h2vAlFiJcQEVJnAvGc30dsKiVv0Mt7Nf
M8Xogku4IyO/DdwoCE29I1s1NEOCUFjoCbXgwFx7oXh4h7uS7FVIXCRYiSBSXHv0wP9zP8I+ADSj
9zB72zDIc9CjwjcJd+69s5/66TiYdKCMLictPGHCj8oW/dHtZ/+HAMcJTUpfl3fXGyP73ctTV5xy
SMRexHMHUplD+m8/Z9Yd1FgpP8PdKYO2gMw8PKSd9dbpXH8icFhWiKmdOpjjiGMkb3NXzXNsWX+M
kqVNbvRoJQ7lzI8qzYbMlXGGBdjA37HkKPSxHZqxNdHz8DGZMhTF8q0Rykz5+2xVXpaEmEdd3zdB
AUTPRJkNt2Zrs6OJNdK12NbmtpshnT1x0o4UZ5wItbDMvjH9EkUN6l0o7ST7V3miyxS8tVEUWPtJ
FwA5yRzT3Mxrg2s4l8324qSEcLuwFR6igFFhdcX6DzZxePwV9lLoG3mIVGQTnK1yqFPNlxCQnKJ0
WON79F9uKirJvmu7Dfr3hf5Cv66wMsXykg3UuQ+lJUv1V0XhriC2e4MxPgqOSw0pLgrYg7TY+K+Y
R/mxglC2rjv4/pTcFEXsi/dmNKUeiJjnWKXd8BR+U1CtirsF98Fw8B+hZYXRV1Ih2tpLoiiy/w7M
21nyf1YzPW9+4hC2pV1YrSvtTH2kPQF15J2JADjsC9ZNmDxCPKT7GWUlhk/p51GMfoMGYKqBBiac
pgcS+G4uA7WoWwOcxRuNykA0uK8+DY6f0e71dzBbH6umIyTam7ZIU6Qq37Q1ctidpjq2A13TpqzI
SrVY7sF2diIsNXwLteyndmvddDM3GC7LxHilX+WLqvU0TgqyTp0B64dbED4JJAyxaPU5Ia2n2Hfp
CoUlRZmv1cSMrE3AM7n6Rcrf1c9HbDMgRO12r2X8MzT/fT/5mTrWbNwgdoZp489ivZcePP3R2Nc2
bDpxgzH6tKRjKKp+js4UOMzpWN/ZjKeBH94xeuWyLaLxbNOmO1vYdpWh23ulgJ+9UArXGBzsjYXR
HoRvApaAuZvdgD7Np1s3NVm5iDAwsY8Jt75yvJ8SDZhcOm7+zAMqMbVka2XGOYVms6f7d+MPZG3l
mpwCW0SRLli3dCN8EOfUbpkZ9SjunTgVJ+UDFH7xq0tn0rEANWUJjeiDPAaqO+4zIwV5gAFbhgGc
s65shPtAhZCQIYFcNwir8J23JVWklFtx4HKRqoiYw8uyP+XlWEkrBTl+PWZPjAwTIqXR/5VxlUmy
zYSXwEl0vFMG8Z0P3lpwdqG9ngqno80lTnnVZroeDjs9eNCjWDYj48JR097r4yss04ZX34F1Dciw
SeIliAtltWKrVZDq6pByKvIfVf7w/Ymlw/LCrYFsf6boI1CqZRQkNqPzzc1ymVt3l0JpHi+6RR4t
phMxhuAKmPWrxYbXM/wSPk4nXTI8wxz9h5vABJVpNUf1pxyCX3yv9AWe9WrygenYf8XLw1NyVPWX
cXvGIxNhv1IPC2+KwgmbJkCAMhqPqQWmM+ueZ8Sz/PUA7kgJs12imvN6EEj3xBt5OVki+Itwc/uc
noLnRCTd0YuVEAMW1+GXqJoReYQ3mPf+VuF+eOZxJqjxbkN07N6AlBcgkFJhTgnAvf4jB6lQr9dK
sIuIHTbV2ptrjlaI02yBQg2yreVrk4DL0Xp2nMG1e4UThjvvCc6uGnTRQyFYuIN60Gka+P3MA9Au
E1Wa01lqql2c50j6Ks4cAl3rYZ2YIcDpW+8NEFMxtQMGS4+ccTCzYOMnVNziwaaBKdmeVCZp3w1p
9Nyo2WtmzgNp4I03bi0RnvRPsDuy2FHG/Um6EL8Na9wmDoT0AOulbqHZQ6hYpH9AR/dZIDHI/oHW
fIYeRagJOHolMDEU7eXeSITzI0zzYqMti2EPlJYWIaUTFSKVnxzmM7cOcCwxzfgWxuF/kmBB1PIp
nt+sBrm/hBHHhgiWkKSWCwn3NidSKg+xbq3VelrPEzwlGX17OEPoaynzf4tUwnCplPXh0Lkb99q4
DQ1z1bnvEL0ENXZN6ag3ejjB0U4Uxt15C5iZJoBZm2qaNH9ZB1cdsCFsU3m/gfakYHBaquxHU1Du
q5rwwl8evAlka3H+h8mA5RXgJh+qV1krYOQngIyJybjtcVkn9nDXAMCIPmC52N2C+Vs2tBAViN1i
SvTfDXyhNnlz1kzMnFOtea4s0Dpsc94Ha7RAf3fqhC5Y7B89THIcnhuCd4ee/fiffIlktu1qGkvI
kTYgzSlbbrL7jlCl86HgHXpNrLpkUBUwNs9ySrmiPjd3veDcuEvoy0tRvJ10E8bt2LV1WgM4TLOr
5FGlitE7aEWUIySgu3MMm6QlCWr+ENOsb1THz+iLeWHmu9F436397Fl01bF6LvQhkSWGn2OyqXIn
8aJCfBkNPss4w2/0bAw06kjDnnlOD2NVNNbOmVFTEwbd5J/CLoOYxSDmyGI07tcJ1TyVSL+I0N1I
rR5I2RqBxGnY6JbhTlFHVJx51hz/bkfILk55mhGG7Y4+Eo9Y5gfbqJONcSjIRRTzkG1oau5rYJM5
iQiwFsikmH1br5V2hstZTP9jW3SdmaH2RzSRPpimkVv6PtWnSrgRyCg20aq3T03hR1SjAY8vc0+n
y8szlwNPu1QxWY7fwx1cPEvP3G0RrlWjjVrHQE62BgYiogBipT8vj8BeA5iKhkcAgsi4hyPm9Oqh
+EzFch8rX+LKFrNTiE2Z88dLRjAmZE9BNa+MY5sKm7v6VPu7c7cZow6U1yVgaYfDk9ijxP082gIv
WRwyUAFksBEVHa4DpE3OROrsvWn4sKkTezAv8mCzjJzZPsdbH6cGVGENpvo5G0wIl+5S/ilm8G7v
5cDxEmNNMcAuSBEmczOBTBnuaG+ti0N8/WGyHbCvj9jT4PoLH8R4AlhmmDb/WThgtZf7cP2IE5sx
5Pa/tpaiYBthQE6Ac7DNbBThBnW+xwUil5389JWq4hOFJB0mofGELw+x/WqZWdthsq1nWPfKDma8
YYfFSGoCdUHmVP9AwqTIdpCLE9s5wJpWQ7r//ZewgBrsSpzmYzygsdGlkFyfog34IZ9PO7x6mJ41
41bLoQGSUYhjrCR1nmJ8xa5zqU+ZIvjQ3eMy0CkUfmIn/b7BaSWnWMAaOia24UxXc9ORbVVfnwEK
IHyE+fJYFR2FBzTVEtiQIQIlzLoaBfJgkM4urw/66lLfTK/fWI2RPuuBWpndFDUO2Hur9K0HZJV6
4EcRTqsHZMtD2kZxSOJ45jaBUulCK3X51fjOaeK5TY2KJFu+nwnqHcB0Sr1kEidUa4jSzNCHIAZx
B+R8ahxBpnGQUXlgGgOJBxMenNnZZiwAcVik1D5yiweOPZ2Pe71ZKJDJxrxje1rjxJuQ9XywJbrV
6R/cWy6PKD1UuxGm5F4XUR02pPw/yLEJn0erqMFuJt3Z6FxAbx8+xv85pzhv5Sxny8zmgHrVKhHy
Yf/9J+2BzPK+kjW+DCjk0/TOUyYXL8kXdpfYMLPSOGUG+8hHKpBxFtAAfNyvqyN10VPlKFbGwQb8
XHoaICnRdLzvAbW8Yo1hk4IMDNzSXbgRz/ovUJWJoV2jPXgstfNfTNOgaHXV7AdyGNbyJEsSEYaX
kuyFxEpdMwtxPkJbQNSVWaLRKPg4Rvu6v/I5QmxZ7dDNIBkn3Z+M8XOUY6UxClyP5efiMZmJzfvj
iAHSbLlfaHC0eRMdPBpW7RFEsYv8iWQKcsmzv9VyzG3cJP0FKfP1Rcx0Z1T5HTHSXJYFu9tZnX6Z
VkIsxwlNiD1h0CQZowvy9pN6hX6J6ur33Bnart9ApBGc+agitJCSoF5mYgc2pJVNMuIu9WI+ho4B
I0dPQb78waFSV/ZN7p4mGpreDdYFFqd8PsRPzKRg4A2GMbVuHBOVY5CykudGzIgRJkvUbgRgnj2/
8sIAJqH2KlIqhVEGiSgAKrkWjsfR2lDNZQXR68LwxJgHiloYIvvn7F3qTTNSudFwvtjQIG+dY67h
Ws05glCEttd2sjU1YcNYVGDweqqeNTmwDxUInSJCq6ry+GaRJedV7z28d0iyAxpCW244ilWSNR3t
GpJyX+r/Gw42BIcmMf2pJRKK9znSYQMP9aBDk+wOqLDu1lmjLCAoV22GFZn2jr3Fo6wOHzaky+p1
9EwLJC4geN8Hm5RTUpY3zwlhXrE/Yg6/+gImdqvQbcqxhC6P39n4NBzafzylYekdTOSync/YZxG/
kOkY1y+JXHOynebttNHMUurQNhERVeeByRNI6hlPaWLCBcerWbhaWGOK8BGhxt97Xratm1NCbX1/
UBFaxqpY0vPcJ467rMihSS6Ua2tjPcdT7Qvp99lPZiqai1eGUKRrRcy3K7gioIArSKYWw0jLn1PT
O9Jp1zq7JZD6bkE5VHLfmUKZNVgOwS5u9RCJSWeAQ3hBiaM5SsPnbmd/7oPW6IWteN4+eIO5IHMR
XVlLMi2/DB4CwG485kLrWL2rymn6spetXK2sB0rxtJQzs4n5IzCc0JKzdw92ZNn7qiLSuKO1ErUF
4n8RUoiP4o0bxioCeSo4KKmMvW2z3tnRrBxU4arJE2m+DXlTgTYRo+Whnn1zbBvPfTm3AyiA8sja
VtaBQWQ2g2enmaVRqNl4XHUApcvqGOy7Hv2xQgnQhjnBt01AchaIoFlsM0EdCpHdqzkd2oIRZ6i9
ymZ8C3hNG85ITgP+q5PofQkL0uKRAfjn9cJMgqb/mTNadBkMZpynD1yW448PDEHAzUlX+RJe5Q70
uoY+fJzPuwMEwnksjaKHUSRVByuq0Ws9TN2EkBsPmX3xoJnyIdN2atZw/YQoJ27T0v5hHpyYbiZg
ypAYScHMtAZd6kY/Deygi6SXah0cyVIL3RkA6QbOTFtqJxDSOo/gH3JiBiK708mTKGNeEpS/Nhtp
H9qUhBT65KVW1gthlYutHGbVzTm5VO2SbHrgSvVazxDnV85zq0FD+8v/g0/ZfgV38Z4j73lKnu/U
XWD7j+GJaVuptsAfKGBeNCAsVjJ5KcHmjEGDbLhF+ng5y85peHVSKFbQTu/cKKhVhRi2S6qwA/9b
5524yFRsvEEYt8Eg8iezlTvE2laXPsKIx3dtv5HCM1CtTxS8yFYQzLqbvoSP41q18R4WDJY3QMWd
os1y/XMw0XhxTV29PCMPI7Q+DUIc405JlR7eOY7A7+/E+LOilPMe29SUsNf1ecUBjxN5eaRTtC+M
lrLQsWkfbf/3dvm4dwy6RjUJ9HrOPnk9GW1P0/F/5YV9M/1jR9mriy7k3MI7p0y0YVDY8IZfjB1b
19WIbzuqYCmEszJmQWm8MzVAbot/2XPioWp4wEoszkUTvrj2HTMniZ0bzg6QT987j3/TH32V914T
mE1m4VZ3J1VeGvygOthuJihzldyM3rPVoamO15zLwV/4jB3ZG/5CETmjqGrB1mzCII6ruOikzr4g
OK7+pzAo1JnmcXp9035h9Z/SJVq5mlmgYK8HM7+L2uoariDHpEcW3QmeTMialJVPPQJM+65JiMOu
YwG2gwUPySN7Z6f2wD03ts/Ahj7NHojIxhv1qsmw6FxALQ7KIcK36XOFL3CeQGljKMmX6imiCHyU
ElTbFOWPywAYlDRok94V5EF9dBfEk00raEAplsh9+iU8EUD4Yh8/4gMpx0PZ+i/qOMktu67jL0LO
rF6jJydK/lu6dgaLVMD34rTViFXwn8UJn0189t5QB0biesmqm6l9qt0Qeeu+/v5glbBo1vofjOi7
A7E/PiUdbzZcObNCFz4E12Hq7lZCjJaI5LZmYtMvTheEdddqfG1t5I/xhNMEZVjDAw0jJMFxkEbF
rZz9Gy3ciaLy0SAygBE06MbCtKlInF3dlq+Qm+ZXLWWHhtHopzvKKVhvYHw49XWp9cyOdGhtWtdJ
aNUK3aG93wlKqE3j9eGe0m41N+g7W3fY8Xwo/uCXQF7Hdf2uBp6N0CUe9UUEt8Z/U+q2Dzb9io0x
TNCt3bhnErBwgiw5Nogja14kHzMpI/GtWESwfcax7K8/+dmv2gjyF31/lLIPqCRl6eS/67t2uu47
z3DUXgfVp92v7H7P40nzSvvJ3IVhkQ6FtZ+jjkM+3tDDwupqkZOhAdtRlhc6RMH4FROYDSfGm6Ph
y4wh6fDAA/6Ire+rSZFqHPet9PFeoZCwd+tJAZ53sz07t5yK5panTPqlViYVG04LxdSXxGDPFKNz
poh6n4KkN7zgFyPk1u960jrG/aOy+bE85VHB1a0F+Iso1XopUk4cav6kfod6yaOor2cLwz9da5I8
CYP/TT2UE9fmHHtL45YnMn3LCxb9sHngeLjv+FQdKczm7LltULpoPr5QhkS36M6gVgP8m9cV3KNy
d8/YqrHvb9OOFvoWo0CwCF8hwXVCRQDgR8ixueY5v36Z3FRTuY71LQ09R6QmsW5fZGssWa5AA/aM
nc3SK8LZLm9L1BLEDfySrkBB65GXf+CmHAYSNAHDKoNQecq7nsFbVtOiYpLfgLOs39YPRBmdO5S8
cq4J0jdr1JQ/tXnESqClIMpDQ63hek6z85muQuHWUwEXx54zcpol3OsjiUV1COA4X0qSUbyUWSKq
erEpGz27ThetSOmIB4irHVXgxFJlIsBBLnn3W68DNIBCoJKprm15PlfHvC1QYV0ln1VMO/IETde2
WsYWar/0qrY0fwJi9JU9VWuLHCbjzLhKj3++A/TkApF5xIpBFNWqgmy8zGwZVvKaiCLf6l+fVd7t
SuKYA3QvM334XR8Nrz3n7bJ7PcP/9kPer5IlrRSP5T0JtHr5hZGtOEGfCaYmMzG0Uwa3Dwcf5Gem
67Oo1VQqk53NeMyBwPl5Fy495TSvDgrH2bJHZeHKsoxgXMicJA0Aihmu1i3Mlw+wrN5P/aQnRSd3
MjmhIJY/uEsCZxkqtKy3nwx1hK9VSEsPNXljgjw6rmVYAkwk06amtPaqiuW9PV0O/m+qIwkFZgoh
EXgr58HLIl9V5+ndNmPTh84Y7ecOALuI6s9PlDYVFMwmlI7MhJHgREMxKbSN8L2GI/7b6X69Phmo
iF/5mVJiGxnuDR1HlmfQYZfLJvCo4z7ZgQrQKno71Eaf+N69xCrAPx5tHrSHfvSHSYs6pCvDHWx0
hNskcniMiW8oQktnDpe8L246NatlqmLTTN0QQd80ClEJxikIdIxgYnSjwaJAV5wFehzpEQT+gMIN
Oxn0BNEdBRlYtmkwIQxxATZ+ddNRbXNboTqoLhAxxFlTvwqz37rRjFNGmVWJHWzkwJpdAX1yfkw7
ulz3TR/vH4LhasqX+TYmg1go6h24iW+iXc2qgDT+qfDfPkjXJnn+Gt1jIKTqAVEBMU5ywoIzjsUk
le1eJoPWQPWoAKprKb+gmIYMo2+3SD1wA9dTPZ4qBiESDdvXeHCl1vyOd7ibrjty+F6/jK5l0I1t
fWRYs+0sVYlD2syIDs5cT+07b92odRyJm6y0t0S8/t1qrCZUZ10QYLIJLadApwIDQztIs9HjbyFn
rrCQma7C9di0YUjVxsIXHA6GAU5/kxFoDD7S22y8Q+p8HwBdtqGuzv1bC/GtxnnrjJErxCnKAhLe
simUC7AkQcvzZ2m2Tsm994hFzc8WoKEj/JWLtye4Rq+5tJNnOrwL35oQ5RRpLajFvBC+VV3AAReq
px6JtxOfySqZIp4t1QHdS6RFxaWgpdQTCfarfMjbV64DCj6pdOkRGQ2bTHGnCLmd9ftt8HhUa+jE
cqBYrgp9UPxhfKqjh1XE5DJVcxLXOI2LLHa7LP0AczflALUlxPEb2XiymyeYuOiyvFeMsPDPnUT1
ZgZfG8RV6RS1SuK0McJrlffdlL25Q2KUq3n+H+c3mxivMrWzv4WTucl5ZEUNyAKQ4mjWJ4kMhg+t
1vkzuRrDYQx/I8Fte4Xf2lmPM0vwnxcJuBAQJA6/Mlv4j19yc0l6B1rW8PL+nUsONgFUfRJpEP2D
6ZAEIXUuUwFlv2vIxz2CiYG0jf/ISS60UAJ4PCst5tRPafGV4vKOqraFLAF10QOPAGa4jnFU8iqj
JXEVmT1SHgFCty4sMWPm0QdGQagTqQxbLAaFQmq0UqnZQbVFsEJ4UGMPHB4XPh8GBDKs7D7EVxOi
ojy8CANLWyG91/m/S1jU9DdU99Nconbcv2hcRy51R7ciw/8CyWSMvW0N6aVBPvGNpr9EdJEb7thi
ouWYvUMW3tMjTCXNRRz7Gyxm+3dOid4HZQmDTYzLyYAYkMpQgqrqDlNiwCYQ8O7kJobQuEyRJWJx
6HgT8BTBeYOtV1fCVASGLJn/tg0Obi9jW3OeD2d6E8bjnNbcGcfAIM7fjwRyvzk6iLLLxhXHqz0J
9ExU50lHNVr5Zu2o4lj1FG/gvWDyYzcij9+rQcmXX57bKVz8B4XgqSbUr7+CtxlqnC3Gi8X/y778
HGyaJtuTbH8LOaKM7JSCck40E8R2vKMa/2REv31zES5Pzmy5f37ITwPov2fVHg4IPqWVOyGXIGkb
1MrY63QTlLZF9XrQrfTRD/4y35b/Ii8vmmmojwFibqK9XQaIlIlrZOF2uObnd6ticDmmwdUz/Ark
KjtcBSJP7nemb02ZI4sZ9GpbeCXjI0s6BWa7LkJhybilc6LTd398bXH8QGM76E1LjNqYCm++KBfe
FG/LbeZQqHawDmfRth1f/zSHvqrK+ON/+FLyZmRCAr34mFIZgCLdBiL/iKiMzqH5o8VY9BGzgTjQ
UegEq3Lwg2AWEzpI3L3XMZrZz8bWoZ/E12TrWMPyCng7095H86o5Lh49wN5T1iUKnp+rV5tlirEc
tacdzaGhISIYiug16Bi3DJq7Tb4M36D+AmxZfXv3NnKDQMGpjEG0ZjAt8iRrWFrnTipjQn4x91NS
Sf+uG6w2xkNIOzUvy1QUmgM4FES+4mBxbJ+C+B7POz9O6zaIoW7Rfd69+IQ8G/CROkKtVhNV17OP
72voTXp48hSOZvSZmrnPyen/K/eeSJZuBH3jaKXJCNv/UTg1okRKGmTvKZ9AF8wR7zgwgw4X93N9
9z8O6LgKC0qVtSeYtbQhq4E/lYluNUDQhPrvq4yeFiG+YwL0BGIdTFmaBgp3q/HjVZQwivj95JPW
b9SiMvnQ4i754/kdDXJWudc9WN7oDm5BHufvoi6sgn76YLM0vz4ONMcCYRbMv/VvMF8F1fZdD/Ch
tgvW2iwGPWEA/6XAQgJOT2U3HumqIy8hs0UT6HOau+cflyEOmhz3Fr2fi+qgoiY94g6Lrx5sVbH0
i+St/ciuqq3k0m+ZjlxirgwqUlOT9UvprCp+NLpBD69YDKBCqkWMVpdEepOkbpkOpRXs4h83RNA9
QixRxIyShHHNDuxHEoiHgNzV8jbe+pzbu9ztZCEf06JcpNkllUuPw5JiPiBL837wbRZ1Oy/u5QZd
kvv1lsrgOVRYZj4aYu4M6J77snmScRzRAqaJgyyBOe/57Pnnz8+SDILAjg8s+ZCPFJzo54k0n1QT
v9MIGtiFXFpAzgOAPc+65xzYTelzo0fKcbmhadMOMhBFnNCbZXZQw2Et4qCJLG7JQPZNiNyNlJMv
FYRq7OfJVAVmercQWgBnx6OSKH7/6SSj0kYr20Q3qW1y3MKuFV9B+LtqSpkgc3bNsH5yrzCO8xps
bjOo9KssK6m+jWOHafFnpbK3IBXhoNMuOJFZFIDcMMUDPJ9yVjRiZefGg8hTFAZTn4Q9DNNn4g39
6fNIYS+OdTbYLOM56jkHlDmYakTsygKwlwngGDMHWHEn7hjhorbfNkdhoBVGxFKXXJY4MyXnNTPq
RIbH/efSz+JbD0fZduB8SFd9DR1GeiPUJLWksD6nD0sRZcdGoTNdo+WPW3xj1qlaywUDrjotchVy
CwEenjcMWvkPwaIS6a1M2CS9vcckD4sG5luhUyOoHgjO3orgoPqD/xdgTtqXfNCPuujCPlaWvYqx
wrvD2jxZH9roiCbdXgJatGK/vhA+v6ZtO0iOLKiqjY6Zz8w232Q4eR/NbiPGJILABiTdbFHE6WrB
GJt5w9aBmgypQgwpkTW8hAWTwR36pT360BGdG9jB34DQOKX4LzGEt+75wZdOsWO0GR44YXH+j2Pi
QW245kHHGMZzIo3ADdIIK+2wl/S06bM7IgbcUN7thiQkNFCfD7U67u3trxPMbQS5/Uu5+BOEuADQ
GfdKU7Q38FpX4ffGjsSji1CHS8sQEpBHpeRYaSBYEIuEQJ/eOV4Sek12LngKsexZ2GFPjY0uKid2
Vt5bi3fwxkZE5Erl36ubqWZ/Tg/ES9jgiejgy4/6eWDzM8GJB6BBUisJM7QsLzsczIQuu7mrTkOP
mxJofLWW8K1JiMlQb/oIHeN3EmMh+l3PGmP0/7NE3on4T4MkoONLh8iE8Z4RVEl34E3NXT5me5cG
z7e4wwlBkg93CBBK6MufTXH2wizUcWN4dcJChEBJUYrBKdD3wrANLOPlRnxf310CuRj9aiOPFwk8
SBqcl5VQgfMsH3ewA4Gw1yV8Ot27qN74jV3hKP8X0nDOywXkNmUFcRqitdQBOKI8Hy/HMvBq2UqG
h+BVTIU4QdIzXxnKfWhDPdsZG2nLOT9jkZQsAq11XLcinQvPvz6udxI3ps3K/pegGXVN+4GNLT5S
6WD9///GkCKnU5yk2J1k4Vi4G4fMhZ0zm/YuxPQ//CkBoEC/4OOYSFlKfMa1PKrI7loSz7H0XFA/
qgT1D+3eVq7aW8AhBXWTl5s2Q/GEZ8WartnDecWe6/YOz4lwZ8HdKqILaBSvXZSX/q0ssa1BsHA5
4GuSrH59iczsRkN43yhciPF8s8WgRq7cvyI8VUdZAJIi7Twb0k8Bez9BC0RAuxyXXf8/DJ1uXOQ6
p4r2Z9yfJxD0waulz9zHlJR5vAWZWTl7DrQyHvVTSQ7MJ8tpdrWxrfgI6rCX4YAwiIZlXEq5fFjI
GRiuPRz+iD00ruWAiruVSIdKIUSCiUyGPflGYIy7lPVibbkEiOFBhs30mir8aWyFtF9Tnq1P74wp
4nj7rF8gydkFwwUOvmk3mq39e+tedFAf+UOIRwSZp24AraCvAv9NzuOvMC8lK8Lt4hjBI0CXj4iN
WVlGSDaGILj8pr3WzcjCvQTIV7WwDHLrcKNTqHXcXxu01Tmzo5Aa+gW9VjDBq6fTzsYiTELWjaNG
W/xlWrzoInUmgaY9gTtUcSLJh1F0onOULxn4OjKzuNivn6Fx4CsbbNiXPDfq/ZYgW1lR1sUf5iMT
Qx7cCSSEp26qNSiqjISBC/cpy00X3x6EHMYDDRyAUKKRt20uxxaF7/fpK+g99lkUMLYOJ1J6e/pu
QWjXdpQC34XfwC4iALULLC3+G2XLrzgo/hYnI7WBVv3tjkU7wpoFjpY0QMmf46pAOSOVB6BHo4M1
gC+qPrROuZxXl4Pqg8owly5tcit0OGIqZfzGGOx2T17wnmspf8uCYvKsMcTak8x+Ws04a/sE3yhN
E9Z00vY8i66+a8oRyyDVUr4Kxxs3nog3/Oi48vSAC7okyL8kI0lbJl3n2cNyDLPmv145hDoOWgSh
iyZtJYwey8FI+PXKRkHi/priLHwvj4F0jMpHYhzhq+54RHbHed8OYw7WAvcdce36WnUfHkdFJ16H
YmSZkMOXKi7I08y7XFf8ZztQ6DJFHXRF2Xj+Gfgp9LL0NeiaBhg4U9k8nsISzYIYXokD+ktV1D3d
SMi2dkZzsHaaXo5rAPgWNY4U/cZOqHAFDTXYKzTxTSr8VPjmU9SBNWUEtYJCeLTT6GThbOCuLu+u
+sk93kqiRNnR0GS0gfCb99CC7fY0hQm4yvhNTLmQeBRAlJmV/yOqXP1o2dPEF9BlunGiCcTTsyc/
vPezPrF15q6s619Z/glnjybEcRjjd0YqULVlMg/2RzPGVdKXcskgn5XyUYtDkOycKx24rlCCckrs
v1rv+3jT0cdMuse+/Q/WHDTCvcGmn2C5icFttUYWJtCLhx+y0BowiRtoc4iF5heqQE7vUfDUCdBF
yJj1cmXCflwWZP/d+SuU0ZdfPVJLZplHq+ALEEM9hkciiFAQZhhweS3rpPtTuQcxQJ8Z9g4oUMg4
hnSFhtmNDpYmYqRjkaQPgO/z25421aakVH/X5DC9gDwxIJvTHWIrKVHxpqUD41CJxVmzhpn9hCfo
mYChdHBiTsE2Xt16/2/Lw4sE/CKuNXkhL8a4OxTYfUIyeDaXQW2Wta0xNg8qCwCwwW3290DTgnDM
8cEd79wILNX374Yra4L9oMorCXBNYo+904XGE7MJO+OsOmRvy0SkymgrxCrVDD9oPHv5BB8jdu7u
mMy1m63e0CObjz1Dm6wuFkrP4BpVjl3HUpj9+MNfx3ADJ9PS7yXCXmuHOv52mB8nL/wA1iCkbKSD
Fkr45PIBfeYu82pqH5ND7X3hyPugHhEKNpzQZoGutGTjZDj2qplG82M8AyAuYh+m0gkBOJRN0yYx
8Aulmcfs6PIRRlBmBZ2Us/lEYr2ehD40PnpWWucIRFJ7Uzekd7iDdFCZ3XAko4ee979ySArkLH/F
ym66ASCeqHQLFxXuubIr49eRVXSPPMe0w1+RCgKc8fXwbOqzlyqXBn+rllX8MZlfbECFraoUgXuk
axnAi6Zf7y8iiCxhZWaVPppzUguj0UijE9FKgBMXfIPFlnr9bOw8oU5VG8y3uBxSgic7uMvyC+j7
MzBK75q/vOKTFoynY6edALNr5kLfA/wsE/GzMjq9Iy54yySlcv1hOuynPFR1DfMXG/JrjacBa2W1
BdKDTq/I9olg+SUBjvFjvi4+mrUuc4L1iSehn+4Gya7GsxlDtGooX/+BXOXL9NS7ij7UYZpZJVmQ
x4YFkap14a1Dg19I3QGNquvz3Fi1VBEwQTFCcH8Y8FsSCfgrgrfhNUUN+QJ+jrJ7rNUq0TVHqZ7i
w9p+4rX8fzMJ08y7rauoZLWWMAJ2f9FUiLJ1cPyo3wPN6uZcK9p+u3thovWtU04VAh4RRCbI3Y7w
AQ4vJPSCg4O8iO0HhogPmn3pFlSgNItRfySufn1xUI9P7bYHNJxV2DqoelU2pG4p24iGxtgmzST7
FZhY6pyraD9XARViX9FTLXhVc8itkfM2oomoRoqrY/6LbV9rBPd5HG7obZvlsGFbBGAkX898iN5Q
pM6A6SSgD/1C5a5Q+dhQhkjQEZYNlxVfuWOa4U4H4gOZr/CSYRWwrnkVRmrjYu9VPS24XpZoS/sy
n33aee2fup4AqmdJPvFaLZaS5uTCuHH5TJUquX49nGeDZi4zDBPOD9OyO+xGUALKRA5mIoygGFC9
wUibq7wR3J0ZGqS4xOXu3hDQ50kc1yEuk3qnnar5VtkOAXUpEdlSheaC/71OaPAGk+wcqsflX1Xj
iQBPpV2LvNLttp1nMA4AefO0kO1T6ccUQkqhCttKXiwpq7S2W7fIL1MmfziWsXapNbiA+iVBuvHE
EMlUavpAp8MPlfB19MaEE41dcEFGIR4z3sXVW/yyQP4ibRSc6mHrnWgG75PIzOFRlO8RmpQ4iRNm
rmVitLSePvTaflRiLVW0jS/QfeHR1g4stAXNdFnJaCRlQB8zJl5mhhKetA8PW7fXxoYizaa48wIP
zNZ4NidrZMcutVW0YKrk6khOzcKXcP/I5JOBtCoKUQ2ANCOCM8mjI6xOO6j82c8MAZQp1ppRbHl7
R3u0IFI8mAC2fHbiyZZiGdGmps0Skn35uVQLNHTySaKcqbK13z0IHRUut3GbtfK39n6NlY4LCqrJ
HWJ0T4+kVV9ksPs9M8GdOZTN7SzsyRlu6S4okfoCeKqaUpBJpH0zAT0bMTlHphE/i0pk6cUFjdcP
73za5CIrBmCfkz73Pmvqku70jYzmEX9vIFk+0MJ7Z9nypTOle/XqEpn6aqnCcgjHWjeNP1rQfrg3
T9hjbCU1s5PC3yv5wLPBk4m/CPd3HMc423xMGYy+FpKlVcqzlPRfByq2GTmkgxViwDI4W/S1U3oD
Ir67a1P1fNC3frPD7JrNbxDGAnSJQlWJ4BNxKUxPvHfuNSHSKHR9WZeAug2S2IjrPNTy3pSW4w2p
7BRGcqgclGnNZqRSNuubeBIYjFktauUxKe9hrMpLfZDxxbzfaPWXoNaxo/wxBetZBODBuXnAxT9Z
C9pAj5b7kPdWtv7jLc3UXXU9XeEH9NP0Ntcvi+tYnqXVnelIxH0rGCzAzKr+k+G/qLLbwlqxzyyG
5xe6FelKT7oaMuH+i034VPXTkMnW3xI7BPqJRzhp6+H1tc1m4ugBgOJI6ncElhpIY4W6R7CsTAJ/
Twi6P+kcTIGNljoMpE5iBQaP32VJnHlMsvlYkKSydVQ/VwwjeV8vF8KxKPfKJk9M4h/Q0NKC2TGc
372s5DdhQMGtNwe8v2X0sJd3A4jpOv/5MM34jOVbWRQEQ8Po0KjdVzGXgZFJFnO4YQO4/Crdqfbm
Q1ZCPLe1jXHJ2b8bFAap52QA2ksTcwXqel8/Ixc+h5bm/LZCvFBFnR4MFgAV7yz+Dsc5AL6c5qyb
VIM0cvX4lGXgzX5YYdiyoG88scyGK+kP+O1YKqQaghyl7Ic48X5BERjnGUxB6VfQbZBoO+/wPhjf
EzaASSP0W1PAtVTRh861H4mhOzJwHISg8LTEiWFSrinvXKsvRDTNydVg76zHidCYi/0pYjiMoNGl
CqUB0bnq26NugItqvpPRYPJVBi3GPIwWLBVvfuGvu1T7ge5R/bfuibvwtaolgerkcqLIr8CLOa6E
GQVEH/XqXvSTl7oVnbcyfkn/fcNLKWh7KTh7eL0BztY8vT+QqN8SMHlbuaQPB4EIDw9SnnKdeEdi
FstIQDnZ8wIL6Ya5ofuOIDi65j1Ua3JY8UW8h6frGOmYTmmdhwNAhR3T4NmrVZ3Ac7TgQliIJN4J
huJn2ohehjzbFXUibOPrBM/3suTv9bxOo02ihp9B21yxpJtRulT5okB8S+iKMngPRv1GcY+W0e49
ELCSbcNkOG01LPkHSacFSw+BdmX79VUirvwiPIgctvYMZaDJ/PSz+Np5nBl4k97bU//EY9G4/c+9
TUs2063AVJWc9qFVPwPw/WqWua49UAsBNTJExnCUzE2T5ipEdfMFUTi5ftZ21Qdbh7WpkZ1V124h
Tz6zUDMezIYPizL7qnW+EjJuO6ZnmRjHWnfRydfJhffjdNB0VAMfVsaak+xQszWyro7rbxt1O24B
Y+CI+Z4hHamRxd5JeiAy1Kxfv6ALaVRnaBFkeb1L1/gwIlaNUWnEMIXQWF7VrRSr6xntZUhzGm8M
rqo3w4B21syUAFbdwuwHSpcbcH7XYCWW6fcJTLpRLvg5Hawdps1pABkW5tJ1GGk2TIUPznzK4FDG
l4sLkXLye1qNcVIPVyiin1mdhRuiBlSkdkfk9zWSYsEG06s4/NxEQ2WAGKg94Y57f7vm5eTeiQB4
xJ8E48P71aDlNuCDmTRZOIOCY6ZnY39eiSMY/pIRVKkIVBCFPcr4YHhv645NCvmtAwBR1x2/GUFK
kKkGQpXskVm3EFB6JSG9XXMUC+neggWxc9sxoByeIrP8Nk7oTvMsTSrjS9IxB+bAqd/e0MHc/H6c
QYKk+ut+xJlljIt0IZbYpWzcJ89h5acB6ls+9mUwO8XjyttSKX4MeeiPvhGk2u0r8RUv58OLcou9
0ojPtlAaJ2HU0p5kBVqd+bfAWhCOjcvYRf/QblXbqWS9oAA30Z2XwP0ryFZfNShl3Y4SgelwfBOi
jt/GtLUJUBIfE8F4/esM36XUCpDf67mLI9r/U0yu5MTwAzdwjItrkwL9stjr0KuGG45S1mK3amI8
ExXznw8zlOwU439ZKHKreX2jFYvUlkTKl/HqhxM7cggW1antI8AWXFhgmNCnjlcB5Sf0dJ8/O4Cj
wu+/oLqlLNQLO6A26NJvCIp4alokKDrJwhenqUNNXUQIrZ+Nof/vfe1iwNFI3XWeCio9TEbceQWB
bbg0aTGDKrLZAPAqB92NrX2sxomofzaX5otaETlz58mRi7AvMlb2SEuguV1oV7SwSFKWjVKsxlv8
4UAKL0f1xcYQuSgUzpNr/MbrQdCYQdyD6KVov23bcWgnZBx5wAGJetRlkgUrSmaUnML+2o14QtLT
8lUEfJTGV+hwApt2pbRQTGSf7EGDAKqJPb3YubDMNzGjLAfSS1ZK2jnsolzjFjThAnWQ1FfOV4Xt
alk+OQGIci4MD244L9oyG9YAuqmcHrDgDqYUUUzKnzGwxZhXCmKjpGrxYzvRkOv1KRw6DxxjAeP5
8B1IbikhFK3XJRuE2An4fZBL7q4jhk57K/NGQ3uy5DkTr3SIT7S28br4D3X9E8nlcEf1OAC1DC2O
399Q6WmsleO8opRxSy9BH0OByYccrNxQGW6oFuFy3+S7/hBHQ3LUHfxmPepBOpFTuMbBepZRMyER
3q1BJ2fS1DIk8Zjpk4KuWrK342Y5Ky9YjwGWgHODayQ5z6h7qXwzlI/FcJiksGsieHGhEMKMWZmZ
tacKOiNSul+1MwIbVdoQzuDUDcY54+50JXee2q/vxnOg/44yZ6LbKlXwj+OrAkV47zpHCynW33pT
9w1sclyQz1v9/F2vdU5qq0acjXWbMmqputB1sNMcu6eO+uVANKUEAmE2PyX4vTADjQPvLZepClKU
X6hjqsAtKkNw2UNEFe3hJDbehCPolnXzzzTOhH9Zz7otZVg5fExXuV0/T/i1aVZGNEAqLpiotiln
JLzqtvN+dtUKUfUHkU9H4qJwWTjtc1eDOdcN35T6VlObsyhty55HuA63nQBN1CB5mumGixIB1Ikg
zYfnfZideILLeoUfN8i3FnRD7GKFauWysNxUJG+7avjIUki8z5fDE/JZPfEA/VIEM3m0QaKqimSR
6aoGqTOr2Ly5Mt/lLQ5xhf3KqHMqgsTE2oUzSEPnpuC3xOn4PqzhxAHgUtSB3/WrO2MdtwctclqD
WNb17TW1Kk2KzONuDZAc34MU++TffxNOppwxPkl57OqbWpftHETJmdX8U/UzU0uG/1zWSTil2nsg
vNFoG/5xw+DsiBBEQgCvDiG3CBoxFyYkyuHgf9anlKEnTqVLB1pR4k3atWbzha+V0UZFBpckbWWI
vohiFpu9fgN5jAaVj52IJPVXdvzueVGxqGpqCsEij+JEXpcytvwahZUt2A9hjZkLQofOYPA+91Yl
NtTsZDM+4JazyNWKOk14WVKEIVMevOG4Qcz/WQTAffMLfa4iDrc5rjMAAUPmt+nlvdjJ7fWAZq2k
kTTa078xa8BTZ+hTwtjb02gAdwt7Icradi2h63khRCapMO71gdq1zq1e4brvFQR95GTEcUD44W+t
FRxOCGEB4yEVGnIpO7MCSuvswK7PqB0KENyRnk5Ye2XPdrX8LeLxzHf+uQlsr958MEnoOkPNRbOv
nKNdYj92qKOQTQU7bBrElq+s50QJDfxQ2CmofUUTsylb0zbUPH2SK6lIDgRJDc96nJGxnic/UET5
vwMnEm4jtHozCBxnCTmhi2DUHr/SfwX06yH68+M74Lq7OzRo1or4+RAYStp89hdsoYbnJVyaghO4
9iNmGxZ0pnbb3eGTk2NZJu+/CjoaGa1b4Xya5aeFv64V+jVdtkz1g7F2LOtSxfDqaEOpgZY2WjYx
QcKI2urhIEURqXwxNNBBM0lec81eyLLZp15VwWHWBpXY+jdF+n8nU1tjXX1vi/hGkUpUzJyWsaZf
6JaT5ITNkPQNsmt4qISMRKoW5e0NwpTiiBFbbaImQSUc324j8zX5ZBcTKU2vbYxedPsBWk4u/qNe
0horpfZfITxHHujZiip1dGO3vq7PxfwWXqFXIyaKOPdVdJxFNEgAcE07L31aSQNxmolWsqjjryfV
EOMiVHmtmJW+kZtbTz2CBPzGjZkvuEpKsxxyRN6MFydpTL811vtn9V/Q+Pi+ZmGH5GT+02ZDOfLP
0iHzeNO/kQXAcK0IFlMR+Yuhg1i8YwCDav2y4dgcnSz9AtzdOpvutCF6QOO1hMKene3uTZK0c2BC
kJkL4QjAS+LCtC0k/+vOQAfUxkUSlWOts4aqwIK2tUWbWzded16MzMXphesT1vJQkfvc4d5EQBrB
kmsKD2kMKFPYlnzfuMNmaLmuiM1kMxGGogJvxM1LGM33xNha+NYSAdmjJ9Ls17XqeA9Kxe0sMTl4
nROzLFq+KXyZYdtSz3shGPThRCU215jvqS7FaOZkbNOqt4XJzQAYujH/07oVuUnoCLmfp0AGg4CS
kv/tUH2vX8/GlSvR694BWdJNenA6TY6HfdfKM87tTkcRUb/fhyiYlErEK0i1elH4nX3E51wAIa0T
M0btlvfQK8hm1WW0mytLVNxjugV6M/zZAhKoaYZ64dqCu5GQE6DRU0CjBSqdUlYGr6vqPiWW3IR2
5mUogQJr+t8t5NtY47OuJWFQWxQesMFaXZEWgJHfZ5wiUtNDGAT8RS+qoLr90ZVyltZS7hcU9D/2
0S9RZLlRp0ngY90zJxQ77jxY7WFRGjrC/dordMJnu/3kh3QHMPQadPGXDZ6Y3Fn97u13+NV5EhCv
JH+r7QS1PWG90xmA2ZE5/WL2tOPUyZvbLInyVgIl3/S6I1e65XsjMe5YHgbc4uVb+J7Kpc4mgGDp
/qF19yehuVBZjzO4qq2RTBF4pG7weOpEcQJ8xLijYnKo/NVzBSGLd0fqan9k/QBW8WnWU5xu95Qx
KG5ZRacVnb3fE80DiyiBk6WhXjGMHExlr2LZnPHEn1RgvSpAO51Pv/AtUZ7BY7O/Ji/KkCQeEhn4
nRoI0upngE2+m4uN6TskJQmi+2m7/UF3kS1ByZbrSBFv8ijP2oxLhgA17ug2HdZ1dhti2umept2z
PnEyhI+FBoJ4+A+n2KJ6nmUmmwOf1n9HSztgCPA5pgybdf33Q7uO9dDtBqp2WCM38+8cOWEsPa4k
Rwu36SRHQYabAEaus2GsfqvYqL51pk6piiJvDQjyat2jqdikZEioWfYitewr+P+wuXFjSf4w4VN5
RwCR7NORTBW9StaCtmVis3Fcn/cmD8QolPmCNEyJFl52VcYFw3lDtILlCsaOAS+fW433W/41ggst
M9dGxOx+xoe54bbeVv1P1cculK4KzjvDGc+teKkVZOcnNrtkMm70pBlVtH394ttyyWbW0KM/kGa3
/4ougDG0lzDG9qLdRrPUwl4EzcH4uIOAIpT4u7UZe3kVpA3RdG4qZe5n40exLaPfjMEpxdOapvJC
V1f03g4FretjEeMsAuUUst+N3DVpq4qurmr8GogeWXkboC3cP2lU9ikcbOhcO/DZ/6QhBNd4xcA8
x4ZcQq6JVNbtw+xfPmrW20uXN1aAGy+8QC2UljbVORlBTJYuMS47Qrbwaoe7ioIeTV6qqW9kjn8v
9gnUbMiL3HSF2Kv2/wyPQX8N53tha7TlCkSms9W2vqKiQNWshZ6AMGAN74anzeLLXX2zC4Si7P2Z
3fh6KZTF7foE+I9WkB7hXtoo7/S5yLxH2+xa66t0vuuc2BSfHymAT5ijjisdFD+NVIcEPc+wikFl
WBkVnVVMv/g+793YW+Fa/xuaQ/kIOhEj8VEPyxjwDqwHBLNDViNind+MJ3vto939qyE363HmQnOb
29gmEgkvNzRVLTq279kzRUO8+Z8TkJuaAwoguega5lyJs37WaE66xauUOjNmmBZQTCEk0rOpyU23
DnUlHIRUB9+KVL3wKzNcPykd9zqP7f/W/bL5A/rBsoQtkWU6oSABqZn8q9vfo22v428RRWvwxsQA
Vygc7B5XHTKLe7uhu/IcgVgziinzEhSCMKEv7vqzMZdK6S5u109Z0+3ps06DQfKm25UDCYv7tA8D
ErW3Ft3NIY1itcmLG0l2W8uu+5RsMipBpeB/bqnw+TfcxZjpHXDNMaxqlsWk21dsVOu6xSEVHPtQ
eJfiPzjfs6VMBBvuW11QqZiKYel8qDs3ADcYl8l1R5njjEtV3XIrTtXlfxEt+z8nogQF8cNgLREe
49L2zoXpfRmfmeQg8Ulmry2BG+qNI2QUEJeUNelrbj6sberOt/t1j/JX7LB75Aj6CFwXFhZvYoRA
XZOjldWgz55PdLnRfMbxfQCNWf84nd2NAQXBgTdsD1jrf3LFaEiwPjmJs8fI0k3umAJdV1ip4rR+
tCDid4cdxcCv3nbzh8I0wU4QpZ0CegD9+LKSsTV6zLXsOkTasbyZ4UqLotqmZLVa/0uAkXkjSXPc
/IBASv1Q0BecUDwFGNnyAyAkjGdXrWhYfDUqAdS1kUv+q7DE2ir1jyGzDGXm2fkdi6WHxp1olX3b
dFlaseJ6TyEp3OTQPIMppYCAaHfIS/JlIowBExkRAc8F9XaNjyK2nlZO/hjo512idNA0RnXopd9w
F4tFtpn4Gs3xpz+T2qynAljWT24/o2qguRGEXE+T7F2ZlGXPjXGtbRO2Ah0bwsd2vyopBGeY2gCl
67qBh5CxiSsiCG2QRF03+hS6y4/ox6uPlMs6/dFez1Hmf3TMh7GPpmxSrvmmC0vl9EU+xHQ/Qezd
5B45H2zzgFlan91b4WJvf9ks1MViKg6sr/EWu4BxrBIKpAUMWoRDSKQEQfFUnDJeuz4NmgizS63L
67vy7kItfUbdTAZfNd/0vskDOKhkx63HuAUNkgcRim8x0VpzPofD50Zj96o2QTwyzV/LLxttnpHv
bgH69WkdIF1Vkjk7EIT8pdm69C0dF2E6EPr9SeFtFdHRmd0YVn+i9h2F2d2K8r9630+wmgWyx4t+
ufa6OqJnumt7MOvZ/3Alo26kKZkH16kmA2zsy6AE8jVzI2Pp1M0vy+zu7camm+KX7i1u5BqC8Qtb
g/rf70UtHBu/G5W8aIe022LsC0vD23d+FZTJC6Fh6RX8C9GNvEaMoLhyuj2zasJc6Oie3DsLBHM/
geuWFJL0H9OrNvgzEL09wJhjvfi1L+L1WwWEZ1W7KX5/q/HBG1PNp9ZSiXuhEBZdNM/+dRvn0iUu
Mzhk1yeMs8vmjhOe+XqONhIF8JXzTK2LaW8nupb4PB9oyjI42x336Nej7t8wUQlJipB02vankHWI
ecTwP9BP22TjB4bMOIIU0NwIz5tsKPICkxz3TQ4ANEKmwHvjnZUyQ0NovPupGA/+HDrsitXHXlyy
xAaVXCtXOBhksDIjPJTII5gXQPozPyyQe6urtaWECQHw+sYSanx/SgpJU7SwwBs0TMCe1IEsDYC6
+S/PU7dvjy4cPwHWbB+3StagDrRZr3Olr3GPmkb1y9jHGvVPsCfA3U7f9892PRDCVHditm+FsvrU
HXBDdsfy8GxTYQXucc1OaQoGmMvvYgBJzI36e+QsSVtuMVnZEwDKlzA1QxN8rdboDbV2ePTNqxWv
0vc8eQvCJdmdE+AvW6x/HebGZIojR+T0U2jAYTFhgrOy+lKcjM/EDBVwlAEf7xtLRsIBj/v97grV
pQfVe8xKzFh0GAUSpe1OdLvMy9tMeYupVIPJMQfzpQux/66MRCRQqqvN1ntuej5OdPR6eB5AvWkC
etxU8Cq8BYTQ7SYxlBQDw6Xzhdf6MxrPvOVMTCsXgzAs6genjJmPr30ebwSrTx5WfsL7ggVHQJrv
o3ZBfQoMs8OorO7ZFdcEYXrX5Mke6Y010L5NYRLtqoeaZCqL4rn56hwU3HgN2MQ+Z04wdwyMlDxx
hTl28pYEU9im4V8Nzh+cwtDAnUoQbBfeK3MsvahbjTxoxea4s7MsyO38OtNvZc62TA6slDW8ZEUa
he+D8uR9COtTjh1BegKCcrD9OXWfAY7XcNj3p1mwCzGhih04ew0fyYqDQ+4n9EDXbe2/dHTimwA7
pOVw2R265bXK8UEqCOoFB39VWc5s3vMa0nUMpEZiVYGcGyMK86GkMBtIzoHYIi4g7brA92twIYee
WiebLImA+83OAjfvAnyQTv+WyrQPRtpX8xPizJcCL1rDPegghinIwcVBJ08QrekRdaWcvdrvLjZf
fmvqvRxiF7M5Gs4qem0Wchasj1nDZsthmrWeMtsXueA7/zcfwu12n3/O9QOPWD06AgXiK4I0ijEO
ZkFJGISXMy49HsR4Iuov8/SV9Jinyj02eojZ3Zb3YDurTbrI6vEgy35c2h2LVybOdGVTPFRyxBXK
3X1uFEJwSxc4gG/DkRQanfrXoweyvwZGWJO6ugcUTijv9UfcOO4I0aS2gQw9s5/DXcKCRFW77T43
lRxIjHs2NGGN9DmvHu5S0RG+haYOiAwlrplg7kRad19k/5OP3vslYjvnR/x+5IMDcK4aJklsNAsn
nfikZA9UWSCDK5+wHp+mMOWwqYLjfC1URH6QhARlybadE0gfPpJnUWdjGLz5XR+6MWSyB+iS5Sbg
nOdEVeG6tDJ/32EdE/dzyKqQbB/2Pw1QfmQYwN/xLgvsba8M5HwGQDjgW4iiS6uUOSIVBfk2Fpdf
deOwAKp/dSFxoL47mAn7DcPkuOZYZ5uHWP5O8arLgI0WswYZKAjwGbCOe7axuYn3xn+RAIDjRL9x
OcPb6d0ieVqMTtVzIjgcG9dydH3d0TJJPIDD8U5oUjCdKbpwa93dOqyR7gzkNZqSfSp+TGtedWnU
hVV3EHLlQdAUJRahpYda2bB+APDJMgrQs3CrpKxoqXekxHy/1tRMffbQnoAeEaWCNC6zHaCzpTBI
bZ0GdRWzThw2jDL+58/xIBNv9X+1j65bupXnZOzxPOjOdMew2tZsseTQxbnpqvhYXTazzAOhA2My
CpjLPiEHVUHMgjJeroGb8XfVsNe9zoUDwVay7CyZienXULaYnJt9wa7BiLd8aO42zAkplBAxBSf/
AA5YI5kuf1qf1uD2Ff2Z40ZoB5aA+MGn/feKwinm3tqozmCDU7ItqGrdMWN/bGNA/vRgJPPVA454
i1nJslKnz+0TfeX3HsgGD7gUnT2z+fth+S5Jb6pIHYEX3MpGOkELu03hDEUWCTcOFzJDD0HLg+zu
8cvI9jI4rhM7OKn1IpixdLw3caKw1smCgwjxetdP58hqYjJW+avNO8DRiPKsi1hPnyPrIbWFFOG+
N07qY4xml5UGANnUZOSlIbE5uU///X2u3GG2FLua7JpYZRXSvWnhUWa8amOjcPvXNdIF7wfOMxfz
gBdqdoF/EQGkmdzvliTy3N1YA/NejXXeL3y+6dictUd46OlwvFgM9AxdAYZByTOaYRswST5TPfJH
WULIRO4CnD9lhXELV4z52AgT29WH4yXe+WIeVwL48w9QBiyphfa0W6VSW9JBGq+5+zubHdfxkXqg
bCELnXP7nUtTBP9SvHaK7VX7LeMyjBoJuAuLBMC6M7722PRiA+MtwazUrSbLSKhz0jbMBPApLChn
dSOAD/O0omtjwEmHjMjNsR+6gNGbvpXl5Xoh9p7iaud1T9A784FFqs38GLWoy5bY2c5hTBCQEsgv
tmcPC2mQ8Bs/aHthSmIVCQhDaxB2HM7uOqS1AOan5+V2cAz2vafcrUhUmWbogFXtmaGNsMflupBs
2kX/M+fit1iUcrR/XnuECYpqFjbXlvVr1ctM0zTd+vD498ABOyXjMFhdf+hkl1lZYgOBilk5R9nd
wbz+PlIr/VSBQ+B3xNjv9oEqbjW8y7zEJPnY8/Xh2+C802E+Y601d0xyf+kPUHBVLSo8V/U0CUDc
b2jHktymafbtgwJzLomZdXP4hUC4YTP6d/rvOoO5tojQZKEAo06EN28o4i1iEJXbuFvsMddGay9w
R8yD8UWzQuHQGKG1/okJAB2wQj8zF6OkCy9eFPwA1avNNEJrG/fJJL8WtOVNT2xM81V/zSA0WkhH
XYpC8P4Fb/vGzI3von9je7jsm4suQrdOWeAu1qmkeIUR9klmuQHQFePTe+ZfdlTNYXzUgzB8zlf1
H15fIXeJAVzZScuzeZtbKAf4/KZPczavVi/n/jZTjOHuluNeB599ukbOearxVaAIgHN3SUkuEzbr
5qVeHUXc4lChQj7RVGnudWRKhU96H8GMAFTebW6knK6vwzAncS78PHmtDZTO+IjkiZN4nPbAPk+h
siqdJbV7cW2pAVQH2rfW6B2+4BS916Gtd0WvEmd4o4WjsfWC1s99XQnowuicz+F3zBBKcsPoqSxn
BwtBej81feZutmRmJT9jwLPn1CIJIoyvO8hxHr0uyKHNkiur04pScU6xyFLMGegMh0k5o6HVQJqq
EJUU9XlY5s/6l/I/86PTfYm5WN6X+mGVG6LHx9rNvR2BD6q3dgL9eWWEgg/0r+STHr7l9qI79fST
OW4bbSgx6dTZbL15R3Tz6dcQqPe5kUKosOeuE9+vWawl5Cn7cqQrtY0rdblG5kQFfSuhULQxsuBE
tcUfIyyICzviDTP1/tYtBVBnPdGfBBd7FGLbHeLyufJUD1wRwhFUyUPAwWSGdMO0mSzIPmDxIqME
aqmbv+cGqZmUj0S3ahLb81Q8hoNL/PH8ICS6NmXCC87JiDLC+QQJPSC3driiJeJ+WmxY5Ke8Zj6z
5PlH897jE1QD6N5yrQyAsuH4U5ts/z/lJ9lkJXdAhFYYUMa1Nd6JCwj0txqLfCaYg+ZSAwgL+f9T
kD7P6NHiNbLACgvoUm1DV9xxYlLQY7D+xNcHCSFhNGj1qdx/5tRwW4bPxAJVKSAAS/hFe+eytKbq
DPjS3kfMHpKGonWRenda+KGYyMF0EtjnUsh66EHWD2+ZRQRYbFe1zDjS9Qiy5fNPhnFMtpHae1T0
w4jGAgbN+XgXVCSJ/i8vyqBqpD/UvoQKTMFxsQ/w9IF3owNTtwSmgkqh3szv6edUXNles1vHwqS3
fpVAG//FKn9x67uJB0Iu2cD4tJwJmxvj4SfpMHiPFdvmTCy3+LuZAClYNBXncDPE2A9eb77nt0BL
fina/nUz15HxHzI/GVgCSv3nWWfQoGmt1oEv6Qlsh+EF5uyNeFuEgNFcXBDb3gRAEcXVS6WThykp
R4uxvn2WadTe7H4dswutiicarAhIZZ0nrBhuU/W4viOF+niAJlqS4XzWiSBeQaRJqGxRfPxgI7DM
9oa1iTTfwwvyK9G8KLuKvn+5XQOREWcjUUVcJrhbOEn2xLqo/TRhrH10wHzNvFcM11FF6xoKCtPk
eSqSP+TLpnO7kQj34SY4nOu0VnIGx6DetuYiDqllUGpVSGDC94pB63tJTAfy09vGGZ8V1UwaRAA+
3ONV0r2SMrScveLiDBbneGBKXjerFwreXjMfykMlaf9lhss/tR7BpeDZYH6G1ic13CJ0srlXKLe4
IwJy/ruQULe/KF7zH4ni62RF33+/2YbEy1zI1Msf9YqN/WhbiScljhy0xlFRSJCHh0iFYXrzfrkI
Ma37MG8pkVik+dOQXsZW7zhowsWwjmX1v7my4YX0Nzc8U3BxIPla+8EAqB3lbdJYLPyttHJAhuZ1
PDM+cNjsAdfl87Zhh7/gjbunu2lxXR98cnnhkALenDG4ZxzItjZYjBa0OZKhdRE+zBKweHQ7egGy
ds5yAZeDQE2OwlHCvS3OSSDFpPWR5IwB1bVLLMui/otkHj31rfyCbgKXIJQ8U6Modf+xcnlyowyC
O2FJjkQEZ0g2VUn1dCG1hg698iQYZVIldiOoVN2DZDE7ZYaYpROuergHqbjLnL1cH3BcKCUG4nDc
waf9yLtGhfMr5K/um6hKgMhqTo/ENDGN+zodFkaesgsay0TMIkss95i5fi8VLoCuu0f7SFAhtNuv
zbuJjjK+01eobnFUytRvlVk2JSQsnLbXXUp9GM+9imRCNYLlKmkh9eRtpXymKNXhLsDPrfkllLjU
1bJ/DDqWZJ3kVPqiKrAD/9bD4eeIhGlTBSD+iR2FGS+SJQ3aXe+Jvn7KDfVnxuYsrU8r1tvYFaTy
IN2GSv5iRoKuiciaCv0UvLPVa2je+T4VgpwccLiFtqNLXc/YM8Kg70NUtP9+A4Tj8OQl2ZM1Irwm
Sk/uOjZjjIExPDPPCOPOUtHHPFUf1IIOiJVaBG7dEPdsa2lbqhKAOwLTUTY0nqf1u4Najg2L9oVX
KZaAOSkJoYtf65EVfJsZGoz7GehnJqfJGIks6xnfW2NzTbWJcsq2g01KIsFKHHO8vjPLQSCKyOs0
t8nc/moPB3YehkHeMSwSvF3LDKTnC44t7NwQX++Sj3MEP2fbPYRonUIZL0CIMP3I8hPr1lTMji/Y
2AHxrwZFQ8XMbU9hhWYBBPkEhQnHpkDMMV8NiR/wO3rcYVZ8qvI+gxfTsDJofLUZoWVcFsVGATDB
pMu/Dm0hQXhl/DVvvfabfGqdOZaOypqDMEWfxkHv1P7ILKHfel2HawkZgaVVeSu9RGyK7GmOR+6s
WF67AB7PxdeIKYVzODq3tM203WfjJctTZsjcokFcXof8hJ3F+k6k/kEZ/k1oPBDYGV3dCYGdf5OL
7K+IqxiffAx6wJy7KuBRfzGL0yVyXM5CsRoE1aSY0pyS4LWEYhgKdqZhdC0CdZHQHKY96LuEMMCn
u64+2OVRPOlukXWRgY5N5T5T8m2FVat2zJHOMmN1eJVdSj2KE+A7WmloaaZdWlmTvW/BdtaSTDMJ
KeOzITW+GLNyMM3MyuD+dCfrVKQUGIkOcnvKyOkx3ObwUAKVGvHCDzjn+e4oJ3S/KPWJoc/LcMt8
i+AL9dvKmL95Qb/kYlF7nwOlQx27lfym/KjQSuWG10o/4m7zdrsjzRd/KqpdeXgbZYd0bOH2/AUq
cE7czafsr0TT5r79OxuPuFP9VtqnhLZWKIjPIN6YZJmM2a7wgyXw3Itrl0ZT+cjzwfi8msE+poaF
rrWy04s1xj/GqVvGwoYV5jxNg6XL91/vy9phAHM33UTup1STIFuOug7eGADkg3lnCG71i3ciXHlf
5ZVtqonmL0TFKdR2+ymu9EbZGrsknGn8TmmPab5KqJvOKyXAmStCUiyxY1LzfE9wYjU/3Ghl95jn
BKKFPcxH3OiB3fXtTVKc4mfQEWDaDuwqMHk3Y+Mt1ATRP2ZzVcwoMBBoft4dI7sOWheeAV9TFnOd
ib0i6KQILHP2wvNKwF228BzmWUk7+zJKIJE0gVPrqxAT1foVgo2nKe+HYD5rNLrxoOCwjZydiwzO
EZ9fBxZv7Ji/AbfAeVJJh95XHqCGsG96d/oR5N0s++s8Xa0H8oMjWgHtFBsPk+Z7T1yOIhpzStu+
A3q7LwoYo/deZfJEJ7BtwIh8QoR3GG7ZH+p4peCCKvO1XrdNEdPPSIdpIw0MAE3cHTD/FsdmNkZ4
E/lNmGUtUmOZSSh8polVHSmQPB/YT/6LZa7uhqvIddmOOmyCulgs85w9ygIJ2FxhaK/74DC8UNrI
cOE6Pz9CfhfAxMsR7T8J/5pq1BxqZd1FYNzNyNUIcOEMbZURolisEnuqOz0azn/JuLaGElZePRUx
jNh5NQEpsuBovPD0TPalVXYajFx2vg9upM0PTXPEblBy5ygXI43JLrbZbYMst4iIombmHhidiBrY
buFpFzJSkRfWdxRHPEz0yLqDQNxMQLFH0VFwkvXud4d6iGEQDzIMGnM8d3G8o0JiP3IT9Tziabde
pzfzFpZ7pQKTBNSDEOx/QCrZ4cSIJaNV7VeOnN4AwqBQmxkz0DuaBUb5+gzW9i8jFBA3/Wda1Kpm
dYPbnLO4dn/r5q7I67cZgGQ1jcr6Eu4aB1RI5eo0oUGj4HAmd/0o7rEhza81JIntRy20iOvq1ryJ
XX7mT9ORsZJoyCW1RU8/AqxJxM3guO9hvSQgI0SaSNu4S+l3CTRWldHw2oWP/KgKebwms2ZQ/hFQ
kQx7iIoorDMX/ASVULP40reoWZpszK2PF1W1m+KDQIS2yuKZCU6eGijhufto1tsTOTL3lCwDIuP+
d4itShHAzuHT8xTBoestxeGRqjKIrpHEqOeWednYCbaW4nEmdRRkUeXniK7hgZ6xj/j/kHp6da8N
F5T1o3UYwMQfXwqishu9sRWTzlchxFjsn+mnvZ1GUxqmNJ6TWzQv9LSsHnW5LAzpY345Pkj2RDSz
Z5hx0Hnp2wPAIpreixPV2iVJlNXT04zomyoE+fhm2ZerACsAyzsiB+Pa70KpqpBgKjst9+h7wuK+
IJK5bLckGmBYZKQnK87omnCztWs9qeORF/1b7QnNFsBDZ8OmWj0/Hz7IXeSjfGN1JMKCMbMk0aJ+
T2E33cCqyD9j0hvq9EgID3rMSuYtv38QVOa6w5rJd0+iazO0hSvr9dDFOwgUaKCG7xs4C/31EeCS
bCIpghTpGPbUWyA5qWH0dO69ZYbU2ZwjPoE4pCtc/1B9PrVqUXKePFzaOcuMeWB1bfGc1nW6PkZq
7yms/VHTXoFUQZin/tFCMeXj5ue/i9ZwaahNGqvY/XzP74iCpJWvnILyrpPMbhvNnpXlzAHbF5Gj
kl8XZ25iQ/99kocya6759heFrMPt/dsJ7w/CODoq2lCDy0Mfhs4NolPPfWDIjyDgH7LM8SEdqCq6
ztUw3y/aSr/5W3PUVD3bztNJTWuVCv64Hwp5NI97eRS5VEczZWen43yrjq4z1smQloj0PKT2VfUx
LC0hQ3gqTBUA2bodBHbc6B4LBjTRHxgtvtoE+kP65ap3GY3uvDSUPI0dfDhWXjcg3NqKnixCAshj
0YliIsTW2+iQlqnWIeYFHJIZy46U38IQIWlFLRcAxsaSyW3GOTQGqaHFC56SNy9AMqfowyF9FDun
czkzQYygThsslKv0WU6BYR8StFMRaxciYvYfGACMRfGmUiPlDIiq92eyL/maEXspTO4OxBZWMty7
02UXmylM1dS6RNRytYXrg8txqHyRI87EABi/fUwgCK2ko8smMYLPXk8TjuAPqIwKNA0KxYG72EHY
mdnaj4hoJo47flxLc5HbCroeRjk0W8jd+snti/9sOAjdHcMTiq9EuNqklxKaA9X+kwC81w3Z6C+o
TVouz6SkbRb8L/WzPNeNBKe4BKBvRKDXKnPxV29LKM9Vnwihe3aKfWCAqxHBBuQclV4qqKQOH7XC
5DlAmM4krz0YcVb0vf9ovWXDXcFsdGclv1L6/xCCeUBy7xUUSMqMTB2vaZNgEYlP8VUOCwlwKwPa
j1Kh+gKt8d2cayhYzC1XQunr5cBh4lkk4Ytakh7AvTz3XJ4YuGS6pl+aLWtw9vNUkzICrb8BGlCN
l/b87p4dVyFFwxQU9VA82BnIRo7/k/rEGyTJiM15O/VwVXp3+zZdBVP//OPZBGBUYylBLL2orKrW
PpKs/N3wnrPy0+D4JX0RFn+4S+/jtPX8Jas7ZQ3ZvRA+EgLFrgkuuGyt9uJxto6bjlj4OrjMAwIK
9PndftZICr+4VolrC8aVbdpLj7P8d6+elOSejbynSfAGu8/KATRGrnHJVDYQ9RbBoXQ4kBcDVM/+
DGr22bjnvtvz48zqdaea6Y7g6Zl/MNXwA2XLJQtYxkASe2mw/Wsly3ECCFMJptmTozRVJGYIlpaP
UQyzxkDZXXXXwrgORsalu1kVoIXa5XdPkvj/61mHjq01OJImqRblFKYPGW+r/VY4xBmc7aknMk7a
EFJZfsaZb1U1GWs0DLl8D6Qv5tFprSBq8KEZokd7vh9dckqGYzQMYYNGox8gKuJP9GM2NVnIRZ5y
WZsCrlVw1wYFss8mIygwjN1BXgRgwUcT3cWdJXWKXqTCgh4LYfOSestJCHIgSv6kPNHP3UrFmPhd
PsrlTIqFl27ApHHMvglAW8UwBIGqpDoqv/wkhFV9HjVJ5nB/U7DB2XSQo7E7ZaRmZHFyzo4D8gg5
59hZiGroSJh2P0sa1mUhY3904o8R+/HSR7R9GeQakJ7q/A4/hfjWJIcxF0l+bSKRiNyBtMnYckiz
iNfY95VfgPaMvVGb8Wh0d5nVQt4oj+pnx8DAoq6Fw4tChawM5ARk7Pr0x6ZYwMo7Bt5kMrNzBYHX
0xJ2sVPiZ7CiTVkjXniU+7muHqRIzMeDjWoE5KVgI/nu5zOevcTuh6gP35aFjqiVK0X4+HjGXwZl
+ne9mrpTNM9RJGc6512XUHpsjBbOIv+MnQ9pWWo5fXYcsUS9y8hKWXYxQICcGJiO7JRxWQSLQzQw
ZrtjZOLDjxZrNMKBqYxTzqOFe4HVANqSDo022Z1Uh6t30xTll0hnAQYERczht3DSAdWHaj4Ld6+Z
L1LgzmyNmAtiKjIr1yqiU8BXuwIVUTZdCo0bJtsG+pcpSbAsaJ71NFzt0BECrd6HPluxSQ7TmuG4
X5ZpR08dolAPQQJBPwuszUmcn2nafdsxVoeUDM2mCAjF2zalHFgghd5t1gwTHzFUPVjdN7Ef2bdW
J5amo8ItuEhEEs81hhJkp1Q32zV/yvscQ7QP/bsA2JsEBml+MbLmzGEB+YWj/9LHtdAPVNW44ApQ
nqzFrJHPs5jgX2qNDXuzfSaGdZRLoWvJZK6zXxEZ0+1cMp2+GlDm0sh8FbBjXFqnLjhd8fdRORvo
8l4zay1ap6ol6Bc5jJwmo5idvk3myzbbliacxijGe6VoEy//fdajq+XICy5pCoZ+GBIRRJdKik87
AOACPvYYosKre0SbMz/oHt/WMRodON8M6wxJNqe0Sc5HlcZogGUuwrbslboTslSSdv6Xc6aVD/lS
zo5toHxJeVHUaTjIFv6pEXFvvTmPIJfiUIu7BF7vz0tjvGkeO5btpc1Ntus1zIWeBfj+AYMPeaQl
NPhp5Xnr+fD/PivgxSBI+EBTiRypUlJYRIukpRMKicYINGJ4j35nkRfSq/S5ND1uhUmnp+18Mnfn
B1vPdwNiRZeVZ7SCFnLYdZHBhp5nOIHypKF/WC7Ajt6lzWHc8vk9dkfHLaY29q8tQOvZ9jgqYkJz
+bdRPtMDg8z9h8zHSFYllKw8kV8TgF+6dVrTtqkMZZbTiXPKht+XLpkHKX7hoDLCclSy7+qZy7Sd
vwLQ3LlDb6HKMJ0YS7ao1+hS9CZvl3zrHQ7xtEyw8sXpX77CMtWg11iME/toe/TwJD0JxEZcBGtA
NPZOJc2cuRzgikjrlcGp+U1xqp6dbEbkn2rrngsrkQklWF6HF6im2HfjRhWOCcrzRZo2sv6m8ReW
yLKxwhV/s4nc4KHHmT33VcJp9xWfHp9OK6l9HauNBITuUZoEFhIqPM95++Pnbdzx2YepZKVxDUvl
4xnNnVZwZnae6B+uvC2DEHF7GnYOqxZYDlRNBNgvvyUXkXgSrvVUouzatagkS66j9bt/Goj5ZM4l
Nfi9QL8XMEPEPzwitPXJ2/1nrU2oFtRbnU0nh5hQJdGbw1tGr7nHj3AEKn6IJW6DApOuJ37FbbTJ
DLRvBXbkT5qk+Cn0xJfxPrVRgz6C6fVR9sSVX9rQcSGsTyXW03Xz7cvxkz+p/++y0lqvWJF4y6gR
lUubJL+4PJCtBD8NpY5RlkHFoR2x1unS1Jmc3pWO5qoPFLDNJrZu1VN1bnSkWnAWLwhZrmaZOGCn
PJHxojH6GmpyTi+fgf9uUW/4SQERl7bPqoms2JU6T+NqQDGJtnWfHIxUrb7fEpqIP+PkTIGtoCdQ
WVNp2Aiwranh8wypHH710lJYvG0sR28U7tL4pwhRkd10eQ+bOqQZ/NntPGua2P6deabCmOzpGaTO
7RhwF5aK6aXWYSfMkPbNyUL2bQav3W51fKny3O+kDRBEfFIUpYhlaW1W8kcBZBjR7AePQNQrVO8C
7rk8DDAwIG3Mhb62L5XCjStHjjx5/nJ6PUN0MeepH6oUyr6aLvBm49EmgRISwVSCPg9F35cD4Dju
K5jo8exaeP8RukDl7PNxWU7pZDEger4oB7zPZS5MzYDaNuIN1dqh1MIWqa/mpaWmP8WfA1QNGrUX
GrOq1kZBfR720q2NVV8E3D8Stv9lJFDyOx4m/Lx3Rwk+qa/KaMVqxGjIioPJbdnnxXCkkre521+2
TJGHBe9mb5uJqn/lf6iw6AivroO1PxOpvdsYrmAhMcJdGIxnUNHawe0ThP5hJPW4xiE08LJbZkCU
j5rM/wEfNVs0JXdpvtjd+GVaETq/oYjVCrVeq0btxzgibCZnp7Ge32O7e4KJ9aGT1Kqx4esPLwBl
KmFQbR65xlBdmnCFzY7zfMbRYK8oKrefmuNZf8vZMpya0pbyvS3QnW7Wdg3ReSSgZXKePEi+tBlT
nsse48yFLuftiOMEkkzk5haH/McuAvPS2jNlnbpb3E9IuTDPOcJBNk+CC9MOyC1DvQniamlJXl5E
fI68fb0gAbbY15a+83GcWdA8dLm57TCe+fGw+/PBQg3rBKPGgbcH/+jQcgLl91VqJQRi/u1CwNJL
wmqOnhdRFchyrcH9iJVCnt+cSnzi+FeM2AJggsWa9VaBYrLMdmhtmmxEkVdzCSOPHwN9qIM81GM9
smJrwFaaqQPG/DXN8HbyKNQKrTFECm5dHBttWuo9QYvSCo/3R9XetlRaAhnhSpS2GvjMReQGY8J1
LsjOnVdsAv5aqfuhQfKIB/9hxCuN+QhTc8F6E2KN1h3ZmIugLNlFJalJRy2ffrdjAMCm18IvFgIB
BXIy0d0pB7mL6z2zYLsf0FaZ1Nq/LHqinh1+Qjzupf5zXoyGAw+SVGN0ePAf/3pkuqsq4QJQ6wy8
87BfIbD5EGv1sI3sPXj5VC9LNLgQ/jbGAVUuL6kkh4YOCsstTMyjA42xVAaySmC0NWOFVIP1TK61
/Ndm4RywJvHhW+lhaEbXm7gxP+ASIuqu4HntIhO1VPQbLPU+TXjJfMCIejkqe+7uSiB/WLgD/HJ6
TZ/k5dEr0RSxLUOf0z8VgRj68pd4RNlBkUGlBZft3PaJsJ2U6DJcqao1po2vh+GdF44IWB4V7qly
hVoyGAHduKtdB694zAlOopjHaZi00jRRTZs1AuKvkG/it56ZnFihuLQ7nU2TdCB98LAztfbj/wq1
eDw0inBuzjRtmA4UtCenyLUcjqwRV2+0Y5Yfd9/ZS7gCRH3VOwntxLZHRLXJQBl7y9XY9OO7GqLD
qT8/ec7jK9d88VpNYF8R5T132svgVaQxCLR3APvndp6jZbYm8WOuwG6/8JaxK1VB1nkDWquJkOkv
yN66LyEiD9d7Ijo/u7kn6CRZAUWI9ZyZWxbIxRWeU02pHUfCXzGqJ5wP07VM9WzzwJhZd+oFKJ2+
4+YYVSUDGytD8iWCbwktmILIxjcfaWl5GC1c689ploNqRCvRRQT7KZf4VidneI+wHj0shFFTG1Wj
8VMh932s6Rm8BvGZzXHZpiBgmEUcGgCmrkkge1nR0z7tG7sOnkM4kPwhYfzApjvYHYbmaubJcGCz
/sUZDayEHq8kPErF2kndGIVXXGMpFWv/yvt1vwjZRMiAmVttI6wUW9Z/pmtmjCc9pdMDfdzQt9dU
J3RzGp43oLJo9vIPXq0RsUXj8kXli4/FWduuDW94TE+FHmAm5n15J2rZBroRlGRE5OeBJ+/u0o+9
hCs7JujyKUQ3yDyqfgdo+GQkOFW7E0LaPDWkpsVufJlnPF1qBBtmY7yiem+C73AvqP5/2yAw4uRL
ZlJVaqo4miV/DnK1CRJCtozWUuyVbfgfgJE1M3jHasxvIOJRBCBVTHmdRmlPf9F5OaOeZK1lw1zs
JpwHWUoLmp1SnzLjEzTPdIER0AybLBF7WQUFVAVfQFM1SiC0tIi0w2cTjL8Z8jyauL3AHq12x9ws
UKp0l6e3BS3syJ3SXE5GADiwDIdEFF2OYWH2EbWMTR7qtzRjmR5VYVJkeD0JO8ZAx4DGwNQHG9cb
RlEfwo34i7Gvv5JKiEmYnWr8WCR7E9jx7qnaAO5jbgFkHIKgK7mSW3t9jiTt64ZnGlUMm86igf60
3TpITTtOoM9Nz9XudSrFT98dlLQGZu28ZE9aPfV5AurNy20wpHsrNAqwa3R8Sz3tR6NMcx08zub7
mO5nXK1YB0gutiv37+eX9Pf/YhGVnsz3s4j3I3gC3dD/yE+iIWDLcvLLfz73e5eHJOu/XtZ8+dyS
5KiyC7hfmR6pPj5i2W0+Bi/zXpLZb3JAgYUV93soxnovSmn6SZEcx7wGIOow2sgaruDDMCdCMf+U
J9kx29h7W1A1lhdV3t7K07U5r4gck11f2lEeVUOpzfGj362Cpe9rm4YyZ7AMBZBLycK/6w3WCqTR
MJXoiPNaMFL0RYHXWVonIQMlOVvcKwKQ2bp6MW0/OXvJgI3KlRgSNihfheMF00XE8TQgIkwBuMVE
RmfV3ykPU4Z+7dbeoVEc7Ug2E81U7TjS49VXim2gJKEvFQgKxfgPyy++ukLjIwShoQ6x1+UMh/rK
ioaMAu8d8f7ScnoA0Jde9xbY7y44Q+4z0lXTR+EBxBvkrlWjHCTdh334vOdNkw5saYFx8OwhJWmN
X+X6yHkPH7O+lEJg9i/h680x3BHgTtgUEnxB0Kj7uIOJgtkdVTumWlMCwlTpfQqRm8r9iBY1D6Om
y8lhs6Nbzs+kO5qiefCDYAs/OMI42fDOcKHNBr603OxzGPLfwkM09rD+0u23YEvJAciXXdHw0eAo
CrVsTxHH99V/jXH+5dvFi0kJo7OXpzqlW13BIaPUPJjJ8wk1CT2hQnMrDRB98dCJT2nnsvjqaDU2
V9R9PydjcGbA1nmtIW3CmYOc7ljtA76KM3JlsPdSs6grYDlkW/SuFSxL9qMcTrCVoXVx6/EQ3odt
sxyIv9mpLXrDuzdfQAW0A9Lev3y/n3lwbAJPzD2MYjHUcQ9wzD4jagSITrGOqKpx/J/VTJ7NKwIL
0j60XYNYOEcbZIJbZtBITLELBe8Fc2PTuMJNoNIItiIVaqSZ2m1A51gMBnJ/ThKLl1k/2mm7m6dl
KKP24q0ZZa5JrAuIWkjMR/fSud8rVU0oxDJZgNP15WNnctiYoCCnICP53iY1tHfAEHm9yUWcsaSL
xL2NOG9MqWJXf1xyIyukf8ZtxduYlVyxjBZL7M/XoiqkWiRLiXZNCIQYV9Kc5Iu35S2LI8wX3UyO
ahoVVv4nUVO1deRb6Z+HDSgMx94DZk8Lq79N3ObIY2OGkk7+S1Wz3xydCIKVgHCPyAhBPqBqmHgA
/e4wBaAlvfXFxkclP/18I/Z/kKL9cxO7BBN8ZiWYa4ai5jhxvDkW937uvSv4EyGcEPmv3L2pkjIb
62V7QbdOQytboUt5SMEnb+5tkilf8tKBwnLdDPxJdQEQ1VJ73+5dus510ZI7nIM5aG/9wHOgLoTg
1yJAC1YBF+atUaic5OUCy4H2L4DffcDm55fCGqMrKbTPwHI7nBp7it/nr591OmBCY6IJFWZwR+Ua
ZDIaawbyJLD/PxfQ+rLv+ICw5+wrpx9S3h87Ap/XXMN/fUhggEvhaz7QmMEtpDwNinKP/s85Qktl
j/LP1bafKzkqMuRBxmCfExQPY+k4kckTMbXpXib/QbRB1Xf6M7HAzUjmbRp2joiJILMTWYZd9NBE
h4BNCqRGJZNwfMkx02rwEkasb2YjQcQ7N69hYsRzVUNc2ypGE989ndyUd8lAsZ4pp6jRXvINYbJn
5bc5LaH7S96lJljvR+PAxE/sd6UBuOuzdIGUXaG91Yiu66FPgs9flc1aWbk6a5GMgJ/wpcfc99zJ
w+Zb15ONl9t676dMG6w3SG+BtNJCWUC+fdDfPAXpFnJc0fNLi150muoLXSYImly0f3Kv6pccaVsL
Z7cPN4wG3DKSrn1ZsCx49HOegoT+kzWGjvcCRVTETpRF8rGY7Wm5kkUXa6gC8tr0Vp508/vbrDzF
nzN5fP5Mp6iv3VVdX34B1TAh59zorPJZozZA+qAIdoBIsxzWqmTlgMMnArQ/s0/yf6d3ToZ3LeiF
bMRkcy+QHbi+sLh6MRU7CR+0z+jpfFHifgDOFtf5AZ3wpDgPP0iLrqJEtt0RGnAo8PmNNEsMHsOF
mTQIl9ClDhVMI9TdGAi+htNIf8l9Hh+jKDJVSpwdTZhz1ZaWa+5d3FME7By9GUCNJivCZM9OOMYU
n7j5nvwH9rYrnlmhdY2TXtZ2W3vW5JZUmWiuPzk4cllxXLbVZ4IpoBoyR0fbtuXNA57IVK8PGtt4
m/AagF/RZIYjsfpzQkSs+2R04J926NkgmpF4ASaPljJZyQe6W+OJSWN4b9B05r4J9zObmpB2XA+8
Lcloc/NVIhej4zlrw8vDd+C9UZmpR5WlStqoNcwAqAdLzhFEZcRxhQGFx4hI9WyUtVigBZNiO69M
NsMrCDrDxpSsJFw6uYXSsAPO5WqBK0iCw49e+bezVblOrzVOM8wkXKLk3hOgjhDOIsdRMCwDZPiH
0fqRqtb2dhea/rtf56Ocfis5CWSUL/F9DFFSSPPkWMpaXuevnj7F/1aQR3LzMVibXttO9znfBx4M
1T/IHZmnmK3jzrmTl0CApzudvY+1OlALCNiCPANeh2cOYjQyauWciJvVe94+kvsLi5BBgHFedFrj
DcQuvHzLNtk6SCMvjlFYa0abmEhM6xtesJfw4wS2W8PjbszHIjxFbjeGLuUaNqGblyTDEUjPwpRS
ciWTD82zJVYX8GDWk+AATexSSq1g04AW1q6kpb+OB7ZNybUbEqFEO5o5Pw6a//WnAfJxMN48sSU+
13E8lGL3K4L0lkRjuIhsLsoCSWnO8/DYBKJ2yW4J5VHoX59ZYMo1LG+AwBNTrLozhPl84m7VIx9Z
t/XsPQAyeO3ZxTaojSTi1/A0PcE9PKUblh0jW3C0CFlQymHVaSdVh15qgLLIPaPmyS59QosUfkJ/
CA9yh/JUPi1alfCduLtlXNNIPvrfrDX4VsXycUMmeo0f3q3SFGKw4rDaLc8Dz+4BCPUkAJ3s4em/
paXaOQTtuRnNlA6h710VcimECQZl2qpuFEdrHFX975vY4lY2tBVjaA5/jnEtw5LEV85Cmo71pM12
3rFhCcziI06KDUJtPkUfED7GiyDUOkTCl1hUX8V62TEVurevfhNFXb0YMzUPolezcL/UBEcIhvOA
aC6WqBZ1cpLTGZdOfVVg7t5/FGFDTdVUWWJmgilUoaiA0/4wT2EN8KCJ1EKIoU4zhI+8tv9QPku7
U34ap92i+7DgvtQRlql7Vxjl4mK/K02ngfbYT3JsorCoKti8YgADMtqPsMzbsSagozhV9XCy48as
54gkJBEqAFj7hp/RNgHpttBt17YVWJnfez/IpJxYY8sufund5asQLpFY3p3ospiilayzj+ERK22P
+R61q3BiWWUo+Kl/xYAe/0OFGOdXR6mw4rXMG+SDqz7hmYrlS2iHFGQbSpln3v0FPB7NmBxNaLGb
0Lq36ry//Xs0hMVScRVip3X2583xDcDYLv+3Umttb+SmOwCybBFL0HSyoF85hnVtRS1ygoeaeBh7
XhpRh1FQuf9ftnLlFQbPeawn2/o8FzvkfndamQR9RBP0obEnT1bvhvYfTTfxjmL5CSxij249mKbL
z0SKEzBhGsE6hXJO70zjaJuTYYjvh1Nn481omqSrAjGri3FmwNd0scBb5qFUOctzmMMRp4Q1au1W
AXfJKAWVzPptCJhpmvsRnJSqtG9HINQpMb/ODE8oLEiDF+1VCuM5GgcYDaKDChTSlCLxSOoEMwRI
W2U+QB/q0uv6j2dvuiPFyqP1OQTdQAJxy45n/hIQUN3aDKQ+f8QR7W6Rjf0DtX2CJ0sH3amKAyHQ
G8ioisqblyL/szX57i+hqIM5ZKUHh8J7sRJ4LcpvSRhniZP8MT8HazgjXVD9338nwwmB4E4XsY5n
e80eu+bsf5Hzdj/Nt46YLjmWYpUF6UP6VQrbP+MrZWjwUaz1+pcfGMs6hDgX3onuIB9Fck04mEMd
mPb2+e1mgL+x4neh1HyyRZO6XE6VdkqRUvWWObhELgsAZvx6DlxBtzCbxN7jcfLPnC5gG+DEGHId
fiUGY4IPSEMEoEhQ+SEWAcQjNtPpF3zAuxTqSoEgJF2zP5J9NDtG2fgWg4AZ4cVQra1UDv0Y9nuW
/Lkry2R5NzRCX7WEzHzd6qRihPg1iKZLZopT2shPMu6LC4Q0Rx7JXiGgdwcRnyiyzZpsnVgbKmYX
uYSa6tOEH5JfHNhcOsgjn8EK9SDFOVLhD8rSw4+nK6Zh+rFxa0ueuHuD6OwPw+v5YU2eh2cJLvnj
zejux2atW+5v4i0Q1hGL8r2WVNFSfXMC6vlA339k0I1O3x/ouFMEjF4lzMsUNKI0X+zle300pNNi
nGGRG/YDFLTvHhPU3kMywtKXULgsYnT2bgfXanf/KJ+I9yw+buvRDe4I0WWytLx3cnpYyIPSjDxF
0WaTaLMzi/txUeuLsdZYuzCBI0FBu0lfC/xptiBnkE9gvmnO/hLIo8GFMWA1CLtdCL5orWbp8ScA
SmsHTyhgPfp8hGgnliTPqRronGKtRL9RPAQynBXSMaKcpn0DGDRwCEsKfly2kRW6KWK4v3O71XdX
wH6v4GdbKUA7LvtMY5MvkTTfcEwI+QXPGmskB+JW9Av42OUV9tLmZnPrSPjpkLnYOoCnorawPohk
9SWBpQ/5oelmaV8fhCoXJrBnz47pkhyPmVqfo5+BUHQrmzsN5BvESws4gmt0AfdpWTj93MkL972V
SrRoIindGVERnWyTqNggBSCAq0soUXbG+pIDwy/tCB8fQ6s7+7IPxcgvymlOHNg4xb8B45PTEams
mpA+Ozgn46735q7cFtmQM/IIBBurI7I4V4N2MWm173+tYWTS+BY3cM4yqx/07+sMVMGueftEFOTz
7TOHhPLeQhSrM7EmW/VIhXhjpzRkbjIic7xFaKryku8OZ18PYw3MqsFLh8Xb7mPtchCCIOYcaBv+
9IxZi5RLJjH29vj1qXKbJytR4DBDuWKzVQRrVPRVlxSq4stt5tLxOrpVVm2fQENlYcdSF8zIgwQ7
MtMn6SPFWMZnq5xHCXjiaVyqKFu9hjmQlMSsQA575kLemb01xvVBf3/hZm5ztjjQUdC9cFHEj0h+
3Zm+9cFGojMhZXlh9CCgwTTs8YBJjQAlaQUMpV5B8vVBCchJtnuPLn5a65+4mEcvPI1f8iPHUm+X
TzNT68fEjw+/sH8o4pmPTDEIAa09dQLb0TJePbeFYYjj4yhq8/nHd1NkaJv8DNZy4Hidbc2HtqbF
vs7JqiSLVObww+ZMmODyba+I0ESGDeo+2NMmjrq4+1AflxLgc29Ckw8irfrxjODYzvYjS9KmB072
Wr0stq5Igf+ofqv6ucQ4cdU5ADl3PiuS3+utkPCcyHw7vwmJg5pdSWzi4oJlnduIHmwO6Y5ap6zL
+29h1TRsnL/FIq/Ozey4WF7oealwC6N/sWR/LUUh61g5xfsifDZ4C8WbRr8O5yAcjjwqXykcSssq
c0NtlrP4m5K/XL++1MeYnEtMigRPdf1M/efro94rb7XoMUQ7HGbIraUSUYFPBGmLR5n9ifs4drqt
7f+nKXkMNbmC8i0oUWmqz5UKWBt2ch11Y5rnyZ/ZrUhnT24ylNZu1W5y3g8ExOXc7Ab/8uFZINqM
17hHFQUJed35Bmpkj6kdkHtwOtDAdGbPHV4SguBYFpEw9DS2oe5pZS1Reroh6NgGNxvqvU2mkgIO
AR1VfBywpSxEc2MgLIWpNgVkUJt4Ct9esrFpwt5CQaVKaeFVlF2sBnvZkQYrSK+uvT45peCSfmkX
ZexnqTcvtt+XMFWVnOF7JXlB5nL5uhqNOF8cYvpoiBgNdJx5sK6qBsc81IsuDit7XuDeK5d2OvZc
08QA5RcW3Vv8vHYOgVr2nX4lIRfpqlz04M42EoQ4xGq7ro0n/0Y8ysXxBKJ4i3rpyjo4wt15bhEG
iSLhvNz4iMG5ujxBrylVSj82yCncsT2AWQmmNEVunXmpX978ZPiQnMw6PlXViHG3iEgiByl5QMM+
v3R/HvW2q6IYjdl1wmCRC/fO5FRT92dFrC9GYKX/gvjVdly0nj5TQarxqD8zJygKLj9/lRRCF0Nz
zFTc3sW3uH5Zsuq+bldrElCKu4UsG6zjOjXnuB0DY91niVgnqMm4BYOinj7Hqfh8idjmL9pX715J
BiQFrx92AiiDpX3Zwu2iLTkUdBdg9+GathVpLf9XqMQQ90V3pfa+x/pt8rO75P1xuJOBQ+5bQR/t
AsoYn43oZj3Ha4a82pK4///6Y5R9/Degfb1WmAoRMZNieKTcaZfxmQ/n/9oDIYoUxN3Nm81liE40
gQ1I3gBVGsqzEevGapi7RjabDOVhKs4Xb0FynzDHopNcYZ+SZMlyeme+dpzNYyyc9/nWwOXgAVh/
7I+AKEQkwdYJ4DGO5pVyij7Rhc1pMlJKhLdGLr36pJqFwunUOmLI+F+jVTk6T8in1AfqoIgRQyvE
O3ufsyLI00S6x15SBBOZ1ztlJduuLsMWCLiSHGTMW2aMe34yPPzj9y07LU6sPx/csO4Wcuu3Dp3C
DR6nNikLiTBrEPXYPX8XudDWNd/t4OCmksetqS0jXYl5NF8YdVfOoYg6eZpweEVc9wS8UagINQZC
HU10rldPyHE+xVHJ2Ug5d/cNWivqMPNlT+dg/4WnU++mfXdKYsYKxp83Wol2AIdTgQG5TVXTcaku
aw6zPDMt0F6FuCLYB49/VsleU4At/bliBSUuT2EYwI2FT4WCDZZkLZyX7WoGT86WcykBQtRXFBPf
lxvuMiO25t0ffqc4zH7ZSa6wYBZoSGLg2SVsIxO8X8YKTKSKMeiWrJLtU1ayVfStJEAIZe1sjuJt
4RjhzUngv0UlsGzJ+kLrMRFYtwqHYyn+hzz6fm++C9CJWlL9uV4pW9HKjXFE2OxUOPkQQD+MNaGv
vCmBwXvYU5pzLWP5l0o441+YHsdzTHSJOGc+sfIvDJVadQ5tJAz3v5OcH4Jn5Pc12f7CYiQDe/BX
otqhCQIrlrK9fZy9BYw++a5QuzUq25mlI/7TT5GwSg1BY1LEA4WUrBXX8qT4lr7gnwP9zIs90iJX
pQ4vVJR6qrAliV96GWWiDGMhHEbQRXkvcXOrzU68TRp2aMPgJpEuj+KSh9uua+gHz9EcCLjXRVRe
RfyWQasMtHioBWpYl7PEGDsJf0cLoFQ0CU8WBdjUbOnHKB6tinFFyzLSwNWwmXFBCuxcEn2TF6wO
Vp2f/NLa6PMN3I/zX2/ph/Vi99GXbQQoFnm1bT8u8N5MuoK+iTOPgJaxTmVA1xeZKYuERO66g99k
DJBnvRmnJTuI1y/w1dXOPtltOYEk7wU/cj9kc6aqdlOvB2WGSz4DawF85muCRTVon5HRedxi56KF
2P+7D5i3kSiJ5XLb0/2deUfhQw3V+R67rWg6sSE9TQ2a3wp43SvbYeubrH+5IW/DgxLqMHoZ3ZyW
nx1n4jBR7kgwJGkuua4FPtE0sE78ay34OMr5z4kN0W+lFtiYailmEumWbDb/wxuK4EWyn/MXky0y
e469YyUWbRpbynEss2RjUFlOKx37sPZTd8uFAnlwgQ+yOHu7d9pt+veiQL2CBVzozsyTzn2ZNOhv
BYvlkuDQ93GG+zVWG4AOulTVDl0f8VLJQZiaUCwLcKOqTemRx4HkyAQFS1kRR5VdF+YvhEN+5YDy
wEqd7yIyXQ2XepHn9LDEp8CcgNEhYhh7gsOZRAuoXtqAO8jsDj9f/iPMiUWxdhXbuXpwjkeNzUha
hrGHSiB1Yld2keid+x1KjVQ0qgzfDgGikyjtA4KxKcg/WVNkj1ex8idwCGLNsUKaGETXI6+D5xEf
Tc6V6LhyW7hba/CmWl+dEvzhcaPVD4tywkoxirKMdujjl+r3TsQJn50WC/gpa66UI1JSqXFFUJlR
RrtLTgl2iOl++VqpjPwmAzmN6AbylEuIXed0SOK5oPIacNBdFyn/FJwUF/6uV+r/jBqg/orKOU3K
fRgxzcr94yEMAI1noqXSIEiZSUG193fyPLup+vj+966ilnI3vpTffW5cfw524TSFDMKVF0y9cKfo
Q8bkVxvNjoox9a4J5f75KEjfjU3KrjncAhYUndPAetw/0ZS4FqNuDcyCXHHNecyhqy3+0es8fzLV
z3WA1dAAVvYGPoEM/SYSJ5fSq/uSapeVYi/cHa2RiZ5IHYTZ6LjhAcw+aY4yHJTqPvPrO93SK2Xz
sZKMGa6S6KP4F7oI1goR+1AyBZyWPNxDmW5uGz7WV3I1mOQJ3UWwbvcn1UjxiPS9V1Fa19Y0bsxo
rSjYjeDIk4bRy5GHGPIoBUGk9rW4gsVPsu6EC6l324iApF1UXpKRA55OGdVgqYEQ5cHHlpzkBqZB
C2s/+bbqtmZZ2zBGC2wDdQLqV+U34766JdRK3kVBpVoD+SfqDz/By5hmBm6Uv14GeIGBr5n0Ola9
x+ZgYNjD4ifuITP8tF43ZfAJoD3OKfviZTEFYlBl9co3JMQd9GvzKxGrxOROAWdqXRHRnqbJnpWj
Q6XIgqaF9fNFSSvq6T19uJ4sBsCcRQqsOA0WX6ThpGyH948xceVw4dwW7vpeSyoXlJTm/w44klif
Z6sW2BDN6pvrHAxzEfDAmBVQ+ixCzGckrRNe6b7uF9CbePH0dhCPxVEt7OzpLtsBpiLLniRWuIuR
Td1jnhYN9Z5No/JMqSHLuY+HqS6iUX47VpRWy0t9bYIv7A5kyYdqbXFlhkrTjx0Wwx25eOvLrl2t
7PwM1NVeCe+99RYgoGUUI8S5Qqw4hk+88hsVOen1DPWWXbNx23uA/7QKJ6GdvdYpVaRy/1ki1cVl
A8AWHvyZwCICpFdzRMpddmMRO1GdNXFLW+TBuoeGg1Mp/Q7wCxv5zyQyN1qoYj1r1gMaGa5nWVax
LRv6Vn24pBQcEiwFTRGXGVAaeK6H/ryJ3gfd0MwnXCRNaBtaygME4+MCvkGTOigUPfSc6HdC8piD
+Uvp4JebjUFM2dPPvOodDwavsWXOQvRc0OIyjBe2OUvM5zdFQ1bO3k9F8sbuhThLaKWz3Ya60oa2
kdgxu22JP9mbwZVnDb5iZTEaUuAr2g65pzX/JWNUggiIqyvqQJrWkSZYhL3vtSsfDkfXj4/fQvwQ
eCsYUNdF057q1jgcXoQZtQ3LPUeBQfwZeU416F1BiDH99pe9nwvVLWG6eI/kDovsVVn/AA+6KEdr
FBagkaLm0iDtkIAjr7sezxx6ZfV7noZ9Oa/MxcKVnbivFqQoohHf4/vpszkJb4X2d57S6SLiimAo
RH5ZUb0zkXz9H3khqF+2hiLnmG3gx4h0e4CxjXFyNWLKUk9jU88e3GukRDhu0zFHPDw2TB/pUYih
u9QjE1kfih7sKNnWFyhpeh/nVLls4i6FGHiX2tD7yN1zZm1tlsH+0rWj0izAYR1DJ6blBiP15nRT
G7Y4V18lcalDAXh2PMedOscMN8VrMKIah8+b5XLoJ55dzZvtKXxrOdzbDUxcK8YCNoRdUWnLvQF3
F9MxMwolJPaz9iLDl/MFQaRYub7a7ivnNXr+pSP7nUbFhEmy2z4uFHuEibnb3mduSPFoQv4/Khqh
DJ1i/3siWNAIdYJzv0yA6DbE804nUgQ7pTbMUyLvprzHMFV3rubGzWPWYHJ22P/Q/V5wdyXXcabu
h4jjq6TA7UVjmhuLK0Sv2JX3yRhg9kLcILbaR3LfJ1+fTRk3V6LLWKJb081BPYnModCadXe7/C9N
ND3u3+uZ95w38w6alV3/f9lo9IbAlBclr848MaCvinNHnCFjOnV3XfXFpg/DZwhW3OK4v3EOAqpr
X9yLkLA0cLIzmAtWWDyW72Uq/qKo6lslqzLGlZqpFq16SEMZfRSd5nQERa4xiwitZeNAxRfHTEYD
TYwQk89RWt5R+dICxqkeGxPLq9R18ZRMQ5MR7CQzIc6mMH4O9KxFSuqcJWAgcqbLWpVCfJBQrepP
W6DcKgrYBjf3uF8XpPJ+pxKTX0fRffIGOOc2ydlKtDaIyVVL+hGPDeVJ97tvzvIsShpgvf6IT0NI
71SyhCzKgBpmf0IeRIULoZuuaEpY0jwvN3R0Oe0T9MhKn2ML+fzM5axxlOeoygI2EhsJt2tPi+W6
BecoJRyZsDd8bSX6mh56Buyw6QtNodUkh34o/oxd9t93IK5JICGtxOdyaYgo3JKtkdPRXFdUElpU
lut7ieWbBbpIBx2ne5/bTDQwU4eZpMwYvvUSyCM895rhuWvX4IF40esE2uUbJiPiLc0HIse0Cn6g
EyPEFCVqraIlqb5p3FCU7UYiwdcJQUUlKIf/xyrgAIAFzjBCuBARsaVzCgbjqjgy370EYicqEBxt
XIe+9h/EDTjJFRebI1DaVTg1Qh4VfSj6nQL+8R/v95QBGF2TRI9AjMYBC89+IZuslqfYf6yxozud
oXJRvxVJ4m8RTaadsrXQA56zqhNpm5v2lyBqDIyVlFYrhxPv+btaAp9VfO2iKukP+R5m+eBfuRRM
mCZwTFlK20J5KROrpH7/7dzKKhHJDaLp8GckbZURTJXkHkqK2J/L8MSzKdqB0FN0BSnETbqXChJs
fhZetLkheafXf/QgZEgEc5UbqxwdzBWAwZE+G3RgxfAvxtdp+xPe1n8jaCmvCGjrJTReMedemjY6
PIPjzwFlllqS4Xk3ka4C8Ou62EPOaIyCym5IJkt+/sZwx7AXUxw1EPE8B9Nd0UVpMLPMM9D9NT3h
od9YxhY4V+1ZnA2zkbGwFANwZsPukKvPF1ExsQTKGOBcBBbjUPsYuffgU8S8/lFCezjeDy5x06Hd
6WNpt3/CJ/Gx4WbsvxDzBAA0OXEQG2MQSO5/XbEUbRAVcfvtGO1aoF5OIvzU3/a1efu6WPYjlCHu
X5WV6SFP07Q6pFCxEOTTu6fMtMYJiVed6E233TfrOUfXc9ngouN/wTl8hcu+j3K7iZBbWNtf0baC
BrtfllBxqrNmxVxOHaIpBZT3mYAOHElbW4eKgDUVYG5J3n3Ez65pWSHtP2MYomaTKPQw8cyzWWER
lP7ZtOZ4ru221hd1ZPajh+w1kaE1+okVCMjfPRBo8OxPZe40HQOhD1BXzL9NYpc5A3TJQJDUS1ar
6KScLmnPxV2uUlWm8lTjn4GOkxy7SvOd/II3EhZu53ru1Ml9LmVtVx0gTSyqdAhvfrSofvImLnrs
V69zws+QCx0sHJWdj5io10FNvVTOC8RsCoYiWtroB+gmPWiKgsAME3YV9sx5gPcOw1IH57WH2ZAO
m6WV4xSLr9kv2RK9y2vvbuSDxVkpUuTzSCOE29VL1e2WyeJHb6QdKl0dL5mD+3QKdkyHDnbGOMgR
c6zWCAPSBBBuyu09E/xB5NkspzwXTWINF6jSSbsE4bAx+fOGEYggP82heBJGswp8IeQ5gwCtNpgY
geltght1RLlochP11c/VnQxK/fk3Hww/zW2R2i38Wqj+dzisGBe5hJSn6BJjsq5vSj21m39tIezs
WuSEkBC+vKG8FqDidJ1Ofj5VM1eZ48et4ZTbz3hfuZGHcDc8qAQP48PGHbOE5ha+4I3GeTLFqElp
7RYolH+0hhnRIMYxPCXoD7Iv6dCyL4p1nXrS1rRyOUk0/uPb7tDF9Y9nADeGK2YZTZmqYKGov1Vv
pOxVwmt0kIU4favabDMyqeljBa5dpmanQpdayvwjJn0pQLpv/PJd4GcXqdTQgwz370U3z92UIwZb
PDWBU8ZJojkbbwJp+uVqZ80T1nC2WUM55fMSbksJQnwWWf/KZBR1lnfXQbdGLjXVwAuEHUfB04yw
RsxIU7jX8oy2i74PBZm1hgOBuTa2bwgQ+elWpipkEZkV04ZvMRn5OCJ7q9/lfpOwEJoiIpZMCR2O
UEwLxk/MzsJb6B3DGTh0OdJqTr6QOoV44F46Beughrr8uoaZfXtdBMx2RAujHVavOI+rno8sfjp0
0oI6dj3y33VWy0fOGIGrL/hq3jC6srDPuc0AoL7HwgxPkTq8ys6b2pkDjl/3KHAsLf07wgZ/PKVB
7NKUzkmxDfl84PjJMRwmXn/uGvxvV+hBk9vfeEIAACQL959DzGGv0NfJ8lpTeejVG/g9SHkoymrj
WpuW8nYUH77AWf20cquMOJE1dAd5fb2ZlsPnHqzkZ/37hi+bURP4y2LZJymcSTqYDsALOH37ikOm
qkwubnNaQfx2xHrN+0JtVfKaaBXbiQT6pB4vy/ziTB0FpT25xkyis0GQyQe7Xsy5V3tWMquKtx9X
1ieVr+GTMojZ7/1GxWpDE2TjNFTTbhtsKXohhlDwIZkTVilwfBxpLQI98XWckAip7yDVTlpQ/kre
TlPAXMJ0hwDdn7PQ39FGo5vS5ZVcYZSxqj8a2pd5YQpejarpBZT3TNUgjH+ZyZ0dJeyMIsxERx2Q
iiJzQBXCZFOm+yuVMMm/kF/gpxQtjfBoIvO2cBRfWeUyzFtZnNqUM1n/wrUUX2/liyo8cB/6OWhV
Xt+lXrimrSHktiELx7DW/JQPQcGX0nZuHhrHYlSbB9QNE5pkXOP93TTzfylzlR8Ruc1M5ucBuUor
eD8Gpd5ZmoLcHJQObFzvWYg87opT3rSX/wqPpVk7oi9MT1hBk1nanjUSI+bfygL1Kfz8GD4P1LkN
f/bsFVkPHhu6O3UfQmjGjYSUK4xijT523P/58sroP+H7ex2PhF91d4NNKjeneQnUlXEJ9c6V8mqG
vQTPVwmRERUEcRvB+nvB0Q6dbRJghtyIJIaBYTNBjhpC/xKGWRJvbJiXF58HsU4YJkKY1Smxf/P3
hhDzmm2cWgNefEN2DZ2aMeVau0jbH1l507xOkIbrJ5YLIb5/dQHIiezPvhdmhiBe15IKIHsl6G3G
ZKG2FOfchYY8lmR4FamXRLa2I8ucOKlMNoTNPqGtgtN+KD8UQoBDCJLc0YX+vPM3QEubdVKZf4xl
LiNFyLal5AgBBhaMK4nKrC0XVtCIyZ82cYkql9bDgOgdVmfwdN0sqO2RL5hdzffpP4jRlGhSAPW5
pGB9KlnuP+Su3dEGS9mw/uiUUkfijBuiIHLMwwd+dCADbSbXFr/CGcKcP/F+u0vCex0bYEld38Mv
ll+R7kCbUCJv5QllpsodFJv7Z3R0u1S2i3UjycOlqo2XjaHWxL/s0Ntz7puid6zD6R/MIpuTUEp3
Ch2hAPrRbh+igjEPI0185rAvVsAOixO7v8rrrqIOE1MGn4nkDdGHdGfSSPZb+ienmKxjeu97eYlw
OtRzf7PxdYx5H9wPqCWjLvPvDlufn8ORXStzG6BFzAWuPIL26fe5HZOdvdlDgZ/FNyWE4YjQJiB9
kt1lt1T/MyARF963S0cbaI/0G7R9u1vbcWlT3mkd2xxRxp4uR/jNBjrtt/nvfnwE0YO/4HBdj+Bc
LBdEIU+lX2mB77UH6P7FpClonp48ct2yg8ruR2OHuoxg0IhNKjX63bjlGzYUoMBY8DSeA/7xNpBr
SDLJu0LQbJDJLmIEM7lbs6bUHs3pz+s//FTUro62LY3Bx8G6o9m3l8ur2p04OAKJqD2LVPjqcxtu
pGDxaxNdsh+jZ33i/R4mTyJv1vMsXcdgFNEBgTbrfEeGmMi/0jCInnOnBCXwKhNL1ZbTa4yO48yR
ATBtyVdAXv2PHccdgNatC0TtDQegRQTUu7hXhlbc/eGnBCeKPVOqmHVdO5+V3petfp1DT+Ravpmd
YiVIIEGICS8no9kKF9CEXbtC+qGX8UFpar12KAdxPmQkwPqNm7X0+T/Tbkx6rpGKFvsqKvHJCgKd
xCkClfQkQNH4h/ORkRYf0rbNqdoVFItUWdDeW1jH/HqTx/F1AYpgcSynUXOOqy1mHRmY9OMtfkke
sa7Ke/1CVwNniAIFkyxa7tCNTF1rlF6lghpbYHODOq6D/pE2hONwDSoan30+DI6bFNr/ETS3oTHS
7Oi9GDtioxSHZ/eMfl9Eqts2gm2d0u8Eo/O/VNlP7EVKxMLO8RdRM6mrP+s+5kWrVZ5eocjz/AhY
opDfTb2qXvkOaNanlnTYlg8/IE8yn45GII3BljpedzLsi1i+xyG2EqmEOh+lXTptAWLcXUB00VWn
+iB9xRcdMgvUYovuWSdGC3p+uEOTU4MoRjptQ9wEXkqHfH+18XspxsvrskrO2zUcdValdOtOJT1L
GLpA/qEC0+h1y9OvPI6Ij0aNpo4ssj/uuzi4u6wxJPQwilWgQrosBkKOccSp4eqkh4kLSAp+pdsV
q4NtJF/r4h6PkwKyM8kKCYqJckXXZK7DO3dUBLVUQiBup2JlToSxcae4MOC+DDcEY+DT9I9+J4dD
QQP9xR//IQhShu7tLwqrVDYBEDY1hzbAfEoTs6c6meK7AA4XGzDYWJ2GoVfcOslcRk5u2NNB0x+P
LrpK31niQRl/dPJDMNyhiH8Itrx7R9VrDlVbk3vImHA4fKMtsMyYrSnzzKDKANmCLV8hsK1MM7MX
/HXGG4SWqqupEZVwxkjnHNh9beOJpNEZ1K49CowUwEzsbFVu+HPdNWzKL5zHYHxBVVxhQsZmZon1
CeerU+FXOuY4m0n/rKevgHHrRFQeg4jeavqnl90W4R6IVQtYPIpWLYy61/dygLm42Mr6nrRMx0or
qHSZGQ/ZZ8EZygn/htdhiott7fL4Exd9EC74GUfu7FIHwmVjvM5DAVp5/tDZS+zMNKdidfUiE20d
TU+D+A/nRCGHr3Xdokk0i9g2GtTAc2fzeFvoy/S8D38yq3GDZWVByu2QE0Tjx7C8p+fxJ7gOYaRr
j+whIPCxsRJWikH9ydcSojMGzyecNI90lrX4eCzmLLlbapJwvOMtshnAnA/rB+YkEww2Yd23tzur
YoA+ESQ4o921/S7ewSDJknOkbZfXbBdKgnCWfsDsnRwJ7cnzo3vryGObLROTpvHZw1AEp+JWH3Du
6sFqA2mG5PvYhBZtO0ZAG8hCb0T/4KFUjZ6NLPuGbEqZJq9YYly/JQ3/Mvv5an1c2ZPr+btGevWn
ULZa1vOk7+EalIRNsfoIHaf6J+NHB9bMgGLmh5Wl6ZxNRLvlQMwl9sf6IprOGMBiqPo+nIakg/BC
amelmxmc7Xl5E3l46nBjch4qunYzsLlS1b0mcQkPdC2ebAIalS7U0+p0XSpLrnG4baulakhKjM+0
f6PAiLpU7+n8WiIYq5pVTGA3gk9Jbh0cBCW9/pJkKCZxKgI+SxKlyEOX9NoV0ePTv1G828dTudAO
OTvaW3EHvkmi6vZQXernjLcFbrQyr+VrYhfFam4KSzsLUn705Ip/iyIKrWDeWKSGxX6fV2XLV1yn
C1rwbSkI9FDi8vQOQ8xTXvZcudSevr4SOL/N3j1haYxW+rnHaaOSuZ0SrBgB62quWhb5aHSNLyxn
401CIp/uqBsWpRF9bxPbtEfT1TRLY2MbQx8BaBjENSToaH00t0GZUPUH2VPfkjDRL1tDQl9ST/ob
LZWGOF5Ct2VHm9rHg50gHkFKbUqcRm3pHlsn++EO9cjK7JdeL6Tisx71pyauZ/80e5vnFk7lV6MW
Pr8NrQmH8MYJQ29TKCDwEOS7Lu6vmPP5+R7eTA1DzQG8cbQcXpMlGkNlEVLCytIoZVD5PqvfKL98
R+opalIUzU7Mi1jsgCqIthRvvt6VLayBa2NeDaHZcEzP+4HvVkzBGiwuh4pvaPSHiK5RbRRm/U4o
mSZjYi0XQ+gP1PX78WfuGcUmjVtJI5c54oQOLGvEcGsrq/Hnw2cHoyqZjWocR8MXLeWP5Rj3cLYM
W/WtQNR6o+un7nD3p/5uvYntS138vfRD5B9E+uOOZg7INt+DBfo4k+0m/W4R2uVTJOTsRqoXSf+i
nF5tUBdFDyFFqwou8f6LT0ULeJO4qzfNS/yS739w7JyVmyzJiBL3n5iIlRPKJlf4yIyVPF3mIz9x
I593TLIBrEQusdzSPiwxAugNS2lSv1DZ/E/msuVEZCFpazvhgfqqFYt1WreiUyqwaB+3XH4BIv9a
AYqOJAhwfk/ZwyMvhHKpN9FGHkP2hmFIBxbfm0DLfCrAVHrnv2Y60adjW6i3WE2jBtqlNXn/jmAt
hvmBMYaydnSD5JJ7VzfJA/GlPD87IJ3VAhe7aayL7vvzcL6Q4uum4ggEv60d15DCkl8LjACzP605
d9OxcoZtInR692GYqMEAnnQ7PE7egaRlyQvG21ZOZ/XQafq3G9gga8VyADeDZ4dSRKxeTJJ9KBzj
8dc2npvlekMWitKQ74+csLZa3EF0kyFUg03WjrXFCRQLXpS1vzaHRbCiB/JeXDYiDHnSwTdfYY+k
gfzGOjWDGx8BOtS2FzFvuSeoQ+rRTN8AeOP0TOa2cnZpImXZGrHe2tg17nYXFBNd4NijmfCGranP
9zzwJjUbwcISmzF7DSujGYu2k0QBZK+sMCw1uyRsXxqFwhxSjaLf+dHw5aCg+DUEqNnd+gqf8a8h
5GTvb4plC+9QAglsUcnJkRak/Q8dChbYgYYT5sIPEe/ehgdE8AysrS4x7lyQynC2xYODG7zQVB5O
n8OeGsq/Z89SrOxkB+Zx782grjyJmfW0MBSS1G69BFqLjp8iuHE8stfk8N1v3A5hIc62ZZYrNbyf
iZwGrlT0ulyzwGPM7uFYXyalQwq9YK6nXKQPkMD/ciXtwLMNVpPGYIUoBpcY+gUNORlq0a7nkKsF
VPZt5xURGrpRq7BzE9RWUwI7/9TS2ZCzzShsp6dkbVPR6WJVaFD/KO18IBefVJOpiH26G85RYMQv
BblYW37/qmZRMDnu3YH6cz4o/iQGcMvzgU2cOS83LOGR1/GWFEfzlkdzmfWLqTnl7TPOkqiCMCZ4
sPrBbN0iIwwXmdl9QoFQvE448H92AwMtBQNQCYnE4I2H9LoW6LsBQhaXtveSWt7jpFw5rLwGq6cT
xbnyZ0TZhDQug/IYstTed0cSQqIzt/+HDKg3kWW3kFFu3nz91F2cqTBvS6A0/1V38P1o/maKah6f
apD/yQVQCbZTAQuH1V6o2rIy+JplAc/s+xigKWGRiVKtPvHrgAVfR3c3qXAoAI1/BSTNmlQ7BLBE
xKT2S66KMxvcgXlMkP0i//h6A407Vj4eMIZqjOoxB5KW7mOSJfnvsOn6N74r0KgUD+fsUF9NelPT
DxSpIwVy2jjtKzh7Exs6GxoUIpkTM7qj4gtyjyuq2iEgApa4bvgniKMn2+/7DLj+LPnrUZQwMX3K
Dpjsbx06E5fxhrhKqO2APY/Gz27GYy96Sj48ae448EuYfNvMDMx/qk7R4iZN2hl128bQGRxU9/UH
mAt5Jg97tPMwDXZjQ+jkUzG+HpYC47nUcdAE5qhpn5Eo7FmjydMIcpKzGVxlu/3+KPeYmyuZhNFh
dukqYOs4/dsl9wroW5GTnZkyvqzPnZjQBbLuwR67xxgdDE8GCBR9ziSLx6L3MtayBClAgHh5hUBv
F7QwhHTflo8N9qlyUSUQQkctpqkXluNghUC/keGEbAMhjGs6bfGam60FyfGEx1jKq+iMVrQ9/I9u
/wkI0UrfnlJXf8211CU4sfe2SBoYlGqsmiwlb2vUk4d68rtxDvZaswM7t4R6DXwhFDpkWd17p4/g
JbkQntw42PwGb/S4IninmuJz/0t4NMBdRTIDOmWbaQm7lxt9Dy4IdX9B4jDfttowKqKnW/NZWtDg
sDhOEvjxFUvgnJ1hOU9TUpycKayGRZEDJmnoM5xaB1kvtem57KLkfKVy4aKRi6hld7yBlXUYpNNd
zA2gKkTddeqtWlf/zp5cqvH8q8v/NPXadCxwcqjBxshtwV0Kx0XQTRHcUpdI7T0FhIxUF9oajIg2
TMAubv5IZSkmfxIAPBBsmClYq+BUTrAmcLAMyEGWv3KwUiJr+wOGFaH8Zef3cVE7/6s2hWsa9ga6
e5ZcsXvqJkVpnRkR6YcCkhDfWIBb/1oaCmWxFZm5HpYXemvcR1kH6xQMsfJnorPvpidya/dyfb2I
tF6SCl1fOTorSr58JFO9rBLHQk0Az4tP7lOmi83FZq9B82heEOsn0PWCEqUYaSMYh7X4WAF7MJhi
uC6XLpg1Z8oPVKNG7gzKvmWDMP8vUwPN+Z3rNVf5hy4Ozi534FNusLJKIN83VjaR9mty99XAvEGw
I0WL7HZdk6SAdanvVZNhwtgJ11GeaaRhiwl9dJpDP/NEa1R053ozuGYBh20wedjcl6SWEnIkWW8d
RAwUK6LgTpzqIP1SZgwQ1sWzFiDuudenefI4eo4CUAR0JnWzYYI66tw4h22SN/t67744HkQ/IwxU
b/XaPhJnAzp9Pz8QsPLga6DVRl099uiqpBajlch+/AX1iZk2XZNbmvCKcLHdm3Gk6MJKGAGWv+3o
IQu2ydZGjlntu2AtWLflm9xwO/ezIfKkTJ89FDG7BmzL9ydMqa90ZL0M3jSD5tvIiFa21zFrh8h/
7keI4/iZY6dpZwEU3/VgdCOeo7BF2h0o683mIF6zOn2WbLf8ntn1rMnpcuAsL1rmxLOGELPlSDj9
dBuk5sdRdczOlvm9jyaj3qbUFPnfIqpDQ6TU7jEU49UAoL4kuAKsYM+75N/mBHdOvF8DTy6T12ZR
Q+dCxUeI1AwgRYxOnAkDc8eP72UHyQ8qiGzMHkCPQgQr/xEleYNwefVboQ0OrBNyeS2qYI6JKYkw
y3IYJ0zly4OyTT3WrzPlyKSZhaFrCrpgvmb+c26ARevi3eGYGumuszyqss1ZzLE521h5Gsb6ucGd
2e+lX5xugvcIyHwZK6ETD0NnbFLe/X1DVGKsgoxyPkzBG7BaqMpOD4xdGNT9STbrJMpwS9/fnoVm
vWQt9It588h8tZ1dkUnm7INIdzgcn2y38+0x0JiUqaIyZ47/Fbjm8huthd4piRgKXL0vQbEoirjI
D9pgwpiHAgRehXmMEYmU0txs7RIdDtiSopWSqEuZScDtkdCcVdG9P/fPudVEVaFHrx/V9Urd1rJf
tEMlfBgIk1voOb0IEa+96pM3T3t1fnWiE2RPphvfisVK9topYUM5llZJf5s0izex0UiFn6ztdqGM
aHDDiZbz9NMv+hGSviW77YJXKhAp9y4MHXKnAKCzAXuRS6qimm6flxnkwJDgGA88Tl+/RDp57a6U
MNwZ+9yfsT5JWghpHl30ceaCClv/7eFL6SvMvVYkIjwiRKtVK/xSvpsXsrTKYocSCw974iYls+2E
0PXBjo3ddZLkKL+IQzqVPdA+V8IbCoQ0TfkbaAKJH3YDqHJtSpD7HOxsLr7LDuwn7xLu/3MsKn+e
5e3di3HCnPNJrAVb9+LQny+kafWIfZQch8U4pqT8/PtdIupTL7zYZXnP1wrV+BEzVijHuGpgKqIZ
7FtNMgSeFgz2wlRjVmBhZH1ecFvyHTOuE9F1SlNXwldA4i2n65KVTzK+xaxh8rAfcS3twZ1PlT88
6mwdniFWFbYaaQVCC2HXkmOER7WkMSHcAaj5mvkKzKx7ZxsUkPhXMXPJV6IEC2HEtztOBzmKM2zR
vhebp3anMwoIyFDAviEuNp5XtL+gtTLsUa9tN+6bzdbovD5YIe1JOf+95qss2bGB7FX/jyMFtQMV
DjZZp9PWNcJzmsBBAIlBHilAjM7kItCKlNXAeSKqDTPCp235Aa1ujCfzFXALlfBPZp5jonIC7CNl
ydbguUaO5kL4wwccdqXne5w4hqMGXzwIHAx4RGzIddIgB0i+POhCxCrNYxo5BW3Xa7v19u6sm5ku
qZ+fG8IFLKh2zalKPnJioP39CtZfiUJ/fPvvsHpb5d6auWrLuAtuRJ5eJmILjEVABEZATRerxxHx
NSxrUsLEGlsgX60nanjuMPVAMdN+dVlQYECgpm1Q0xO90+KsbjQZERtL7tW6FO6TMLZWwNpAtfoy
tUN6pwTliDhVaBO/Fes8huaDiGzqVINJcJgSwTDAaoYgase4katqz7dMk+wJTiDz+fqK26kvpm9R
0IMa8BhLECUL/ED08g9g0zWV/4d0HWSjlc+o+k1aBaJbly+13srNkPcy73XA2KZRLfY7Ij/3BVqk
kZXLcg2crtvp60H4dMZEwILQZ90fzQ+F1qDalSf4XYzKvf1hdDcXF58QoF79LgzvJOis7lcdV3WP
V3UbVaNbrophYcAgfHFUPm4Tr6OnfSxNOPRGLr6KnKkdBHVP+ckOOfjKoWgMxgJI6F1NJQZPKgZb
H/CjAqc9SgRr4DhD5n/Z74Tu/1TNlrTOJ5cb9T5SeeNpUnvQI7eLNO3XqND9oUBoLDZ8ib6tFLAh
G7PY7GO5a/axv/rsXgO6C3iB6Veu+5lHJyVyDuIvTGgsZPW4zCdRXkinD9bO6UbfPdgYc6mDw8dy
xj797LBecha096tV2t7kvThp6BU/g+6ICfDVpbuZj016Lw/wOm9KqQUMeWbl12p4iH9QwH0+ke0t
PTLSpceLKhy0aTnALMvzb0SLS72A8hJLL4A/0odA76svKKCQMZpFkzAUE6RKZ02hsqiNyxkKZMkg
hfgKLNMMNsCu/gX9v6ViOkzdISwNjmILGn0ScRbkXAaxTWimgfZiDiRGXTR38T4n1dEY2Qo/0lxg
vESUlNapfbXAelV/7M9AhNWdHxEosfEZkjkVijITtBVnls61pAVU16cFvwOsWr05ftGPiOSMQU9b
A8RPh15Bgl0cSkwfiav+TJT5L74EsJ18gu1ylNs9INWuoZn5e63bheeIOovohk19+WPuawohvgT/
OEGRSecGGgpgGo1pb2lUILu3JD0jKWjXVpw7Iad1vAblTAf0Wjmqxt8QG2TR4mGGA0SO80VqxTA7
lbvtzj4H7wYEQYnnRzwmJyZ7BQu4HudxSi5+3JMws0Ic4AShSmF3UvCBMQRzzb89LqXbfSfaM153
qA/eKYs/ujvYppMeTvYidmPgqhbwec7M3Xgixch5E5ndME2zdQ/q3d6eq3Dodk0YfWM1hkaFQX8C
lJzvg9JESbPrimqRtw6ivMdzpGrxXkYZuezretYMLAKwyExHBI/WCc4WKmMKMeppz4YEEzMqogC+
0HJY0oH3XJaILk3kmbkm24bx4TjAgr5B1CmOQK+4yO+QJAJdbDVdBxeJqtws2A6C5pFQHaYSyx8G
2nQQyane9uZkzwnUTqruFECP+MY5c2q5yLC46nJww9LUKlYId5mZ125eABzAw4Cct5DMlDFi4N4H
IOBkYJvUGtaQMO3+cysnuMahJTx8TH8m5+VRN9Mx3lRFjDswtNZt95NrfizLy5ym6LQD7XsWYQXD
aRB/EWlaRXDNRsPvmAemh8XQJvgMz5qRFyft99Zrp/1p+jRtkXkn/1S+2WPX3EHybV2mnn8+SuvE
0ABmVzn5OFJXKdkmFDZmlb2LXp9ms7AudD9QDHqv6yhFllamp89Y41LzaQTE6irD5mQBltspdcjh
v1hXZxmipDDsFbfn3ukHT6vaI01TicI967Oq7bmInYiHoYqkO+qD9pVarKGRIFXLwLEKCqvqQBbI
MYuvreuqjn4TEDxwz1xKxMT2EKR64GHIBQVC6MdiF6BD2hmz+UwfqCyL71cZHeyFL9sS81suIncu
HZXUjtAGxyQLM/AQj9B3Q67lKCugDwaUPQ/qBXwJlExZzhmo/b59Bx+HCg8fQN775/x/7s3TqoAc
VgF2tMYOAIDPfFPA1lKKL/fIsl48Rc0uOtiBKJxdTcWRT9ivgfUgZ3uFdi/BE+R8L/4Ia08XOcBE
ohpVeDYU8HNyFtX9y1qvn8cWyQuW8X44M2YmFLeIZDCj4x8TCvHTeJnVZnEPr9C3+UqQaNS2tX9W
0QVxcYJblCdIJNzU2CGRSSpzmDMnf+vzsb7Qpp43nsbbRyj9gqY8aompXeV0mkjPqPB5DoRSBg9s
yhEieJRFGGaWjT6EvDjI3pynLL7jXdbtlJAAWbjkka3ENH5jn1nYn/lRNQ7tVqepkDlPYDFXBgvo
rJcy1+9bB2Xe99I/HY73pGi9RoYU7J93vsKPekzjT5wLx9F/sDhM/q2met11PzB85ErV6w/HByO1
vdLyS7GzqMfPErt7wH9UqjGIMiy2SzwN7+vKVNC2NMgLxzPA8V6szICfBKwlp1md9eYRhZX3Xptv
AgdfUr/NlwfF3C1AYtU/Myhi49THEUnoLF6Cef0KgN/3k+RUaGK2JF7DybmiEYHHmTcst9fu+g+J
lb7q8+h4rsBy8WiwtWqM/cZ33hfXw5qIr2oJbCkB1vYIu2xlCwk7a+DEA/CmshYomSVf8nShO1Ze
vwSPXgLSDtPSf6AKT3vY/k75qkar04LSLDSvenZQRXUH3+OJ0r9uR5/9NJ+09ZCGlub91SDCw+V/
KYNkXaClATia7ZTzOAqLEvFSUNCKuX1zDxs4vhp6hLDjgruXkSv2tDeqUFXTBHQW6fW6Nb4hOwka
DWKHAXHgBsgVlh+mqh4UBvwnwzGYEyNCwjQKpL2M1UqQQw8/lFgpQ2oFRGulOucNakXxsJGjD31+
cGN6iNx0/G2V/nWgoBKIP2atLin2vzBsQ8Buj0O2JZnJ71r4+qdePS9FnMWtHarnmQgac9g/X9pK
Us90Z+k9SUJ344KEWEffDFQp+oT+vZqEkWh7VHwH5br4dEd5l6a18DcGt0Rdr3h7Qt6cGScYfvhi
6ryrA0hiNPu2+UjvVVgavBHn5Be4WvEl0awXyU7owJSyoP0Aa+PnryqwBEbG2BpyOaI46E+xlcf9
32ln7vexOoCdxn+tyR6QDTZeB3K+vHGOu3HNeoG/USBn+Pwz+dMFRL4Ng8+sdRAxFu/81UtoeWVI
m32gKQ7lIXL8ujGheYGXxAAH5fNnhqG4ESiqd8OoVxZDKGbv6oo2dlxqaoTdAagu0y0mwm6Z/owU
B/f9YsMjBx0EJWXGr317V5rlmWcORQHcauKsnXzfUWjxl2s1mfRCICBVS4Sy0VNmaSmj2a2u0syk
TKbje+T8lKpEdvhRotNYBEwuAjsXR9itX+JIELiVuYZE7J1YQeKuAOgpnDeufBcByCiVmt6Q//AL
TzYGN8O9SnjXA7Q7hEVCwhYg9opVSEn219EfBqGq1JuJi2BJv4FUFXOo3ZbGNY3P59WyQiRpnISq
dJIXsmulQRSTgPBpU/B5MyElvlCqbOAWoC01/nXBIe2QnDmzaI0+ZvMB3LLKzqSS+JdBnK/Tfj7F
jATpRjWI7F+Ha7bTVZu3W3BTfUqOez7RYq0Oq/fS+E8BbiZoPJg0oiuxBCe+PZJQvTcBoq+yIebq
+NlDnevK7BFLrPY02ahTMTxJuOykVKXBL7ZdlNVlmuY6Htphqn5H0QwST54YLbmNUKsA+dL7ujvj
7+fdYaHqHVfGKPKxV8yEcqX8+jxSnrtcMY9pqVCPBGEeeukJn/ZfC8ieUNEulbjQFzWo3+8SKTVl
iGArGIcolE6ZyxXYuD5CHOtMHL8FU7dlkJgLtW+zSF3Fjqm0quFbxMNarnxxlvqrcRQzmtP5fR4x
Dnqp0Vyq1Gs1cnLvY0lSv3GJ+1XL1xZuaE7CVctb9vhExM72LQPNiRbsZNaYMZpRNW73bTETQJxH
J7tfk1NFqohAy1cRkC6bsBqHlR43hz7w+DBXz6unLZho+qjDec7iRaSD7OQfADe3BJ5i0tR8fJNS
PCbY2DgNYdgU0wBmQ6mi8t6/uBIhlyuwoF/YJB+tzqbMr940NXXqNmU0zcF0qh8a4aNpjgz3p1ZO
wj/M/H5WFH75/PpkVlXuEUiEj3db4Qws5WjoxrGou+RdqV8H1Ux08bYcaw7+Hvuwk6rslo8ZhCag
ofsd4Cbjd5IjWnM5SCNeJODWeYGOz9MxDY0sEL2lC/FehClWMEuWX+Q1iKMBVGSQhaAI+gM5Uoma
TcripylTkmMND5GoabLoi43EwR3p8LpA6e6h22VHtuVQhi3QuwQlExM5CpzXS7lANfT/MoferPMp
8ec7ZBjzENx0/p7PaMmOaLI2UnY1onkvZYKWTNtdCr+x3+OoFWBSSJVLIr4LgZOky/bd33pe59Xy
7eUr/UfyUCdvj9HSyPNpVN+fCBgjxqmZBkyGURsWtauhzQ2BDMYitopYD39YygP0Z3ipddToZDyy
1vwgU/H1bAAYDFZso6ncPIg/087Fq+6Miuc0CJQXFgwdZr6M0YjYntodoobmp+IjWvykB/Nbfawt
+KoIydL+0HdrEjwK5NAPDMbZPo8Wwra2MdYAj3NW7D8LPeeSmyU4FqEQhKTz4mHTF5y6KuQtJoKT
nynykIJ2MH21qkQJUTY04z6KmfOzdQXpp/96A6v43s9fO0vqhMF7izlSQSt2+0ISOZfDlGdkQNUn
GOjvJru/FXWzsJwgIMwUUrp/iNmFKM8sLiIavzt5HqDoJR5zd6mtudSYuiN8ft08QJjxQVv5BX+s
sy7+JGblqwXNmd0KEz1j5JjVhS4TdK4qIgzYoxLspEEPJnu36pG+4Kp1F3sRn2CI952OSYihoCmq
KamPXQiITpnZqQ1UoiRt0VhLPcL5TkI4p4SZIvjQnl4+p0AGL1CQoNEQJfp3o001LyFfVVjCtDC5
3oVwBY85gQThd7RLqtHbx5JJ4pPCLfKMwcoXFNiUpjUlRGYpO6+FmpF1DQ6OxfmgzOQ1W1swC3PP
GBGqnJDIcBl7M3P4cfacmu7oYJZKSr80YvjR0KKSr1EdAvz0b7UGyfX9k/lWX2j1cgFlJpye6LNF
pp7g1wnPhL/+5Cx3KjBfZi0+w+8m3Ni81kV5F9Uc/6RlHLoEuzr0p8AYyeLMwNEwT0w/g2cdSCFU
D40m7MvskRijfnvja6KA7XRJi9bOSfQ4v1v9eYAz8eUG0A5Y0MhHDJv5ArKeAZZyr5bKnW9WFuT5
E4I7BSDBsY75k6bzjleVM4FfVu21zc7UMyNuUZ5nwmrt5gq6/AGZfHzrLoy0hyLd/lYQ5E7XvyzM
R3g4RFDxYSzQqpJESCOoKpkaYFIFrpv3aI11/DeA3gpre7cDJ3jY7eXd2dv+Cp2vlwJaZ+8KYsTm
XqEesrSC2Ikh5E2xPEt206j4zKwVF/0sGXjamAYRepWfqlRs5r6vuRmvDqlxwGpujVANb838pyVB
k3MHvOVKO30YjFZ7kVMwSm3dYWKUjYFK+LehK/023INg+E4dStstzeV8icsSA2o8LJPvy4A2I4RH
lECYtE3HjpFIzkftI7uzCTLVJLDB4d98Bfb5CmtB6HZaL1fRo0O7ehgFS2UbH8qTNqTLoCXff7qu
2WKJOnhdqFsJkba/9kh7H1RuatuxD3ryOM+NN2EJCTMYL+20/vKY6o/1VlqSGuCQrFM6sqzqMi4z
ashA1NF85FuPO04m8X840y+kRpGt3r8pO8YCmcyitmu1L2BHYQUqvmzbuXXTmO+J8NSss1qut1SM
GnxDHtwD7jlR3YWVlgS1jo72nn25dYz6wPf3RmtPbNbDu/J5SKwoKBQfNTJWRUMuFV1U9O7ATJUZ
4BZLjaHIuWuYwRsigsmpRLnr23AUOoiieQER/M/Tx9nn1pzKDk/AQGDNUyVlTdBHKi5gXF4KJdUs
vs9uInpzkQVan4qVhYKijERrnLQy8oaQYQym5hFhMqbtwEx1F4Nvlb/l5XBOU5CXvbSXL6r1edT7
rk3lxjeiVt8ppfacqmd1sQnBiqY33oZWQJuFy66OL5QOLJ0HLzQLzzdVbCbsVy4IYdPa6Lrv3iGW
lyxA6KVXYF4rtxQUNFqyFVXeg3NO2VEE65E3BNfs3rWkY/kZFLFpIXpuhZ26gKld/hrWRAUQcd6U
K3hLGN/Eh62I2akgql2nvKx6HKqwEQVVvj6lf1/6dWZI/hGIZt5zZm/5cmGo/5WWxr31WGv5jTht
rPlnXxPBjLARoETQEiFr01u0w43WEUDq2katO8tWsfDBWwjmhBpwVebD9+8gEQ7xa6/scjtDLjoB
jMd+RnSb0DJN7i+Qs59pHdbaK92JJRszPhuH+EDzznHa9ZOKMCBZ+zdDKFmOFo7DGTJgrzqOfb5B
GFQpM8tDt7GbGV5yU25SaJm5xXuzXDsREfb604bPO+hO8perQwqXZs4cppdTI7SP0k+KBFndR1QQ
PzwXZH06Umtx9mX7E0htRmf3jgJEyI2PdGdQpyiE38PPXhoTFlQknfxFezoMeHD/l5ZXXUayxh9y
DXUkX+LVHD3Z4YIjeh5217PTHbEJ1oXIAMGNiHbdY2m1w+xfvEY+iaBjtGikJVQ6BI3Jkb1kpvQN
6JXjsBNWlw24klEZm9MzWhlwZNdPA5GgrYTzHooooyZHLbBjf6LnT3c2JwbcEHpKS1/7X6gi1533
apYnA0JBlWJH10sLbHShWkKx5LNic9FN0lgPKNjX9Bz5tlvcA5vO9MuUuZWwIA605jLTsNfrTFp0
jm/r8t5E0aGMZaLxJwGqjuQjYsFtjuAQb+0jA+RQoShVmGQNtTuC0EMCqcv3VKObszcGnzc2XB2w
a6YWL5TyPBxYM7Gf0h7bWgpm6DPfts5Inva2Y3O7hJY7lPAwxj2KjPHb3DoTjUGqx32qdwyA0+Io
NbINLL4Rdl2lxSPlhtOee+XIYPZxDDdgvI81zHk4Le/phcBtL4La+jiBkfJNupK4KS9KH96lZrct
biUVO0KUuYcMsYE3ZnTXYQqr/p/twEdMoa1ktvyJgfcBOVxyQEtSnEMtSDTgQgUwZn9CwxPSfFsS
gb9kocp+Fq2+510mftnqO7cIw+ZX29+MH7xKoE7ydrRaS3nFlaliYlLZbzoeQX1NFJpnTLGzAhMI
MXETI1h9+SzMZ5CIvgj58kjB7u3RX63pci5IssfDLBJGG24uNuL3i754MWUsX++cCgrAybLEIXS5
U02idplUDbKqOSsjuOrzXepvwohSJwptHz4Fo8WJq4N/hJ4hr1mmjZiG540mfkTdzILiwBJ4yKjn
HbygwDVAL5Fxx/Cv5C/baJIKgSVZWjnKx9EpKM1WJhVXL1SLzgkzxEYxSB/o8nJphaE+tFpTUEhI
EMsBe2CXpmdw5i52SAJnKg74HEQDDLpLgmXVzx7JRO2yoYLGXZkedHW4BUNYEeXTcyV7i9B6SIzq
wgNljQMzzb82UGzQgNYD1h+5ROqeHXKL+gqxd54pLTnczuGHV7qNSePlZCwPXtmE3Lk4WV/rkrVz
UUGS2OoE3aPrtdIsDO33BQ+nd3t6sJgstoDn2aWo6goq0kkBw2oEVCGFA6BxaNXs8zOZtZuatZNC
GQ0PB3lI0pChzJtowM1aXsaRZqLWBqbxf8Alh7BhmgQ2U0KFK6xtaG4q4+4w2IlEkg+bRM2pr3Nj
iE5AFIOxAk6BBOBkIGKGGKazQfIdvQinii3KA2mU3FDoHjqNwoW+Y6byD6LC/4vBP6STGPZtcGmZ
NxGClVDa7L78Zdck0zGTkp/Yfk0NwnsqAUfYQnFAeEjsXEUXpXTi9q87U82XVrvma5h7dz2DbqzD
H0SNpNiT4/NVmgGvuh4nwf8HK9gOmLyTz9NnZsvZ7WwPEVIAszUti08LOaLUa+0t6tABlWJtDU5y
HHA0wgINqGYJwggZo13vYsq5e0pyTMoQSKdPldXZcWv9FIv+Gdu2hSpfdCKeRcUvgsbRtv0kLgAX
Y/SZfcHrLN8/3z8xRE1iJrvMrTPVheiXiWen/OOvUvy4n474TNLTWrOZxwNDsFNXB69jWnyG3WCO
w/tEyVMESL0orgDH54Z7Y0/W8Iy3yHBImXJoIjXmT1WACvZbIvd9qvXJ421VOri2aT/I+LQ0KvA7
W90bh5MQElGhzzgszHIVlA/bdpcbp/dKrNbLR2GhmfGYRLiEeGL9FHYF/Fp/eq78LgTxuHEDQctJ
sHWC1cW5UiAq4G1AUiGvYNMJlIiS9HSohOY3Uwl6yGPt8EZTwJzOcr5bnE6N0INR7rQ6j+nIUpQq
bAmgAj5mOfFa36nGJ1L9LmvWrSXigXtVIVzut6iaD3tGrHXC/PSJmOSigDFLmF2B7X877l4STv4g
KD0ThwsX7yudElzF3Afk63brTq60Ooog8yz2Ax7p0U+I84pXqZ1y5ULMNRhuKJnFeRAAwybjCa5h
6JwUckHoazPw2K7nsfXLCc3ArnGQb9cm7G1dI8hmxO6Edi1URYiQr6jk4AwjoMHrRElbSnT7oiwt
8JELRMb40Vkp9uAOqy6BK8qyIHh85CQbUpwncuKSbtK7c6VszAM4xsTKtyzGqQXuOhuMa9X0IydT
U/3pTbyoLDA6wZLPqrVCRsjVIHD3VeIXDiA3wQ5hvU48vy6tnT9yq2CY/YeTebkxdkAgWYjgnLez
v8z8oqzY1CHZCWGecT0djh0RcF8AUg9+SSA06BfXnWkTfjDWEr5ZqckWOccfdMjIMfB7INUiP/1K
qf7A20LecK5tw4cF1kzU8LGHhoJT3ls78rl7O+r4TGZjx3Zt4MIZTyPhko7askWKhjHAr3hpFVM0
zq9j48mjh85ZxjcJy+KIiG84A/5gQTR5eGrqtiJWExytgnEoyFm4JHWtsNs6IK4vBbpvbrpTSqb6
rwx96rtGarxK+wjsatJJaJGlzENbc5HaXFrpvzanNCfvIatWFnm7Epnvb0KKvSnUlRUcDSXSbVdX
v63PLI5H+oCTQibi8KdadqsMmSWmbHTIm2c2QMK0wIC3A02WC3XWhqeCoHhVygSvKDAx0JoPbkMF
Snt+bSCKREJ/nwbpPCC1m4apkrRhBPOPuI+HdyBvJGmrEnMu0ughucSpFFPy9aww1+v6K679/5zs
T5FdyIEJC26DaQgtcpM8NsURdExFM+T1zRGYi5CYL+JpNmc19IsnjvoWbX+6rNo/iYXXC5S4Blx4
riUql27FPV0lnVsoIEta+ZnB0RKDNTBt9c20NGBAV1rlBNdFM+44F782lEZk7PXim7NtDuPNqohl
nQvIQFOUedAj79dL/C620mFOMsppBzz1mV8jzwuDVNewF7r/L1aBg5tGCQ44E9/CRPojp+DgacM2
YBzVxZ09PpOYaIupFmWboOqZupDY+KA463Re+KyUXEAguceMtGPd2J64MiykSU5sGBvoBPPlNWEf
wlhkDRSKsYLk8CR/pe1DM6EzGOcoocIGy7yu90U2rnRv4KK83R0XUvQZsTCp3Cz9wWW7plUcjKUp
pdriMU7KqiApn71HZhTe6N52SnXVeevFZ2ahmk6ihevhNOL8kFs+I9vSL1bReYWYsV4uvo0Xj2Zs
b+aO+nHUD7vd1DXbp5pkW748KQeclMa11S4oLLFSEHi9k1ide1c6jpitqxiZABydgMwKko0LZ02e
m4dnBk5jDRvBG3pVkpUrAKStecIlcBHv/JHgp0IcOu29uWdbYfRzvS5UgPj8pCaHfbcfjB2NyttK
wCtSETpK+YgapjV5Xp5XrOZUHDRmnUz4RHLzMFlioJBr6Z00uI6wJzbN9BAfspfZejgj+b1QpLPW
9Xh10x8rV2mj+RtsXIDzF84zAXScdq12vDqG/f3VjK2GMU6CLcWsM0MXSNnCdPfA6JK7SU1t9QcL
Zzscq5tHlDCszsqYEtBzt2F6X6hnr5lWUNXHzeWFjQT5Bvc3HY5adiZ8q5k3/LoPbroOGA66Co1e
LshKvC9BezF3bktbaYuT7pKggidlB8Kz+qwCW6qzUdUsNe5HYnVeag7METd5v6NKIBDUi/FK4g/w
MhW8UBi98pAKrVi/jxqkRayCvpWNds81VGCw+pVRQEfsVkEOeo1A+NzsBmNsnNYqxhOY8iwpeMht
GUQOtlSYTtJru6Y6cCQO9vwR14hkN1mRvSU3G/VOykU0tO9jbyrVTUQfvGBBD1jNv26v94XsT2su
C7/ZiBEbQZiuxAAM5nEx2wmpQJUe8Z1t3rjI6xQ8H46+lyi0jpSPyQM3UORC2coVeAvxQk6K1qOp
IS8gQa/KF8ovt5hqGTZ6E3qpuDei1do4DZ4u/P9t2vGP9Db5v6VaxsTBFOKZmwsS6kwIShx+W/Ft
rSD3K3WMU2EAyivwdsyIgMAW6vujzJJtVWm+TQHWFWdDbalS8SLkFQeUuFuOZ75koZ3Bi6+EWGzJ
WkJsMNjgQqcIAdkX43Wklr4+rLh6pfitD7zh+QkV01DtrW1yacmdnn2DQIY0zq4I1VSwVbBnXTjZ
9fBcZ2gdYodmXuZeXG6enaEPeIVfr2OhZbasNBE43AkMI4SgSrhiTk3Nd2VTbC7Z9y/L/UtZoo4r
Kx0QIfcceGi2jlHAax1fLoTu3lHGm5lJnKA/5tpOKPVyJYjwV5Psk1cxTSRG4AZD31WE+eHcZg4v
CYYsK3/68wH7bf43vUa0TmK1EWOoHg7Dgyf1WnfuNXP7aKWUbBdAvzXoyWIuA9Lnp91uviXmmCU+
O8rlS/BjOguwhhTYvYUvAbKiGz97S3jPky0vtCH0jaiNEQiJ0KG/ZtUNE0EbwvNEVAzses/4gsn5
gU4nxDgEPyCs50LXipEj0W1U26iYr2eqFdP8AbH0bQOPB2c0dbI9u9f+kna4GfyLBammeoSUG+gz
dOsmMlJTfbaFDLhg8jlsMVhgAN56EMx3cHic5KEjoggOEn3pBOkAbKD+nITH4U1DsYWD1ErR+eq3
M9OO+viiky+MKkRgiz2uVlnjjo4sYCg34g+Q7WuqZCDhUjW83IO5nzhXdgVoPunPJJBmOIyM3ul/
Y5BWzXcJMa4DeV1IQEiMd2nmnoeMOhDktcualAo/dbglXZaWLc2W5b1gUq12wfAjogzZD6S7Epwr
HXXH7DHucyePmlv1BqW8zxQ4vuke4EDqzoOCcq0sh94Qwy9Wfxf/uJNgWMT2fjVK+GFVhh6j7x5F
Qliw0MUqa64dPvqyn0D1LjvzPr21X8wQn1PE4JF8zAhPw02Dd031d9qZDgvTgfaG6iLB7V3mHsld
aRFMAFYG9Ijdmd0hAyNJ1CqNQz4+TIypXw82LJvsy2+CPGkdRdzHcjYyTQxVJXlgE2sL15sgvUYg
BoFtHJPb7iKDxsz/nR55m1Z8BVVmx1ENUVIkZ7caWmB1npw/xUC/DvuK7qSUl7y3HOJI58cZYVAy
uu9lXBtjAUhRGen5w1UR9s8oBWBjl30wv+6OUznvUoIjYA4MJQdyw5DpndHfhCBRnvTAk0ieeWjh
amRSDxwygmQ7OtM02hAL6BCBNTRwd8n2IvphsNGFHG3+t4IavqL0m4TffvhbEkHaNc8HdZ34egB1
1dupysCXI2+juwgmB/7mRelbQd5vMICMLK1sFCgVJyZWB2E/kG5OwMYNjtJJLFnotdUbL4XpXWhy
04fDOJLR2C0mWOqPKzpjtZAAlZaY2lx8CH/3rAZUpdgQGbp+HewkmyY6/bG8fvy41av1x2Qwlx0C
OyLyVQMWj/29N9lqloxu++BLiUz8TRuQaGllfdM8Fj8K5L+R7quXtlXI4bBEZRmTFqskWTUP0nN1
BGXw+5U20sFjE+nKB0DpeDcbcRln56HcyUGiXgy/osTcyGF0WOP/gi76x9LFfFY8Da4S77ygEmNx
ultvosyIGDZiWXiL3RI2DHsPXlSCM5XUTyeoECwvdypHf9wDLZxgn5LneU7vHS7lo1+AaeHt/mPT
kLVF50BpAF2MbVjFMJt3qkmCPiwaz98pp4O+HsMHITZkooiu3vVgSomuNGU3vpTGZ0jC+kN9lLkh
yk+TTyaGcTlDDbFhrtDILuPkG248nis81jZ51bQgqliuF/qSNnPr3kxtu8LzSOuU3IfQj8BNmJwI
ifHE5bX85YKukEOwHwvgRsyqnSANLo1TH4N6j42Aw/NW9Bjbe9NA3RR58wA8YmW++bpkxwGvqEec
out7/etmPADB3/WNXkcHdxS7jfwDvsrTcML14icehzNi8QuF0hKICSPrCvTm74fZLDUGX7Dfv3G/
Wt1OneDaOcbZu7qhnv6u1Pf/380vYpiQBWQe93ovD0rOxou+j/8BB2buR2LIS3kPrwywEOqvMQ9g
USIDz2mD4n7XONmlddEBipXhIy4+N8zTk1QeLJvvCdiNUrd0Ws+HBtXt+cV5VfrvuAiXEyUswicx
8mhNvuL/55EIfYKaqmZK6hyScrAWlFohNyB7oU02DuBadk0yrhnhxHrQ9RntAzYs+NDZq1lFaO/m
lsA1Q75tyMQlq+4YJJWmwlmXVtHT+RskgwdJRUJWnSG7tks/oAtDWR0jBXCWena3lsdI8NR7Qkfh
2YId1DCl42Wl/GNp1VtePwJ7qeyl3RTHBcDHMftFAN3p+JL6gI/8/RpfxjrCtEvnkKtVc1/nNKf/
07AvhmbzYG1dIhFbIgpvmYOdgqQApsgMNjJ5Z1gl3iZI0OV65pWTp+N2bhMp33dKsrqe1Q7EgJjp
rkvcMmAP6yK7GLhQJuyhgi+zTfTrrwdPutzUKkVJ8cc6qQysXNWEqaLxMcV36+FLbSOxBMhrS4Y5
3mVYvOpXCVecxbyuwuO+ryPSslImc6K+rEJmjCx1nEHg7dj9lb0ULOlF7TwNscWdOpZwibkTQblw
lnlFlYXOaBWk/Y07PsSQ5QsXzSOm5kWksCuSMxpdcm4+kRM1O7z7LrFw+UHikZVqOxer960rC+/8
P4t+n7pPmbqerU7SiKpRERZ1ibeYu4B7qKsI3PJJc6qnIbVzrTyKZAh2n1dW68F9jdo+/sCuOprp
DUcHhdgQ1FB7rn1pbs4DokWSLmS77oUNJPOKXGKf8wFmVKZpHHhosn5kLOyXnXs/BH2GCxF+SWT8
LLN6G9E/aTJHg3V8B2Qxla4UZvb4P7uknTFKjnkzwmYFWIdbXApeUFbSTzBBSVfOz0YUzTn0Kllk
l0+LhxizW9Ot62z2lqS+soHBWHUe3PlOUmDc869UFMylGj9yjXpXKLth6tXqNmZw18slw1btpTon
CtoGajHa/mSu7e9V+Ou/5CXW5p3/k7DS+2SBTaXB0gSRA2cjjBfBwDsuyBN1Rk3Hz+PkTzE/PIZ4
98utdg33E3SDID5BwzfupvQkwmGgXUNc7Yl0ILN2cHFBRgxRJoY++0HUna5nS3pIlT8bZd4rPVN4
WEuXg7M7KuE++XsJJf0rwmuwjXB4Mgm97aLn5P85QcNEwqDJ9FQaZ6FQ3kjwvryg6g0LRR4ZfLqi
kioTx3M39Aw4dv6ktuH9AB/0F5xB80de//WoxXoKEZKxILRzewJMNvgxX1DKTMa8Kos1EdfMfolR
FqObbYEXG1mcIw+wGeZQF3AxiDcNy76ZHhh0CiIWhEKTpjZva7y5yg9/c6ARj+t2lpXnWFHnMogP
qEj9uO9KwT7yqkOwn1HwUSBBVX4e2z21qoP8AbrgtSVQywbBRJXhBqhGANkWTUEPvZVeKcm1m52y
sVRLZSqcA7b2vk7AwqcWTlQARSTQ3D5/aKeTSe8FJAJBzejKUYghUJTEOrAiPby2tkxAjpfRtJKD
QHyQh0oLJ7e19T8Qpmf9CSF8w8kESXK1NsF5sdos9n1NzYTRriW8zDc2VnAW0h64lWpx1LBKfhWS
pU0MX/3TV083TGdlRt+mRoNBMbgzZSp2ZpxABpm4GCcg5PPLKkb0nGrvqpVIUzyAH9VIFzeKZAGY
AgZmdcWn8+E9mR2Y85hrGoUpfL/oi9Py1VxtYE/NOOQh7YWezGSEngk3fyy3k58UsQbFN+hJsK80
ycxvUJyN4NNrsfLfKrx5dT9P/TUh6MjeVAeIz1hgP0MGYXWGQvSWvAuahSzDTaSus6cqEiw01/7S
fpQc5jH7xaGbls2GXsieKa9Lwo928N9M42XdpCMBkAUfrMjPHI0FBtxnHydBL9flJuvbqNN0sEzU
ejQSVAlvhDs0E6i2uV+PeOi2Wwp6MFxF9MODojZCpA4lYvDM22etJIQEq8muiXq5rTphaeINXnAi
RM8F85HyQ+yon7gdJqyY77v3lcmEWqjSy45nu30OX6EJOby9i4lcSGPHZ1pCLID5t0qdLsrSVlLI
99qL1FtlLEBaVVmKAomsWa17o5Yybe/AfPd1m4F/Qm0X9f6rKG6jKuFEq8Px8PdO1FURQ6SYho08
7UsrDXBv+g+KYwxkKc53lM6Xh567UYWr3xRuZZRv8f6snFY2LuOjKPDgEjIxs312/k0Rwat2PtYt
UmxWtpy7OW8c8xryrjrbwBWuLaAM8QT49jDMc1afEyqEQepY0FgBlvRAu5bIhDgpiJbOyqotjCdR
6ByKs76cngV7fLaQH4qtInlfMBPYtFMupFqUYkGxIcdzZbkQLafGZQcZqLQibuHAXSAGBhIE+eka
r8RzsZMQwd/aW3t8pawKFWxQj9qBulUJgFsSoGFmrUquwMMBvvOYOTUXVtKcT/1j6tIHYOjEqm8/
viRRK1x1KAiGlp1W4DDfA0h/CEcrtWNhJLMbJr6LFrTVeHWyYdXW6JlMUXeIWfp8QBperiukGxAs
vp0YGq5wmMG6hodmapq/gwaP+eJhii4cgXFBGx3ocaMW6yGwMlqxV2dSabwz5MS0JzL+ZpkCv7rT
TI1B4qeCN/sOZXoAh0lBt51e8qrJ2tydHQiqKTA7870HunXFp5/0iuawLLSvoQL0C3rJ4maqUL4p
wrxh1nxDRfp3E5XdnDLr+q4JxDX4R9PSa3r9esZEIvRjlgDZWEu6AUOu0OVTeR3nOWvo3GA8vDWZ
hrrGTxkI68CG5OhAXClqaSDX7CEAa2XWnlDz5mUNARNPyR+O5f6h5RM4dNftdW+GuN55wr+Qvaga
P9d3Ro9cyxBVGyphvTGNR2wHCrAH4W6fiGbp+1gNL9LBnfnq9k2SoK6nvL4QJhlO3VV26A8u5xgK
qX61QZnwGbx8iVx6otTKN1llpw1SLkVAu8AhG0gtFKVqubVHfonNITJ94fGNEE7V20DTPiLuRPIx
e3MXkN6WkcrgNyZ9XybzBFu6EeWFhps0jUwblMC0ydCjVWNYme+0+WL/CSoRtW3YynqgX82AF/j7
PZkw7XDgLmZ1YSwcqj4NlZFQDrKkYcnl5qvZT7gOA8gZxC8o7CEzPrCX1mR3zLr2t2xmrB8ZL0C2
JO8n9uzedHMef7lh+D3UudN06NtBx2/NekiWBeNXTTLSJKoZNBknoLGqt+ILo2Jn1cX1fKbw8NGy
2Y8w3iPb1O4NWSxvoALGrVIyQaOznXFarkCZagANcox5KwyvBHXVOx9EXHYceh1BpHuxqCqGNLCV
rXLB3N70H7O42enMmGhNvGjlxKIetm49akUQUSH78J8/Z0JVbKUzattJIAxiS5nRgHUI5HJSxjsH
B4fHDVJYOP8oPJ39Yf3gfiQrYdN38OlH+Cl/FYS8+ShiA2yWBHGIPhN9sR8i4KGjf3bVWb86y5fR
RKXp7rH/ym8m0qKtMX4OnE2DOMAfYkca0msUMeS7H7r+mWGQW0xx4cJnJ7h3abEyuaQbZq/Mk+rd
vod7s6VRPNrW832HvwjRmF8gmjg/G6vidzBoPte/mkNGgOCdBhAg5VyAeGNMK5maFtEfRcCnpXp+
ObWDu4RcvJwgVhHuiilYiAD5sbpr8FlfwXjYLFW7jRSZWoHSdzYBa4hV4aRLc7INCMyYro4dnC2o
4iUhUg/HajUo8YTMCy3gxs6wKE83Wz5MV8UWNUkgUMxBtPV23N9vY1t8OB02GyfhxNnuGIReubkG
IUKJiSfgO7S6HmvCTdg+0RypObLI22mivPlHDCm0rNCIcMhP/568+zpuR7DTxwp9qdq6czbQZYcJ
ll0mVboTxbha6ABU44MgF11c5G5qtlWiS62UXH0zTAdtWWRs4CtMEC4iFxCgDPKgc+0ysovISwEU
wG5VYQm5fxHPmHopA9YFbCalnw890udNDrlIRuoIGGhILi5JcvbOpx574LalYuuZpXNlDBd0WA3l
u7fsfR5RvmnrnMTCZjuaIe1uNhrbo9TbIIyF7oNpXbrWZmAY1LUnaXvIn5i0kuc6Dwg0DMb4JVKe
nRn6VseE4n5+NSK1wq72LuC3w3HjQwx900rEfY0AGlSvvQoEDHczeommSL7fCGYZnZdz5Ui/KJuq
EtyTXiR0qC3V//Wu3pCrbUp/tVgTzF+T3ojSPRabki5/xp2Kg2j6NtnbcrEg8QWU+F0ftWWtiaR6
FtBwmnddH6kpyPQMMTOYLKsVfwBPqyMhjj0YfoD3D/FxwyFHCeaiYYWkGUACbGhSLi/vUtsyjd2b
KMHuVHukHZItBbyKrBgflxRV42cSKdppt6WueJNww6m6Vl+n1YdA3KN6lYuuaPJQNv7VGX1csFhV
NbnuYSKcelrknyBL691IoTe/Doo/ENpBiuydwQ2YpgOENjpJodWnnYUGguZfno2C2ryQMWkWXyt/
OsBRrbXCS6lCEeQJcpr7nmRku4XlQaPdGFFAuQL0q6fke6pEAEXP+WrMlrr4rRPUyDUOuYUoL4pj
BRc2EknkRk66QqHiGEqejdhpgt1nWaCycc3BXG/vkhTftDwjSdjVGuxpGgZrL3yqw+wlAR4+vwp4
U9/FvSYG80R/wORptiWR8RDYsc6+IT77SbXTX5KAhs7q7IijxlZ26TjEiWuFJjWbgY2HgtI2P8Fp
2AM3rOsuxPykPTasnJg0bfZFoOmCtaRViOR0bcKNTtXpCwK0PuKg0b4vsQQAUlp9ucAPsuSywa+Q
BGjl8D/e/4Ujrz6WTqdXUTtz6L/2GNtZqUNrxWTUN1JXjes7kLiMjSyRaVva8ZPNXBkK9pdzYMUA
JcOxdLgK91IFdmWtMlw6ZuVWAvJaaOrnxMoTjw9gdTok3L9z61bRF8Zmnx99epfZdzG3mjw5TIO5
0BihcSVdKTBdciRXgN/sT7UyU1+Yt3GNvL6EBLHGItOeAYkacKF0aRHiGAnOrJAOfKQ+N1WTmUJh
fgYDQdnBemO36O2A5eDxeubkDWyJX3OtH2iwssrmsitvyuqVL+LkwsTamYOTa72DwVOIpNYBGYvd
h5H+f94Lhi5No8UfY5U79QqFWd28NeO6bKuDRy+uXsBSsCp6q/g1vj0G2I5dkmiHY/nOaSRY7EML
7YtgeVIbOQzHCeSXKXe3x8OXK//jyJb9Jom15bKSE36krdbYOyB7Vz/ksnXDYxyazPdtBDn1O6pD
s37mKbyVMUUrczo8L/d7J6+5LpKlA8BI0EGtdGBKTFoZMGqnnvhhG0uosVs8Ga54JJkoIvBevqgE
CGxKv9jQMLogpX2204jyumtxk8VDkP0tYcxqS8bdmH81vnSX7adTYEefjjvIzG7mRxKaUjZEzjo+
EPQ7V52efVPAXgq1SVxhU7gjvPJJPci8HpSjBo/TVBF11xp/ZKMg/oc5AJZAdVv8tGwIOCQP83W0
QhrDI8S0DCBEVvklq/PRyLS5N9/TqufP6waCTP9xw4Dt3IVNm5wZE017KalLZHKKi+z+lQl9BhgQ
Wq4/YJkI/h91m7NwBovOQzh3mz+ra/pYjl48pioyN9vpcl41UW5UqcEQYOrx4MZXRwV93USPrZ8C
+PXEynyCtp2ml0kO20dfxYrGkXqYsXyH/ULAQ5YgD/cZuQEcwmJUAG3EHc0LjE2QdBjZLTw7fImN
Zs3oH9EGNKC6gumkv/ZCULRFGUzzPo1Uo7zS/+5qlcp//zmDU/yBSEXv29AYZMtsSryKujKl7Rp3
rtoe/yUzihYGmKxWIBRqRc62vpxIBRNpfdhbqxZhA72a9Z2nK8xRR2N+TiZBOQzDvmDKI+Mw5N5w
Eycn3d6F0NrF4BwoH/9YnrzRqgYLfYbABhtiuJGqnkVVs7ubm95fZpJIAIi5DAEb1zHFSCeGOz0B
EGGnqji2qv72crB6Vh8MDJShXwyqVst8X+26ULQk0YBuOLOcX7RuIS8X623O3saZJNgihtpu7R57
Hfy/5NBybuLK/K1QPTCykoK35elBDf7cgPFk6AENdorf541DutAePXvn2OmyCR94bV7xCrWKkiBk
QYVGhzCYR57ERUgKfn4GBS+3MoPtilQS+GhxbpcwHPRFN8DAmGW+geb/mRqvilv5tlMw7VBtu0Fm
EFSQtMTOc8+PWeZll6tV2u6o4fFO6oW2ahtTOMlf1YsSLKp+hcxIMsDv+AWRuICDXIAhkf2SOYak
hHRu+X93UfLDdvkBjQySk2oNsh3sLNGJ9wqHh+8vjuYuhiIcX8ULRL2Aj18BDbeK6Y07RqPLD+cy
dGqgkf/X7001kpdWrguOgNlADGQiba8i8TVjZ05rvbsDS5UAyxk8n39Llf+qi6eliG2lFHZCOzxk
z1RSxl8GM/1sa14bSF2dGVQuraXQz4ylCNshN6vnrLK6nFtTO3q4axIzeeuW5N/GIRAguIefV3Ep
G5F3kmxlRy74Pu+UuLA9H+xt3irMioooghpd2cEazlvtaWp/gzR93dzHjRy8hfnwWkyTr+Xssxja
E+5gxwd6fR6LBQf4+Xa48IK4rjH7w3f+NkS1gfb2AiaZITDI9WN8HgmRPI4t0At6LpVEXVcHAUFz
1tWiExx6bDITZVuNqnveuW9qiKYxr3XMUapTIk15voGvNfsvWAlExgWyBLlZbwjDrQGcJvyU0zJD
0Brqwqvo5+UN7y/bcim0FqKZIeA3sRME+I6WFQ1kEJfK4p3xTIX2bXUo0ZBOmeAVRQCyqQ1DQfHN
kNlY1/jvvurtdIe5i9nGpUtkxuML1L8TdjgCeWRY6rlxWO8Vqn6u9tGvtDSKXhjgDDEMqXlzjlXS
VPTGd9BMNCZrjPxXKiQ0kxKJ1vQnJyCyaV2J/VsT+6T5i9fPTFtnGKGxyAQ+BeNTcv3m1ONR7qf4
Th1oKEEF5aEHOy1wjkFyK6xrvbS+o9Hh98PwbsxSXEiUDRbvC/zHcvCszEaHXaPTwxLj0UhDG3GG
iq6PKkT/ZspvYy7cKKJlhBk9SB3Y6ggcwNVBvyhNtuFokonqjLn8iK2fN3EHQUTr26e/RE4QtREI
PovJbDBXqQkwimJOzHrDO4lXIFUDexsMbg7vLKzS95fBU/Vl48DHXfQkXzOxHVa2cP2mZDSdxGQ2
20Rh0N7BjGZ3E5AxT8J2JAHYuufRNBF6mb8l8mQuk3A3U+SYUAyEeGFxImbbpLW+n5f4flWbDthb
L5WBx5l/wJrq2tNJEF9ekHXOcKDncNfyd6QO3258wXUCO3L6gDuypwevX9ucCWXcJ4fRxk5iXW4D
pZvlyznNSmjicjblT1+nF88DAaKpabal8rqz9Iix7zOLS3ADKxr7C++gtT/9IByGPwiQ9ldT/tX6
sRhv7nwvacJEpcLzBojEyUZ1dElukg6GVxASFNM1BU4HM4+tq1bsrifiaNUDusI1QmGY99QLIHtY
woSTUBlunMDPu//Bw+LiijryVKEAf9IiUJZpSodbR15PLqeIz0Us5ScBhw3vCK/gyVz8Sh1mU9Mi
fwEjxM0krW3phItuk4F7PqiAn7pEpZItHDFJlhDkEvZ2iwKmBrpPqFi1qhBVcepqQcGVXgzsYnrc
2MDnF+DknBrfHsPaF9JF3Z3rZqigV+LHNBEl6+hueVsaYMDbX7y9bS8JlNhRA0ujwx+5vWvWNyY3
833i4LAk9TRm2IFMzeYsDyWFRMfKN2KKmzCFddDBLHzb9P/OLe0Kb4rH2xzophHnbbYiFA56GYo1
c6/170wD8zQtgtC6dUeQE9qFLgCSlX0HEC07XrYMQyMfagVEA2lOYiID5r0MuCfsF7zqGZhqOxF2
IU12iButBISlmYO55/Oq4gTchAMNiSqpDkxOfFkqy0RdgnfuTkcOcJMV31wp71Nb/ISM72bOaRls
3mYA11KaOjqAUjuQJESnL7QqxZ2PL1ItK9t6zlOyleGBe8lZVS0BpeU19teoJTkqWyq3hUZeG9wM
d5RXJICpU03RSySM/mShOKBGIMsOwklm/4BWDh+iWJXGoo8WsE1KVdZIOhn8QDK3GT/PXsxFVwHP
aI7EM4BNtqqXUO1N6sqD/CXcbBK8u3hT17zeBsOHd2rp5J0ojrnaKCGVwvLGOE8rGql5UgyuDZSg
KCViz/wCtTgRUrJx9iVEMZviuelPHady3vO9L9VUE5v+cPt/TrfS24NNEMdtFsBLKhxk0mnokFZk
yU/SlE4mWe45CKAENjye3ibC0zkaJ+O/2h6tlXXgDYU0g0cJD1TySeWQ5QrPXUt4hhhvKr921kWc
9W8XeC+d5b4UfJNFx37m/wauU0rrymXWGaODiqFdalc9YHtqb56BN2tcKFX9RDyNOc/K+Wqm5Rlz
uXcuGTQEwJiUwGuEZgudcHzgDSKP+oSDm2ZFZY358BFsGKZxxCv//QDOY62CjcvEg9X9Xy6ZR+0x
u76wSgOXOOiyxXshpP70cCavXxTnp+mY5HdKuvj1ttzV5Rx0IFbU4UktkzDn19rYpkRcTivji4BF
L1vEq1FY/ofyZXj6h2EsNqOULQzIaDq20rIi6V4dVtsvAfJPdNJSUgTEr7TSN963V0O2Q5yc6r8t
UxN6GRGvyhNZQmr/EepDdFvKbDHpy+nrgOIJe6wp2MRJbd3SdKcLLAT4vVz+3V+x8tMPRujyf46z
ghEw8oAYGB4cG0X6Sb45rZrLz4lTd6Ar+jMPvV0ADPI9JXjoF9hDmt2o199ZbQi95+28wy06BkXX
Nrwz3g8Rw8OVN7p/rTcPC3iVC2SFHvit7f0F73r1aIEASpe8lggdTAul3vIcThFBPVl3NpYP3xip
dTXxRQytwKOlG8WpkMRTqaNbEsaPgAz0mBz5d9MkjOn/d074q5819xA8YIuU6mUSdn3c7uvm1e1w
c8+hqTgo1RkMPM6dHvUVlWq6qpBoTcPoD5V9RV4iX7e1hJFlS/lBOgDAQWAVkS7G4ylb5kKi1Ylb
dgRAe9u2VjqsLWQIRON2UVJAqRAUd3UWdYT/kktNYjl3VIIDv67DP81VCkM4zdWP3ZnHusCVXguu
iughACnX8AIPMCq0HBEniIwj8LHhdO3gE1JX/lyuEk69/f8zYUVxFcpXwZcI05gd1xJXm4TLb+eB
GDzqTg+FQGmuv/iT/Sp42wReD+PM8rgjI5Auxt0ak/QXMsiGYvuYO/Qs/o/9jGm/ZV6mJZEMMU/n
zl43ezFdXMwE5gWUR/WvVh2Bz7OB3gZ7wbjgDx3RyXFfucsdb+hfrMmjLYCUjB7IdEZOrqCnX8dI
4r6ty1yyzhm2rc/qcmKA4s1UqFe2Vyn0ajmZLnyPP/hf4IFAeSus1yLmM8A1GcLtF6H8QoZWIBj/
rKNJ1sNLyCiItE+LZ1mzFYXl5qxL5Y1FJa+J/D3yd6zxpopkusSIvWljA1z3stqm3Phup5fM77fe
EhThQfyg+kXJoRlG+If3PkSipv/ib//i3rAIHO1ScYzm7GOyObo/s6XEYECxW4vE9kcmXg2D4kgP
T5CvhyzYNSvhU7jAC0ZJBNq55CX0SAwKtg7fV/qgl0rwJ95yJve3/eI1uKmfWuaIDd3ZC+1Nfsvt
9yTvK273L89RnJkWlJbtCuT01L/XZkeQRwXX7dLmLzbtopL1XilaDlix+2gsjQT0tyRXFMzY+Xn7
GrQrD0aYRNGFar9qy6328Odczh8NgdhrIrVRoymxn/zS7NZkeS5XeVGXfAETCK5ZMe6WsHqMabaJ
pC27R9qJLHm8hb6siezogvl0Wpq/aRxFa1U5AIhlSZfKcW16biUU38foG+Nj2yBM7pENOG9K/eNE
BW7r6ub+IrI8uLE4Q7giLXjmBjCOsrzIIB/tGE48Oz/FquwT8Llkhtp2ERbAWhl8jT35z6EOrLB9
Lgxydh8ymP69qlF4nz6irljI+ubrKJfXmdp2LRPt0QCzKILdq38xCTtq5U9M9ub5B+Ug0VKK0VTE
X2CNVMmzoA/chuLvWPt2NAvb+g/ba6TgaO+fTpB/ToBRvGoOZM3WVAAeGA1OaJgtFBAVORVwpt+M
jfFE71c7XBVEg0gXH42VXK9W8rSqfzBTaAoYscjYmK4NGS16+YTTeJITdjowr82p16cRM3vF9pss
1mik5P2AHiAqZ30XUkAzrayZ7jJnmMAe8AaLm8dL4zoNUUag2QFv6Q3k/hD/0QbbF3zqQterDRmX
/9pmmj80/LZh9ZBUMvHQff7kmYSp6N7waIxspVsth+6qONU52diyk3uXEQb42xJJws474RCFq3E4
D1fj7KxiBuAz/0Er15cye/kvtvZm3y2Mpk/KTYP7K4tLGI/9R2lvxsd2z31DA95S2ttwIxP5dfXS
yEn+qaEBArxB/L2QzuKDB53UGjqIlua8hxYoVgTl4qbwDip2f0KeD9DJVLhRIaUyrI2QgJlkQrhC
O1zohu10NoLhZ/7+Xzl5keXIrW73+vLlMHgL5RSaaqkOnin/RJ+cyH/mOLt1jY+iKHuy7bH8XFeq
XkKGnhRmpuFR5qS2eqCmoWZ4+RHHjrEnCbiA5bYLBUffyeJH7iS9djmWZ2Zhs+5ISz5zdD3pxVsN
+a0e6YANSeSCXeTZ3dcdSNP/Tyj4epodwhbZRn9d0EgIHucg8Pnm7i8nq6L+VHAYTsBx3POnbGmo
lXfM28JgZspG7omc5fCqCesag+iht19cA++LqIfbBmbAIGu5XFLxosyg8pCAwaL0IIXPZcocVoXy
u4/37tkKAxo2Vv4Y7ufiBCSHxgTVgN3Byu7GNgRhEeuvHhTaZuCwwHvr0Tc22kgccgLxROC9yyMY
TonNG4uibeWOZ51PGBClV3vq1uuHOcmWujhpqoxNGIqKINEdBMu8e3TaL8S9KkVmzlcEk48O57so
Kn+rJ9ByPUl35aT3PMhfAHOqYkL4feMQ3iVzbnzkzgRXw3lOZNjmSs4gwjlIHPYUj+pGqxZrkcqF
UqKOThROTd5tnL2dy9N9MzvrQ/hWo7lbPfW+dNZHio323vEKTR9sTHa7TSR+kJ3xAUdQaCuqfw0s
dg/dARMgs0rPJ7J2GnNis+6sWLDEO6EsOT0338CRpmo50M7pybh16nB2HgmoMilV5szIUTBpb6F4
HQ/XB8bsIBM3GSmpaWcWGTxUdPJtnh767xxsyd2XyChWqHpeEs78CNLO65iv73K04CFhXPnu0ubP
vtu2b18+qdU6jYaThpbcSg5R/HmnOJsweorDSgNo0uzBQppyvucAZhoZTEpB3TSFJ57AqQCSbTmA
3r/KwBUdEg6beXQw2ISHzrs2B6ykSSxeaSBTRNZFAD6V4mdk7sQyQCURw4gGUuRdflcZcaezABc8
dCWeamZUymwyKzB2hHye6/kt5VY7a6624Jf1FOULEpcQl0amaJ/auUBjfrIzy0oLgxB6MbDZ3G+4
TmlZCQopJYURTmdUKwiUPWF4Fw+m95CWjLn168O5gppTmTtUAblX3lrCTwaQxtVfnAXSDHnAgPsq
1tv3CdJmkG1XrIDfGBKFSjDbpIZw3jI2n6bHXEv2Os8EuSuIVIFzXaBeMmBR2YrUdoXd2Qk58Y4W
mKR8ioIdKaadE/boiqIHpEK3bxMiNHuaycFZG4hZ9XHJ7OVGYorrVrxv+JKQhkiySUb9kEOQf37/
SpYx7fQEnnXQDIWnohhbLBKT83qibZqTBdMCkabFh3B0K0YCIVzya/YyeuixmHpWCltyD5Wlmgm8
XrInxhJSE/mBrHj/J1de3109buB3yTokJVYF3jV6rF0vO9mOTR10IWofV6KsAq3qJBtzKSnixpKz
4veKVmy26L40KggtMEmMisoIb15LVc0Jr7A033XlAQJSyxd9NbCwRnDfCx+bjtO7LLJ9ErG3C4pb
zXmTdboOCKLvMt6FHVaS+6NcgLqaL0RPeOoriwsaVBTqLpusk1INb2cVKhLDLt7Bms93mEfnAoVc
AOn4esF1SeGPwOXee/jGh6TUXJlzb+MjJoT7+Of3dFRvxqFCT71Nqik0ojSCuZaA6Sqq+g1crq5c
VnSa910bP+wFpjJcuUrSXV2/bdrVVrkr7tTq+6u/J9eSwYL6suz9Bz56WnrB178keXg0ADMHxaQk
fzUna5yiWAHH0Xm5K4rsFQE5hPXFof9Kxjoxdl9YiNa4v/0qu+OstUFOSBhbN9VD7uMqCB+dvwAx
B5JCd+/5K4qtNiedjDgQutxFSrrcyhDwyAI7f+ZOod+v5um8UbVZ6rve+Mov3719goh3mZ86HRKS
6ZHBSD1xS+KI3POFwAAKQZ9n+HmleFtu76TAopRpaes3Um6+ao0TCU09/9GpwPyybqUCud+fEO9+
MgSYDCv3PFsx7rGlSyiqf+EpWtghqAQMrhVdW0xCZ3EJssas5mY6Ojl1VweKmZfa81t5jYGzV0jv
zR9mcfWR9cOMY5ek4aWMKBC0dXyZKXBnRhTOHZmUX1sDgbIwvQsuriKsi984MfFdK4hkd3xs4Dni
XUz09sbtZYNHBl/WnNOzo2Q/elXLQU8NfJDLFDA7wwhQ25YlcuDaO+ok9BJgjoFrl4JcK7z7YwAN
hyxEhzIY3bFlVsWZFyYqZ8nzckcAu+FfGGQBYJcIP6PetEO9A/s253ABA8752hEPNJ2YJ+sLaIHn
nmNQXdOf0lInbFv6dHvj7q0A2iFL8a4ECrCUz91fGHHE4TFmmyBH2hDgWYJrcmwgvVSGV4A4kJBg
mYtsdyxskUKOIwXP1l147nvfY074suTSfuMFyCfGag1MfGjMDvxnk7slcIl4wazmFlRji5VH43oq
5oaKlhR4ktxpdH5VeGUEX7tUkDCH/zua+Neb+xs+ka6HrboT71uA/UXAVmXiqy3vEdbqRP2QCJai
2npB1Sw3iCLKOrW3J54vs8/5IhD2wUfholJGK06DEPy+oQ9qsEddiy8qd5f8AykLHD/oe3voV0md
H92/9+/6DgQE/vbrB3plX5vSMcWKv3ZqFGsZmsljL0Ly8lsctY/NjdfOAnStCo0jMQRDkJMO6bJH
vFaf4RMPwnYm5UQBP5bBS8hHi3X1qIaI/Gfyggrt44eo4kpqVBTLic9egB8rs3QJFXMxJ6/bGuvA
mcNdGJO7DoHSgqnz56+NnKqMbuQi7EhKaGocGvt7MvtImnhtJ3CL2/bPYIeqdjHtccyR7AqUxESE
Vj5n2UrzGmGiu0MuweMBpJfrRhB38bDlIgY6Ao52d+fUwVVK+oeC3m3TfzZXNCUkPCRfuxf/mFsA
jXmfcZQOHSrBNkl1BaZ//gIseUmtQqXffodfUaE4bozS6+TNusdY0IfL6oFupe3lm7+99ZlHNJj4
FTuX8YrrUhsOcrd/GN+jpQIet1EK3sfbM6IhPIIUDKKnnbNw5CPXoUTzDDdCBJvAX5wwml5v9are
xhV7t/bQV2rFQHoSSOTrOqxmsdXoOfn4+GIiEMjAVDNfqzJnV68xFvQxT4D6bD1P9ZzHnPF9zW0O
KRkg6wbtBm3KRD6fd++K8eYEnVhqwPKGjC/8LTEOXhKftgdRlAcfDeRQGMPY5g45UQhdrq8M7C0y
1Po7/lVA2Oc63yQPtpsk8e4yvYEqwybYx5Xkl6CY3Xo+GWm8u/ab0IgTc1qvyDIc7y9DGch2l/ka
dCWmyPsrz0PkYK1aAzY45tnWxZbczAiyqq9vmf7Qzuw1bqpuBYUdiBrxmAR99n/RAoXdM8vB6s5J
Pk0z+LC549A7fqJPaq8faX3VZmj9ev+CM+qAJk2Vdpc8GvT1b4BZGLvGh/XZQDggF3V+2/jb790s
8ozi966wDqHF1c58Ogt2sa8pgj9CScj2ms5n25yjg1ngrWhPNQSAYlGmkUuQfXzzHQdQ81cCNUEO
LPEUc/3gcw0YgBmHT+0vmaiP67W2spWu7C9s3Ei8tAuaNz/b9e3lXPtHXoQ9SFA8zpYg3MzXv6VP
/dUko/zlFVVz17bJ/WaycVJCwaNIADKNd3gsrO+Q6wkCGZ04vNcmbKYrzATLX11NLrZpTRnhwTDW
E5L3WBuAws14lWqLdIMYm+HqKYRJucMMpR8/tPp1YdSaszn4LYnwR5LglzALcM2scV+vyD13xvQ1
PVoHWZGTifM31yQmfhWgwHT5WoU/FaTE2hcN7yvqQCrN6q4GP9AZCnbtlITr40lmtNL3kL5gDWSb
NUn1YeaxlJjx7z/TRUGLA7D/FovIYe/EYIT6bIySnKpeYRtOPoxrL8+YJL0mrNbII98mKost+aED
XSIBKHyf4sYjil4zUa4/mrKxPtoBK56GlryslkCPOdKMuTKOotDNmk3lLOu5FEs2jxLRVJz5ddtp
FP1pghOQHUVDxiHTgtLVrr7AR9fMoHGzo/XGFT31WfcQs2gv2x7KRd1YB6CnASlr8GlIwvHp3RyW
c/S4zOg5V324K9UAZap0m7pB1HgJPMW8oJNn+oKfpll2J40qggPNtLrUI19Ockxl0IOXw3TKSvPO
v6OrYe8o38w31HxSm8zBTNRN5dNYll8ipDIdW3G+NuHhsFaj0U2KSHBt1Ea0y8YR7UmHUOMTMr/Z
CIavBIHtMRoqs2np6zHm1hR0CULi2fcBOT/QdKt+KCPJclt1QZ6BxcCcrqwKR7QEW0+hwI0TXOaE
1kC91L9tebP/AqM71fvggwsvV1NAJDQy7dIn7XyqjujHM44k/53pv1xl002+s7wUczZbOJPLKO6Z
sDN3HIhDG/cSl8VuLRahBFlpaeRDrZZjSituhPl91mVf2WJpFhFvT5nA7v4VVRmRu7QvHXutVUMm
jex5qoWjRSmU3bcD/FR+TQPIb7QaMYEDYr8cGFi7CJmvZl4nOWycyggtcFMQBKKlEUhTWPrK4fnJ
T/4W7ycQpMXIieJMb1tV5XeHQRJFbwtIbRxqGa1hDAr5kbF9T6uXJaXzo7JA37KZQEA4k5VCDAVi
cKuzXAl9uVaeWMxut+2rqf7TZU+T2bwBFITMbDzO5SBQ1nD4sYNW7W4p3LSTvT6BhF2tgQWtLyhG
sSXWzkh5PjFwyN2+4wjF6UHJGP0vnQIe1Ew49H8/j99u8gvFaPUKQHrzK8HbkxMYADFQWJ1eXL6h
syNpegB1q6jLUolVIDXrBSOkvf9n4SVCovWrZzQnfjEA+lG6zmAeU71IQzJhlAcg0/1DGpQ9yg8U
MoiCniXLOY24reL3XkXCbkLZBevgwBl2onc7ThxFREa7qC031kYpV+SudCGnibJhW7LJK2/0rAw8
xcH7BrXYHEnMUcyw1D0KKKrzjvb9LGHEnw9cLn4tWuDKRv7+i/jHUEix61yvLoHmqojkRgBTVCr2
JxNR5LuZoaTTJXu8B3tvbhuyOlw3DRfrvzVB9d3llu3X9fBOdRHmbgo7D9mZshIoCSoZ7+kCsPEb
Ia99VL9K/EvydlPQgo7w0IliEuHIuBq9LAq6cC5REX43AVRPkW+4cJKiOxoDESn08Fy4lUcClrWi
Xp5JiYBjU9k9A6Kl19Nm2+Jb5oi762kq9udYUoOPAQPQVI44vmGkJDPdjw2jfn82gT7jRozxrpmW
3w4Sj2BRVdI0zz3/2vikRj1+kn+nMmweps15U1sC2no1Vc0aZBpaIQDHr/cG1ka9nEm9vvbtnLfp
MgPWFkpMAegkFjlDl9ZOxPs7Qq+K3eO4UrEwxs73ObUG5ooG1rJnQpYlLWWHUqeO/SOXRlM3gK6s
WLbPzdldl5ewvUV5YwfQ77wVAhcZzJPkdDbduG6u/pRlyPhgALkD2eMA7UrFkfEMLfhV9uQ6umLy
bWBzUyWHsast7ZJvoeEqbuvmPfMxVo+KzM+3Vibu14TVAIFQqHldq4hym2rNeyESQW9D+fdlcZCd
ylfNtdwBEJgZ1oEpN+RV7GU8Ja86bIAVMXx6+FZjYlxg98y4BvkbdY8Yry3dTcAa7Fnz/HWjy2KQ
7JgDFyNS/RPdEVtd/dsPdCG6APHc896zR4asbIZ+Sqg+R7QeMS9jMBtF3etZ7YpFTMGYlAyj4JY0
H7JhiFrU56Ypmo2nCpFRodglEifXxxMxnw/9ca9ILU3W5BYkMlUkeHV8FZKCX32HOLmMvaOeYEdG
Oe7xuc5QXXTnJCcqtS/9pd8gpCHrBc6XjBmcEp7wdsJTaX6yDr+5UEZ8WDKTDmC06rs09LAG1xTw
Iy0dk7CkmQ2F+URUBjDEbuJL/xapkHuJ7AT+KSy7E5DI1l6jsFipJDZHP08EAtzH3lVNpq7QGN6e
QG6pZ5OzrGvAMdJZAIkeiyu8ceiK4GZdJGczqOEV5/ir9Cpfs0Emc5PHHYK7TsD1Tt8dCbfXQ5e4
HI8poyzTOgfGdoUQlp4UoaA04YEsWPW1cHP//sGsidhZlx9gKfvcpQZsIV+0bHuKjzD4leduIDID
SKQb6ynRRFBTVVRCaPcR/vXBTN/HIsoMAxXh9vZiUVBE9f672V68PpPvo6rXLd6wboKl7TfoYT5P
bGylGNkSLrSsfvGihWhyHdLPeUZmgMT5edpc+kQKGgblB/QvvEh72CogAbiOKSq1zF6oHzejmD+N
bVH/0LAcSKwTwFWsgTQ6VlSHEmQXrRdvwBI4bbWMMxNKwFWDKSH4Ip4gOvxBF4rzecqH2BumK2P7
XGc3zS42tQXwOvp3bFE67V+/TDSvN7dxBVDOP9Uetc0KjxqSu1zZKQBh45PCwFuWmdKbpxIM77/6
COdy51lFrTabmZQOgopTspLdyA61rP1R2q9cErkACQ6/W8hqaMD0NBpW8BNq8v011xppu2Zr+DNm
h8eOk2uiW1GPyDMmFZiseqHy5RguCc1rQGQ3YjjVKFSqOTmlIcuXGgGSIRhSuUBzuk3zwyYr048U
+6j21L8u7disvoYP2hvMSahiCa/SpqrLBcoaJXRV3fgu6wTy4YRZ0RM5hyGWnn7EbXArhhzbUg9w
wVMyBC5J0fumaaqKAO1FO2f9Pi1rD6+YerlMmmodR+kEeBY18dnzZseYFH07mAGaCrWbiNGcBJoY
BoHxP3O1EjforsNmXseFyvSbUkAvtwCbBqemFaDZmbRUP2lfiZMyi6V1+e+eM4gG5mHIfTzGThC2
ere+YWhGSbiZDj1H1GEVC7K/6o5Z9ClgkNgqUS6HTGBOIGyBDWEYmcpK2EnN31E04KT/imn7t6wI
Faz3oMSHU5fLZIKP7Z9O21zk+vqZeL7dEKcQki3Pj5xy36/TLy3qKg06srJe4OGFCAeve4+uEYsd
bNZz6cm4vwsDS4B2wfUTtpH0i44dB5TtkzJHgn1FzAZsJm/SntPUzmu4O+eEaAju3/i6jUAO8OJm
ItfPWCGI3Rkjfjsqo25CEUPLmaOg01lkJ0Zw3ikee+3mgellbDx/63k2GBDc297BtezhU6zksnE1
iSO4oQQ0QjVGKV3Oz7eYUC1gbmdja8iM1UPy3rRzFhyGzZy6Ch0Tv+Y57Ybil4eRo2Z93A5NXhq/
mmjAT2mNJCaZrFAnnOhFm4CLDe9W9DUHTf7oTCWeyC1eAKoBxQWXzyCNRcoAdKCZ+2O/rVGC7yb2
WhXOUj0VzbhKA0pPYx1lutPAcUDllgg0kxMXqDl+hBlJcCxNAZod3NihnTE5+GiH1ZMNOQ9YuE82
58+H7q6ziTjun/tnv7vnHAky9zwEhqotfxWisoZYmoob+0aU1iN22sZQ+/EF0gqIMmdZ9pwO7Vxo
LMHoWLbsxodE6M3oXT1bZVBao2ZgOrjzy+moolLGs5bnRh8fba4hJHb5Pl0XybxCxJzfdnM0INC9
3vKB/sgLkY7edpGEmhR0WoIFWnd038/lqR1rw3iVIQPwv3YXruO4s8O1OEpPVLdbfpfaPGsL5AGc
fRm+ZEXOO5aw1VZrjcme18i3SWjpcnGLlKR2M532v3s5Empw1oaSer5Q0NryXfAtVDGYpGLwVS85
FdDjPxZbIhX8IzL9F9+tqgtS1oTaYWPgtwa5RHuR0aQAMEKhgzdYOOOETMnDdNuKVNLLCae0pPtt
NMdrytXco46LiFLGShgV40ombDdn2WiOfiGyBvJ7cOwWAXFrNb4zx8UrhEgJn8Zd78ocBlmiVw8b
Fiyn69AA0mkHO/wN+3Fd3rVsfv5kNeL1mLxMA+sw+c026rqii2leq7HG/1kMfenmAo75y9xADI0A
abSZ2BfdEqHe/taPefyP9ScI40s9aW0Itm/eG5j3Skf7aGgQHUpUf1UxiSIqx81G+YHXSiRF96d0
/tf1iXWEQa85J40oWodgvwzjXVyhSe3FqkLVcdJFE1dhDNU1WAvTRncw5oNh9qpiQDCUsMG+bU69
fbDKFd9gC+vsTHw0yU7wCC5p7MpDycBoKeeTJmM/vZ8IlQJ7zcm0MEiH2RbOnP7s2kF4Hz9SfWC8
/6PZzjILoKwjKE7TalBKpLL46GC98FKGU+Fw8C3AXnYYUBPwBq9KgxwmE+LMccG+4JEthtwv/pJm
TIVH3grNC1B6g0e9wphfC9dbwqUG+A10EJn+Cmco8f0Qx9d3zjxcxnHLD3Sf+E04yAJFu3mB5pPE
JWnsxsfSN1zx70Fh4BoR3Vd7qgrKMRJVbsrqBSwFHdvam3YsLT9GeNhFi5FO9GveXQgeALhP/TWe
ukCOhL12W1rNBoLiHynVqUntV7SoJMZretrE/Zc9QhclVG9dkdl70SnfyJkKrI1NPmo5xchtwHiS
qTKGnyj1OXtE1kqZ9kmMnv4/tVLR/ysaVAHfk+pDYw7ZYNvSXAm/gn+6Zb5itfWVmBg7UBlkjoE3
8FT83lMi7MYo7JRqgHF3tRQ4pNzVW2bGhk6emMiqs7ngzhUS+8fP3fDmcnsG55qEU1mW0c7RNiOH
qSaJ/oIiEUKDUTtYFpoEq+WAenPppb6QGnsiO4r56Q230kIjb86bIhLYAlBpMDm3yHJa+AKaNwWJ
WbKMgrj81wTEyZYlc3hII8Wx8eHcRfvHbm0CMU4beIq/fhPPHqsiWjrIicLyux/mgdkvXmGqYk+X
Uolm8VqmxINE0wN6MhBk2dgtDG5Lstb3fp4fJJHCvy0RiLTTViA/e0VoPXwYJkwJzIo44NISZ7cv
KlLUv5+YiyxyHemHfAbpFSUEopEl9xICA+aSyA09zL0c05asxI+2C5AThY+OOa7QPdRETLAauuTR
Yoyrbw83nGnpq8LSkAtivhwtiVk1WepIIzW0/xt5UfEFYdi8Arik81mQcW+KjtdX/hK8v92QRjrD
vrKT/emwlRcP70g5q5mdjaxF4dUpmir0+mKrWO+bvRjngobVK0rvU4cLoJzfnhzFf3B033EK/mbC
gpuFOXz53rN2bM+CBZpkYekDEp44eX5n+FaDYGRtYDK5UgtnF/pIgxhK+rLOfhycUptk3kscOo72
B5zHoSLGi3sxJkc2h8mWyDNLHzJIhM5kfcC6ZKzEiWoWXZek8vtfZ8WRwcq/i44vgQdqYGY/gfuC
HHJeY3SrIcxXQGLThONtujlyJV3O25dXVB7ONNPZxtC3Py0Q6oGR8O5dXh3nqBufM8wKj/n0Rem0
abyojHtj29oN9hvXxATgfGWBW0JcLO3YPSWJguUnUjxyD2XM9FRn95UfZKc5GqSO6broos0LWUsJ
uNCLKrV1D8UucNQGoeEXeyYIxLHx8Q1UE8wh3ApOn/BPGm+06CMtN15lgmmo+MBOeBujIYvC9Mx5
QcAAZEAv4SHXWVOMk+8p8HndxP9Q+QNwGyY36KSshOc9MH6dAKVF9nPL8nCj228zLKIbXCXbQRiq
r6l7soNwynFJa0bcgjHLirrqjtqq2wJwoFwKIxYIaF8dMn8860No66fW3rrKLtgwp4BZGjAHCG1U
ieinlPUVkNH48RN+gCoQaCBuPvzems1YJAhM+A4NGIFbGRieTL/bM+ZBtaUF/QnZMmgIB0eJi9Y+
pgpfs5U8FxfBMKlimfDnw0BftmV1J+lGhYSLIZwJrVLH21O7MVj/LOkRJEV6+CPejkJ0DTVaxj2Q
nLMF2ZyAmPmD6aJ4YfEmJjb6zxp4hsfJyEeB8ia3aVJZh/47SC4/Ed0Yf48vjHjOB2JI1I8xwa14
YnjarKSlLzwhQ6F6fUQ0CnDqkAe9M/g+z0Y8N2eqwa/EEfRsMzWsd6ybUJt99XmkgDmx7uafUhvy
2Nt6aoATkSboQR3NYwLSpmCVbUuy+yNcjW9lz2eAgO+Boez9dpLs1TN2gdmO6jrzYtpOtQKJaTdu
SdixRW+ez5oK4wP2QVHquMAoMcyur5/obO+MWDBtSaIgIOpM9imRgkwxFvjmCnVkm+8mGoEIBsWz
/FpHr94N29Gr/rcAgkDXDCceUNLA2uBq0iItKw4IyImpmeVJbs6bkTvy+U5AYekwGjJPEP3NyiUh
uJ2BB+yRotkIDTm3VMMye/yG4N0+TaudRWYJLb4j7w8iDpLAXkXO7XSngLZ/B5NYY1vOxxDn9nPe
1vWkUvfmAJxBE0qF/bRFRVNFwIniWYqFeGeMDKNZU8lrtRSQjomIuOznPy7sA1b9A4BavXC4cgKe
o4hzyv+qz4nlwSdQSz9cRxWXa6yU6Qe09HMDZcWw/mlTtYV/Q3PmeBwQUOA70i35egjOBzivtDwA
czQKesmbzkDZViHsWtbYB4hlIDR35zd5C5PtKf5LCHTEKbvZUufC6NY7BF9KAh7sXXHcsUOAuuSu
yqWHAq2l1NF4GM8B6j8enzY4g54qQwQ1njHIys3geMCnXVMFTXRYFa6oE+FohWEufuw4rsvegSdn
3QsCLUw7cW7NBFp9ZlH8XGurAH/uMHdG3OnVl6YxY9IkGs84UxiktPEAoBcqsRw7GCVYejN+3hUX
gZUm4VPAM6gaUQGGRDnFHGZye/DRPzmlfgaJN4O0aehKPxkdNTQVhfFl0tbpZG0SOdyCHTb4M3Sf
FedpNARbT60uuCRKtOqmfXBCpWpv6jYEa5FOYe4rVg4Hcb1AmW0LuDt6couvSyMJr5M6HreKMP7r
UCTT3edZ/6AQM+WVCl8ekJPZ0t0uQ7ZSgXXtwN6iHNtU5OW46Cw7aj2fmFI4wSHGwi8Tpxv5+JUm
/tHKIN+PBa+HDPj7MkyQAUIL0MrYtdTpSium0figY9Bnm7A73j7GFolsMi9PKIltvF22dnWjVBZb
OL+fQE9y+MDKXe6Xe61mz/XNtHzX1v9PZMkbBicQ7rJKOAamcgxRQMKkhak3GTsqkH4r8tg6UB0d
+gAiyR0brRoau4v6LDL0qmLZs57J81THVcXrL0+bsKLNLmWQ4POnRcPN+koreuoUkwVcTuMg1MLl
+cqyDgIyleHoTYkdA9g3RIqT3+LBOhD/mFI81cyszsabV3bpABDTOgy8VM9R3vrgnCoWfUcBRsUy
iC6BqSbYRvVbzu8dljIlY8y0RFDjNvkEePjY4zV/8R5UbkbI4w9wB8F6BXl74xvf5t+e1ZJIYHbe
HYObDJOn734HfTWU+9ueAsQlKrnPnbKoSFWFfgAEUfZ0rQKmJ5xSMckq4PkTims47XU7omsagq70
Vul9XrJN5ixrzh/m6CGlwWcfB1yXsOjEqY4DJYz3+F69KEeKnpaXqYhrouKpsJsVjU3Om4VJ9ibG
j35MxP4PIxJLv5CQqiQJ1sPlLGr/Til9m/R4aIvi6tx4uzeBYiTqzrVn/peNeGPJUYxUiwqUPQHv
P9k2rsqMiCgs+Z7uixjxhhq+HkRNWfvgTrJNdnEdTFIsnR086TsdHrQl9pMHavJlpiP7eeG1QI9U
TSDF0hwTQfZAmbd9W64dCqt0epIvISub37JfbbsVj5gtXzWuHPo3gFrhFTHnEWned1DtHOB2a7Zm
jFfG9ACUlYK90HS6Wb9vMw9viS247ck0gmsHtpFR6Ocb7qFe26udcpSBv/9NumrMSnpbeFgcx+bM
iy31SkhHpQhnw9x2RhnK2O5QW97XIqah/hIHRZH8/fR5+nsGGiQmdqmhayMheHIS5dlW75LtNu/d
ikj9j+UYetOQHbDCu9c9SXmkeja9WUAiL8JnGPy60LoxMeyKcQp8b2xprE/D9mvahiGly+Xl0AEB
njP3PC4JbRGGeyaM+sJRMHff/3wCf8Jj011dIpEt1nBae7Opf7Zi2aEaqusXo9ZgoDGtBDXMmBpz
0XexnzMvN0UTKm6RXxSSPrv5ctJcWSUwgWicvAHJ3d+YOgnYJMcAS3ene75AT0tDVI3f7Xyf7I+M
5ECv7vMCnBhihz/BUq1U+UEW61SzT98TE9UWwkxgavSj2SGInn8FIujChZ6kuGSTI8yFdV3jUQW1
4UXEd+EcClaqxpi0Hap+oGl3UV5QgjoAF8eOqLlLyVAbRVnfTlF0/o04Ne0nmbW6b6H/p77WYCjC
b10VyxeSZR5dQAMvg5UUhypdeqg9tD23tcRb4TQxzGgQIKDrdN9R0HIzMuabmG6HPsTYqLzCsIJa
6Qgp1CqUAgNIJV02/OZkUCFuHswQH/gHi20+EkkaFADX2wFl2iOhRtxTJxVMk9lYfF5S561WhZef
KkRjbeeVeJEHnsIjMI9OIMekJ6uuUXK6XLBsoZkRE0/VeDnarYMJn52D92DUhDpSw6dPL35jgFCS
UuvT/cr8fJnUQXkapuRfLFAxyCttFzjUjxZen6XlqTEWVNw0iQB/T0YqxJyiHg9iMlJGrlwLpKr2
L284iUmXKuiQOFQzmsnD7e4EerOgDQCEM+yTWXbrwStPPaeI75y86F/xgjoCEShUxFPiVUcLtoxC
vyjS/OJylF1gTJv+xzHRrMxmhEttIuhrkcnZEOUNHo6/6OwuiGO9/XHWLTA5EuM84yB5Ish4zorF
h9MsKrHzDDgDjup88K4ZrjPluowddfoKvgofu6SnxIlxXDJsBZkrKfLWLssULb9ynPE1ZO4O9nHB
AjawouvaconK+9XkxHncSPtyhmolW6x04N1Bp1tkTmSU3Xry3ppVRFpHFAjqzH2c6hv7nN7uFttM
KoS0PaNNbUBP2PdJyUEmV2pAqQmPjXLKUAHXQhuNVkhI4kK/wxDERYRoGvZK+huZE9BeIzsL0wP4
c55BnZ4uU9VPztOojHOIYTYFH1xECf671rq4JCqfaHMlKzDCabJ1MFbDc3kwd1HoeAleMZv9jx+E
Q7IgE6vf4OEkZLJmssvtUv3i+GbYLDdtb/77ldpuwweAZK0n/qMaikfdegZGtpkIDH2DDF9Gxq+1
M01UIDoFc3mnAvZdUYj8DZD0FAWnvQv+eCqY+/wefq5487jrE/0Ltrv2C1D0DcFbnaLaJGlUYRgM
q9SPD16v92EsrGayblp2YGQowecIRIMjLkkk5lGo6qrl8gj4l23i4FYTdsfYd8BS+QCQeZJQ7Fz3
1eEo+KSICg3jIURMz979nnVLbClgzbtal34Tbl8ugKTbUvhUlJSQwPIVC2io4Ag622O8m9sdWZwk
8uVu9Y4/PtEy9mFWF7XflpwvH0c3Q9eFP5fsoJ7jcTJSPXer/I5PCrZZmuvVUUOVwL/r7tQdXWP4
qwVGSdsYGmYIr0blUKdRy5niuClkCncyia6d6OGYV/f0xtcOl8QCNrYDpWc7OVhjhu1zyXmZuZTR
69epq/5YVW3Z0JRJro9cj5zT3H0VNTdjU2VzeiF3Z/yIPSpD/jgl2+1mXYWbkH42002tydAM3En9
3Y1c8wpKA21jnnLDchO6WIrXzdf+i7rCgZECHAXfjdTFTaQu7EwPY1f3L9Teee/1n3Vw2ZdAZeeR
QT+Xmvy1g4LEKMl8R+C3rgu4G+B9EO2DIfOLdi3E68u/4wTvaMsfs2lYgh4s6sMfMaHgU8ifAxA4
clJYLrdN+IL1koS9ESca/MMhNldm5yC3EAUNns2ZtkT5vzZB87ZM3NzNVZFjtW87MzDEZjjlN4lh
jk53OOEpB0u5g5mHs1QpFpNrF4Pk5dwfW5dnZBoeat+TvbrPUFZmtalV1NgE8QW4h0OwfHiBC2Kk
ZOchJcZSI4s66pGC8tXb+vLsY7llXu5nW56MLXiBzCljdqL9GXENj44PPNOJgpPfK+VKu+HL5Rtf
LEzfyVh5PwYwHhOE7OeeQ/qRzbTLz9AkKIL1lSLVbj6YNDWv/tA1m7hO5uYV+EJtwu6M5BmNhMzr
RzDeU254CD1Y97d51hK+agSydrr9fYFboD5HU9FmFO0vdAHodS6Ec2puxDTkApr3y2b2Y7hdDTav
Rb490JuBjunr0ZvVLBj+H893KPWEugeA5XgexkIoiNjs4EwZskbyb1Gtmu7PmmRDonzr2FtcCpDs
chWI38K4Tv9cf52bitMV1FLTUidRc4L1QnnCWgltQ2ELhoR+rQml6wD0HhI4zp817cHc11WbjZGb
/L15B29ogjn8VqXsLO8URiRDMwmqQGfnGt0Jy39x8ydC29RDV0dtMi70+UmrQYNIRkcbJO3Joph5
esA92ny4KPGi7E0Td+5OoGRFRQirPvZpNzNez5im4V6cueikX0YP0RwBGz/IIhQbmFOI2MDDvRbN
1zsVzplA5VKjIAC0XET4M0OgphZQKTCkHkd073m5qn4IMC6qzeJxWRmoAQchclyNyOWlkrSjp0NP
GMeSXtaUmAfn3BWc4NhUsq1X9fArqukmD0n6A5DsbL9JD8ln5vWC8mj5jSnsY+ddhkLXJejQGZaA
3oti0fxcN8KPwXa4p6v2XP4J1VXZwzfoQxDlCQSPuzdYQsMKfnhg3wCDe3wuMQ7c5/IyNZUM2+Uv
gT7kgFuZiNyVOVWCqw2hk8JFfsevs8ZjSPI6cPpzfslNDYzPdwKkmcsw9jmgWO+ZuwGYpCpiUyTH
3glVtVw0gVWKdDOJPo00Hkq0Bje4n3jGlOqiwEZT0uSX5//hRLtopFDPBV/nNLvZK9E4rfjcQYgx
VJvf6XxoK3taeVgDXdjVGwKUdpqt443K6N+oE8IJ3TOaIRiBjoY3QkMLrCl6yX31rkGTyNW3Uwqd
axj2WeVGco70j9YY6Ubizwrhf2ZRzNvr57sFiuCYhD/XD0f1b7dJpbt4SMWHUjvYjNsWId+3iXm9
MW71stdMfZmxZ9LHfMcY2WX/pqCvosPZJP9uwV6LJuyxSuKE04pNhmYDxQCfY9+mdIBbSq34054c
8j8JYSoN8Ye81O3vUZiS6ig7vXpsQlFUN48FKGDe8uyHra9ensSgxuhPVyNnjyMoQsKFejwVO7qz
ogt25H79mi+j645sg9KGfUbYYB+5LVjZnzIM4rhFgL2D7ec4K4EXXpOukmy5/E3yY8NV4oLiddh1
9Nho7R+ZROV6s1AHIWtz2ym8Ii9m6uIkMsuQ2Q6e9h6OP2xnNQSm8NLJrCRwpYwl2DyfviJucz9c
KGz4OkuSUAvThTafnWtLilEFIhjJ5xaf7E2AsbZY3X5TMfOxidDJraUFcTb5TYAnnikgPy0yyDht
dxOAFu/UQI6jaMatlAFWVNuU94oHS5FU9KxtMNGaIpQsv7a3mHivkoWHIdy/J7Zy416h/ucllkeu
K6EjML0IHFDSqESds3MgboiAGuqfUooNVXDYJpRo3Wd83PKYLU3jMk8gKd1K5J8L0E0G0tG26JQ/
hHXwIRY/WMhRnmTGe4UurjrRtKb+U7AHj1VdIrC8zPoO7rhVA2r0wDWxlK7M46VrNBi6eJ6lnx4F
RIlNtEM1IfxyniJQI752Q2stsL3VXIeNx5GRmKkIRMdMe64fvVBDboCdBahfkSmT/V5GkaLb7+VF
Vdfkng+fE27w0fkQ0sk9ii4oHxyS/J/wyqG2jKXqlD8ENJzb/NrlmteimXYcKrcbx0OKM8hljb9q
qPO6e0v6CETcEc6UAzdjbcQZH7/fhEwetNDEmLBMOwnsN+psBcieOd+OxVjuIO4cndzuYcIlO4kU
z2mtNKBVqyMf7PoR/RnXRxdlpYOOrnDDv19CIxMcU8+quqPfSX0SXU4S4bjF9w4hGeGMy404tT50
OXimRH6iIVdit6mqsl/5l1zb8SyScJbyEWBXuftJa26EKVw7Xs0H+rYq0a5u4pI/35lpaCarBDZ/
FYkJ+4DDXFZ3pYFQc724sXusJkOmXqDnB1xHzUSvq4hExDShvQegVYEoxupXPA+ohVchKqBtK7wR
/ZtrtAHHszeqHcqI7x5HoLErJbhbGYBzGDtcr6t2hinkGpSw5XB3OTlujW3hMv6N3bhs0+54SPRu
FR2cw/tqEon5LS7bBWIJQI1P12FQWBIsC+HFu7ACBpwQAjZYoFkZ9ls1VcW8k+3qcepDZUHI+/Jy
8ZUbB/J9UxxPm9ZNSqjJHvV9ZhClMfFM6yxwONKEWR/Yo8ZWImW5A+GKzS7h3/GHQKDQhzRY2urx
KWIQcVgWZ1azl4EroLXUS4NIj51l0RvuerCR1LKyk77BW8s/u36ViaN7IJedEBaM9a5bGwhnaVMi
f3v549NPvKjzwzzJv/s6NXEOcNddo0G8rXqC2PrjId9SMbKjIZFOz1ZQD4oX3/NdVJqnlR3pjaN+
EF3Ty5DTYss/g4crihqeMLHNnNTAdZ4S3BV7hVLYCnCCws0Nf5lS2/dXHm9ybW7Fhdz9AxJns6hK
cGHcJMQKH7rcyU1kNSKYdY12mbXb8SMvbkpOjULexfjf476EnZl0VxbMthInhsA3vG5WARIevFZX
tzafWRhjfMrJ1q9XiI9v3w+SZbsDWJFMjC6kVvG+xdXgYTeAdzTHrYc1aNMuhc4pBPspxvvA7IKd
4SeGb9fyrspogG8bQa0sys0wxY8Kw4ZP4XakMc+28NZXG/MxyHOug+jkBwLR1h0Vky2bsHdvodA4
Oy3T4stAp9WqitzWfXxxNNQ3K+dGg2VsexeQrdjHBANsvytGRBPSYZbqm0d1cTS9W5pfg2/3bWcF
2gmX6iIR1NqQmfqaYDB+1m8DR3VyGxVhm34Kuy/aEGhBOkh88c8WjPgsRHQKOwJsC15OwzzDAVy6
1esUzkdzypJJRa5Us7O5dzOo6vqYqGfpTAagR4C/rpCGMs8B8t3gKdc/fmXcx2nAJq6rzvr7wcPq
TkLr0xkxwie5ZnB6Xu9cOTx7ZRBY5qQb3tWLvw791tdx0oR6tMMfAlI4CqN2Xs/xMCCQFLows89k
kQzQkbJKF5b5a9q803ito0R8DkIyWbaiUU2T8Clm4iSXfiMOU5NWzRaHJIWNlLdnC5vnV20sf+0u
63b/Tlq/BEd6cX9Yv97BW1FH/fB0TO/ez96bHSb1dd8jyPYlN9SsDJCpB3ez/+vg8CyfTb4Mcraf
fsgV0IH3YP3O8fvUG/LAoun0RWntZqOJEwEi2F+jij8HrhzXqDDorggflu1/rx06VzzglfO/BH8k
CAdt+LzllMfBsE5WfzSAX9t8R/Y+X0OYCru9O6qKuUzfqsyg9x8+YPI/T84LU/yc15peZkVSwZy4
qVGiZSDSpGsQYJ6zTZ49LaKFqNoJV2/yzGw/+8aKbRYzQCviFoQR2/A7o7SVPNqtpLga81nttDQJ
VkenDFt16eXgm21+/MVm1QXhtVTIb66d6PhL+aEfhxi0D6hc4NPjma7cRHMKg6qL4bUBbbXzZyps
IATQrSCYGiUenFhFdRXxzlMwqer+FOdalE9UfAY0JbhsidfXmpTXcXvaXx0MXy5ZIXXnDgRPN/Nq
Bf+sZPWtBpC+4tU4B3LaJQnNjpFwVoVHpCDLdph822amujuNxoj4ilgwKGR1kyuolJ3xZqVnkPFN
lMHsRbj0IEGGrxv/Hz+DwX/3oV2s04eq9h2NsbdTUFsHzRidUT08ddnB1n2skZHELPJ7tnTzMrJQ
04/a5fTO1X2KX2XeSSAO7qwDWkHFhNGH0T1oL8QCE4RJseRYnheO21N/IDiTKmfUXfFGnIOqxTQx
fqsB+/7FqoayEvg+NdToBosyr+8l//gP3e3oPcpbn26cK5UYREkneej47CXC95wupYxeI//P5uCq
2b8Iav+L+LxJaeaTVrZttovyrxYhjfB/J8Sviw/1qvVck91tivOVQyLY8LzM7SYhzkIEFR5aSdU0
iPzaE5Fx5fuady/XZSUy5jc5c0//aXqmeEo2GS/xUXhTQFaBboS9Kfh2VRaEsgrJ55TNCoDIRu95
3QONBk36vLnGWU7AmwG4sw/wvg+kY5kBD3zqGHNiUEG5o8UyYe3LQw5HMEbDlpBgS7Yytzrr/hMg
TzySAV+iya/izYV5UA0STlmdfz/vX56myDxs+bK0pJu9Avqhl0gMcEPAP8BT4R9uFjx3Zc/mPWG0
bm2+1/qineD6FtqVGsDpOar7AnEXILquuu31Mw0BwLWnaKlRa1uW1B+1Hbhqg2NYf+99rrHl5e0k
YyQvZwMBtkBGW7dK4eHgp1sAk3ulprUU9+L5Yh5FQEuom+nr/Nx2mR+7fsxjMDrSTxOnJbgsGz7Z
rjR5WNJQgRjALxIQWdUljt8LGA2Twd57lw4xXJaCMBUgqTz6jWCBnhfZruAFGy4VoG7220v5jGw0
JcHVNtmYZm9NFIHy8v8RJAwUdw+TQB7jbkVgpBQwxsBSLBD28cFyVLW/XeRJTdQwORLBNnEEj2S1
xG0aM6dJ+x2dKmTIIyX3x2FGRvUM42xDBZOkJhVyWOh3DU12RzTJw5+ZNOit15zikluUcjouo50p
pMcm0i6k9ub9gHLepF17sbeHV+4CKnQLYCg0Xn0CJ0EZQqV3SkFlzuclrt0AHCxt4n0+An2B23FF
/gRgY68ixvhw4v38pi7IvnfvAx5ukxRTgboxSwHTG5ONdbqJ3AMssAkSQot2LPUr3HbpnKHCoHz9
/OJEQbWooXmx8w5Rk2wob0cn+FiyKUUPWKZ0blQcU5jgE+q+Xp4IFPPitVRrgQCtws9UsdJNGsr6
LY0bx2Kqtsg59DM2Un+iWq8J45IVvNGZAoKWlDJ0hJ7MnggqPeWtU26oHJUlH7SyedPKFgiosE8/
zrBjitVGEuF8LNGW4t7JcQv/BeWKTPzB1lsD3YOZDYgsX+DaqtKJC93VfSGpdui6xufc3cZ32WGk
p2KklpOngyojahnue00ZiqBhOawzTQg/3CDdYuS3sjMP4fLByK/uo/fIqWijPaGoSHGAq45voTW9
qN10wW5GChY2nhH8azEaZiAPmLVIEHSraPJVGlmUmPt0qaNzaXwrc2kslyGdcHvSiHNdJDHuguzj
rEU4BF5lLVjnGy/ltbFyDa016RIrjyK209J9ABu50Nr1A3zzonokOHtTBouvlJBZqFMrhFTnCQH9
++iY4Y/B30dhis6XmedwN8RtcrDESI8/tcysTdV/SUD2EjrXzVgdUfBuXdM0uOUpyUpFbmXi40Wx
TTYfkQLSY6cccFrwFN0dR7OiyIdYO9UsOivoTUADBV+rG8uZNBTICwiijapVkZmfhWw5+6laqgK1
JClmUq3GhHFh2QGwaE1GhFQnpS02FHBg51nkO9NIQn6MPMrsiIFBtx3tvxnHmoHrUG2Ze06SMNl0
Owton/yCboBttH5910horJjIDNUXnlK4ooSZVdrdC5O6ya+JoEQYIqCNPHRQCDWfmm8nrK0Ucts4
dJnpoEFsyQ7KeVVvyyLlc+ZTYTaxZsH4R27nP4j0dukqSrQSIaq7aHWaxZw6mcq5kXfyVQmQLiny
cTpjV5ijSXwcJk7/elQi1+ufDYiTSTmmWzESrIBaGvhdVOgApU/vKMEhnreat9JYneKK4HiRc5AB
x4uFTZqIDkrFoDm1zg80ooHBtVBehmB+op+8yBIzb8EqFT6IRg3UwIlB2TEunYrMa0Ge1qQH8ov0
AQcR8zqM7WTZAZFwdoL+GcfMAKsRU2Gxt9LBF7ItZ3YVuIXnoumjWuYVpyc43PqCcSraKeV64WRs
CnVeUE8jV2bYBVPkmOsnNNzjLNA9LHqC/idfCjeuvHbQzomtrgWD3ftU+LXvCtOv74MfGb4jlp6A
Qz3GYzQs9+j/6t1nG0bQJFAuTcTxPtLV5TBWtZtJo9ZgZOJYAevLiF7F8kyOjTUPIpOQVaubKtNv
urWPQS+5n+3tGwh1OsR/2xcE05bOYNthTiN8SVgX/XtD26uzfpdaBehWL1MB7tOqVsPsaEKzxO0n
n2Z06dElrW/8LOJyJTC7LU2zl6P+xRiISLtqKts4OXvLNgAydwl8jOy4UYLttUU3UeZp4m5iJzK4
WnenCQIRKTafmttVNwXo0U4SGCvDBSnHl2o6/8cpvsHZJc6m7ng1e5dly95uFhWbMqZ0v02917Kx
SuWNGu6xVYBOfWtczLlSmhcM+ljlxRcpKkxNqNa888WNk2Vt+3IRmPEPkbhfURsd/oZMbbfL7JuO
zGmXYjuwppHzqXsqj0RUfg6hHcZh3h1TrwCurmqUM8YtOaOxF7ewwJhsbxoTRi4gQMFO6+wCe44d
FL2vkO/q/VZY4hYBtVwJzK9nqn02KRQkP+sRPGKYMV4GQOG07Xv7EWFalDMtzddHUpRVI0/idX8M
kqvjiCrfDxByNJ/GxZQJ83mSLN+4rxBS7wSFvAGpCmsrwny3NkNezQ3rqVJCHFP6sMc09oXOJ5gS
n2MowVSbXHZyBHtjWgxfezAzu7D2Sp4kBOBDUpWLMeMUci1Xk22BYKILWeO/8vaY5dXNzDHtT8HR
TsnUBwb05qw/TgNBE3M1fe/KN/jTj5uYxCTMOb/XzWXGK5sbSWXbRL39IwMhjaJQnoIx/Qms2EOP
uLKc23Cc8gjSorczAIH8/lAHk4CxyLsoQ/gXMLGlCvUkpiQt1qxpKBBRS+M1K+rJw2VP4dKn7vXl
MPKkcGBeAJRSiOQCqtQ90SJAEFApngydjVY7r8rJpBqt+8e3ZFmkTz6gsiU/QTcgI+KTEFFIATXZ
TFaEUZRja68kuaYAKmuC+D7vi5b8Szj+xguRr50M2ze6LXKvYFu+rAWHqGBLhE4qembHv/9CSmVp
hfle3LTJ4l6hEPw4fp2ak8H41bCO5eaGHGrAmF6aTDoBA1+ARyjkUcbFoW88S3n/wMBJLhpXDnj7
slB6avYuEYKGw+ph5oimI/FAwiSvaO7AAXCJA0CmZdG1TOZVhJW+2colAAXUQEAxeyPWQp14db++
gSe0ssJ4ym/Sp/f9AWeYSv0UGNAh3qk0zn1Ch1q9y/mnjt8Gvr7ZxSXgKoZIEL6P8tc20hoItzBy
JyyJTkhSNwUSM5+kAxW/yG9I2DYI9IoLV/5y6I9uPPaUsMFBpRkFipT98H+ncY4gB9a80iiLlITO
8dtWfJpi2iuGwkPDdkYf9ZvY1jMA4O4lO1M0qOrBAk+wHWXUwo38O45z/KxBjsLzAirQXsPvPlWm
IADD7D4J5PT775KdRBR+inf3E531bgIbHuFruhDD2PqZkH3GqrOSnvwnzg07zzh+80nCnsiTPkU6
uepXRWvUIvJpKLiHGKIB6+SODavy72kuOVuWg0cAlicu1I1AgMOek8xCzUku1vgzRl0VBe+tcmF2
eGhhPRp9lFXKGFwPiR3eGT8FfKXYZ41kuVdRHzcn/rk2nxYj3ufkjsp0h370waoMJr47sOozu9EZ
rwp/YdL3/cjtzYNYxXhrdw7TGp++2jYIW6Ti7cf4BoxY6GryPHC59HCuSnopmjJq06BLUQkRKMm2
uie5XpRYY/bydnz9aXhR4+qUxgPiGDnyIWDMXaKZ/zjutYiLuWv9H0O6+7SM+W8PY8xlgOLn6xl4
P8qiDk6an2wpsK/CQp9JxfHH9fRBjj0OvG3tWKv5PqWTqwM0zezSNGKmUvsXLr/hysJTN3onm0oi
EBbOQ7P1th12sCnovXpSluXON4ONagyQ4nyHswlhEcf/w722+wDNTYIYVymgjxetNz73s3dI0jww
haFzYAxmzRc+iyhaUbiNBRw2nJs3CrY7o1kF4NzJgNKLeVQhVvIDLwEk96H1ubd3BfVrm0biCYlX
UOjAkJAuQrYMiLu6zKaNjT7VzR11IvkQjI0OsWwM5BGORSnpg3ONegb/nIw04a8cK93eTQCh102o
vBq6Lxu5YRCLdpllJB84W6R/ZLAsDaxN1fIJteaqmz6NFeEgt3oe3KR/XrKtg1Y2e8Oo6WiD2HEn
MBheK8t0pdcnY/zoD7DJ5pBmYU7f9zuX3ZMFb2hIqS33cuwHQTGuot0maXF9zdJL8Ge8Bq4Mc+JP
gfxmyz2iHjtNkb+p6qbkwaqLn6vA1BuXDqob408A0XRFz3l5SvICintugx1jTk++PdLmYiD0D8Sa
JmHNEoDNACzlNiBbWYlmcYTuMsVxe8BffzdnU/cAYX9dPpmYC59oHZRQ2CT5VgDwX5+zPfv1lq0z
d/2S/hr2FL52E61vO08J77F+cWnq7nLLRzqWKjSDpFMBuPkcathA/ovpggQ5LrBeV2sy1Rtm374f
PtLPF9eRY40KEFz3Ev6quLBSxQ5ycrVMnLaEFKUIzkeutnid8xsvi14ZDfFgociwgiz51LUQXaTI
hYNappHl1Teo7HH5WCRPTpgixFACI5/YxPqrcBM9qF979SUwU4TcM0ZkyqiHZyjly4MkPEri2oGF
0gVbpRKhkMpSRsk+nic+pabsNcXARs2j8Wrqs0e9ZJ7aP9tPEHFb84HldoToTeKAgkPKimZ1aZr9
IPGD8jACZiAHxwFTDE5e+9d3tWl2YH/MrxEfaoOgNh+q9mJwwCkQaMQJoTsXIAtHHOQCMJ5btz4w
/UJ96XOHl3//+GjHgC9RsnJCwecsKTFFYxwgD1x6hPcr8RwjARx5T6Beu6pfm/6XgtsnIJhqC88q
zocli9L8ruGOnmJc4RV2Zh+f/fUBrAcQj88ag59zYkTxRJ9P0da8pLq03BWqj0lDUwXMIUonXADu
3fwHwTtX9XLKQicPmY3sPuE4y0ylg6ApMIuQGWLU7oCwfblLARlOl4WGBZjsKPM+nBXAuAvJJaIT
miuE4ElJQ0+tcRfT40fB4KgnKdkh/xUYn5XbEPibZjiWWuyrqVXmqXOFwb9GCC1AOt0sg4utTpol
k3662Hvr+JnXCJyyr+gp9HrprskHDNHzfIGH43kKIZsnAcF22GJFrfd2t3YemXNpxNndESmwFqhb
x1L4M80EXumhKBcfaax7g5f35n0YSkd5SeFgfshUnZ63uziSO4OJAiPcRWZYu+ge4oB6VcLSP0Kj
GjAqnwbrU4LI5vqeF1wv0BkcT//OuyIiP9CM28rDEsdysDm3NKcDnif8O6DR2V5lpp6dD1SicDE4
uaa3o+1IpIGOdP7AOUrkLsyZCXdGyuUAreB4J6ZDkDACSlf/HMnLWHvNN1KRZA5hTgwcP83GpNwc
hR1qHVWXADimN5HeiJJW8r9AF2av5R301Nbl0Ij6Fw1FxyrKksuksjZgM2VoSzsvzdjLkevAOSES
pASkhAetMtlQlOgogwuwUBr30p5TotYIgji8HZ0BT/NeKGMPerqA6gWwPUpHT9b0cRWtzqxKLX1n
WagGoQWj8uJzBFvg1n/YlGSH1LlxdjeXABQ5GOLO74SZC4pbVhR2ieOHwrZQmNmLL4w90ISIeQYr
65cxmp8NaYxBTF2SuccgFCWPt3/IoqCyf0KYCjZa9fW09zslC81atBCgo9eRveSeXh/PhfFBC21i
fK5yyqAOYd+Ha05yMnzcG3SqH2efW2f53x59wfrgP7/imJ07oraRuGtLTr5PmDmhyvNYWgM96Ink
UodGOOVPfk9L0RXU46GhBm42SdpQreZ5QtnsDjoXq32umAjLSlEpfLIkvXc5ziBudW8V8JjuSs35
REBU2+qsR9Hdj0n2Do9NCeWQjMQVk9wA5w4nV2aVyOcMihsfDO/6pGer4ZSEacKfTc+fl8UZIdoy
Mc8LQMlg+r0+adcXUhAmkjdUR5phrLwRHpAfIYO4gE4pQXRHlN9IYu7PzYPmFJgeKLKvI8B71vlT
rTTKtneENBg/27zNwcP8xu7DDYMiX0muvUNZxd/3ElBu4Bt/pvAV4SyZlHrRWgFNLLy2BXLj6UCs
/D6rSDBQQYaiezyvwPue/xa7aS6vPfLbep/MP7XLtNastKwrv9qquFfMNawsjbf5W7CPUlVNWSXH
CY4EM60zbWYSi1+C83QKRuIFZrISTGK4lbtq2of/TwrttBzQg6pN4XtN3HqD2OTczLfSlxSOOtxz
1KdZ1MV5A40LdY9OZGovaLS05ZW4tJKWMEKkUsReOJ0Y2T6EtXwpcoAPlh0/pbDGPR1oEtXwVcT+
GLuJzuZB8GZHz+XyMQ28cLh9SFU7lgL3wUcHnTLO12UurgSSQ7WCLu+duyjknP9bQ8EiFi2w8p/r
FtrLrDq9jWqJ9vMhujOlpuNZblEwY9NGBoUHlzIGj4MUEEsq+06crAkzT2Yq7CYm29Dc952BLq0n
3EQWtdXKHFfi7A/mDshxH7G02XJ9i1S8SO+xetv0zmqGZvuYMRmuRYp3dLlL0mNGbunhfYyldsKC
g/SJF7btToRw43l89GeWxpDAm/muz6pUmxX5bzId9rZjhhsjQ6u2UiuGXFC3S1bcASq0MK+kZdMj
3Py+UnpYFe+tcxsAJi8YsZN3f2jDjPqeuy1KhGmzpRjWiJbT/hU17JxVoIy2razDXAB9yiAIXVSs
IaBZDKkONjBcJAeWZl8BcbHjWxT2b/26J8qGSNGnqOeCt9WCAvFO5maWiM7DaYFFvibur1nNvrCI
CbJ71DQtl9zOMsW3J1N7O9KshwGv+NmlzWFftvW+5Ql0nLsJjmlU8Znzc9sGu9qgAF55BE8I4Khc
CmcUhCu+oF+gYgmJzvolf9sDWhGKCPbt3O9cMbIl4lzqbZQhrsV5vayu5Wnj+y1iwPUrcaLHiSUI
b7U0qB8O8snaFac6HYoMz/Dd5aF+iIaWbU9kf8tSBXNzCEK9Bqr+vvAfQHDeNCRRib4kumETn0ka
2g1kpVxhIuWYAyl+GXKW/jpgCOce/y2WNTH3eT4GEtePbDdm4ZhE0b6di8lv/b9pV2byckgacvoE
1XR+bC8H2mHsTvjgttBo6Lms9dBc5b28gF8fPU3025WIfjiyVrXMMNg8iUnnTgDf15aS3htnKdCv
Btm1wePtotcqfi6HTzmUCd4I8x3ToJnZiyCI7L1r+yZ7bALh8Tt5CTfso64v2FI2IRipfyIbHbnJ
7JkoECZ9fGuaY76rzUwsAw5LzdpYzSEl8VHCGwUt2RL2B35TZiZ/y2z+fdE+e+iHrzr6cEepHdio
HOK2Sg5WiPtZrkQ/746hfk1DKA02bqss2VVfcaaaA7TM4b0SVNvnbtCdoM50NhFTJiJlULZCoOXK
Kt+WnnYJPlagKT/XI/2l1P1Es59jy3ySo0qtajv1akg7toGU+nXqAVweKcLjlYZwJSZoOm7P2q4w
U1BaQou0amoy874EIUN7OYis91jzeTKbepnAGWf5cv27xMBStf0GQsd8aC3pw+oNrXDO6W+uR/s9
b1pBpdITOLeJc243jHkbElSh+MsEHafDoyuQy+UBlZA7bjdb4Ti4SE6y2msva/oEOr46dYs9rC1v
CUyA7ovqNS7WEpzBn04801BARe1VSLfD+wKa3tSyTC91o3Shx5TCXXL7Eyppi8rRpKdclwut9Zt7
aBGY2viAYSk+1iHVwAaBgEKQkGfcBDHmyhMa9qHfCZ/xhRaCX0KRbhxZ3pWZMPKRZhhwIN1FZoXn
Ds0ycLXqC0asSzDOp1+ElzDeQ0vXuMfFfd9JZ0UC26HY0HbSaoLYXve0RcnTEauvzJkWJsnRQeCV
S7WMYnXuw4V1MTrxIasiaIrdCuoRHJ7H79xfWE030VdTzMg2X2JtFX0UDLpCn7ELw+jCsDXAok+a
d7H3C0BfNITpSdeU9R8bQRKA02pqmj5x40tRE1YVPbn/nAkXdji5o+t7wtyclwdy5QCd9WArFibu
ETLI5/ES+4cOEooPMENRx1nKXxOsJ/yPKJq4BX0Rw2BNvY0QGpXu/9UsGz/9oSevZv68F5GLg/mD
GRF7MjIojsf2b33XWaJZf4JPNSXBZT2ccyIpqzCjvQIo9g3e6d7SF0WXm8sUjKyPtP6/DVbZcFnd
KVaj8MCuoeVLQoqQEybGg0XfuSxz4E2+vYj8DCKkb2v5SUeq29ygXkfxrCGsxntWjRDjBaFbp3yA
9Dl6WK14z9HFBsC+ysy1vjLzHKDpsqhj0NbWDzr+46CBmltMaw1EPO53vWOfogLq6UU3HQnMpVE5
nu53pZxHh2f5ioJIeq2kUUFZJ1PW03FccDK+4+8ZkS3Nj792wvQqFWlt6wJ9MRFB7XPWMVCSQ3P3
FW2n2XXgVDWJbT2dkqiIslRiqgIkPneFJWH0IFD9bW/Z0JQGCJYy12t8AbYqrYvm8JxS3+3XEMGr
q5iBvmkHBckZQqRoBKYQQPnSJ9N7opdA9hdwQKycMiJkuWXZ6VjX2Dhg6ttGQjKNsUk7pWPxnjvd
V2ZTLZ3GtOBlvhnMiHPSldEOVqDldc2xvLrZoowFIerlc9hkqxeKQ7kXoCmbNyWk51yG81Y9Ep9G
8dAGKYtZWTZz76cMkT5rPqVr32G99MHOmfaeS13EOe1nCJt8VN3vYNM6F0X/bx3QQNIkMF6/xGXZ
PqEbY/zB8w5jzJoaFBs0cR7YJSbJRHQLdO82I3I76JvFbX4aTsOzmsm7Nc53JW2xIb8pWX2p1VNL
TmVDjSGreJjm9P20TH95ynz+AQQw09GGh5jGVbrKW8fiiwkPBJdTHLlrCowbufUCCEpkIoA5z+G+
t01Tu8o6zo+PE/LvUQk53xbTDEvpsUglHzaVLnOc/oV4U+iT0mY9v4pl0aJdtkCIvOCUEjo/Vd4h
vEDOJsftbUGhxaeq+ZkgybvOHou/wsCDHT9Mv5WS7lCCs6ANfvFdfqGQKneJpYXqdhK15YGRIp5L
XEXekd2n1p3xTI4lCeayEFT517zmK2qF7wddw7F0D9c0muva2MZLbsLzIYwvRBBO/UhGyNK4+Y/m
K9Ma2b4U/lRvnWChJM3ADh7LIH3L0d8eNTP2oB6fPWrNwwwIFHz+6/aDAH/ZMP/azFMXCNf23u0L
vpbQ6DsrNuciwWFXzAKMQZNFqmeErk847y00u60XjMRKFfDWdOndglQ3llOLc9SG8ATxntEaLjy9
/5Mncv72cFygXsDO7fKNEBOzV0whWHZBP7Ns+4RQsDsRcOoEf/BzgNcq4c7FvD6o+BllEn2XhlEZ
sfa4HXzID9ln8MXlxkYU2+XxnXHFndCVmeYFljGubb6fvtSegQbBRobwbSVxysD2L+/EH7R+5Xsr
qH8aDTP/CVeNY/xT3KUoJquZTdv18k6a/Ey8Ha0qlSa8sM5t8NJui+nm9y17lJVISvKYVZaYkEDB
xYi+32yLfeYXhIDWj9C6uolOLEbkaPaGrkFL5B5PZq6Raq/BEIEId1aIpleoyHW2DkCRSfKTh0QI
Jd3gR7aoqwLXfX02ydeIrp7/sDJZkRnfcw7k4nAZbZtXpSzOUja/mCBECsK2iKUGp4wbVaaLqpIa
6aKr3mOhACjxdnQN5ffDrjndeW1atX+FnQdlzjAdGSe7quAUPwyVpJvj4WxvRv1ViSf37pd3hzGg
aWQvRGuX02H1fVZ9GkV98n/4xDJOUHLH7hKx8g4Rb3YaKQjNqUTK9l1pG9KuwJT3azSaGoIr0xVt
geBp/Rfo+F5LOt9tuixoVr4ftlz5u1bOr/5BbQ2uDYiyX2RqcOf+t2A5DMaXEACmF/Ig4YvmnRD5
cSJnxvJYNfVe/fEMa5tAMjd8ASVaz3yZbwfXllUiY9kb3Y2fWGBIYW1yEs6EaafQ22CCMYGSQAxY
Oo2jeVn7lGvtPqjjhVAfXCcq8W/G4ugAA4FG1yUZBNPB6aWxOYkl9f/QDwelZTrko2lpliCDniKx
qkY2U1xnafMwpKOMBuR0KVtNfQQm+qmoM2zb2KeR4s4iZm4BYxAYL0Qo3D3e5hfxp6RDqHQynq/m
V/UCDjwhb13XupHj0FkUNp4VKqRyrTXOU1fuZ8eK+IdfKHi+K61xA5Al37glkGd98YM4eibAoxQv
P92q4/Xq3PYmWYfDdmVFgygXZSAh9TzLJ+XZ6aYhWuM2m4ggIWwyUKKZveiaGMHqiGbAfxe3TTwT
KMUuaVxO4+h4EaFC53oSrK5RztMeTcbtqckuZLdTLMnwWjZmqs4CpXgCbpEjNlAEkaceG6F8Py7O
vZI6Ag6ccDo6tTcGzBd0N6FBDvOvSA1xAG9vtXIFurp8xJ+3eeebQUGcc3lbor4s4CY/Zv78kShx
NC+eUuIshRoY42qapxOZBV0bbikZDPcK2fp+QB7v3+EDn4ipK8qZNOMDCTwcfeGUQJ4e4BuKbLbm
ZQg5MMvRbf4rQMyey+CNBKnjlIPwfuDEPam7oZFgjEp1fkf/Sp3uhXvFv0e0PxRGl5lB5/j3IJud
Az/lZpdOISdWmkbLZPU23UEd7AxWv1Qu30Q+gye0Hk7lmHWDP/ZKBJ/SERGIsy5PGT9jkjD0Jsjv
l+Se1FfqQzGgyT2KubvzkTH+FvkhJrWpeNF/wVw0jOUQGrcIO7WLczNsSyPMfB25nM6IBMThaZVf
+Uu/9aWbaSas8QKSUZy6voFfD8p25r6FwfxwzY882sHeKRz5Ak2KTRl0g412A9SPqijrWACyCD6l
1U+I6jbE4mFrATIqBLrfoRJ6jXbbDxQtbv9QSGZo+L3auHGjABf0a7IJayV0TwHJz3R3qKE9HKf4
jPFoCCL1RHZgoeO5eqHiT8USR5Ueu83CbUSIfpXZVwHwxnx6Ps7zmtruk/xS4KYTDHu7/FLOsZFt
OnRJkjUw9MIqftAAiouLIC/tHxJASaUbEfIssrb6uK2nU/t6LWJLBvfIjbb8BjgIlOMvPDZavD5G
5X9fHn6vAA1Q/085WIzK1EmCZ6mxDnTVSQmfAJb3kSgwdPN8aX3p4zhJJ8Xhkg4jKTqx7/8FXT8b
htS9EkUcfxVgYSvPFw2z7RW+fjWiHIl/415ydKByhnk2wZq9YzvvJN9O+RyidLOijEXygrY7a/Bf
dOVNvXMriqtzSWYb8U+95Xdsuyl48fhLfOZ3hY8vcG4oacEhETH2tkUX6s8hwuAzdzEWKrPc243X
B16p6JjoX70VH6a51v0beeHg5lhlK7gvtFUgXWyeOuF9HR3lruc+BmPOPZ5YtgxgMRPIu8RTp+X9
j7yn7PU0n7ymqBGVjerq9QTPVZTuM3YYVuZviWfNnQNVgVBDRON3MhMwK0kOwUGyQ5iAaxXBkkB6
4DNz9W1y99968B+o6tAKt0NUY3n8NnRp/gw9XiMkBs0JABhAjF/0NirsqEZbOFrNhyGr7Ohvft6d
7/fEDdIskQQ1zwvWtrPEmZkmjTcD5AawHMqBFjXaIJicTlejADFRoacH4zSuyRUdFU+F4dWFuSZG
HLaycCXFryPISIrKBb3tHtSAq9oVH5pRE4bK4f/cDsxK0GpGxFOxK8U2weDPpq6GNHgYHoo5qE1M
3vtrjW0jGSGo7uNNLPmCsCdPNHK35zG6dvFO0EijQ19HVhFbl42nQas64RhdBmoRb1wob+iMq/3I
ypIW0MVwa99GW8rYxy5fi2JBgLovVngxSWWXq8GFWS55Sic5BcCjfI0JsjOMA72haMHG8+zqiSrw
V4MfitGrNRcX59fjbw5yLUwTHupTgwapjSfXVkgtN2CioH+pULnBC1S4cgiiCfB3mXc6M/WVBK4l
eIIeatHuLAiLiWwXvj9nwlRszMNM3esGyHYhQ66/S14e7hWCHdFg7SQlqoKLcNh8AEvZQlPzvZJR
i4xBzYBDzN9030tXQm4HM3Y7fkodwpiPdYeVwhvzYqOSQ2IyyrIGXl9UuJkMqKX03vsMkWM5hQi1
maP8YEzJ9Y7n4OEOK6gshisrTMKtI/7ukgqgh5Wg+pEA/fmdpFUlx8c3IlH7IUgLEDECWfERPfFi
kszfPTx9h860QFLrXHZZbMxIFco3DHIn7mNUCpzjNdtZmoh/mjJxZHItotxZrtJqJAdVhBMtOWG7
InsuyN8t8de5S0V7wfY2UdCEraBUr5eIyfxpcq/A1Jv3ERHSjpw9DcGZfT/BMmdLC0YEHatWGUX4
OapmGUrjBVK7tnuCKCpf8k6Ki8uSwbGkgOR/r/tMjQ0cYGu062Wqkiv+78+LGt+GrpgZtIVRwj6v
9lrfZV9rRA0WnYNYJeat1VvgZ/nwKTUiH1MGEt2QB6NPq8frhBYEVRBhnOg97IHdUJXMw1LH/gem
N3xDu/FvmNqiSUj2GM0x1F3Jwai3lrqsFkZBhjgFACq0a6sf5huEbOEFE5fmQv/6VE9Qizd+ZFiC
9DGjcftzN1NwxpUgvfSaQJABammx5R/Y2kSWjWW8ppWP1tp1uOKngSmWZD5UQ3cX/bWvJJ7FVBlk
fiBfU74VMu2yJZdZI3RHKis4kGUv/Jb9seFVmGircyV5SdGBI7A6z0Fl2YaMQZ33en0SlTbK7Jg6
MiWwfCPIg34o7qnMGTXkcIXCBsCmyK7P7s9G3gvNyth+UpwSUxC/0Ghc/ZkDGZZjdJVd3M6Z+0TR
IvSm4TgxD4mjamPsLm9/QDypNG3bc0HYUyWavT9H7Lznb32vzVAmYfOqHnDGmYV/fezq62RKdUJD
/3wIECyRHkHC30UvU4+S70Adh3JOvdk3WmdEfUPIdtupETGPRG5ZJKOSG1NaN2IcyikPPKuoOREu
agLexbY0pFEg4uHaUtfIQ3048nqVYKo9aSRB4jX81bQP0d0gjv7aUKNYV8VlB5WW6h0vm+qRSKOh
ML/aC+weXkUDiZ8fSDPM1yEnW1OYAgqaA/qOVJhAwXozRsrHKQzu6JVfDjWL/OqNoWQNlKvPaUtn
rtA+4E95fATmJSGQJ2LDXyJF+22y2Kn0qZXfRQXS+2fLqGB2jYqokegAqAi34Bg10d4F0eMTHtgE
M9HqgFfTQAg5hgnB0cj0mgWmfjaawLiPCDmFlcrl0MeolNrAH5Ebu0+cspjvKAJNS4Avcf/uf+wP
012BtMSI00499j7l8VocW+7sed5v/GOpHHQ5K1HCW4z/TvewVviGIF2Uo2t2EsbYB3DvvAkZMZbR
ThgYcDN7onDor7kF0o5zRYQzPzNTbRLpquC0ajQJoBWhFB2ThWgNwR9geqlpTXybM/vOjzkO/pys
TUFwFAddE4FVaKgYatC5UgR83RqRfsVvRYt9UCymASY7sQ84atMQ3WS1gMUhmOY1IzJDRQiEMJUj
dhRaa+bQ955TdXBxVh1qcmh9w9uVHjwYrK5qtNhfzcmJz8bJD/4Q3OQNEIZH5GgoJjfo6cfQ42ai
yWLhBtf4/h+qKvw3Mn/53tfqjm7VDCaN3/2KFkQMx7TXQMVK5ME/Mua176cTinNQ9Pkt84CSdKWQ
RdEobHrARmowLrGXUGGTjyu8+niRhFYfLz1vC+/dveUdsjbcGrce3XFL8Wz57ruz4L77xZC1TG/7
oW10EPaSNj1G3Hw5KWQcJkHt7etSYteCHHy+YvdcV5AXRCUA/aDXanWnZeAkrMcDo6FjOp+Ywspe
KdQYfoWGLh+s9+5HdJUCRPY/l65hZOy9XbmVZDescTMnDNVA26nJhRPcjHeCe8fZNfYLDGrm0kb/
UOwCumTfVP60JTrZvXAwWgRaVt2RXRHHbgQBfpq9Atnl3VZzgmajbbYtQ2Lfra1xE2cfvThWgkYB
9gKSG55bOkukzvngXU7uWe//ke17VScrRdsL/JmclmUfTe0l7p+RHUHyiZUTcatRmPvx91BygUPd
lTEb/xRu1Nqopx9df4rcRYrCVDJnBrARn8KRGym6Ky8nH2KCMWUVRZgGe5kmdQ6VvF5yfAIdcz4+
EXiN2NsMQsbDh4VIzNDdiCBTGE04x/o/qTUTF0CcDEXKRbjTHHxHFbQ8XcMSg6cEcnZuVvi/9aj/
AgSxZ+ZgzovrhS/6ZnjArw+tG8Qme+rIn2Aw6jW36imwZXx07K85Egmq2wixTGCyktmSA6mSUhV4
/Pa25VaR4quzOfMtkYj5bRdD4Xq1KpV7SFurOQ2mt1o3pL64fg/UZqgh6JJTl9Lf87jbSt5R1rpV
XmTjrw6V+s0XJ6v2aNYH6Yy/+cWTVZmGl/ZnDeTxIJn2jWPltNSi4HTqbH5iG2vOIaW4REl8UHSz
el4pXifB8wnNODqo9i2hNdyQg/0hvf8A60JCR9pGBne6W8G2k8ltvL6qwJEjU2Nw28pHmCuFkr8T
ikr+VaAE77YMIGZpabhoHz1WzcLX9ey8pVyQ5fV3Fx+L6/ppPAxqQ0jDKsKOTePl1cP2wAG+LOKY
YL9ujufvUlhYbdZ+3T8Zo2ShqzpHIZzguDO1PgtofxrBEQOHRhFrOVjdBWmfDM/DbijPD2nGUW4w
bqgZzVUQZSE4BHyfatrv7szb5GNcH3TxEMVPW8/KbPjimfDzDy6J/QQOHgGHJUk2Dra3oTGT8w7M
I6WT63+Ucyh3NGtq+Mznl6XR9DK4UvZ7VB3rJpsnD4ZeUcJfzbganwq7bIjXDg4kBu7ePRTrV2UK
OF1NcRB3yKwGJdQwKi3WuXpVtGxly4f3w/0FTfpRlZXWR9iexqny9/4DSyu1eivoYy4OUOQTbgtC
jXimFPXHvaFjM3pYvNwx+57aQWIQhmui+jE75uB8/MJJw6UqCNWf9ArvIREr0BCCNrBp57cyQYNy
a7EyO/H8f/zcUAFE5fEMdyhZd6UrUm7Iv6q5/tGYfbYwhz1VKdcZIqr4ZSjlCNFTEKRxw2cmyzep
wwmdOGmodECWbKyvFLneMKOmbEfcN8ddI+pQ+EkZ1MpWjY/DKD+/byB9P6pGBWI35PNwFigF5jbn
Rl9maH/FX3dQGYopZJmZR+t903xSj/p3de9qZJpkqHLQBuA6/DpJe+7pW9zrURZEuYqYAaTLoMM9
qIr/aW333/y4KSM1dbNh4Z6Sdx2vVgyI8mT1MQmJxorg77rK5u9+9ZYgKflk4nFWQGxfb2BmiNvG
xLxtpO456r51nejyxPhJvQ2RBfGTtGn3GJ6to91/BLQaACUPyAMdbLeWwzNrjYuhyXje2f8DXH2u
c+ECQQFXt24ClQfj8xGB3q0ioj84O8JZclyb7tbUJedJqdPRXSlQHDeWFiQ61SaZUB0mfUYULHUh
qv13aITmvY1iotRj9He4ffQ5UUurLkBp6TLm23uOzYkVoJDHub21GCv5aYEcG4omyEftHnIwpf/1
6lNUpGUF+20/XEGNVb98E3/tpyWmOUOVeB9SggMjuI+sksXfKFA9NHcYjRKfk5kYFARl4etVdlVB
fdwtu1BMHyH312t++R75tVh0CqMdbJafT5DjL8MntwlT+r8M8O7HO47yvaCpZQr0SEK74Q3196pr
fbPmWg9w57AhYWLfXU5qC5JDHecDoz0v3xFxb4EdNOTPYnexo0JDPUNBrue1ypFPF1wJwO+IgmgK
uvBQpVZ7QEAbtpDv8nBaANoNIl/SJTn39u45xJvUzFgIzsZmcu9WNnFZ0NmXLTiBmn1hAEdL2wnJ
0ZzStK5ZqmPD/2nEq0s+iJdmorkMBSdM2Grq4lP9taH0MqZ6qd8DFINvA837ZVFeFbuY2KlFpr98
TNRjBrPR9cyqLNHSYTVfc/Sj0b5f7sNQsCiTnNRJXgEJS0pB0vjY8D96pGLJTj56fP1LR4zniV+X
jfpSAqzNs6n037peFYVeFPiI/dSOlfT23fYaRO+Cmf0VgtVU3wdTY4+Rx+tkBZ+bDA5e0ga8oKLy
0A7jH/vvOnr7dp4dfZ891c9ECgNkvFAHheYmwCyGakRX7Cs0+n4A8GeKOyun1HBBWXkKfFVU9c21
H5LymzQvgJDaMKOz+SoDxVNQtUZnWX0NuHO/8rgzcPQJIZMs1nmWYFLx0qJF2M53hGghdBsisF0X
aAolKfK0ZyfNENTolpPgR3wxP8KjuVeksJaaIBbipdlYmdPjsbocetcgozUpOCBg8jJPakJeRnB4
+quN/PoCqWx/e5XJazNHkbdlJnIVrspupMMnyy2Cie09Z/xd8NrUdGw2NXKyf26a1QuRhixfwrId
aAPFwJtT9uYcOUBBtT+KKIxybc1mVwnqRycs9TfF7gDNgdZ2zhPOrrQK7+UPGf50wqqADVL/LEJW
k36I/ORQjhBQ8M4UVOc1O57jj+8lyklTlci39AnTr+Vs4JzdzwO1oPp2hi5PpuqiSxSdRZWw4GiO
mPagWZeUh8i2UJF/xu+0rrJ+NZFW8Nd9mwQYDuQ9/F7dos7xROMIb37japujBwCwzVJTfw1vSXSB
C9V+sl1luVBW+P0dphgbe5kShGiBCW4TgGzeoWYqjXeSI5C6er7uE4Qo3gmqqgzycGU8FG1oUMtV
I0pgLxR32VZ723yI2GgwL1dLAG/IU2dFcR6VSJJI5OSLYscenzeHFilq0ARNwOEAeiK5ICj03Xi8
L5ubZTOv6Mr7mU1xelq6qPagzBxrtF3NkKVxZ7LznLp4BPy264atRS6MW7MBfMjCNjLKTUE2g6sc
6sfDXhArc4zslL01cQ50JRjdJ1Gb/6VvLnghQsgV+UboHDf8ix8TsjIOgztLR1zJqqGBSIaictnl
5mO+yFt5LUFgf0dvdH3ojNFDN5/Fmnygzif5gGS+5rCl3C3B04H0DQ6/speIbUpMS0huH2SYyUt9
BU+eK0i/PcafyEJCKjJPZuMFNVtfBmpIZOYbg8NZeGzVcclUIRH+/yHWsQ84AG97Qmy/rEUnyQBT
Y20gmzb2NOMAlArBxSf3JBsEfIqX12oDpGEJmzxKw8WaqJKund0rhEytpmFJIOOqFL06iAeWglwr
P/Tlb59wMNfNwcUF8zRm6dpDP0PCjutaBmVlaYF5PCcWltL5Es9/IJB5ploHRddQbZw0+CJ+Al09
H8PCecTXjN3CHG6cIs9fcllvSDR/qVJoeeuUV91sie2ZbmJgYIX39RgaZk/nrQLW6NzdNd6+VDvC
1FMvqHkoZnoepyiyNyQi0JIxF71ccYI4JTmGX2j2eLlQokTadgbgJawNcRlojqLEptY6KwIgkdTe
JtTKXYVprbhQmdAJdyfO+j9PYUs2VPFCe0O/ZGS84pWLY9aM7RWDwDA1l9Z13hZNY2zHWJezDMYH
fr7WYgXt/7YQUmIhO2hB4u4df+Wk2kBY260tD14hRy1EjAthYHYCHpQJZ1cEO7DmoKDPmTeut4Yr
De9Hisi1BvLQk2jKapT3X3ksSTbs/YjCgvMS5WphGqmVBm+L406ZWd4FeHzJCLhJfy2iuMLOvWW5
TyaOnFZwDvDhE8ltSldD2S+jeGT+BMIRgoGYkWYeT2nCHwr+AqHtj0i9Bx6HlNrb84sFZgUqYf62
wA788zoUIo/rH/ahGcv/Zxm4si4ud26trrE1QZ0L3ABQVCQYgu1VcLvk9arykv2X5gXpbCsJvW0S
GjSPBtFIt7iVIPQUXJRp0BGJVAvCtLEPEJTSaFOEF/ZKeafYOkoWNxWfWbC6L7vj42W5C2KR5bGa
DNYrg6nA1Jlp4q0r6Otu5d7ouhZFNLC8ruB8fFlThUpZBBAuKqHpceJCiQeDDOLzKNukfi2EmRXe
pn+Bm7D/ODM/6fErUnhvmVodTlgtIslcQ/XcCfAeEJX0aO6yEb/CdLPGw1ia6r6vTd8OxRyustRN
KNC+70E71i0Foz1MiLhmVbYA08nOF5bF2RO4f/OadsEEzi517GwciJMLEfUwFdrDMSdqdISvL/n4
6zaXf1pmAHKmRilwAUj2JTmtCj83T3hbYcvVIZ3yVes/vZeQ6eLTHZScU3n84FGvnPuH3XttKI1I
nRnXiFyyixHlkrEpcTqIPKSFlwEFj+FKbL9zQLhVUv4Xma3El9IIqrhJ8bkRZXKq1L9Rq9Yr5aOi
272Aqs6kgOW/64GeNWkaDGdm4WfCU4VUuXqJ0ZAWNjRvWvB0yQ4F6fckOrH91bqZuP5S+eK79kkR
D6rxRLkoErnJkbErcOUfkwHyf49HEM9RMtRgIhZcDfyMppS3UcKLU0Fo+66oW46xLObwS1Hk53NK
UfMBtNpsmDetUNYQ15Oa9lC/+kXBEeBNuUBE2KDLiS3krI1LOh41zRWzg3q5LT/M90YVETUu7U31
acDzoYK4dLE3L8VXWGvebvyR9i23V4TnIf3LnvU9LNMiVEWWka6ohPvu+FNo1eRVqwH5RCCIjFpB
P8cFNT6A/0oZTLoXtkm040rFVyJk+oBLd5r5DrTwmiP+qj2vXuFPJVw5XOYZ64mYEXr85ixVdGHe
ozDkUpuNmQXQK6m9hBROAoVJ5vw4/+QoUHzoTgWBM0Z/Jw6Jm3Fm3DTOOlnrG0LYWrZiNyvCHPca
ohm4jqQ89U3pUSasuIMoHtcGJOvYhmPphKDrYaQKG1PdKgiVYz1lgosp69SEZUXA7/YuKzZ9HveS
1j3ysrZ/zFmNQOWx0DlTn1LXXErSWj9j4nmyuz9SXoaO+MnqAEI4vwVJawbCrOok7D/+mLbJJwNm
GpWhtVuNfYb46oX5Nb1L4ML3FP9h+JHD1zWXi9wGiCAn3xIiiimdYGp54/FidebzzLrI05UAQL6o
zck8IlP2la3sEl3qAikWiaH5gbr6JszfaYRIPEDYs4P8xDw8vuEvPTz62VNwBN54X/4uSBmaIjTn
W8r7jMAfKPuh6WCh/DvEO3Y1kdMD4ZeAhFSyE8+1gP8sPd/IfhRqUH3YsJnJywjk3ABb0zmHWrCm
36jmwNYgwCL77KFV+RlwOaS7RclQPlPblahQx9qwrd2eQ4fk2A7AgmZaR8aphV4akKCcTVk4l11w
Vpl7mPLMWBncaUyzb0mHO5lX5cOz9y+JjdQVKgT5rkqIYBvxXibtp1U4jfvDxYZH1uS/DLbDDOAe
zEqs5kEdI5k3Z97y/rRQO1QOdxUqoCDNJpeXSTfwRRN5D/6apxAOyTcFgRJ2/rKnwiT5dqoor7BV
WKzgxhfMKYHhTkYGAIpxULrbbLkg5/Svs8s1zgDl4+qUPdHHGoBhQNzajiRbzusHWTj1fErE+b6g
psvh0zZdZylvRyU/PhE/459raYmjGIXYDrGiY8pmVNgb00Z0uW5IKD7MyBff5DzDggOyri9zqZyn
rkMVT3DQJ+JZIScpfuFLieNELsOZ6ISWZN0HSBA57wxxG3m8ZCmhPoP1CqxDwbKcllyB8KABREDf
pIqmJNRekdkeb4prDfQTE0hoP9nhYJ6Cj9cnWgS/dCOI8uz7xvVcf6eEmMsAL16St67Ba23p6Lwl
AYstW1J5PhJ193kiPENfeqz6GFdZzjwnJbv2niNQ8V2BKbPNjd+jmNgc5QNn/VkpL8qrP9DvwEt5
kbzQyqWAgijcb1fGwyTfPgr8boqldLduPZ1Ib+m8jq2VewTeRhJMPPWrQKNODwhBQg1YoOPjS2WU
Owgouq3og+fMCTGCnovI1zCeqDpXk/jIq8xvJCT/wDlt76biTQTUXoRqwQWbdQRduL6mwjfhctAb
NGdPQZS8vpxEHlTMo7IOBiI0Jegn0wqM1E4UfsdPxHlY22Lh6uXT6crGngL6BzsBZX7fN1huStzI
VtfrKQ00OhjSlvQ+AH1cfgvKD/U/zpbGQlIPqEN5rHLGkOuhtmXRI9g0ED4SdWiOBXvpoVhBE7Ju
PmaG3mo0LqeS/lrpu6221MjeuH2byymjX/HKjHKLDsXRJkwtmawGzWu+MCLosxSnJdcnWqiGo8BY
3LS+CXTOkocZmzNNtPbWoKpu6eLw3K/WsRhWXx6/Yjvi0aGvgg90HQZ2bDDxwrsIqtxTR0ckQBEq
fCXFEFLmr3ne5KgkZ8SEMbbBgmINAa7xecQ89inu0a3sKqmvgb7wCpFvIzD//yw9ElJAoblXWZtu
3Y2YiDO388WqPMlBMsFo+IaqMx+UFLlN5yhODUFJfwhAPlxckJ4IKEkTy/V2IhllTqPN+nSKMd4o
r6YzHeQIWeFyedPGzW9PkR0YP/BjF6yvoTBxCs7/RlJ4QaphKII+BC6hm75Lo6GycJBwaGO/VmyO
qkk/s8tviYlMNcSVAmDF+A5DhgLdD1iKqVAg4AjLt0JgreN2UNroY57csrS9Brmqe7tZp0g2vthc
fydexZ+Vzezhzm5gYRNKteJ4+OlrgPBPlkHSKjG+SD8PCWBop6ENv++tYJ+pn2YLC4ON6dS9NXl6
KRQFvDOaBJibtiGEi9yE5XhtgN7ivFY8B/Glns7XeUCoabQ6WBOZmh0kfeOuzpOuDLLuu4mQmoZs
/yIXmf15G9bVjldDNl7IeIPhxnnQaeSF8Wqav2Q1pxKX8RzO1bhbB1vyN8HdRVUpE9XfjxiKMvts
R3tIMPr8/tMHcRUIixW5RRD2EAQK2Ncm5slshjADZH5Bdsdp1FW5Rvla40UKWcm9V6LCxU7vAlgn
O6bAI5TaWJGnqOJzTc/LhBLIl/mFOBOVJoDkfNhUMziQUu5eyWk4AIplNZZpubB7LMrEVej4tcqf
VSyrjWX/eMryPxmw35aczbCdA/41wcpK1XE05ebyc8ZuMrEXgLvPAZ1Y4F0RF8uLhYh2r7tY2Lgz
lhRuJgwb8DNubPhcTLzvnwYMXwKKCS3EP1SUqLD0q683Bn6NmStIK/LcqOv40KlZ+TnC2e32lDDd
I/UbV3hAwU4gItx3+hB9vCBvlw7Xehjh/jLhTejxx0rqovN14dHiblrIaraEGOkmd+o+KtQfmwaj
l4uB/Qqpt1D6YNrt4enV8Xfqt64fS4wb4Jqf4SllvV49qhdBU4BPY63XjCMRIpg7Ht4CZaC36aCQ
/rR98LbP4SOOd3uQCf8wo+ltDAmSx3p1hmN6V9AQUeGLCBoIX7piIXuUZhmgQ5YGQYPziQ+TNIUy
5VRTg3xvDyTI4zdI99n0x9UoAf1nbGIjTnLTag1DJd78JY7woman+OLGSspuhPCJ7ze11PNvlkM0
Dui/7nCxdf7jOSgWce4j0lL8hHOEgS2EjIKFcWgL05jsRYMdl4bhLuw8JBfoJ5fAo98v96eGgDn8
37pUetUsnXPxVOvsvYZIFQGWVK8vzYjlmkTzeNk2VxiL/S+uYfo6DDUqIsN9D7txRpWVwWK+Cu0i
6v/UTLl7aO0/1qsiyEt/FrT4ajWyUiiHfAxw6yKSIKmFXtEF7BzROpXL0g4tyDENxPTvVgp8xwTL
rK/MF/dyllQ4NLgfgByfXKGJK42QJaJNOEis51kt8R7fSoo97nuHhY2zhbdQB4nd3CflzC5WFdjb
xf49tWNL+1h5nC7KvPioU+CYBeMNZ3avuxpaDZOrUqRGhamNwAc10zPaZPLbACwhZZJHJd7uhTTY
ATt6L+VBt4Vdfr23NsVP3K6xvFKZ8H4IMxZExozGOoZGekW0PL9+zpD+qQlAZlnUmCz3MKhiWei7
ihf/MM7NV95SPctQy9bEqxMn5/wMl3b1DzTbykhbTfyTknzzOJAC1P0+ixyDolchE/N7VusP1B4h
PCHTQrQgFceXpY5drV8IdlbJHdE+Q5QIORC9KsYoNnePhZrBQZjhSE8xZbackpElKy/JEk3712Xc
aQbh/U5LhALqBK08CiKTlthSx/oNxoCWyDZQ0Lagh2+PsSsuvm70obZuz4kbKElCJGReBQkAhLpA
sMYtN4OgLany3tQOgd91W3CZEg5oj/QXJC017GPu0+FuHfPVM86qnfhz32USRaEhRrppOtpJYoeP
ar6ePRatfvv4MVRVjGwzhbtqwEwrcxzwAKRCAPSL43mqHN5lMMYDiQ4Ay/EkD7XgeL5vD/SG+qVj
1T61J9ax5w4hhtp6XqqX4pUjnssXJPB+KQ60OAZtd4fJSv3Xc+BCyXXvRwKNg+2hTLwnTf+65nzI
fumBPL+GskfznhE6l++SJTxpzl0uzyfLeL1xBChRdySyASvP5f73aZakNOe5FcoI23kWgxd1jzqZ
edNCa8uaTBQBwcwMRKyTRn8OW79I/z/CYlOk0s8ywYeiGOIV/y4KpDDbgfWPR5UXcGxonvJQX5MP
y0qnJnp5XCBnsNoXRGn96xqCrPuXMEcy067CzSYfGaUuXuO0fUuhpmi5KwjRQPTQFGzV3NUGr6za
sTyfBzpZaYhF8Kq19df7up6Ot1J1NMINhnFPxYV6bpLUpiSwfNxLjii0y8jDqz5AwCL87qASMfGh
WVHWp47PmgRBE/iWIT+v1heLshogL2WiEy3nkhRJvtIEYmUP/xVqOiq9rF+wdNj2UrzT15WHZs9I
nHrhCuBQgKvStFroqKdOQ1JkAFiSfubWiUt9f+Bg1qK/YJloIA4ugg8kyEsx/zUXD/mCklIqB33v
9fmqlxVPnTEt4b2mMqjItuMJtDow3bL+SJ+gr6B3cLz3998YoAaGKCW/jFEcFgMKPOvcKrotP9p2
7Fxq4m8jdoEgwoLiWgu7ADR2TFvRwb91xDmmXyFYA9/Gh/R/68Ep01evtjNVgJXqWJ2L+OMMN3WG
VUijGs23DXAxwJ4Xo9d6pEWdhE2fCQrK9g+U2lzteUHsLP5Nqyw/CUw1mCZxnJuVjJVyHCwfI64t
z4h1OVCSci5KHQ0RIFDChY594ci1hLLsi1J8jdVwRFJFCs87lGbMVo0oAzalt3jhPedGsBz6m/IV
a1IGMIaM8xRiFatENixi5Adn2s4Y/F1HPhCJ5ju9/W6+vdwb764dSvDXpJBcxj5LDc94oXcrKcN2
z2TA07CCE9TMUcJwT5qhNSiJz7y7a5YZNZV6iohzmf0gNySAvP7xvkvGyP70g9gCxpa3TNQ38Wcp
L9tDqgQG3kJC9EpLlm1s5UeqwSW9uX054fqUyQ8HmET+lZZCcp1vK61gDokiUGU19IDadaTOIggX
BkHEwOjBaQ/DbJqavEBn/Au1j4E2g1SYEUS1who+U5CgUErXzHW5D52jtHDIQsEHD9DuzI6PMfPV
Ge6x+laMvl5S2K7LrnJxYkeEtFRauTVrTzhAeMMrxhAR0RT2kDISRXN+nTdz9ReYsBtCOfpKURbd
+RITkmwf4wv05rTq8eoDn6ciSkx8WyBDrFAwOSQ+FxbGiv69LCkiEFriw8CsopdIqCMYmrgHLzTS
+AWHunn9Is2uieUH+Kz+vVO7FLt0l3cEFCQDQWlgcIk9cAtg/iKMQk+x+3zAaMtVa0uAKjV6qn7a
a6i7ybwVwJYq8JK1Gl3QRQ882UUb1flPlK9JumKv81MeqCsxvTZ4wu+8Mi4d8dJFSOuM+Q/QgaaW
lsWztlvYtAsKVQoxj6f5qlcj1mRPecASTDyIjUnDwaMpCXrbSon95HQ14786/MkvYft8spmEHjiD
CwOom1wI7an+Xb7hfDi22CYcF32yEgl0vf5jQLR3NZEHYFq3/Zz3fa/P80nuSKdFMw2mRoaQTTeq
T28JxLl7PGcae4osSHuFAI0pVAHzh8x+zBYsiMzLM9Uiydpn3Avf5L300HteUR58uxK4uJ43vXkP
L7tnkvNgDriPpFekMRxBp7+rHfJAkA1s/y4RTYvJXURxZGUvEZb8xX5b+eB7IgoYREmaIoCfyAws
clciU/lqr9/Pc0/bTRsBxiZ+gn7RQsnida3jJKsQBxK7N9bnqKU+32PkdIr3n45bkKtBx8AxjK63
JYTQbGp0sxMM7IdVG/SxKb2veigcQ2bf9gcFnGCDYazRymqsoSZe8B+++ha4OknqHeTON0LXb9e+
DBecNarWAMUJxY3yiQniQJxiSTzlMRtU8lOfxDiroj4Zyxc5IWiE2TdtR6Xni4ZzpR+GZKLNqf4n
THY6X14UgYVMrgEY2v9QX9xU//mB6+alCskO1xjTa0lrX5bcFlUGSnHfeTpIyXlEbmGYRWFZn44Y
7vmdFG/YVqNZzPBzc7UsaHehYS8UOn2iLmOZTkxgWKfkWndSrJdTnnsPJ5w1xgzhxAqeUpgX68yb
t+TbvxmohLkCpqwFg+BOcUkz83ygx0ODDMk6ZKim4ynDCnqhs3p9c30UXQFiQi0cMBBAvsTI8eLb
3hnsHMA9q0jnoCWihq/taz2EX9wv31UothwMqp0lOV/1YLAYL62ojKF+wiIMA8+VCqX8jQpgVmEw
PJb1VPaPfdJi0gh359rpgXoS3WgE9xAzRKj6iDcd8it4OEwD13WJ5vxd43TnVqnabkGlELTttlzu
A4Tph9/rf+RqU8Wc5R27EE7MASOTv6EFFHOV9xlZGsCM5nG17RqIDemEhybXlVd6b++xVHCqJ+5Z
SwtujT9eenxmxtMjroBuTSZfuHpgDwv9r/4zGfvyydBRLPBnQ6P8dTOXLj+bBArW+TTDTH/LSSpN
doi7cNb2xmjmyUOwY912DvEUZT7HlFw+lFHPRmvSshsR5Ce2enT+dMuGIXY/PlK64mKfJjxULXVO
y7KtxHgIv/PNeOGy5qhpK7ALydeZ7ET+hjbNnBmJEBsWGJaVUSGqLkNMKYz4nk+Y0v9k64veZQid
5PGMq2gbn8Ae+hO9MXa9BGlQCi7or7SVLZQ1cvTKtBY8wu6cukRcjX9S9xpUsrP6/JYGn/Jd4tST
l3iVBTKb4Zsnq4a9iQ+vQzLfE3Vnaia1jVMZC8jPUV3s/bLLByhLiD38UuOULpjG7Z1NkMGC5uvE
7uHEtKpHTP+yHk27nbEpyeG06/57QkLcm6Qg6JdhmyDbpamAe4jXji0kuKk2vNR7baQvhOi58C5l
amlNrJOkgirL0fK/iyVOUbhq/3juExW7sw8/mN8KvgQn3o8RkA6s2kC9Wx3BMllOYG/mr8lY+cXL
tZxSUFNxWDTUanxrAnT5m3LWPHzK4LMBS306LQgS5rtfqZ+1eIZNJ/bcMyFbms6Ncb3v8ndlUDUG
cjouZbAJs7FyNk04nTL5NIczGBie5s0wQQ3hpf3YO6w3+GM21pFnMYfNCxx9ESExPmVKOu30NxN1
I3XiqWp2Thbb/Sha1MW8SszObcXhm0qunW6eSqmilPsBHW2c/4xq1VJ5Mpr0IKEsiY3M+rKNSV17
BxiRW9sQXUlyGABJ2aVr4N1bihA6a703CuwQ574g0FGOf5jG/MVRqGHoZAcEAejxJfvidHxnyzDK
X/KkeyWTN3JUUolwL5RzBfHWprSx3GSkOu9HKIfgL3IkZCobOz9Fnk6y1ZgXw3eglbxhxALEe8NG
2CqPH17IYPuTUqqw2idd39Ll0M/5i7pA+7A0g5cbbnu5sCocXOwn9wb2sFvlPtYSBv5Tbs3wXxz5
b6TS3TuFV/41zr28ezia1sOV7DeybdAqwPERszCmi8fLjITRCh1REW/C+y57S5dls2DS/8flLr6L
fMs7vkBlGH8mPB3tiGoDlXR+EnY6V9fvO58LfO6X3s4lO/prirxWzHxbPjWG5FIKn4b8OJ8ednS2
D2up28VEhBm1qSTva8twFAMXfIsGPSa7kCnxtCjrVrZ+RbKGwGe+IU7W8lxi6lHQbP3+CdXUU8at
bJJL3e4jlFTz/EaXHFIgGL1zFSey9QdIcyQZNLpjC4lebbZ4QdX0R6fv8AN/a9m40cT0J5CGGjTH
eq5Oh+ZhH8bRS/Dnj9P0hqDOQifiM/vBmQgSlgwf1UhVe/H/uYirSYRUSghcbi//rMx0lzTfkLIw
nX8cuNf30lpGs5KfXjk9VTGuSHB0nz8YdpMvM0L2MP4gghL7KTdmCmOeHwihwNZJLjBzlJjDwH8l
RiK3o2U6sO7k/PXTJILBolWyCgxazjPf+nBIwxlZw80sU9WGT1El3UggbroT59WEWM18UylgAFx4
d3lucv3P5jbkhef7cLZv8znzHjRtPIY8thBEy6i4Tk+yDtwG2oF2NcxpPlI5hSMFRPXdXi4x4UBa
IBQmxMzEmxyK1GWY8GF3+vG5gpT+t9TNFwB4/qd944jZxSONWmkux7jzl+BVQLGbekHRRJ6A1oql
DdCDjkUylazonbk4uKDs/YeGjtiKmR4Gfax3T/Ewpzcil098mv7vZuvRVUZJu8rdT6x+3jmoA2x3
ia2xDPy7DRqi85bl+krmIAGcLEwC2wNpjOYgowinnNLt05QzkFJbhFIPLVnT0ssqrH9K/3uJ0GY6
WeeCBDwCaDTZoMa3NQfpsvdJE16TnchFVbnzPtNxAofTp6gNfDrrX1c/vaOPFpQEN94YLpFa0VDT
pmPaxmYqqdaxW1aeVIkmR2bAjBa0wptn7llYvj8d1CqPHTaXnKR86WxNjXJdbkboQSbT0ILSkq/f
fsXRM8NtDkCkUjnLae3XwaizkDK9FAmQD295mgqwfyZXREvJxtSxbYQYvfu91Xw3Cg1y0yI36bz8
KE0s98sIS4SsA3H9ipTcawMclgIpbADUE39Ap0Bk9PUy9GflhW0aeiml1siN8W/VXZYisOgx+sLo
dFVe8TF+AzrF0yNJKLPq1cE/xFhFurN9L2UinGzhEhu7iDmJPn2e7nuL7vA7DtnjkdcKS6QUgH+S
1WUes4xaSOH8dTArYf7Cw9prUjXxQ/mjUaDu6NinyN2WLOH1m2YasujZ4GuNcWNZB3p2g8+IoefC
zTv+xTtXrRCnr+TCCOuXcPZ1apB3G5rmKO4ebdsoIU8mAKy/hDdUyZ0QzWJYbKuDNp9CxNJgIf4L
RKdOTcBqEcILGRhk8ds9o8w6B/LuhHdX1X4W+JaS1lkfSLtUWdfZzjY/540w70znw7YtXh3SYIoW
tFXmck+rAYO+rH0bZVh9U5nPn0ovcp7DmSRBV4AF06ZwYk+J6ZNXdraLeXTTzH9XfqkZT+Wv6MYI
0hJ5S11sXbO0WpRK2vyqDpyvnJPLgv5zvWt54iiq386c8NyG+SyZ3gvPVFeY2Dhq72Kaw90HjA05
KsU28BdoA1yWVlMdIeSyRvtgHU2yjBEDy4BK1yu98Su1JWn6v87HJn8geGxMGndxs2NvajBgzHUn
HPEvtbD/pYzqAArlLlcTOEEiMOqFb+WjKYbxAxBlGW3DMN5k65JjqGlH3DnG8KOeR3+PnLHkZbrd
vYXiAaw0VtOt2Hbgthcn38NzgMLNlndoleOHQpzWdvZMJnXbwWBdEQaDNbfwxVp98KVdZXGlP9yd
aukr7oc3rbDrs4sVQXJjlVGYWhCpH29zJeV+c605SiJrI7CKWiU9IMNy83u+mdgEk04roGUVqp4x
R3aPrfAtzAAtPFzC2vfKmfjr7CrSgC+8QlpjYBKIy8erlA8cSpBZL2Tyz3NTi2UVRPf8eST1gksE
kuHydVuJeD9e0Ga7YI4GFm+3V7EMRkvHnaMXW2PtiYOY7YALDpHAE1jGW9pLNApap6o58hzt3MUN
HwZZ73KtG6wuynGmXBB1nZ55of7iRLWrC8sp8zri7FdnQH/NuBN/A/zVbbGCH1IAhOXUrCj/s9t2
gQNRBV40JQvgf110Vr1vS+BOLpwnwCCgidH+xsxe5KGpaMsX+GNLLDbV1pVd0PWfxetACJW7jqXC
xUTiT7zdiAory1V4WUUIiFxe9Pp+rjK+tWo03el6MwbEtg2QKWqcX/dthH6n99SLKzt6py2mhsMO
hOhXfCcb+p3vocNld5ZP0clFY8gRp6lYMsZTRQu4IZ5eZs0s4q54X4/B3JfItoEKaZw6vS776r8l
aecHRVinpJEFxUkdmgUT8i6QMuK860xMAutNxoFN8tJuJeDrWwcy/ujV8A90TL+zqr0voFHdiHRx
R4pRpVQuckyqsLYtL6FfEqPUvjtEWixVdLbjtu1Rr9GZ0SIpil0t63vmDlLBgfwsEcTvS4NM9unY
SeQEFB0hU31vhK+Z1CmC+xf8hQGo388M+ukOsCMOMaL0vAoWp4yNVR0cJHW6GVNWc6zhsaiJ/4Og
xytiRPqb4hIHDUYltN/H62h4UPtE/9kvcv6H9a62eYUE/kajBXNY2JEFpLcEZkc60GuB0OTThzuj
8O9ubrC/A+pqn9ndwtwpIb43b2vd7sMBEGHWOMinCmVgMBK82OCBECZPY8Kg8yWkgZaafo00rmFr
UU/QGys633Ks0Kz5L9TeDA6Nz8SmdHT67ffZpJjzI+fEao6FjTbpLpAldz9yg4x4lNQCmdw4Zyfz
X0g0AvOUyjI/my/bkb+L01nBFQDpYl9CMTnqX37/9D5wkKCcDt+omqZsHlLsC/VWYhXM993hoCER
aFLflbQu8e2e1zj6t9HKzRD8FBgfMWS0zAYaA+KWSeOiSXX1Y1/XgbU5n3ZHYyFRER8yXAoUOezQ
84PGC1WY0LYqlyPcl6l8QhUk7I0yTHSOfguWIke41xuOFBGeYHgqKVSAXE0zi5LuUKzuy/w6hdej
bJ7eTD10ZLXMNWN2FqRxVr8uRBY9XQlnJ6XktXDQYZYBTa/M0lqLLaodU7qJHdGbDL+cPyJ1p+A9
G9RjDVyBLoXW46Jo+wG6BfSQc4K7n09zwVz/Pc9kY6ruvMIkXvXwY2z/MEgNefn1kBWba0FwvyDj
vahfiAekd8vZdhZTY+8bUAKjzyamBlQpd5JvECsBUYMLFnejafmNmqqgF6719Blo4VJkwywW+jmL
SUptBI0qROX30T/4IJHedlAtomi7YKvVZqDWbsITrg5nhxtC1hxxEFhnUps11PCPmHZNanwWyTFG
pAQ01uYVcVVcDvTAkEJeoU9fNzIwJpOQhuZ1drjxBwO19d00efgM6q4CRMe1FGqfiGx7C/V+9iGV
arXXd+fesN/A/vPD52mlbYmnrKkvUY9LnaF8KLBcffTWYPtHEBq1adqysOZNe7/xwT4qgYr52X59
Qv10UcJ7LgAoADvppdBpJ4VuNqZ4NWkazw7fQrG5qHySFXN2eOYrjSPbZ02z0ml5UDgFarb/LioB
Als42Sv6//8nuQc4LFnFggrK562FsF7h1316dqo6qbkEl4zSyVVHMoLvzmEfaFsIC0kV03/8mmWu
VYhjlBl75eBHxwPHfhSMrprgvbR6m5au6Xwfipal0urFqDy/rY9oeQU815gr7IDDjjwNu1gKfc3+
mAe8pWu8EAr54OBlvMS+SV9C+NUBES16F+pFY/Jq/D3XKnqE2v27HX62/ckvpfD4k3DMD819X1lt
Yhou+AzIVKLjnT9PehhWmvb2kss2uQto/JziF+sp4HpE8vZW+DO4x0k0NpWpzMJN0JWtpJYCo2AG
d0u8KbIQtiD2Ig0ekJbDoMYRDZc0DVsmvLEqk1AF9TBw6fie4WtIAg7MTYG1OOB8l/Fxt3foF7b7
AnARE/93NXHVO3OYHQW3sw6IDWO237um6EOhIle0t7KIaKD2bI94givIa1+SnL5maJcEuxRBUZ+c
Zi2H3DCV2S6GfaD7XkeKS4TLJoBmBL26d4PPJV0ZRE8mKXcfn4GQBeriOKGNbM2EPb1Ua2N2GgiI
4x0etr9L4ncGXDHuQfyaQwwuxxXLcDiVtdpkDPBTesdZHxYFz+MU3jYTLxsDkeAEqnEX49VANR8V
HPJo3GWZ70gZTSFGnTdzGS0UPXXyXx6fD08CRaMZ5z5Vxa/8DsG1SjQASunpf9ceajAqoDW6QWwx
ZMLl8NWQ6vFKxNziDWe+bgK7y27sr4BRdXRLQx3JqQ02ljhnbHogyjDAHbV4WiuDDwq9qGHfEwFH
VEQDp/WIVb1r6FBoW44WCmgYgD4Kge72Mtaq5Fymv3ZKuUUCrQzEXf8f7CYpwfkUUfEdnk7E3j+E
o0XQ0qQKEiMgiV3rSOmcb590eYcEDZ7Y2cfSKp+8/bPNSy0DNvrnENWG9qB/qVcn9vkdWF1hbBh0
e1+qiCIhQ06ncD+O+nMTt0PY5f2/GgCq6uQbNnObP747+UpoGRRpYtc2doz4HIiXYitOdzqAukA9
nfpWvAeGUp7fbc5kHMP4UtOGdOGSHcYh+hM51RIo/igRfQJy8gc7MBk5ghBE37yK4JZcuhg1iCqY
JlCAQdHF+lIRPPaBmHaEuJ9Uw3T7gAJv05c4mBeduqIZB/zsd6yG6/OUE80LgsNnuJnJKuvbc43y
cSjyEmMP5hHm/rjt318hHhWS7nWp0agV0ut/qiIcOPFoSgDidgIx360ILCCiSARb8hf2TJ6KXFbJ
bQOUq5et9RXu+nV7wamge0LxoXZKa0pz205UsMfw5mbJMz51HSeB7NaBvcc2qGsqbyQcaHiKW0/n
4qljGhSv6s/EZ4HyO0+GCnNezf9qcb/hJkv8nP2wZh8b+HSGmM78BexB+LGcoiAQD17tzAd+Y7wP
2xyMZM8IuoFlwxzBcj9SHbq1g875XSwMCoVpw3P+EErullf54FF9MFfM2/82+bkCq1gliWAv0+SN
FC3yy64tYxIn8zR2mS6b5Ej8YufyHi65gwh+1cFBeMsYmedOCQavt4SdEdjZ3h/BZCnzRGADK3rB
0r+Fe2FOSFpVIl7f6mKOIUB2g8JkY66u6X5NkybtyWbnLTWapRprQrNIP20oSZb9jjgrODVyh4vW
v2BItUMB8k9ohjwnuOOmVCIfL6xK2+te/aRtoduo9kIqoeh8prBVFVvwFdV/vPQVAwb16w4BCjMS
iuSJJdsZNWRmFc8zrFpkuBVc+aghcFyvDPB1JtbMpyDuiuRcOD6/VLMEpT7Zsf1OtWou85ywhNmV
FBYM6oNcwp3L/FG5V0ew1XyqBZkhS+9j79I0yHQh06X8EJm8NiGRHShHgzgWsZSdZF9oYH28D/kK
qgUQGP5qVojZjPKds6M3CVdkRoXAD1Ci0UmuPt9C4Nfm2LPBsyhhFYOzywo28P/6JJgY/oSKSRLk
UYKKOGrp5lRmov+FazoBG0VbyjMVDJGCZuvWdz2GE43XYJdgJP8IjGJzWjjViyEogWK8BWQFduPv
yEeyJcZkEFxsRnFeIXYsZ7T1tIZMghBBPlHkhjkeHTgNL+k2uo7GStq6aTR7nff4A+2bON13lq6x
/sbfGTXcKnpaCHzGgMPWaLcPocH5syyLk08Oc5Xx1uh+5HZ0Pv7fyeh++b6Q37yxrtSahPsE2BZI
nN/WuBFuq0/MF8JqTSIsXYp7GjZkM0+/rqVwzkkGi+KtK7BP6p+HZeA0Eg8to3fGt0jsL8D/wEF9
z99vGnRvxoZeK/wFRJ933b3BAaKL+KhszkBf0rhUfhkNqCWI7QA7ek7pH05Pnppf2oqOBcN1lP3x
iQBbN1qrLluy1k+oG6CZtQ18ftfsy2EZmxJpG/weMXmm9kE0GrhNoM1ETbbGwQMNhQ5/GdFQn1Yl
ZwLqd8NDS4q99XgW+4SqoTB1JvVZPiVzyasLu75wdjbFXTn13Q6jsNb4MN3w1LvnqvXVtDsGObxu
HYJ3hI2f1XDkJ+mo2Gy7gzJeBLp8rI3ob9mLv/EZiT7xHnqSotLod9l7gWQNAFuAuNn5m2XJ41b9
IKN5Qq8WmwJmoxC5+rYtnNy74YEQzXZS1yneBkWZm07uLPWaLQVFVTz9kstrPWgeNvZF7ia7+qHz
bJlFfU5qi6768nq3DosX81h944F8FtSSISplBiPOe1Am/gxPEtuJcpt9Sb18nBDmcLZxenJff9+3
imsnugltHhkX/SkgMVbKYNb60tIL1QjFeZzc7wzmsfPN23Tcc3A40PtqCPbyqwNO1jvd6Vss+mnA
ategKbXZ2CJzA7c0aCGK9abEMGWaklebSuHuHqhLL8r34U38ARsfE8vul9pSZaTWZ2e5d5KB0rQ4
IPmE5bUDNvmLS4MHZw214Y75prWIw1mtsoL5IUQ8jRpcSSd9hy8dprDoRhDZLLk2VbOPNYbT5AXZ
szcHmwZtPphjonb0p/Nm8DAMFsSeFUJRimCPRC10r4hgpHN4Yhhbb3l3qW/GT9SQg1n6NQXGw7VR
5o6JrRzgvRWlwXZPrp+t5ujxUH4LFCv3Eq3bUkQkBOmZSBujcHdgL3AnXi+PJl2E85VdLPlVkpfh
cZwOe9659ddFfNlGE5EcIO9hYuV4DF+eMdv6DtSE2AvycOzklRVuNogHWLa+lMByUGso9rGa61Tb
vjR4FRi6Qc8KqvqOSfwIZoNAbVm3sEjbtaNis7YB5N08nolRkORTd5dK8NINOWwb7Z0253EvB/xg
Sr4FKVO1B17FWOh0nLs2eXbG+8hk9l/DIRzkiVS2dfc0X+X4SVslKBIZDqO14t/d6jhpFI5HGlv7
VzZ8w7YVGTkmmZ6dTGjRJivJ2ZAqzYr2COgYgKEB6MH9C2PuSJytDXZK8BaZaFgIWs6EKCEjUzW1
OXtyuBo2t5GfiPYsa54JueyYzNSSRq0EvEde1y9nFTefg+am9pMPtR5f6z5i91iLAH5UpFgz/2T7
TajXWSmtLpnW+DIAFWaqryXOmqpyXBu69RcnhOywN2OfN1MZx1Pe15WeCIpelPAnWz332gEcMH3L
r9i8FtChxuvM9mDsYKKmTnWy48ayChG5JdlBkA0IYNM7fKBTmkwWQZt1diMJlHOevLQPsqBpqifN
3jbfKxDttf9z9N2I6jCq/tDSTCH6x8YiGBjY9hrafRTZmsMRAY4nkIYg8/lLdLVzTlR9LuMO5ViS
kItTCqaBtaouMQd77SwQFcmeNc128V338z7NdXTsDWtZ+ZwWZ4JZOuLxn14Gv8U+ncV2zmYc3Zc4
+zEemWlImHpmyj+g9MU325hU+Qi3wN3TrBqYpkuHad9kOR/cB2LSFYWL0ixCBsYdFnZcEmAfnM9Y
Nzb+NJXf3FZkb8gQ4KF+jbqvaQevPx2KaSmWyFufEgepsHZr7kmi4ZiSW1FD0JiBzi0l6rxEQR47
viB0Ei+myqgvB4VlXuhVfT5lTZiKAR/30QuXgMqoRnSMN0wdbj6MuKJd3oL2x8fbHFdlWQRbjip7
rlef69+KwxtlCB2E7Ui6lOCbtO5siQajpfb66Iut75/Lfj/q5S8UDetAlhwRLGMJgcgMojwbFlQG
Oze9OhU3rme4UJYJwPJCKNKEoktPtEGy/1+TlfD2P9lqk4+3I7Yio98qi47B2aAcDB5UUO7AISy6
njd7Ut5TJCKku3gv5mAOS1j7lBU58FfBPH0XC0WAZ8cAsOQCxMq6s3STWB6/VKoarkkvdtriVPfu
cx8RTjTVAzXMyCf2ZMZRsTNS5wUFo1UPchPE0xTlXFAyS5LaDXj41HiuiPHHwbmjIoqpi5q9QC8c
ATyOPo9GhEcxZrjCbKQvG/8K22TxREskzDNdzBGh2EnThwTZD57rAAyEM80EOe9RJirjKpifPz1F
bsbF/Yk6+S4SvcaxlNvsjh0ijg6/UfRpRfGVWrKZNnXXj3SXTYrHVFZrrJleoufz+wDU8GKSHWO3
drz7N3NK+PMKHdVKYMei9IoBwLItdNie2MdJTc+jsLBv2/8UrE3LlKBIDB40oAiVXS91u9lbqpCo
kFo6gxkxtEmGEEZYcilsg/PDYz7jAbAhjGpMpJT8BPSaZXgzn9ctiS9aasfH/rmpFNVONJwE+L6v
JEE3tSpknkksn620LmG1cJJ+MfWIo6l8Z/j+1PyD1+k3BYLtNN93iGmAfTuhQ5tcVRG2a56u1ucD
ZDMnUXXD9AhaR3QrHtMC9jYeimlEeQacVrt6dsAWdiJfVzU9jCjGMh5qqs6cTSsopPachJI/13G/
2fZcapCrcMJdG8k91RKQAnZjYCxVVAgYfVaxLwSUBnkEVWIvZ57OEQWTeUts/Zp8/p5xCFVh5qEQ
mWnMETmPHNoM+Sn9HeSPBZmsCgPtVftR3lgb98nrT8wNraLOeTlm44uBejRhyHw5SoCKfqVuHS9i
EHUKkUHpICvJbKr8ALSruWToszMSgFPMIWyg7dRPKOhVT2JTiNrsZ6UDpTg75/REUyT71YcP5LoR
jySWfHF9wjxYqTV4GaxlwNM63XFDzqxflKPlR1WtqSPPo7S9op0q6/bFvUDzlnVm3z9wcggn/biU
DAbXd2Lo/4h9n3S/g5wXFowYo9IHIx26ZAe3Vo+b3rDGHfb417c5YIu+qAtoqFNsFojqjhRQOZmR
P+TM/w4TzeNd7CR2QyFR+8GWW+JP+OjvO6O14+uLr8yGnNYMS6EG6mALKgCXcXCKq/dDJPNqFJB6
o1KZHoRBga3tYV1ymUJLhihHfLy5YmD7WHqm1tWGTmAcQON2uRmY5JnRiShuYrqV/Hf1QdlLD03a
JvQRsELb1/nCxMTXfZjke8MkbjpKiq3qWDgmdriAL5tSLHtyAlnWxXdn3RH+k+xgQhSfOY0R9YPf
5kivYupk7HQEn3dpCkra6JFWY+MtnZkk6g7HjgtI2Q0WT7F/r3wViBe1/1mJVVerGTpSvbc9zTmx
XBdXHVUc3K9S/6lq0blSIZFwPuydH8n9RJzmG57WSs+yKBHLMXl97f33nvc7Clf6kRXm1NxVOSuV
NC5iuvdDaR+8RP5f22VOpk2MoiH1C9TsAi7vRHtPFCmDzCHuuI1iGCjB24xzNWo2ny8WmNWqrrcl
h7X07W569TUIinYHGZNwVsGZo+OJAs4LFFhP89DRRcEerDjmKEtTQl7duAsha3IQub1U8Uu5rjYu
3JYUE5oNDci7RRcu0CJFuRwzYn03He24wccYfHibmHL5oLjqV52ck6cL/iQAaZPXWSpONFe8d5UK
16w5PYKanjIuQY6t96Raghm7tkokUgBbu0OnpS0iqqBu7FwGrEFzJndwKi0GwuJCTFNFNR3ygUNF
UlX0iTJJinchhvBfAZVsu9m6voHk9qjqhNVzwJTu2BaoxACN0cAVqtjx9HPJ+k9+8tZ6z/a2kbyB
qtS/bzgVNySlfuox3FJcNbt4JMO0HAhVKvXaozB5JB62p0nTVBFQw1UioOfshDc/i/+slU6TRsvp
JDavEiRPA/WeYAt6t+Ejm8LyLXh/hG8fmG/tth9tJamxdG5FGp5ZIXetQmFbG02CZeTwjOKHxLQO
I4eflNB0l6ZvJAoxPgDtomYB1CLQpfswQEencc3nZ2Gvv0/xUo3UOJS2gC/mCVgd158Al8VmfjN3
bOlbC09V3AK/gBiiSEoV5QiRD8CTzvbyywZdfRGCC5b02PUHbi6OA8CfgRtc9JV2u+ondz76wo0B
x4YQvcXaqTBEvVHSwks+cG5mmzZ8k516LhuvJBMRQmM0M6W4QmsNf5dbYwGxkWacZS+ayOaxvCsx
pEQ493SoqoImGv9bKth6OQgXP59ieblT1WT1bs9/uiHFr1lV9RYyno9fJJ5OtN9YTUJl/Dj02xvb
RbqanGW/JZXGUn8RCB+g5orlDLwMZsPbi6Fmr4UfKF7+GxmeSs/dorA7FK39ZjbpWSCL0hOPPRXk
89Or4HmGrUoJXH1tfJY05bBkyRA21rp1hy8xPbPg03cNAW191QvrB//sty/vA9xw8+lsID9TUiC3
ICEc0V3YodsXkpM0rYehADSOE0FrtqqUwpF690XTZOfTyB+0DzQBFDxQ0nKrOOxksqPkGiDBJIUA
BDKdm3+mjWk5ZWA1br5sydNGDwjcYerVwBGJzN8LfiaDy9nB1u41LPitcBeOoTzXKXD/yVkhoO7i
7uvNhYS0KLkjq6dzBcqJZQsb+tbH7mT7zK7J3X11j8oKWXex4BZjDV5evVM6V3cfQrojulvKd/SF
K1T/hcAEcpcv2OVHx+4jKZKU3wkQnwIGh2TO8/E02Bk2IdeZIi6L26RPrSCULng26SE7QaqcanV4
yrN8hYNdynEn0Ard/vC1U7vMgKK3I2BfGCM+vCp2C33WAXwnttEahlnPrhKfwZ0R9d6S4q1ABdCx
ctlkVjFCKmhfrxIb7Q+CZFq7vwEZl/xigNwFePRvShcvM+cFncQU1yYe7TTf6mg62lyiJEiJ9Syx
xPbO7C7al/LrWuP6kEhuFlE29S2qNAntyD5px+ZZh0rLWHGlS4oS9hfLBmm6CEyaLN+UDFqteA+s
4LVpmrSgzHQPBbJM/T/m0Qn3WMQ1VCZUaUtexYEEgYlfzJLcRrn34VYmdiW6x5s6dPjhmKfhBg+N
G59hL7b+duTj5GDN5r+MB+CyvntHQMWELBlDB02N1fEb/nvg8oO+9ZNmItgRSOIeXEdBJDfSa9gN
0xbIA5i6EqGvTuzyTpevJVpZziazQva4x/ru90hiRAYnWH17d11COxDLGqPiGQu0ss9MIQNIL6PQ
DWG0YR3yIdD+Pt+Aj7j8B9Kqsssbcyzq4+m/7To5F3ULe+H26KpmVFHZaceLFdXNfkIHdjTKd8+f
idbkYnN43fa7uY00SbPE7RVTalpJOQt4pkiHCXwE5hN/iUKbEZUdgo/Z73KK4oZsEUYh18ck/8xD
FR9aMOq6uH8Kv36VcpbpH2WhiNM0hDVfHSctytk8Mjum/5iHqlId2BZWL3iJGMZy6eqEk6ifFyfa
gVFy/IXYLm1+7O/auT0m4Z82sK6g3iQV2FHz3lswsHE3VRNOij9YbQtgnNp90aTRcMYg9KRH/9eb
H5vediBWIOrgAbBPKGTePZtTwnM5u/s2Ya8v3wLCuEgqplZp3C+AOazy+tB1T6nUkECtxBOt4FCp
mfzK8z/nw4F+KKWVxxwVji19UW9HlBumXgnmrTMBRXe6ShbouRLq/YSfoWPpXFd+ku2rF21aBMP2
Nd3ZgBLoiEPyv6V07N3m0H55gj+RlMv9uFNrpJ5lA3xpmSdK20o3jKefOXVSMPd6+t5vzj32v/EZ
UxFxPK7v6xycZxZrgfUVbqMkn4J7Wn6HiMp/mD6l4H+kRadiHQpxrBHCfh6ErsKvEtKeOzOhAkOe
0mJzjuuGkSmhj78KqtM6/oJydKBccsD8XpMMlYeOmndvuVbnQ4klkkzzOO0LsbTUS0yS8Izk+7Un
++4J3rFNay9wY0ehz5CX0jBLU9Bvd+F6k/CICd0dbUXwIb4IIqA/UL3Q2MMmfBIuENNrpvbAZLNs
5hyPGIZxpgRSdeCHDuoo2b4P/iwelW4tX+sHk4JTovZWelPDqQinpn8qKkLy8S3C3ThqfUov9NNN
UP24zPzSx9msGBreCdzC7ErVXPWPSunDa8s9f82ZrKV2Pbv8YBTsEIBrMPU8KiKBmjkyTAYhbBZ4
T/pHGuMZbA40YXxTA9Ibj34qevrqqjGsfcarkdVY5LUmqTPsOvN9HCyUlZHXa+wN9zbXIqucZKul
mAZBZBYhj5tt58DJaTL3cmRXe/pqM33CdmU2Yhr4Xj4tmFQxnXSd0xkEUDGNmrQFlfJeGN7YTXA/
NS56L3IrAoHNX2ZEei48r3ed0yl1KgcdSu0jexTCtt/FmIXvigU4pow3tLABT2+Kb9ZXgR7nwUzU
NTJNA5ycGc/IxANr9PGu9hpbiCY5h1oj001/CUj6xxj+Oilcf7hx5SBVQAG7gozLVz5kDPGGevQc
SQUfjHqudWWZavqgAnEAUzilgLCzoDhH+EnPIHeCxPv8jc/JnXhaJVw1aTZ0+oN0l+bCyIRgWu6L
UXWFiMU5+SngVG7LXUT2m10H+VtzKrizr4EyLyB1RYWOCDi+Axg2a210vYnJPxzsYpjPBMee5DwV
v2OqdOw74V1iK+aEYGnc5gdIvHFEBmyfEPBKyAcYsTZQf48FMaOZXOy85/8ftlxvKq7kf7VQqKON
GkrNu715favZs4WlOlciJ2FAD5W5k6ZEpvxcUePamIxXlbTQt//jIYwdvNNbVHDDExvr046jwOye
Bqs878A8hFYMfbgmPFbFCBEd4SkwOAGh/b69y1S+ct1fauCvws9ZfHdNg7gx+x/IuGrrWHIrjcn6
MYgIsFGXEQiHf93K4H9ilqkj6grRT8LY3aB0CRbx1IktNP10oDEoYTCJr7xNGiAHjuP8EJhZzwaR
0aaPu4BasgOPmfX5jpyEvZkuxOXulMh7SOfZhioLObbbIPLy9I+3LNZgmuVrV6A8S7m51iMkQpI/
Mm3NC94jbxgUEIifzBjW2AC+zNvJkOR9ArDrgKVABhbcN5mnKNUNEDtXBQU2pLgbqRzFllmP4UdT
TGaqjwbxJ9U+KkV3iTEi9cKJpDzLEisHdpK1xly0sPpbV6w+AUWFag3fyHCokv7yxJBcIopq59Em
woLkVyizkoBcaI5y3ji/+iyurN7TWBIQR5mG1gSbAPCBpOsmBOsKHvgMv2leSrWwTo+typLARIR0
quszbwxyuDWbk0DBcLwmQI3IsjjuA0CNnHoyW16UmRSqKZpLd49Fuw7iPOP/TV7y08WI/WwTjPKE
EjjHiNvivZX3fn/HNo544CH881hvVdPTlvDFpR5rwtQgcHcp+hiI5pKCXVHja3O6SH36nUlEQ2HT
FWnCM62Bzl5PZfgnZbWfYsLWfQ2BbJSwW0YhBnKJoW7kLVezkvDSNssZKvuRW5J9MUp5xn58YrFZ
1w7TRjA/6O2fovAP/nLAlj2qpCZK8inLnds1y38QdZc7wbzG8/jL//RucxldBvWVRpAY//f248vu
+pNBjzViqQ1sLGAKSv7dJ0cfQHqLM7lMJQgdUHWZYIMdEdF+vvnTWpXfQBOQ5C3Yrm62LOivtMYU
2+pEwQ49Rf+ZvWv/qOilN0J0IzbXuf7RgDiXIBO+O2TMX60fU/SXl0TGkeMjAXj1qeqvmo14TI+m
8nggSjVg86VQ5hcvTQA8z59+hSfJieLQrFRE1ic0n+kgg0J5e7kzXuEOJZq/QUvY4ifTfE4O9T1O
S79zGDsTjGrcGHfq+T/3dGlToTthO6Uzd2fpWeVyaTNC5KMA2WB4e8TQY0aEiXqvoM8XGYJAoox4
K1go8ASEAe29jCg9DaKote0WvGvjRNls5dSLSrqKJiiBax8fDjifgx2lnECKTMtjwnWXPb0CnxTX
QFRsXXqdnJoUSJz/qHdzDjeLpbR1dSejYrwCBeXXC4EIMj7EPK2LhMRP0WNoTxhZ9dy0YkAqoZkp
ALYn2pWL9c92cbFcvKe2dMjclR/a4f208n4CdyvKVAohvegvV4yYqPiim8KeS0IlCknML81fkbcF
PqFOO5A4ATY7WTwNWeH3SjvQeDudVlz7+hVzjHqKQIBAFtpdBrCxP7S8sw3S3zPg4hbHJ6yjv/6u
vxkD7CbRuMf5r2Pfnu5WVNnzZuUDraTwQXv1fVwuQV4a90fd+VWzF5QNCgSvRlG65iAmvZ20jxbL
5mb7T1JffF3uBNIavJpkKT/wH0a35r6c4tyT2ABLvhKSQhvVWIpTNIc4zBcbjhgRNn5NOfI0x3nN
CgWqG3AB8tM7U6s+z43Lidlvz6crRKyDXR8FMO3SqsC91YI/DGX6MxOn8dhQnSpHEoTZUjv6TomY
Fe47YlIg9XAMBa9lzUrmtVZ8OnGm7C/pxwwWpHHjGB6MxyF2AVCi+6Nzos9kq9WNODmB6by7dhHm
/6NUchlYlhcGM+pn11AoKDaXKhM5AX2gcivW/rLB7AOTNmEsUmPd4l8r5XvD3kHbxGf/7fiyMZFO
5Yq7MDaakxe9FZwG6nTRmuoIdFgaZoQHX7k8RQ2gk+JOBfz8+0Th95cxLsA4VRlt/kBr/8rjRt8c
AAnE9YQXJzW71OR3UZQUf3GkaYKtks78MK9FoXlVlaopG73Nw4mUBT0ZG1HWYSkOH7I1QaDuSMeR
iU//obja6GhF2inAAjdJYY4svCnkyUcbnYgUzhaATiY0ApgYsRDmI29JIImfTi2GHkIsFSPcY9k0
pA3o6k7J/4dWCoPNK0p70Bkq7C4gSqMUDIJjXCs9VKFa3nUPQt5pDBoeUlAE6lHoToKEUWpyYsOt
cg4PoLduNYLQq0gALmn+lVDb05Fh3A7OzEptc3tkUM5+eloDMGjUF4a1S2C71aOhLOWB9HLT1TXc
j1UoZlSajtmBs0Jr43p1X+kygvVHrhK9YWOosLcP5EgJr/KNyCfGqc1a0R70WjY4TzNimWFcEHl/
Y+wusl67orEsTPYb57PAEVB+k7I9LiX8h7jBcqau6hm1hb7CtNTu34ix/N10N0cx5kuIDLMYFe4F
ehShqrUIss3R9qlJNevsjvVHVmhubX+Yq/ESVcpEX3Xefx93BHF8oBDluAVnDe8NHBb1+PJzW8Wx
cBf0X6vITKgqxMvNfoumcCvCLp04/MW1lQRkaFna3n6sJSnSYe1uaZKau+ztoZBAGyEeVItZc1jb
uvvOly0rosaZ+N/6paTW7RaIPW8E4ghhYXIrYBM9VFg4ddPSfphOGpDW8GUEiyba+4/BHnU56O2N
z2DO4BC/0cfhtRp/mxjQ3wTu77r9YxOIoicDdmczJLuRcTdM4PqMj79EKIOBYecAJPb2UdPDq2Lz
tTa7iHJcLHNgGUcfXfolaWG8S/uUS2ystSQXCAtWWiPvScH908fJhkQRgIvPHsfC/zsl81vH1MlA
tNeLVLO2TkIrYKQdJYN64LKpYleLYyEQXctsdoqteqRfaqGvRBvX8U2QX/Osh5paxx3TgOZ+pYP3
nBja6HnoZQdNqEKgUbTxyu9IPYvEp4hZFrtvQkqlAKUP0i3el3yn08TSfKKlcoad2idi7FoO8jMm
CRcNfZxJoA1L05ecRea2nvl2snr0ujtQVr5Hj11+85yOACUv9cyHWcKG8zwOyoWs+3dVajWRP0jY
UtOMu/GzosTb04TL7M6bEqhYDysZoviI+NVSCkDzCoC9WMM2sU3pQdF2EyURngvWoMPvfjILAM7b
vhSUqT6RlAV4USBtdv1LzemG0nvuw+OtRDLKm3nBbF7PR6N6ugpfvocq7n4JDn6x1v7YREQTROG9
TM6qo0dSfIaDypSNwXfaC68v5B5vK60M2dUyQjOahOhBGx8+W4I09S+5dJrMOEl/2UbHAYYDXx7B
qFoYa4DTwiUvQqdzGinih6zQZrJmVTAZs2etRAEqsxyVgMO+kLvlMpXjdqM8aM+64psx0PHdf42k
NxO/LE/n3KvOEs9uFpzhO5PcZNiYoPt0nZ7PpCL+VLufzjtrgaqk+SI1a5gSjfEjomr8nyDAo9yh
T27GsAp+CNQeBCmpiO1c8FQMFYR5JPUn6anz6ywkc0nh9ZQ/+6cp7NL/Ppe9DxvrpRqISLNVGaLC
o0ESIvPoU4VG8ZryS8sIrNJxHq9zoTmwVPOgmrRqZ8rqoyzCgNnKSV38j/TGFFMIsjNUGwa6bGi0
+NAFMAQWTyfmmHt3BBRH+aM9wwWfKbWj+TAlCeSpcadg+h1g21GBE0USiyW4AbkD3QKJ8Q5ui19U
+16SUR8SNfAS3bNfncI+6IWw1O1yuu8LtpQYhekOJ2ZGP/e5K0CmXAw+jk+BgCPC3+NqKRXoYDNj
E0gaLyyAlbDHTLYTzDiMUIXQOm7j/pJrR1pt/8x+ePfAj0qECsri6ZFnx2YorlOu3gk7LCVFN6TH
vd55PxxDqzmYKrVHY9eq1aWHdoVWJ+niim/VM62xShMMKMWM3Oy7qy08XAmSzYG3tvfhGi9zW3s+
E81xWqceGpXsfptG9QHcigcX7FznJGHJyOkZGqDiiyVnSC70pFvS+443vVYBQGpkqHdnG8tWddmZ
aLd7tcm3i43wTiuBFcswLofKDveX/FjR9/ISJw6CSCrIsNHgDCin8yxPMON7Ylevzyznt5UM+YKf
cBl0DgCL/XIwlOLC/kgLA0pL/6QFoAXZto1Nti4upqUQJuE77OkKP68I5UvGO0CCPOVaF8zbdiv8
LcSh/kmmqf3q1ijI4RTHSmHQQ4GeQg6Uy96wddw9TkMGhlFL6hU9FLmeTmO0d0vHsO0OgzyhwKpJ
L8zIsV2mWKGDkkXt3yJLHBkaf7eMIVeMIFug9xtgP5EllL2T21fczH12ApF7X6Y/g3K43348MQCj
W5/V2EGE6HpJbUwMc7RPznSSHs/UtOU5GaXIUJ71X4JQzQ/LucxNJgg+wOmaBQ2IMrTSMX1slXeS
82NY9WFoKu1+GjIUabDea1nDAY567r8Z7umYsdvqVFCWQ6nri2YOSjgVsyq/tVqu9zwOkfj+QXWq
pYO13CipCO3rbTZNv9DlRKLnM9l9Rz8UzSszyGq87GsEflZ8/KAj6U5VkqCOg7NF9I7o81wlux9H
A88ioqxL5D2GKpds/A0KKjR4/0p5IQHtBFhSmLh6Szcj+93Ihfh0A/CE7PcFvhhqguaxgmdqAq5W
cceXITpnfhwq7JOoTySeHscUeaXgBt5V4S3CsoNor4QV1qyu/VnF1I9dsaIXDKZN+ACoHkL8ge9q
NbgxZE1m+tjbDVRcjPQ9NAe7pU8pxvw/K4IQhQ07SpOh5CodFjvqMXllImMYEpnqz+HQmdbtKpDv
e9Dsyv1WLiZIvNEcqGiDhCEbu/E4K8cSRsCM4ChgTyWpGie2qCzWtlQlYbDPQHhHVZOC1fg7gOKk
aqEI5Z5m3ZyzeSW4fbztMQmsf+T7FTfvr9/VTD4l0hZEDh42awCUUMCqnokcooQRSC/Y5fFFRkyh
xTLRvhe+yeWCz9nTun56L1PKzZML9RN6uiOUwuDUnS9WFT4O9KhOUUd+0ZhrlhUuKoHUmvH+M7a3
3ZgkTIaVYi383ALqUJfM7IVBxv5a573wvHOy9PkLQbi6sW2pUeuHwlR1SuUV0gzMWQMjiZ2drdoT
raqO74HPA+uvOJ9BBPbM6qGVTVBA76u89mxVGHvIuaavEh2bD8joulFCZpfKGu3O37hD92+VzFvX
w5Cx+59PM3vfwIIh/RfAhPMQZUkKwKjWS1Q0Fp47Q1pRIko+NdE89Yvpi3QakWxLjkyf9J8AB2SC
Pe9WgWXuAI6PqgLaZ/4MqTMhCXND9Z7RNUD/RUj9Yf/J+C6ME/7/bfL5rb2HExnzuPNNxR26wzJz
BLWJguwCAW/p1P6r96WyUwfxrxoebMl0/dQv2ZnlGMcsZjTLPrEQJ6P95U0XS+f4ZhsmhXcEBb3G
KuNBfyIfKa+hNOxEVlcONpz97JfPOt7WcCc+/b2pjzTHd25V+c9Pexe2qiZA5/syb0vAsh75OdHZ
0zOhTS2fdNR9JTN5Efw4TscLYmpmkwzNLJNIXhl6h9Iw8aqIv9hNksRQGb5YFKba1k/HB2Xe0Qez
KZRQYrU7i2Bg3OYZavBhTbRWqI9pTvZNaQKDv+FcflBLtXRZNWl063dvbKqyADMkjCzTkggBfxgH
iqqAofuSUIsHhDEc1P2etFcyJaCoznQ6EuUDXCOAiJbvxFD12Qc8bz1E84HCCq6stuN7Her7fOQs
tg9maepcxc3vY2WA2Ltj1ZGmz5IvgQ2jyfTMrMRnXonpHnxQTmh1KXqKwV1DCeV1lBIz+mKi9C4i
zyv/OS6+VCMt7HNPLf8e/CLQalGh6Ek9d0LS3TtaGTe7v80lFgsYvLGJfJvQa99jVs6cmLFKXPsq
sLKeGl1x/pvTUql2OaZ8RIaZEAARDOvPHkjsEr4jUs7DnhHtkGLMgy60JhUSyh/7eNQqZLHlw+uX
PdJj71QX9EJl1Ge8GFGydF36INC9mdrSj46/32WH4n1sfAlwmMqjCCdGsVUp9GEhZ0GHoI/yvqp/
0wH61WFEXb4EfEjo1S5lg5hublPs8iNwiFtipr3po4o8Pu87k6CAEaRFGsBp09ELvikEa5yI0/xq
paASCx8HKp9V5TjLyS+hskiv/zghhvbGPDQPUY2SrSYV2ROOtVN02R+92rT5QQPsrxCXAfO7Lxfc
cxkcjvwJseS1B6uoXgMKZlCRwexfAmZOZLJplM7QutJCtklV/TbM+/dE3V7JAWjtzIidZ5LMVRPC
y98JD7G9HnmXKQT1Ffx4DMpgGZMxvlDYp7QMLgyTTeENZVSNOIfGy0OVxTnPOl/+fueUZ+JUmFE2
FVZ/JlDdq56wA8jniWRiCOxfe0lFhtDjOUde6+ST2Db4+vXo9ePYX3BevIqes+oTx0ZB+js/C06N
VAiPNfRJASVG4nzFD+CDyzphN53yj4usiBDVD+ZoUGvuUDLBfubcXWxDr+MghBvuztsma9GBpjxV
+iMPWrekEst35B3YHjXM3mrBGURBqjDMC5yEdwwRZvtBwDp6EMNPCpqWoyMMHAhxMtgAkUSDV+A8
+oRrhdAcDAH67VC5oeyqbXoXBTwt+Amvo4oOiIWrt0Bl7/QNtG/xlNryQUZJ+HhzVFLaZzit76St
5HvaGAB8B0ljZbEVlZyIXgpyl4oIcgFB2q1lPlLDG4B7hsfHy+2fcvIvrEqDVdwg9gc9qmbTcosp
9VrnmJfUxpPxdf4kd/02/Ye4BYa4Ic8y/zntbrHYcpHXOU6/4egqCLExN0+waLIQ8DqRS6TB4oNd
GYtBOqzHyIwxej2X9zeupTD5QnNsu+L+5f8WK1guW1vaIelK9GQIAF26/T7j2W9H+by/DeNTohEU
w/O9D6QsRNLQ+lwhOcS9e3iU+bVGtdDHXmQa5T6n8fIjb6Lc9QqtGHzHWTFZxBu1ZB9/pkXpSjWw
tyrNJ6LUs72hfqpYchjCfmFKCCMx1+mPRNk+eJrJgDAN6JUyeYElxztj+6ArCrjvCuj8+Ks+i9qW
FfYWBTSi5UGnrqrKVNNbB+wr6TIGISOE07sqSl8OPFTyidE5ld0Yes8ZmqtXPvfEzBc8AU0SC1/x
/CA0FTuE47UOoKQY9VUopHN3frhEp2I6SVjgNW/Ul5bdfLSy7yryPo/+vXHS9qHjpHest9r/WNgn
T+X7lR1pR2qr3JK07yD+iJB47k8+9Bucx0HCq5WsaRwQHAhuMZdBDDYhk4tNbIvwyR1q3erOkHtt
jHHoQepgTjeu1yGxgAKfqxUd84BX6KERNuNfr9WlhH0tketQ4ZnCUwO5TCf2YqWDA3RY+H/uog9i
R2oCLp5IcukE292uQIOaP7aDhqzM+428slmXiO/vjWZ3N/9kclYZUrE7w0NV8wFMGPWw9N0LjvWN
FojL23JXWUnF9ZfDT1V20vT6s//rE/evtBvxUeKT0CXT6yuYxAp0pyk79A1BTFh5t5h+ZSIDNJja
zB749zyeZOTB2UgA+tNAQLskvhyZEAU8v67cMhoE/kI8Sjp/Rs16VInnWMh3qvxKY4Zow3rWRDkL
M+N0wcivp7JtgN1X+ZCRLPJPLJAtZ9J1RVKixJi80D6QgQgFPQI41KJGT1CJmp7UXFOz+/rtykC7
FJUlZzGQFUvV35agxq49Dy3o0lI2bQCmnh6P3irdPQkL/Jtywg2HXdyXAloc0dX/QfBpctJbTvf3
7OUY0of3jXKwNmnQWm14oZaRmslA29smg6sSd6FB9tgGUkFFdaUv3Bs6IA34DEWpVmx6Dtf95GHT
VgaKaIEGF48HfzaQEGtMh0hzn/j4w0WZ7SNWvhkag1PESRFCJNcoNbvZX/7S//G4P2Ku0upUPIWt
FfW5l5q7q9QmNDkfPxSx8Se8sG0XJgyEwkVLPx3rORS6pu9ElPLd0HrRtAXaDlsK17x2h7ZhPNiY
Iq3TIoJdXSUw1tMpD4FtMs+ZTxfG1RI5HavGCDeyQHAcb9yGR5hlU5xFn+D0vi1YqNlv8UA+efCq
2oAamwU78quDXDewT86GbSk9B6hoN1gPzQBZ1OO5PEF0xOaxnUzkKRvM/FRpINUxlwbSfnMAQii7
Cg0lQRuvTZhO6X+vUDkH7H1mUvgF30aZgUf5MQeEn8YGlIHBLUm1RQYTy3m3VcPoQCXCCdckc/Rv
1kIdGqIvWPCgokwSM5j+qHVvTeUZIxtuYw5MMInsHcSX8vxiKXXIxCkgj1E2rrbyx3fbQKbZPoqU
R8lB5znPWsISRyvTIlp3LKIOtrZDeGpZVTRHsyzSLj3PAWj6BV9PPzalLq+cQFsX9MMWAYL1Yj4O
LUmVTfR1dfm/s0p6zG7Li6g9niLMeRz5exTv7TRv/W0j+a+3VD1uNj0RanCAtKHAZa8RnMUhzYzt
+bs8xKrSzTmA2McZnUUTwtOoDbX7G3e7/CFzgK+dEjRYViyVDyvHe+10qRDjtUGiyW31UT+jpcKc
tl8ia1D71ALg41bdlTSlqr52ZfyN8oqJ64uOSLnWuwZNCb0Gs9fq0MZtiG1fRkfSQgsjg1hs3Ihx
1eGehbDzVAfQuMEPq1+i+p23EJl77BNLCwoZSYbw8puSSI1O9npL4OibHjOpCyRPfWMXH/ybNZYp
eKa8HRg8xeca9qBTN3NT7uA2cODgF/b6hSbWhWtKhgBR+umZNJibum0hCEKejQaUICGQ3ApqSyPM
lQKstEqfnQoEvRpE/Q/PyRCq8uGkDSOBn4rtl+2cVbVxsmId7QjdL8oKyxQ2jPRyhOcxwzR4FpRP
c/uGN549+hrY/Y61W+1jQSaDmp7mKqxM8SGuUDcJSiViwCn2kSCcGV4DkHE+U1CrUyiTplI2kVkG
V9CCoIZ2YcQfsK+sd5k2ZMuCWAOl/6leFbnJehpnTYDGS6CT3ROE+zCHHPgRgTAOCl9xoO3UMqeE
wLtcPwv1CFmHNzZWf9yPIuILK6fCdPudz7k4wxE5+YJObbQygJ3YYFVfbltvKT+yT3/IdWBlGu8H
z6S4DzBZYzbx/hnBr9EKXbf1tUGejdKTBtcPcanbwO/SxJ7OmHzg8NSbhHK5NhvvGnTq6bIqH5gx
v59T0VWvd3XCkQ69FBUCUtcAFJbCtMCP+PvJ6zXZEEhs+1+JnKrURbeY2L+7pcKs3S6V8PvMVr4Y
IzN12St6ly8zFP1g9mG1w0DcOHw2XOv//L8g397qymDFzmfvaCSL1VWADdaDVedr1s/Pov1jnaCb
9zdFkQmX52s81b3KTY0FwXLTUHreX62LjfY5rsaY0RYN1iGEVP4lqKSZg78quG2Yx4sj+ZcfCdjU
2S5lM0GXIz0MO5y0qqw71EJzLZAhQrlUj97XOdOCqa9lW8Q4oND8ajIfw/C5YEDlPAFGeNNXzJ3I
Q9QyiBXmj3/r2NahxAPTCYEz9kOgxOAcJ5iNaiOnCQ6kDtuDhAJ904FjuzUbZA/eP8PCtWURfDGT
/XyyZT+LixxJjddOmy8hLN2b+netrtx1+j/LCf2u7v7/3/pze3IYl3VJ5BLdJc9/dsO6I6tp2Ej6
FhHoMUxsxgnA2RptTo/42wPR+dPb5D4iMQy/SnCj6HCOgHptrLb90GpkwObVefnaPsKzgp4wAFFF
opzWdyRc81o1URhPFVt4kuqRWncv1vPwWrDDUQ0dL1lY5+2r7/ID1a1SPDUySWVeueNZ+fuCeFC3
le4jNdQXZFctwH2mw585fiwyz4YLv/D6pkVrPKA7vikJR95/f/8cNykBn8YiEP12PeT0VUrVpQ0K
23JkQnK01ziLnXa4yPnzjZXLtcjJzouHn6NXt1+KwcGih588XIkwpHb1oEpyQMnm5fW9rh2Qx5E1
pydgUM7hemm6MmrhceC+c3LrHEk339o6ImJ2UmTdigZnjOTd4dYNsNl7yu0sJb2uKUiQOPtElH1u
H+bSZKoWuSQoJU11oGWoAWbsPCEiEwHaqzWvOm4Uhqnml+dJY1QKdlwVFgpYcpkeQr1SB80GZ55r
2Sqxxa3LCArVTExFdC8kJHC1CzUytT7S+uidtqFUP6pRmjO50SuPy7/Xtp7jIr+pBjiZwvzKiFo1
SVyWORA18ahiAKdWaWMElUY7E2+lVcc+mhBGb0hNebstvuITubSRx0mnxgWH8TSPfCtiaAnbwbq+
neFeE9falXBgnh3t9DO8C2cUKkAcK9ra35SfIjOrOOvWj8xNJ1xPG0TMFAMOlGiqpPN9+bQX/VOQ
ilfghRdK9+QxoINTFix/7dZlmCx47MHCPyXdyZhyevqFa/bHuXRaGWCm4aGiUkjdFJ3pC+DEB4GB
6H8WyCPT3lFpWFzEGCZdfZPI1Yy+edrEh7tEWF0pqg348chvbRB1jkcep8tvcEcXAAGoA8nc8qtW
nYuQw/PhqHShelZZ6f1smL2teJIP8mKuD9OUPjYjAWZhwcLy07FsEixDecRMflRsQ8DgslKv/ke3
14vvOYecgu7qTch4PdgoFVUQqDHwSE83ZD7G6Q/mFC6X7I0K/dN994ozGfBCTPePQCJaVmiGTZk+
5WoAzMSYBWiwaW/eYsdqc8MZDFcs+kbRVaGoBFc0fnpYdFfksRld5jJqq7Cr1qZkyt8IKvLtOa9e
YkJnANJgAVOfHdWQoTJtuaSCYgOaFvXvtblM35hMqbwfWoo7wbw6XXkQIKJlRppmViIosWsUuHd/
kJKtJPAnoHTPffnCBGmdvv/TUVlxFtej8SCP6gV7pZwEWogKqnPb/Vy9WrB7pli6WVCIcZ8SfEyn
KvBJJjIbqMTKHj8Naux2iD34yRVTB2NxOw6CWOpXD420hWUNFs6K1YhwSrm1jNXNX0ki5ssydxHF
tjx92yEGOeu+5LVLxaMug+Rdr0C88LVD8hbyAe1I8mFGN9Fnegp1vwhmd+Pid7h5zWSnFghuXmjW
gjkAPyGq9p+kTdPL+h4qjP4m6gD8ELrj7YDp77h+TgA1U1itmUTTRcBgGg3ntFpIsYZIzoHpqh2o
VTSzC1nG9HixiqaGs9Ha5vGalB1LgbkF3u8iBEFs9Xv8vaSRtYf+h07/hbMpPcR5PnwG50Z9hHkq
tqYAGRvVEkSWQ+Z3SnNf1ub+9wCUAzjXrFx70UEEbrguNCYbl+06rxNirzCkM/mo18Y8SdG6rG0i
GAogfO6DJNbwbc6Z1iXSkEopftKGIKQLfwbiZHw6Y0WLnpbWdwK2JMUkfrDT+8+dfe/bcp3ihgzp
146Q/vxbf3N4st8jZcMEthSMsGPDC7E7pD1ADnLUBce+1pW1FcIrnc52x5DA0ijNFvphvk43Q3oJ
HyQZEPgupGhm8l6uFjrcB68w2HpIRSvCytvgL5xa3wLKUGJI21BI9nvEd2FGPbCnj/XuAKZvMoN+
l6bkitqftsl4Sb+SUXDPjl8rLj6oqQ32E79mQhA92QOlvoKbn5IgLZGZgTavWGUxKD1OpbLwANk5
TWoDEdA+ogZHCvOwh5OwJTSerr7P5a9pcMOQF8RyrlfWBBDVUL8TmAlzkgqvvHIKoFK5XYPeOaZg
6ou2vdafSkqZJSdOlcvGWPYRjjqH2aw1dtmO3Yy4dyfn01Cy5uon16U5EanbtwDZy8PuzgwRWwui
xwQ+G+9QKHuUWyauAM6Fds/JGF1Y20IeRnHbjIKn1EYj605bqknszSDTwq8oA2/cJc0xUKOmX5oA
NyXhEmBPe2Te1h94n3CSaM58lijzpc2fTbHhxGRo/6UbvZaQiTyqazHOAqiquntagUNWsyDTzt2o
CpP2lXaFTty4iXbqHdd/nHngIGlKZeazM7Gu+1I88khcyHM+hnvntP4fS4RbQiSmL1Qv92NslYAN
1X0yQbjYDch6M7f9qTsPGnOgPd3BW2wZ3/vwN7djl4Mdv+ztdsz1HFQluRfskYO5v1mnPisN58TL
UxM8WIS9NEENLPs1N4lU074m7TKb/a70PRHUCatqSSYWw61RxWpFH/e41wMjypuIes8qJpkBHxdT
PZRK7xn3tX/vTpaDWMM8kJ9QCnmPmf+q9IoBnfZSR6JTP7eXIuT+Qzhurb6zWWe1ChksWFVH0qBS
dOBVAOMUtjIUnbi5RmOK9wwAhMintbgSUbUjkxdYCu16CNwOw6DlCALAGp/YkOT6iOLtFvzgx5Gl
9tbxhGPGV7ptj+sMffeyJeyWx0dQupdlmUevF7DSQuniCHAlNmODxcj8wJqZhxob3dLnTneKzvrT
Ta7KINrFzCPrFp2XjwDG7Ce656+T5ic/8UT5sT6k+CX9kcqFlYJcE2VMXI05CQdgOSe7kammJqcA
Zsp5S3FS2kytONVytH2CX/pwVZziTNl6UyiQNYqhXUDufPovsBb5JtiivQfHgi9MuvCcUTeX5Wlo
5clEXBLwcz5nRpR0R/TrWFDuLGHYZv2i7u99c/IXj7KBhoz1Ehjc7LmoOrHS9GSvp/s1IbhHJ8u4
/85BzJplv/N1Xefp9unfFxPzzlX9JI9NLmtZCB8+ohPLqcZE7mTnHnYckygLrwrDoeRcJNnVJuAt
4K7YqvxWK/Pc87c12xezUNGnIrZ5SK9YFj8ULfxRvIrb5aFap2q2mR76bAnqkt0uLLdQBFkrhm+G
7Y4nVFdByE1f8hWAacLPgLeN4EwGkB86qt29igGX1WzuTKwf81pcMlyxj6Vlly//dp9HgkKOuVYt
EF1b18K/6LJyYFT3vO31rkpdruzSdqQnCb/UhVzbt2Bjovgz05isnYA/1PZX8ZsHGj3fNfSDuuSI
0cHHpU6PO7VO4eTTE+H7qh+lcJy8VxNceokq+ZJ6dux6ahFkMGpnLozyFTYWg79Q5w2jJJH+FlvR
SKwKXHaUsqBcXo6Y3e4aTethah5wvUyaevRuqFT/ewzqb9ZJHRXhdBxENByJ+0T5J1I8TFVo8kTf
h18ib1yvg49pehVBaMwko4l2xyacLJ5Iw5+uevQVHf7+TFRm1OuwESBJTlBA4Lu4fwE1X3Il62nI
oiSuIKb0Q2kzi37dYtvSD1WfAj2XGJXgabnYOtA9lWXRegVWd/PGtEGj0TtauSKvw8DgmxnAfYi3
fBqpOCrA+RP3oDWP7sP7XPA1ZjHjONqiiGeyI6IOdSTSF39kNTvn04AukrfuPCchbhW8l9W8xKk6
h/Y8Pr4Fe3+KyzTHVU2kZnQ1zKCx9Yi5mlSukOx3SOlTUKOiq6fq1URsMFSwdRXLmGEYp3c7d5L+
Vcu+mqTcRa7pgajd2f6rAN4DwHpjQAE+tvy2m5SpPCm6/eQbQywHm3O8EvFpJAHi73nRHszJePrm
+Ow/2a/2ZvCd8nyHck7q9iknakW1gXJ2ys2ebY9GM0d84+PrVTSakUt8gvURNDEqaJm5YDBbY9GC
WSkbhS9SIyvdlAjoIfCTi3C9maPSs45/EXUOp3PhvNN8VtCKQGsn4BYhiB42yTaExIQpmE+0edIs
1Bg06HaEXbwFRsie0DMA0uSJyb8cSLmFl/wXE++js7cw6i8ig7kEIXNl7OPD8k0URBwMkIr2pkQr
CTrXHJwgT/ykOpOIAvL8TTL6JO+KvikCmZJhC8kMDxcpnyV8ZzCbQMWwVZlL8guGDkP3sOpsodjQ
XE2GZvBW72w7Vd9m3+IT7oc7uzJNbjNs7arQLja0Kdjp3EcA5pdXDhJF35XXb5Kkg4nTvFg5C++9
AD9MTPudrjHg+7x/kg76kwM1lwxDnypziQSwOjlKAdWECDL4ySb2OYSuqiNBiMK3veFyl8WznxsK
PcguBki8jFxnSvZPdWp2jvWCnb5whZHFx4OI04s5khF7e8Gd9A6ri3GmUNoiOL/PjnO/kDsHieq7
XQUkdQhAl7PUjdokfBapjaa93Bs4hcziI1uAQfT7/ZTje2CvveunCxfKzoGrctrkDnAWgQpmRGtO
Iy2pMCH5URVTl63jidSLahDsdsIIkoucynXbBUVLIDeY0+8EHT9gBeT5sx3jf0XGZbNVR4LTNhJp
7I1oLo1zrMlu3IMDVpc4VIHeLb/6kMvqCgCyN1pOPVTOxYJUDWb8nTMYLbRDrQz7XM4Idj4ivHXb
MR98WppWtCOYzj3tGbf6fJ0jFDgzII27tiNFwohNXyofs/L+3XMIC/LvtusU3ksqHiLHXrKn6Xsg
w+PvE+xUNsSG3T2QKemy+3rAmrQda1AEnMQlt/YbXCiprtkq5pRaXt5TjD6GbZJIeDMoG67tFINX
P/6/gUmFJ/5x1+Up/7Uwuv36aQUGjbcuWF3nygYmsdECunx7lKqO8rk1pE5aBWcry7EjaW9ePc2f
njJRI76zQJs3eayvaNZzExJmnVfYzsct8uxVE0o4O6JAZF/Xip0zvuPkrs9y6iam9mgU8tCFIc7h
8HAq/Q654PE/9beoPCfshqGvemR/Wp93+sLRmBa0QAv6Vg4NnVLZXNuWPHsZPU8tiMSXEvP4lg8U
I0ts46Dr7mRewHbS6kFrsE0oEl6LcFf8cSe1xnuwRqU94RPUxVphD+rcZwQaso5fspg76HavRX4h
vLI4UVhT1xVY453bwqJmNDHdfLAXnmFyQLHt3jIdOHTfK8EArz38/XPRLYZCNpLGajRzZkpMESfy
Agyv0Lm2tQhuMCR2ckWraetJHC3mkD2hlkfM9HC7JYlFNR02JuC/nrcrQbWhyzCAP86l1wqXtVnr
XfW+1oe8527nzp9cslmcz+1/U79sBlRga5DWyvFiSW8HtVYVfzQfT7sIZVVtkyILoBYuJJWdbPLD
STmMqzwWJS8MQ5p0qH6j7Jw65yVVXBiA5F2w8KqpLj1X88aMcdJ9w5tGcYHZ9Dt79p7brLFA7ZAA
E34X97m1PL25ZD40fEqrDSf6/vfab+o75x0wzHo0BbDGi3OqW9dvdUrZSbRPtlqzzRCgT+BQk/Xf
mvufKGF/WSvpeZkqJ528NCsBggql2L0QqTvW8L3b3FF0E6FirMn/5Lsl8tBJHkQV14vUoKpsK3uS
I44qPVUf5lhsFDpOqY9xaAjXZ07eTtPzNWk24O8+GF5JflQmk7v7aCWEEzgfhcGciGJ2w41+GK9M
aki3O8OMubhdW4G5Q3BGccWgL3bxGUtuWAryt2LoYJylja+aLfVowx5YLeoGMsSKXFHvz8Ht6PyR
ti6Rpxs1h//dAvh6FdfPRSlSP9Xnqn3OCoBQYWsO9sxfAq18P5LyK1sBN+LIGI1plQ0eLzugm6K8
xuNfdaLePQI+LuuVoAfbw/6grJkRmvXeGZSzj6lYIJtzK3B8AFtNlf7iuMrDXCbpiueagKvfeiLl
haCi9WQzqfxs7dYuwFI1J26Rm/ZUZ47nSg6VwU4/p1Obael/RA+yhY4pBsJboTQWcsRnhP8IvyKm
mPHcTw/hY127sFModoTV3UAn+pKt7oXWT2EP42bw6ap1rwga5PXlq6RGu0uRBSnUZwrXaGByM2IJ
D2xtbTO5B3ccwvREk3/0rpHBovAcGf6O1cJJwWnxPYXwf0QYjQVfVt9M8qwoWfdAOx8lHlonPSNE
aBByjRkUD3rU9KsZL7/Pi+O9sevmqPBHgRCCaxNGER210v84JcGm6N0eQHBloytaJBhJZkrDr+6o
krE51cadp1sQ4DI9dtrh78kESNwtKtl0UZTe9hMw/CWyutTvFYreX09wn7Auj4nyHH/XewMySRxG
Flxld5o8hq0KGoNgovjL//scEYPiQ0rDAYVzui2sd1BjVMTMpYgDGgkL5HaKsalacwTsnk7R5L32
Fp+m7UYVj54GW0k57BAIQtwF3bvqlf5b6hI/nXo2gzqraS2AJw9mTy1VUy92luXU+drzcbuEuo+9
IiWY5CSsVmLqFPC+BR4goIej8v1LR3bLIqnfxwD3XIf5Juz+Qzch8aUcQ4hYyJAj/veLd+drKkQW
W0a8lOE8oJtCgYjGQkk+gOm7TOzXcIgLeppAQSGQ+1PbZeAH98GBMItsid8AW6zw+SVFIafGDLTj
OlrT34U50HPxVCpc04YHJD/xdGSzgy5cDOI6bgN+YSNAX0hqj2Iz+XK/+G7VWoCRQj1d9yLLnfyF
DkkemZImvMYTUr2vSC2y4orx8owOA011EfYnLJ+tMc6NaFYA4fCX+gyNX2k9s9n4P4nh71zeJ66d
gRuY7QTUys1692smbH24Mjo47VjxRipTmYyHmxrld3oCZpYqMs0ImiL1XQneltoqlBohu7p0J/qS
bQ0NcDYWEYF3EmDJOKoJxPIhBXkLOW4cYx8rV9VxzzOp52aVDeDlWgeoq/LaV+OTgajLRTXTSeXc
iw88mfO2TZnTiYcxBT+KhNmjDBdP5Gu55Vxm98nj61P3ABFNmxPUROi8q3sUJkvCZoLLHlRDxZNw
fKgLGGV7S8YMxUoMVLUBjVD4vwCUXESZdklrcrSmpbJm3vt8EsknvVxUEOOHnyIooOWZQnUsBbIU
yRfrkLkWTlkaMiEhHOLfPpmTv44jUpHlXIsRBW0m5R2weO81oWZdu27mouo3NXX8Mpmltj87l/WD
aew6Zv7D3jjGl8zhdqh4cUZiSB5NkKpuJuBUKAU1Me4H2MRRmCV+VqP+HKqq1FXFFkdRM3AmjI6K
HiSosdBH+B81y5wcnTMuxwUzXNhsDV+I0hATr4KKtFDxHR/ULNO5yvGoItoZtzrD5+gQKXp5TvV9
9RtSDIhXxmHkrxEmTvrvDoOYv6saKNMGoIKq1xPIDNfpHf6ko/xqqIBdDYmWEoGyZQQA/IlewH4l
TytwxqjFKkeNnjOlWMXcZmP3wZG65gI4ONLjRR1dhaqj8scJDLJUwkTJ9oraUqcGIwx6VDLKYA/d
Q4Rp90XTGNQ6aQD9WGP8ZoqrJDXINWUDIAC6JsmsUhj6I6n0YgUkD6jjLrmTORX419Puq2K8hX1X
nEnU50BriEDzhpbMXKs+IprnPngWrVm/vcO43HSns9y5CFhHA3xwCaoZGJpyQMXHevUkVcyyBDYS
hrHRTDTQ5C2OBloKDoT9hXPBgGihkl+YBK5qctw6iJKZu2FCUcpwflD5PE8LXY4w5CFx8+vWcUoj
tpoB5KA2lm6KiAf3O5XMjViNDc0eFM01iVgpG1f3xURlFCGabXnM5kp/gN2tl+Q0GM+n5KoKdyFw
D0GH33nxDDawlsvycp0my2TnEQaYLBZ8bA9hOS+dLOxjzcdtRSUUsOo8vWkR4/L090lVGSvI/4CK
AyJSobIMkKhAY7v1AQWx/mBnmDoQMjiBcgAwo5hu8zPqZx/5G+ei/b5TH/xzXVLYFWUNkwme/mpk
176YnJ3T2iIrCDCo/u+VK0wObRrb7p78ylnpdoBxcdd4kpdynT9mnoMlgFuX0AKBSC0+8qgeQ6o9
6eCPdBnrNVQu/zN8q/iLRwPyvrIiJgRxeBfvY6acITxO+P27XE0gkCKvuc5IFTcfbYAZrTXNGAed
/D9/JkbYcVmq2yogykQu8Z4AR8dZ6AbZmRgogStpSPuSqmjC/9iHX5opRCBhG7omcLAphkPKBYAU
0Z2LUZyi3CQx/aAIYVWK4fTkv8NTed4+/31su2IO8xSOAtLafszD7/4JHzZ/9IjeU9xxJLsT8aQF
juyMTq0TtxN2kL3h1muFoXtL9M9lbnO8zUdEP0DoEG1XyT+0vVRrnK8BpKpVCNKCML6ZpaeuhLBC
g87XEmFa3qpfCGQWls8KZZeBTGBkf8KUCjyIPbC3kcC/Qw41Cn/kwL8Pu3Ya/BDC2SLz2PfYsqS9
Kf9PvS1BLSxirhxewgr5amkc6gcMhH4Cw+m2hqXmx+43L1vKmzGxGD0Jj93HyQDw4emneOLNRt63
iv+tfRfKSNDxx/eUEFWAKwcNVU8oy/2XjceqtEOmwvOkaxwnmpHtE0tTQzCkx8FhAxlpF8W4X8sA
+2Ib2uYiq8Faif82e4+NoE5/ggpjhk3COSfsQ77Ugzw4199ApOWNSb0gjS+YmTwCS8PIBWObn9DJ
3SSmRYQwtLdLz8wyLsrhcJb+Li/s0fFIBjNHHj3MUxjuS6mPDPV2p+HKCmEHRqii6yKb11O0K2Qm
YW++yRrB0d209N6Z1oOe0T41PbFYtQGOiM72egOeNfWglnxckRKQ8bQq+0Jtgl10W4GgQfHqr06j
82MYtvLiARbJuMyPcOpwVhrCVgl7uF7C5/scO1jBiRl0WFkgzmbeyJnXtmRC+LfC+jeXuwCYTn/t
a/PkO+HUpwn3tbrGP/tmRUxa1TZmInyJSovE5Ud6fX6RZKyqhXSM1gVgRgKbC7P4Snismo5m0ToL
WXasJ7Y8dWF3serZJeCgScBU4KYylDs7WDsza8I797FgQRR80jLy/TvVurB+nT36wZ/g8WT5TC35
MkYO4qY1baQcnEdmMa8iZaeJe29NFsBsP+sKTZGZHT7qDupgX0NzALHoSlwsXdCmtXqo9rrsqyrn
/3E6jXPKwmMI5/Ea74aEylzgxF23mc3kqYuk19Ythn3j7HWXksTRTYfvwk4WIJ+SZn0rc/MoUOe/
VXWeTYcuzcWhiTiTWssJJBGvbp/i7YxlV+TuRs0H7V8k6XR0wrW3WPCLWWJ4HlYto+QU4FOnl+tc
eEMngDeZzsmMSPfgeY3IksM2Qx8nmNzNatVCIpE2LKyQJZ+fbtrXpoUXxxHJKWMMAG4x+4y5aoe3
UbSJ4AKolxlpIuvxrFf7F5NSw6/CvGOB1aEbDToxAHcwaDMiXERs+C9RZ6Y6e5v6xEcCXqeU1YHr
XapzCJYcldsYzap9HVQAO9UkwW5x7JPMIuovKri1qUKKlmKG9OAiu3ahtkvOOmtn8E/5ZykS0qo+
qgqZ3tVLb3j+KahtXZ4ZVGZfZrRs4RWYP9Scdzwj3BlOxgSM4rdCdWwgD9iOWEcqqSYU1bDF8mMs
phuuNioe+P/3S8+XTf5sqRNXX2qoiDBnIl/0soX3eArDHiqZTq/nbCj5BJ/YAOxSyljjvKQpUENk
2j6AUDQyIByPYaOIURLjqhxh34hHw1M7YBLpL/OG1HPLL/YBGLkV2BAqWAYbQ+wgJPeArhO2nbGL
fYoUAs+A3AHhOIot1qBLHpRKqgjMGYjUXYD+8VLQPJVbCiLHwOG6RFE0lfT/YaX/sV4NSVy7O8i7
xfXoypz6g0++xxUnD/tqd9BJ8RVHbPpQgcyavzzksZ60k5yYwLUsbgiKcleqbQ5k7X3sxEPZzBwW
qmxC+uEKoD2XZnzjQ4XMLlqeZN9NL0x9vGYPqlSrZRcHxgcbTGn226/l4jwh3ShUZsO3DLltYq25
aZQRgCw9qok3CJ0b42RSs4sk6OzcSu2OK5Cy55aoSod/bPhqaLv6Etzs74zvAkFY6JezBZtk9ITe
SKexGXJeEfZNf+zJVC2Apu1i8tQRG9MP+6ML76lOGhzf62pLroyDW6j0hAkDeghEXZppA2xdmo/z
TsZIukmrzCXori2gavwlgWjPk/273r0QMJeSvZMqroy+dCldCdAny35Ljsw9TOdFWjVXsLWwmzbh
+vztXIvyCN87gcgjOAQ03h6rc5ww6v91uimZ2NUfAaEgSqeT8+AUKEs3HBVi7t5JIbvAVJOE/u0z
2dlV/k8BDBpZb6R99rMF9qf9dvka9bgJ6RGIEVtediDfL1vp8xJzoy4/uvhbGV3KF4DdRikqW1U/
f1T/EDl+nG+0odYXVSUFBf6oFXuTFMhf/Pl1jj1lAmdv+a0C/8zVibQZGtFAroOYaVGSkT8bU15s
muqcMoJSrhJq3Qr4UYm4JJrrr4D02eR5WlYWR5DhMyDhXHll9G04/fB77S4QJanjC/1UU03TRqA8
ptlbon+bIZkzSATc/r4da9Am6GMTvtgGuip4a8MnyMNq2y11YTARVO2yJ2vS7bKPG2lg4aRYK6Hv
Xk7sAVCRIhY7H+p/VLAEggvgeN7oOt/zFLGnfuaZpktQhcIMqcGQ7bKHbh2x5PgXRh28MjbBLOKj
SSaIshOx1T4s73hLKgRpQiB4sINUZVrjsARfAP9N4bJbS3vpLAJKXCxSoR1NkBWQ5xz9oFm5Vnxx
ajkbktu9kE3RSRa+OPo0def68MEpxMAaQFP+MfBPtRjMnBbkXDBbbuGiEWCsBSuw+Uknss6eCp/P
JpnazWEdBs2HlwKPxpS9eR1g6NQ8PqlxyzC6wwX+lMLF0vF8QHQlFS5mAmJwIrm+C8deYu2jdYXa
b8ABB6B3vCp2kfuMKYPRGnFRw8A+dDuQHr/F2Ebu329F3oQS77SA1NJnDn5V90RHZWQQ0ne/Qo4T
fZ9gBCC4ryqcx8LogT8QMLwSfxgNMIb+KnDZNaQbQgDbUVKKLHXvBJii+H8CZ+LHPZ5owKJ1ew8a
wW/EqMR6KCoJTOIbDfrCXgzxcRPxyeGhW8WfKhgBgF8uyBiq+ARYiMlbaXctgABGkWwaBdxTTLUb
BfMpgzhPdhg5Kme1cePTbQhAAUpS6GKi6V7tahMZr1e4ckG7G+WNJeVF9ovP9g5/tCpVu4jwuW76
6ZHbiy6UsrKmQdGTlHpzJ3ngBAfxvcwwq7LsAgtrpE2sUOYsjwznrDDl5WKXm7edhWKjsYCept49
7RylWpV6fXYrHd8SZP+b9PL4ToQnvc6F1MZaMKzYuuSVS5SdR23cxQ6xQfFTE07BBi04YsdTCW4S
QpHwJ4gWfYOfRl/TUvivJLNKJFrPwQX8PiaNlQWFWBLSPIZs/mhx1i+mHV4y3m6itkr7wX62budA
vZfQiAG8TYvs09mabyvChjxxcYpL8DgeIbhxM0lyW8++cZYMksgyrLJPdr6GcH/EaN3dmR/nXDLJ
JSc5bIya0z/J97zuZ5/FZ5d3CqyiBeDz1WuS1PhljoozAywcGZj/3gFnPtfAIqO5skpV49M0Q96s
Cro/NB0nYHxr8x1Ci2jdayLM04xnELVMEiPF8DeT4jNTXDsA/0y1+cNvuQfRXHLbrlFWcJDsoJi7
iO1T30iubBhWz2IEUyPZIcXiCogCLPWSz6SrplZqBVRETKoRWbLKMOk6LRQQBZe0r39j6smoj6tl
5qciJIhR2+IlnDBtGq8x4n+lPX6Dtt79LRulTdwlhjife8suxV2KJG2sYTlHKSD3bHaZNf8iGOH1
MzQito3LEDHYIRNVwHTtoL9nzcstQ5NV+eZG/Iu+ty68lxGzXkSl96iEeGmi51QPGI24Gcd+DfmZ
ahUamqvn7hveTpIXLucFZ3Bg6/cOjpVyeklBg2Q3Etgjsxcaa1+Qct8gut3pAJSbR5tnnvTr4qw3
XkPO4USobyF5kc5pEqRaHFkwu+cBYkTdBoeQwiwZ13qXrWj+hXVbvR48kaCYdMr7nD5DLyajbjr2
0IP/fd9RKcx/zeTrNxm0AuvfSNlWdGaj98Ic8HaTfs72Z9iVwldKwlTR0KRlceJmTmv5W5fZji4V
WaOul8hrsJSrq8wkRLKjH6GAJrpL5TyezZRvp/eLr9fzWFzeQ93WDpB0CjwVnpkdJlCwFbkbdqjT
l/Tmb23T+bWVM/+nPVlgwDbG5bgBOJV9z6m2H1RZ9tC+53/pHqOVrdan5jD/tI3Zf6UqMJxNqgZC
eeAsuuAKKofP2r0001I/2O/avOVt7XCWX3lnkzwzZDju9glsnT6BqB5F/pYY3yuGIXSUDrB3zOFa
zm6PqELGUmJIyoyOPD6mqlCbnuMdTgxQvC0WvKoxk97B901ggwxogjVpRu6QZEqLRXYV+UFemglX
q/Sc9WZl2HQ1ZiRBenw65Lk14WvLOIBzFm71Uy/W0GgtwY8GvpyFuvvcEseUMhYvyRGNF95Wytd+
jWRL/rD/8A27xE4FhszxByInPPn8ucjGU6TPlWt0y3faugURenHZaim1xJMf1SllHPSpfN2Dt8Cp
3KHxd5pxwZPH8/MSGCOaxwIZTDw+1knk5x2EcxzVw6gLIre6OPwnzpJlchAoe9mUO8ZwGhlG95Qa
QGsCcQvmmgHT8bCq8mfof/JmrAnSCR0BP9i3NGRLV+sRoEeL+mWTwHW6ACqZo0P16ZdN1pKJAwHF
VLEwReKn1yYjaAJMZcpI6y2ACQ1vDeedK/eHjguehOics/M6viBnSFwPLvMX0JoB9dW0GB3505oz
+B1Vlh4SgDJ9BC6kEFLGzaOkMqr9A01hWaJbXHYSXqTp4Mh1xhjeX3bQobxxsAkqZBAoztzsAzRb
qz4fX5zRJPdBDv49Mx3bZfx7lLwHTJsNUjaJNJNKQaa++d9V7OlSOCQnjGAnOYHzGJcmYuS5UR2u
AQn7df7NBIOUwfed7/eaEuklw0BWO4xIl6SqAXTNSiqL1uXziQL2yozKOsxUC4VGgQMQ7sEMHw2U
fbJAlu/CrPD4KgWD+80SGaOGFiwlhuGSL8QjYZkKc899DWgqO8SWTeLzrwW05hcz5GMHhJUhmYLB
QRHR3CD1h+CPAFGBF01jHyLeEZCGudVDsZzGI3yFUig9axQpG+afwqUA9ZUBzyhEtB9Yxtjk4Y4c
4S/e3zvd+yQT6p646Z666xBJ+fyPplae9ucoaklSEreX55bFrCyeJJil/diqr+zIcJDf1KNl6igw
Zw9Q65wkCR9yU7tLzjfkrZd+PKjyzDm406Mlvem03tffAAGRtOIBBGJnnvYgN8F3iavp2huHH7uB
5tkA2r+pRUnKAUlEieRptWWYMaZg4aOmDO2/61my5j6mInIZ17l8mTN30PJj1nMjsrzUMCaArk9a
/KYRT+HJyoY4s4TyKaNQBeHyJTxhgG34BEmatvNNZU4irO988o2ObhUIjJVxP9RGpJFe1YZrh5/p
05jp5GrWkcwoqE9hmXd4yFg02kLRq1qWLhExaNIPbB2d4GYuuXeJnM77P3W6UGdhXZV12Zoum9vT
oxVxLjduUe230Tluaouu3yesrBRVHxUH3RU9ywLqW2ZExaHNqjaAG57kg88FaTwaQ1WI6pJ+GPW7
ALs+z+3EbfNKM8ejrFQjyvN3Clun6jGnx4cdrHD8l5u0hrzHyHwoIPEp7g/gOh9omhbGYU9IXagL
GNvcznYGDWusGDCSP+jnD962QCun+sCAGaYtEZPoz6QR171W+fmW+Y8vIbTltEdHbHvQ+tjNicD8
xMlnIO6kkVjIh2QcjHu81ydjGGTsAJjnIS0/Mezfuoed0ZJrZtx0tcl1TEdSlrtpytCUd5KaZ9vm
bL+M9JoaUwUWhnzaiOFYn3oVXyNSDSXIqtgke9WWkf0K7xJ9FOxPtBmRzrRt5wl/OfEkaSbu+iHM
v1w2eQShKqWbUgbj5Um9vwFA6aqpVwSzcJOs3N4Z4TpWcofgDluHa9QmHQtBmDOMlDI08C0S8CJD
xc3DkGxCXLqt2GUXlPHH20M2erMeCZ5KuZLOsL4M4S4qXxTOb1I69Y1ClHQmPrCiiQcuSvncvo0A
xj1NYRo2DpjIt/IdnHvuk/XjX2lMlfA/H8Bmw4C/S+UGhVJru8HOefgoKZYhyCJoeMTWLYpTIKT9
gWMzTNkBHAUw7gA3Eu+6OiKyb3bzehfYmXMYPFWjgfuvoqqlncOhW69y/gLut4EhBJLxRA7KH1GD
HPH04UjyWg1rn0xCq8QrpXltDhGLyMVXw+Pz06yHGaJTzP1TNq6ANCY6WtUaBND5VHNX7ERHKfZI
RAsmYiitVP6dUTx/pjAGmy5+uJgbfAQ8aJGcQ/37dmJwe5iBdfFokRwZZw3pv4ZPSmS7rsTlsIdU
brv3pmy9bmbGW1zFSX6/zheACIdIVFcF5bRQDCmucQ1s5mKvJk2ab5NREHMoUplhqMBPKiMr4HnI
OqWM/K99GR1Qp9mqwYgiH2qD+dBvEtlzDhiM0RHsxUQiJqOWwmBuFlwhjef2xsr6h4L9/xHyHd6y
nGnWxFkoEfZLwktjns5BceCEDo68RDiV9ZT2PQYjgwgaLim4G/FydqkyMUvFfNC6D87EqtnzdQvo
mxlbjRlO0hj1x/pg7Dlivgu5Z7dToP34SUTWdFIa19GBrnbbYNcMFKKMH+Z+3EzZVctioo+OMexi
U5gMNqO4Kqb/vcKAxU1O3QzDHyjzX06Fyz3se2RaqnerZrcV20RlU66hO/oixwecUpG380o2rpPk
2hizE2ccH1GK7oiFGeK3FS6U2vaInBulnjHI2jRZyGCZhTLmrFzb/jfLQn54goTeE8koadOVpgyz
CT8MXtFiR0o+9giIghTnJGWiJsot9VdYkcZz5m9/k9/BcHrwaC5HvToaRGCJE5OHvNt87xU8wD+n
mO2sElgAj5TCkXmiGkD+teFbB5H8q9F/bXIYTjA42D8/51FOixw8JmF02fOtWDAAY1NT9lxpzbK1
ZzdtlKBceSjdPGQZstrxqu76NWeXDvkCP60EFT5T7mLwuzgkXEgi0YzdJE8OTnnYdpGXYICUz+gb
PmWwPEUOELEZvhEagwRTpuKISVMHdjirzKbsRW+VGMnsgzPUVxwub4VSR+SrKuA475m1VYJjF9TE
x3e+NF/ho1n+tSC/w4aGO1qLEBnWHUbABq0G0/EMqng3B9sbP2F0dlo3xDEis89NR9T8M0qIFLcM
MyNqsxJ5AtG9jkFw4t87Bg9Ap0/89i17+LXRk3yyRv5arCk6pkRG5XLIDo0LjPMzAktmH6iOJT+x
ShTgjZqvGGLjMODlBPJWWUX9YHf+VdmnedJFU+DzXeuQi0W0d59/eZLUpO6e/eYS8t4syWIvzaTh
h+da65WUYhj1+6GyJynVi+4orfnKtA5Ydu7LERRKwAV89mOOTLWKPYu2Lb9K72lLyTCbPummZv4j
UkM5QyGhXQB7RDrMvt4Udp9RZ4hUu8IrVSuBlKe7Alvgmp2jWGSUnOlILJUzxK1JZKYk9NKVMziy
tS1T4oGYlT6W+uW7/dnNaQs1TjXFOlzLJKattOrRXCh9yMYvVnGO9/+qsY/NfcHaV6opuS5PR8Ba
60TFtXECMohfuxvb3u7A3nLpI+Y8co2maFYDrgogSkYPtAjHlqE871352MZQSI+JhgAp2HeHEqmc
z3u4m6RkMOOXoDuaBqGfmx6mZc4iOBamLstpB3GA01jrgiHMCcBEQ573/JvsWUbR5KO6F6XdSslq
XcsHen7D6+rTWW+m4t2iUKuWLiksaVANpidBRYztnOy5Rm4AsXPuognZS95igybVf7Lo7nCgUy18
qjrIoHpqAmV27fvDY9PjZLm90Lrqqcv1pMFl8G+94q1cEez3LeH2ma+cEMJWykGSkaHlFhAG7Bd5
mahYX7M4oajFNW786nu3XWFzCXy4BYcXBTxDsjdoJ3bCl4zd0cbOkaLq/g/FSGSMKipIiY32DmqC
pvN5KaopipIA1Hb6TVGIVXm4ZbQ3aOu+k3pXacJ619DPjmXy6zCnzbwW5VQ79CZVSin4Yf68cvyP
iMAQL6xt8lIeGmloPJayicPLtJr+wWJeQx60EayLlmhWdnnfiP93pdUCocp/ZH/6Nos+Lh9BqB1x
S7P17Z/ACIBGSTdQbpIn8VLq/xIBoYY5fX84ZVpPPlnlWizQWlqp6I0WM/RznODV3YsCjN4oFKw9
MDuecaiwye8HIqpGynPMbpJTiFwarfMU7rYE0edz5QaimHiG6MIk7WlSXXVls7YRg2FMDA8Q5Cc0
rqPh/vOI5tmUVhnBv2JzFvPCyFwPjH1cNr5KKaia9rSIyXGs+wKTBcRji5bnrSckRh/Pkj/tXYlH
TcWhulcXfZDIPkeWz4xB0c/5yNsaYx9Gzlgb9Tv1utV1K9z18ffOH5iJZ8Lu+pLGvOxzw8G6w6SC
jGaHpzkLKc6egd9qqOSXoummDAf5DsydKU16h033p97OT1B1eJKgJJgZjlOEClpzNN722r/cBTOh
b623JawUJKGce3/TcKGAs3Vu6rDdmIQQeJ0s12KQPwzfa9dOdMbAy05OAIcSrG+/lFZWLR/JwV4f
Up9UFV+43UybkdsJdQ0q7JgFbp8V2DGvMkQo24jYDB3r31YamXXau50plG+7yHCPA0TqXtmKMUXc
b/O5MAmEmaFQozpTU/YLS15DpUKdjI56H9bOw1KUONjtz3VITXRYWllDd6JuSA/wBOCnNJw3/V0A
GvUbsmlrktoQ1hAGKRIeaKuVEVGH48x6zGHBvZquyA0ijEYgT3jUI2MwlJUbbY9McWRbg10vvF8g
Cy5SJq7smC4vs/Q0zPlN/oYdihZOJ5rgbKME14AjOWMLa+Zau5v8DbRoSbIVTRavc/nEKWcyc+nR
OGmEb6Lj9r/14R5ehtoupDlbGdOfsNvA1aga1R6gsHPy9QlItOlhGGdvAC1EOsXfvFPjHZkz70jG
A3yMm/3DdScKSjjsSsvLugp8EDkoG63sm3rrF9QC+GyLMUqEdyT/1JuD+AFv6Ta0VC3biyjyhQ7J
fdrue97YKt0G+4l/FbDj8rX14ADMxeowY1+zsQFTIloRzgNnKCA9EDrWNMPPp5DyCF3W/1nuQstg
lb8BVNt1JNdyvRXqWnr/ZGQkzcpHjUFUv0d5XYPUO0Un4tPrTo/SdbMlmVEXuI773XOf2HWdGRP5
Z3KIk9S/2GTVWSjXm14uhxJMLTcnIKJSZgUgbKYRyb02unkGuKw9lS278du4hkcKxhZIroLj9W4z
AjTN2/7ZjlZjzTOG+VIIx+Al/dTesPvdXeh37VyW4iVoyxzCCMctf5MkS1Z65lThBPYujBcEOnTi
xD2BiX3iaIazgurrSm+sUqgUhquB9T5p9IO0ekvgr5nmhyGkXSHc5hECw8oD2iQd751xR2hpODuq
91p4GBMx0fWSi7xmHlHZJ+sq3gYSHeFJwy6XuVpDhWoDmENyHis/3BPt2d4bf2/M6nspQ1ACCVx0
KQJYfLdBkRw28CfRvEpIC6EXMw76civAc7RxMxt1zaenDuABLyks35C+lsMZRq5HZUJQvOdV01Ec
3eBCPbc6e3eplQSnS4+swf9IeOxo6aT/ak+fKyYUjL9U9x3KpRSjGD65Z5H0Ns6JURjpHJOIIKH/
YloqdxS3bKAEu2X9v39KQVgSB34SY8LkrAvueMEcFhV7FDjjVaT/oOLNCLr67MjsfEJPsvl0Sm0G
4UTw3eewbGE/rZkuzpssnzfA1sFcmIAz5DLkxscDbxBO+qX0GpFwH5oxntB5UqPipSRwLhTbROQu
F2VtkIsMAoxvHhE63fxkEKa+9DWSKrOSgjg3CvvMsIXmqaPxG8Ilo2l2YKGLRPUPCbMid9xhn3ug
6Xm0ESkBxU7XI9ny0O60UQ22+38NYLYZlgJ6g3CLfp7ZqxYe/fLDtOM3B98VG5kkVEhU5rQx439R
NS9RUkbgx/HE3bmirSRwSTpdr/SSF7vmSk8wPlimDhZZf2Pc8RonZXedg1HRz0JHaTqQjTqrZQCN
p+P5ZjQOPEpDLD1plE5CwxZHwVc8mrQsNRrP4JyT4N9xoR+W0EIBlJuA5+EN5jdkREfaE8g3ie24
Q/TA+tqGru5kJ+Uq1Na+5vfpDzEN4q2gEJ5aSFNK0L0r7sQlpnOoBuTuU/zTRR/++RU+9y8dnfn1
6vv/uR0KGV3uUuYaSXXDxRjZn+Zx6Dkl2z4PpZB9qfs09INmHJ5BqwG929aDnPbWGVnQOfiTHYyV
XW8gZ0UMVkL05Jt3i0kUPzzUtsPRb5HtJaTFI2bFWtWTOxxY4LlyviDQePMWZR9sNBaZ0tjM/PDy
GnqJJZ+RdkENte2zI2JA4m3xzufvoDzw1q0BGbAVtuL/kanl3sGZhCgYOHdr+I3sRha2sxIdU9um
TufoNQmDDrVXWUVZO19q/abixHTJgM06qoxQ2CmVioA2IneS5YurPtl/EE9A8jCCW8lVIqGhwQHA
f3ciMc+sE+9a/GQUkJvXTtz6FY2p5+cqAiWtWSLFLWBz5FotrWgCHGaV51nSNH0CN8YXjQuxXc8E
y7sWVRL96Yw+IiqdgdGwTcb1csbUZo6KgQQD6Yt2z+sppup+s697jgvJWUuhVG3I2SyycCc+71l0
obrCLejQjTofPfg9Ldq6P5coohdnWGcJp+2Xg5XIUYEhzZb2neOtLmmZHN5YkIkd9v97CgoUq3H7
5aUVCjLpuByBWZlPk9eo62U6y9dD5vg9IGOPwzEiyzm5K1pDhSaCcSsgENohadFsQAeHlVzofxIe
yyMK/z6mwMml7gC5CqYgyys8lqZ3IbVLOu3GJRaUI4ag0JNarux+VDv95wO/VoUMyasNCcxlFPLP
YcSpG0fZEa3ciHFIYLiB9xgLCSi/1rJcDaroJbGOYhEUqPKr/GEpcZ+QtRd4S3gAluwn8Q+GrVW3
B52BuFXZXwq9VpBZRjhrpLoXzKcpZppHVXwed8xzS7QYSj6J/RRsKPDnx/yztew29+2mhZEe6Xa4
n9jq7QS1W2XIaenSpIgA5hr0CUXqwVig3gLq26xa0LFlUwUgGSDG/2HOhjeQHbTUuOs/OP5OEB3k
MYkFefA=

`protect end_protected
