`protect begin_protected
`protect version=1
`protect encrypt_agent="FMSH Encrypt Tool"
`protect encrypt_agent_info="FMSH Encrypt Version 1.0"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2017_05", key_method="rsa"
`protect key_block
WszABqHa//glMsTTgJQLvTDO3OP++Amiiy5Whrr0M0s5V4LiRzgZFqkTLWVTQ1uMLoCg1rJrY+h+
ESr57q28LsHQXFEYaYbZWqa+gnqtlV1+gfZB+ettpTgB+RGeHU12XpPVVs6P/rxnd0mLYSn7qAiX
QYLM3xAeHRvz0WvXwsemxVxtvbQ+Hhphd87iBMWYhVHXscz1TDXNlz0qMWGCMVD2GcFTjxJs6IVp
QAIUlwcbQEiefs5D9RW+Feiwzne9voN3xp5TJhNPrc4KrexWkMBdcFMzFBPQMymZaBu75Y3AVTod
P19WL/KLROz5jmY+IQW7Cw4U2zlOeFOJifo9cw==

`protect data_method="aes256-cbc"
`protect encoding=(enctype="base64", line_length=76, bytes=71360)
`protect data_block
kx8teV4EWn14ABd8bHKoJ8CMrQEtLAdobabrdwKyRYYAWjoKexkLKszZuBQodItj24C/ONGlb9Qj
19D1fPxS6H0Lh5QmjIYVItN4jgSchPDW/GHdnmISLCjQyUbLXuP6iLVb93R9iQxOFweGZyneNsRP
xUYIJfG7m5KrfylfmwNSodczK88AnRsL8lrNhDxTXTLHo//19nP/A5Dzn64FtB0DKIZn+ZKbZXqm
cGdxuWMa9aEnoc0DygjoZeF4hKrkZlePfrBpzw2lp9X0e4oF+jeP8NiWvKjYvLzsPCnu8KeqSuFy
tWs67EkZYuLtZZQK2OqxaUhtBliAXeF5HsmAT+wbb87fj5BUu/+siTWZbkXKIU1VlMjIkmF1sw5V
YhncPcUtOgaiPfANVGFzo0Iu92YJd2/XEWBDQ7NLZuAOtH4lDO1dFIsPPI14YkuBdL47BtuNzSSf
xg6hTF+zy59tbA4UaZ81XoKMvGRpu0TqpDiqw0Hi8RB8DniWUCdwkgvLujcpunGs6D5fyDqsVQhF
pGFyg3ojtnPNF+q0u8+hf9GdHguUSKvI/SmfxanhHWViuMUv17QekErbYTKiieLA806uGPJ9QqIg
sex8UFVPegIV+e+eA62WkMT86m4VvWea/vkgValNxZDoOn3nr9AK3XvevWSn0fQuE8O9sGpBXwGz
i4F0fjQhkAT1kaxo1GJPmceS5oVdvS3QBbozjsdGk01JgAdvXo/H7H4wVnqHn+BXsowTg4bdEwj2
QUWp/XTFBxBG3ZXR0FAFsjoYMMNeJA1aGNeULPIyJ5OUeD8adxld8h7ucahee3wHCls7F6t553tm
Nq8dflKunQ0fTadUJfOumdJbjhr2DoB8J1rLETzf2v0Tl3FNY0scQCTwSow9HhC+cCGIt8wvXh++
SbkSBqU8alkUwGP584WLGWAEK4H5hDBksFjM4hlFumAEi8NwyUMqMaAbKGextJoD2S4LNtHq19BE
pe3xRRZnHAVzWw9aDQu1PgRB1YuNAu/efRoTTKqHICj2XQk0Sc5I/h5vp/fWQxorjwnALhSsvfsr
qk19o9gjICO8jjEA3OnKjjDDbJiOc7qbKIllqk79tvs+IXKDVZMDwjq2E0s25JWoelkE1rrQRW8r
GHhjID7EjD5uOLVEEl5sVsa2Iatrm1JqT3g6nCIQJyEWvGpicj0EO5qE8mGJMIIAD4FqN8Xr4ovr
04rxfkJNt0PbGJ5YjM3X5D/q8XBgIf/xbxGSf1cRCgvv0GfLpJV3Si1MwBKOSURK1ADUaxxAD6e3
Yj6fEu+YNUejkm97A5IMUyqpFIhLspK9fvN+lBf/cZ1t9ocb6lSBJaJkHZSPrenkry7BS3YJKyFw
x1ykYirt9fYvOVqf/xHH4/oZ7L/wVS8rpTvrXOkG219O8d+AJ4zVwjcQN44+vLfT9CHqkajqbR3m
Y0Q3LxiyZek5V1qvnd1iDSLcYl15LafV3QqJCM/3XAURk2pnIL2oVDi6HTzzgMy5kfSGFt9U9d4t
ukfPMnU2i91DnU3olU1Hz3vTKuvWOub3fKnV0EsWcIBcv98P7A+3eSDCcZnGD+f5anH924YuULcp
QaMsVjEzdGrOm72YqfCyvEi8B/WGsw2jzhlo9IJdoZ8l5rCUhuUNmdn03wkj8ow4CDzSlpdpz/Q/
nrCp5dJS6UNon0Y2qPWSHmqKlJQNQznoPzwJsPiVpaWivUJnf5tamxA46TXb4chK5fnxvu9jzUTK
lbSz6Jzyvv/juyLCqCEoVbuydWWWb3n9XuuQd1R4Xgej7cv3kuNbyvZudhooVBimVtwNfucy0A7N
wNvNuC/bCtB2fcBdnYU8D+CmO0WQj6axoXKmQ0T28jXcFsnfWeAObabLQJ+es45yBtHJIfSOKgXP
4zevV6giNs4g/xqUg6LVV8MesYZGQzfVV/cgj5EHTqZ+scBvdhdo6JVuIVkcw1YCa/t1hRqgZlxn
0aLnKb2pawdJdafzcZIJ9r/AUt1Xxz/SbOcTRuP0RXerwVVq0nh8L854R30F/Gal8Imgy8YfsRvq
hyUr4u2+zURu3qonYNNhQc9JwOlZYuAwh+Wwww4yfaDLbI7UjG1cXTnWBNqZf4Rp8UhUdo8WZhzn
gnH5VYzssc/vcaPyv4vqLkQdUCmdyM0ueox6Oziv/M9LkVq6lwVdPJKDmxBsDhug6OUdEnEwIZv+
fXR6FcHvVgmzZSiZIvyg9sVisszk5/RI6fnX3CqC7MBVYcdVl3ImJ1fCrU5jYDGfDTRCgIuziyPe
TSYW9IGFgRnVn/5HP8G2+ZmWWRQ4QV/GTaXQsvvfkSAAuVOXgcZm6L9Hu6zHnyfw5WMdPKyOe2nT
zOeklT/wN0aYnB3nCUB+IS6gqfoPMouzevBuQgYNlMatcCbqPSPZ7m2iQ0+9xB39RyOnI7XGjoXQ
pvfLxdH70KLSDLJOrBHG8cTh24eZBneExvxbE5cK0/2DtAu2Oz56x/8O3ns3SfVBZ9aHUkyCwvDr
k+JtszajY6qp5a3sKuVYVUBACmdieRfvCe4zCborGbcXtjpQfgzfAsh0mKu+MHRsMCADysjda6Ar
I0fppfmiTWzT4p93JiaJgqrgboDJumKLBGgDljqBH+JB9xRJWRy/BtoG24DlrZwTzQIqrWDaQOAT
fPbQcQ+IEM1rbc3HH6EaZ+l72NPmM9lIs8Qg877mj43ABjtLZGAPc/A5Y5mP+BCbOCDeY2akXaY/
9kybCSlWnNd0UrcrhOG/AS8vE5K2+xbcgCT1hOyaI6okZCQQx/gAW/bSK7CngQqucFeALFSTNPyI
prCXhjiTOZxcQUMCLXhoNV0137yiv1LkZYhovDk7nKJBcRGyNqtyTezB+HAauyh2DZ313OA5cMhJ
LnzeGTff53qa0UutHBluO5B9z9b1YWxUds3yXfcRMS2fsDuJzlbkDmUGmh60AonSgaYw1qhkrwPL
IZzo9EP3Jvlf2CW8XWcd+GFnBUjKD1Rct0J7SZuZkR9NzSFUE6CLFTxCLrWwK/5O53hM05f/RsjR
O1I/K3v43TiCkkBBvrP2oIRvlmxFen0iMFVBLf9+ef880J2Aclrw9zvBKSeM4EF/xLaVdJyyawdf
VvCrOtj/Kt9lo/43yhClKP04ynQEBe9+mw0HAYGnVmAOJkfXI/eZEkWx+L+9t8qYFoCT67uc649F
ibvQLx8GoFeTiYNdER75xvBvCfezGHqc3V2LbWKethrBblm2akAzcT1zGdn1BkGmeBmrkKaAby0k
esfIHGaw/iPCFjoCaBf/S6OdRgHvlYQMLT+mu68oCxiwithwPNRr5vv0793xkvQlohMZV+47JB/k
WKdC65Ec2Q6kKw5RGrLOLyMzLshyZk61LItrp+cusrNe0BmCHX58n3KFdkC7X6vbUAXv9Rkp3Dke
RnA5d+Om92rr7E/kegyal6PljdvAp91xprs56yQu7KRzFLkw40POpX80ExshubcpF2Lubu0u3FaJ
n4xzKg8A9mn6ppXBKfCW7OTYvBqIhpt6UHLYkqP8LynWj4l293OWRobGcw8PA6fHkPW7APM8yZQz
W+liaRyC7Kv2ECzipiQYIuN8Tl94WbAlV80cbqdz6+R/1givpZS/Z2NxtyRVO3vJTuSs6BQPTOXG
f4v1/oXnjaiyDQLCLshEJUTPqxpW3kDK/KOiuqmGXEYoacqtQcfSy3puBVK+hChNpvZDZwwgbM8j
RjwCbrl4OIMRbVzFv+7O3E85gFcRETMkM7KGC4gwnZxk2uDEIWlP+Wao1E3pKwPciceuAyZ5BqMW
aI0VokeECEcGjMyUY/LUrXbfVOBnL+9+LoBnoOWe8vLvvC8xLqJb3t+y1kZrBJNFqzDyRdYUH+L1
d1Zxf3yQbyEIRD8RBuFlDwtZnwYcwJ8Yy/jCmddbnt6vSxBGyMv+2fpbSZ16ycsgY4B0Eg0RRRa6
N/k6QNYdiAX9u8PMZk4RWgxrKZ7mfQ6RBBipSEEbiyY5KqRyy5OrrRDWvrVuSLnxMRGQapZcV6uV
v9Eg0XOrVLgSZmoBgAn931wR1Ko672oPU/8r4i+tlpA/iY6O9KxT4H5EWDLfCJe4dVji2BNMGFd2
Vi4wF+RvWAFK59AnjRlg1M4IEnwoAB1AXkauqsS2aSOTn6TmEyOnRgGNE0VCAEg84k0nQeo4bXSO
cRqJqJoobFSSLRYLa1oI6NbLZlU2XetgNQEUMXIrnzCEYugXhu4nEhXaUtfwXXM4hVx/zjewrRgZ
79xA9ZJ4tWG69Tu6/i0XI4mlWIdwOkjmoYEuDp0GKg8R3rkRgSve3w41NF/i8oJHV/lVLD7YLAgU
Ae4DdRfYZPgHrSNVfVTOHte8mWTjEaz0aZG26IgFZwdxRSTb8qDLM58KnNV9sz8Kg7ank7B+/Irc
2VJZ5Nd4R4XpM9wRlbxhYvZV/eaOgSB+plnGB007DPlMy+yvzhecf4qP62wacoyrqsIM9Ie27t4q
YpJ/YZLHjRkz3kvFS7GGcQ6CmWATBjfrAmu3NVkW9V9Xl8iHqxBRArxhLe/pig0pzrTSsKlTsLTs
y+BlvVGcCmIEcQcKtJx60aKMUFCtPcjWcIUvKTw/kI+HBD0p5kdSs/StiOhnOL1gSvmlmWtFTjfW
9+R9Sm9KL15feqGFRTXD0w4ubE2dnGEeSW7eMv+2HpVaP4i1nGxmBiC6Idigc5Y1AmvfH/pdu6jH
590F2CgaqhCG5riaGFJ3etGm9Rjbi9dWq3r7+rPCHxJzXSixN3QdithGDRk7xLRO8LSZcM6Gq0Zs
lL8bB05JvpKk/xsI0W9kOJ35pTzGdE/bwOxJ4OiW1iy9FmXs+Bzu8l6hJ7sFUYlFXrvm9RvoKC/A
cC2wzlo/WAjrjb4a41erHIRTxwDf9LduuLAtIv3OSZAZnC5g+I2l//Zl93iZ1U02+6dYAgoYp+OR
vYtNmqZiXUUqR/79SjuwpZMojU269KwRBNrnBTTKKheLMzXvKQobFWBv0YkWyB+APG9hJQWFPUl4
QHDoD9805qKzAp3/AE4+HcsT2n/tncIomeSsCgdXlTCjDhNPZh+hSZf5hL09VKR2hWpN+zAGAgaE
BC8kMlEXR6R9sH3RRQ0uY5k0l+o6hkd2Pj4CkzKVpH6W/y3PtFszpJ7tTQUtOf9iblfoAOheB1cM
CYGqCFsrQrkWuOSZ/emhCuqd1P2UtVpJel5SUJYuWP+qrQU0D4ombgawIBxojUrfoo6N0M5EYpNm
yn5otOHCjFIQ04hTgQhUsGrjUzaRGhEhC71VBa2YoarvIIn3hV8KDW3zgJpJgU4IvgJOWyrvQye8
iNNn3VwDTJXwbKQApZ8Nf8rntKOjeNJ5XQXlXC+6RxSnzIesVmFiOKqbY8+Ws2nnd9fD1aVUw/6k
hEMMJUAN0ehwiwRed9Tbolx2j7fxONSRxEQ/7aOIEBDOq6DYgjKEwGH+pDhLE6tRwvTXYmdjQUTs
zaA45M0b1FFZbqzBVWQkvi081aktqtBN/ZChkMrdoqSAH5MI4/vyXRkSUnLgH7jFdI8uS6VaGX3G
uH7ay+M3FKO/+gUHB5XuwP2/5cx8cFS8f0GHQrOKEK0xnW0NJCVurJewOzKWi1BU58mtbgw/KDE1
mKE6D04l8Z6CwiIhBMCGzWdLHEGZNwNz2llA+l6fWcvKL43cnvaOWNxIOyn+FpqsoO8bW8QNSYtl
0S5U8sbLXPGswn07CbB0TAcnAyMVX7u64C6SxFBbKee43a4UGLuT84ZeleKIyPejV9UGOaFnh8gH
KJ5i6elGZZLBa1JL2bqbUBoACwhh/NXrScXVklTLTBhMKHd7Py5GVq+nRN3Qr9q6dl/dCS3Bso0M
zux0BynknbQKOkoR/BNF0vv55vBooWe1hWMHh2bJ30lfWuGpMDeyB71YGA8TGGtzzG9AKj0fCRQ0
tyaUFCklD+0pgYZ2pw2cNcQ71mah4UD+n9DhgmrSVgzgtAEL4r3dDkLWGwtKCMQ8BIvrwfUy2PzS
BX2nDep5vLWklwnAShjCzZkpsUovhlvJaAJo2+LPkai6b6Kf0uOWZuNCcuBYEeN8l5RmYdlG9RXy
lwMDiC6XS8iaoR3gEyaJopzPlLgAqhh/KSt0egCHH2+K35fYMv5YcjECUftsTcEu8txDUAoQJajM
ovuoOLjo7DCfky0IUnTUBVU9KAnzlyglFM4cbDKywEXQiUQGV41kIwFbIDCl22/mocvaXLpwaX+6
6hiCj1w671c6I7k81EVchY0/9Qx1heX0xTBoyTpxD7xu3u17R8gW5i9ElSh1ph749XoLH3uoZ6x+
epFglKiC6mfDnxOX1n+VfabcTcuWvlYcQpYT8n9Zr5J8EuhKkj3+euHAXs0X8n5Vefr42Y34foNl
PLSup0JLuT5phd/e5XHvOZneIVL8Dlz7AH39uP3AworpBX3BduISRlwiM/2T5v7BV8VUctqNIIR6
cUvAgbph67o6AjKSKfkk3ao/lUzi6cUnSuHBejxzPz9CVfVk+YSVoG75QgvA7qKOuUKiO17HCRgN
PfczEwQUugytD0HYgduiDOcPUAE2ZpSWuZ44PvIdyJeCwG4sSTl9fCW73PqOZPx0jPP7hNat83UK
ixywpkDrF5urCdzCvPjZfMsqW8D9I2hslC6mOJwLe8oI/cQyS2gH5RQBGdqkZ29ZoScIErKtV1Bp
pd30fL+HoFKkh5PfIXSse17ZdzGc7lX/uCZlsY5r/eLeJLszPDASDtiSU9emxQzDa/+dv0nu7FlF
62dn+Zr/g1L9wjQOLz9IJDCtEmbzLfTdvcqYAZ5c4xl7Ap79nNvX/HHWDM42fDvp9xGSXwoCS7nb
9meUk4CWN653mEzV7mLRg/hfIqEAANhHdCHUVwoeGd/G9N7Plun8e4vbszuuTFTvmF0YdL3Jy3h2
nsaMVhf1/MoM5qXm8OaaWSh2XOkA6jEcLfekrZSRjqaEOWYUPL7T5Z/9P68d5dRHoT+qbIOxJqVi
VdoIZyqdQLGpgiJzFRiQ4Uu89BScyGsFKOuvw8zK9Mp0QNi0Fb7Ol2+mPvWWXE9fwX5jvLGcQBXo
ooIBAbs+K34WRDRDCE0yY6Ad2Z2XNJrQFpRugxyo2aF+PvC/XWEVGAudEgAui+YGAb+f4AjWvY0Z
7DnSz360siJzAimiGz8kYYdWtDUt+qiX8OvLko2ekQFZaRaT8tvyCcwY11PYj95mdE043NsRgVPz
O4VVv05HzPLnGPJT+59650GHzhT6UJKLzANEvTwIoOt+ajqIFunaC1h4seFc8BdkjjkwfgGuOwMv
CuO9aR5fcrhRbg8iteURihKzCLe8u+mzNyxA+zYaG+5TCWOtsIppTYP2B4lI1jQEiXaz3SJq5pW+
UGeyca+fkjgX4VOdszCIEoqiYX0vdgcsmCkTGkQZ2yVlvQMrvzwc/Oi9RPCRBJWuL65538i6hEem
iOrvuA4TTj0rLUi/FfOTKCVYvSgAnKMAVTwNDMfAlRgLicvXUI9MBcUYjzfuz2ry7GFlzCCpG4yw
yrkv8tNM0Fcq4oDkQ4ZFcUsjr9zKwZmDEDB0bqX/HjobTFVDZKg00pM2tHRU/3MC4TKHABWHhJ//
EbQyiKYP0dSeuUbgdZbbHcB0PfLDFEkIAhHJy1TX5FR7WUiv0G094LCXyHlcXc6X02K8sr/hQ7wA
VZmda+I7nz7wcFiM/hCvF/wAm2e5U9deB9qfVhCPTAap7WS7r0N3ULXxanjcaBlFm+RNfvN/ao1J
t5Fhn2xN5XY4ic5Cxnmu0UDkJjhC0im4DN5hXA5MF04tGnvE40iOxFQmlSTHnxBP5GO6qVK1EFYt
fXA59cVH5NuA7mRQZKZTpCIiQDUZUVi4yOvWbYWOTDSsr8YlU+MblcXyoY1dYs4Q41WhANLupHtp
+p3TS2J/zlJx1TNhPHqgfCXgdYNqzxkEV207Czc65lRA9qt+RRjhEydfh3flgxv1Bn5L0fl55oVw
i+56F3sCbVj0xAi6RCr1asFrkxqCh6cOLiXeX2JH/VeacsUbC++bdrZ22w+W8E3kojyv03zuG+hv
urraL3yGWG6KkBnQsFhaYJxziV1j4hjSzKPk5dPnEt54ySLmKXWPiGxDQw1zHB3quIHDtKM9A9s5
vTRt3Dn+Ysqtwi+3O07rg82Wt7D/LlAx/u4cxAl2pZqU9MQibsGuubZTS1j19US2gGsgX85o9Jhl
HCE5jVGazXS/IPjCjEc9MeOh6tqcC7ELF3CwEa3CCzM+PPH+TSWmjVg2TCa3TTXp/lSAKWUXm2oS
u3TH+dcVTC+P9fkLxMt/Vq9xvVCdEkPZ8Xf7lVBHw3Ens53bWwzUKmwQnPC4Vw8S+gXuA+SH4EgR
Q4zlJTFPqJLtfutsVWH8wQPgRXPFpsZyZHkSidWbjZ4ivEpqQOLBAYZQSVi01wmmiNqd+FPabkhh
GiEo0Yi+MwvBuAMcGqQvj1JQDHWGFKdqIYzsE7yadaWp6vEeArJtSnzuEZPxxf7eO9NprSFy1tLa
39s2lCNTvd2f9tdFGAsvbj9blJeGMXmLmxZYxVooDjFyrHBGOFxjwTYbp2Eyo5bp9dIHFC+w+7Vy
fUvnlk+qBB3AvGPg68G4w0L+71deVBj26og0GqAwgic0ugyKhOB6Dub5mDBsecwrM2WPdXdjroQZ
4om6HSrp4mnFjvhECFai0LQWkVarJTVLFs5RdHHymjoCDSo4aAwpK9E3vzrk03/nUnFcMeeL/B6/
yiZlgRu31L6oELCqllfAsiK4uo/kso8xVl1nt8jAkHRxuYayPr11kYdmQqoQt5W6ZTv2ZB1DwLLH
ki5bWpgr5/puWeEOcMVhBK4T9e9c4SQ96ZT/EE7IDpQEBRQr/RxiZJ/3n6Xp04vjS0DpousTGJdu
y6PLyI4lDf6ksATlwGEGXpUTuIbc+Y5i8zeD9/0hTE5l0sHV/LWgv1s0d09Y/ppyuVgEYbUDc1HA
UWy+KthgD69hdsEO0qzIaVWegCmx4/Y7g5NgcgFzUpu6Yn74SQ2DoM3IpRixrKHTuXgx+i5iF3GB
lwEWF21lFdEO/ET5wxmt3PmrsunsoHVzt6pHy07ddZbMx+2/Za98HdF+qwt142s82acmuBgiHq2y
Fq2OXZFO4exNNlfn5ND+EoHwdOrcjqylBwBwec+bMfSI/S4KsaXU+mbijr9L/osjSN2OmY6jPgyM
2AVzkmTgiXF9GgKyaamndOyuAQGYDIoAKybWU9fLMRXZ9Q0WnZyXxHa48NMZlaajFx3P07nQ3BnW
jdRditzynmw/3XZth5n884Ur9sLbpA6obe6adgmwRhzOHoYqQZUSTmHZblz4IvFnb0nZZK/jO2kl
54UdOqOC+PYKzvDHE8jEGT4D+X7NciPiuxYRpMMmAOXuw1OMitmhBM9Pv2gXdpq5gvwdGZx4o8xN
ZuxzM0qrEWbn+1ustqJyyelwiA5DwjT25xXPFjkZVsrpFHwPDFWMbF2Bm9FsNJLJFV/M54kH1olg
5pIczXV6Rh4KRREbhB83DsIt0GGp7ua7AU2ma1mHYw+OwW1RIiVSfEBQdEIN/Y7lBSaqjePcDrjm
RZ1zje1MpL/dRgrOJxmJlpeFItaQ2ubp+wGV+gZM1lOmtF13elfsfERtCaYSCbRRmLVw6XF7XXnJ
z1yjNbxa+NZOPTpP3eAbV/g0SOQhka68EDJSt1ITWenvvkfp1F17KgIZLFb4pm1oAbov2wK/DW9g
ZgFIN9PtCUOQJgcnmXuTyxIssPUsZl4kr7t8eVEXbCt5h4Rte8FquzTO5y6z0FUOp3wp/nTb23sU
bRFajNLlE0RzKJ1gwG2H0CFDRzMd2HtZjZvEs/nRKhmmZPFkRx5Z5qgRRuTjabUru5vRBCiuaI3s
4z7r8TN+1xPeqs6e6BM4tV2ym7dzPTw7XsN5XWiTxltHqpByKw/r7W2H8Bvzd/nhALLaHrEWCh87
Xsq9FTq0a6r5lT+NG01X0Anbv3oUfwJ6iCT3GbMszWsXJKiLf15w3C6+IXF6l8Dq4RUJvNIQXM8w
ubZQ2gkLOrOifULPvp8rDjCSw/2NEyYa1DCih/h4ZeR2wcG8D74WBdIx04agdVrmzcwkZth1FCLQ
guBMqxaVp/OTbypksOTDAmBSQLZc8lt5tp4Ka3BOgPSydA5ozkrMhC9dScgxdZzKJv7x2oegjbZu
sr/vbtRgmSYTnUnekzMn+hxxTPpI8l1bK7jVIci/l0Pc6kQiWSfrJjBYm9+2bfRzvMNqxdIw2hxo
JFVEKPzQRRP5gFK+p/kSp1kuMEKU/wPBQEfeWpgqoiFMa8RkniWqkZnv11z3pUKsHCPehbBDiWeD
y7cP8aSM4w0nxT5Wy97AUq/N53ruQ1cypiPp2IIZ/dyJU34k5yZRGErY73YSdF7BQbiKZRn2/GUQ
W/hqFASjGRtkgBHUKc/3InIoWq36TIE2PKPXc20KfQXC1L1UsgIf3+te51w5lIrHlwARwFW98BWo
odPO77hshlyaykjfydvf94wvcd5QCn85RvG93bXMIRcyfO9jVdHvnC1M7rADkYdk+jeYVU98TRoQ
v3FKlAjYid6CJZ+VZI+cMaXDcD6rfGr3k4O27B4H+0cJl/i4AzybM4DmLnEUH9/6QvggPjl0Bj3n
9VlfDo5ukU9ieqw87ZXGEYcQ3SbFq2qpAru/MT7hcr252fvHGDa14XEppMv7aVFkbgK6E+2T5iwU
uTAmRYu8DGTl93BADw9j8YEhcsz7nGiszPtf4o6CYxkP3zN+VfzGMSyz960SzI7r7XdU5OUbW3d6
nYnexA//dR/OczZgSh7bSRQB++TXP0MdGiZoMI8G5NRzDmjeNfdu6eMfsqW67pf4Bd7jXIRZ/QKh
PgDM52VzPaJkUXLYL5pqJQX+rBNd0LJQnkHDmLMZrOZIku2+wILbdkoAIJlLPBk7utd3aQjtWD6D
AmMrpvrWiNdOsf84ajW/ERkOKMzlmwpVDk/hKQBvx5IELngk85ssdl4KBtSVv2p+Yx6zCGBkhV3W
rO3+pmm98Ac6ybVuaGtiwpr9lv1fgvX9bjYo7OM2NpzoEBc/NxrBfKRefwiG8dDse7kpqSPWXJr7
ffMwM3TNBOTx+dPvDA9vDBsOqikF7Fqoje0tH81/0QJ6MsfPxtconOFuxtYvmhDApUPqptmuEvKl
YKXph5MV/cTZt1LDTGUgEbSuQ8+adRlTmcPTqMpaVodxgQi1vHFk29UaZi8Uv07NyP+Vniz03iUz
GjfMacvbGkm16Osat6jTAGlk/Lxb8Ge3pOrwoGBN/PUsHTkh5uXhWxnDFoABGyQXKVbp8sbm/bLN
Ahd8/Fi3Bab/WHiJAt3jyqYBtiho43ojgS4rn88zZR9fhKTiRHrbog9LlzqiDTP+my4EwibnxtW2
ABIfOVT+ayo4lLu3NY/qbtRBwJXK8i6kj9+cNTo2LDg+jQH7LgBrd0uZrzoj0v/Xo4fU/1gAXf9b
drgaImlL7Z1gb4Wffc/XML00SKOopwz2vyLNnxdt1aXigdZ4zWRVenGwvjQs01PkFVLSQylP915p
2eJMjf7EdVnYug5EAtQhkf4eUx9DpcMZqGC4lrC8LkS1kfMOvsZ5l2VVktTf4YM6QPFREJ8+qI1g
l7UZmUh171qokJKhQu5fNEQYuVIrB1ZkJ2cC/kox0/opi149IP4ywldB90minnGHXLhqiJfIfTaO
xs+D3Gq70olTV6n01reYdrpW/C3JsLYNRZyUg4jsqTpik/NNPt5EZM4vYWtv7sHOEAhcBg/G4uG9
qbQWF3HkLfEGwMilp8DbCLGTMd5Vcs26j9Rlxh1bmIAVtjCPODHS9+BDDzre8xQwpw6WmuWKAnlu
ANdBdonuNruv3pO4oz70RuJWPPyuIVbN5G9PRkQhtcH5zRURRVvJiGtyKpGCn7EmjdYIal4y2uMf
u+oK/1QaOrzmtwhbXuP2R46C9yXhLckYPeINsKJoXwnNm4oEsdsCopRnd0amoGSb1+1DuTCqD3nS
YTnZ+zOmUvDVOSASNs3zZZkodjlAP7VX2DYzHkFQF29KD7Ol5ScYLFmMERsNInkTUg5a/wjmlYO0
Cs27NW7dmb3wvsGf3z6q/8k2Jui/iGTjKXatsORuQoqmXPK7QKuh/hOIcRL2/8P+VYCOWiAnTOtc
IF/rmnbD/A/QrHKpwqqSjLvUaFbI5WLwQlLts/GhFU3G3uC70OeW4pA8DcTxwPpExIJIzW7rWEMy
hJuLE4/wyn6sFbXPnSb4Ss1FbEGMF0c24VjnmXMRleHxcrZvz5D1vYDNv8vMchbHIvKBwZIjXcct
dr8zSR3LENphN/LpW/2AulgSvJRX9+jG/BPy+IsWe3tu7te4eLfJhbi526C0guVXNb/7xkA/Ex3d
LHpU8q7ccBO/OZ6CZcHQb2qvHrjqv2WItrtzX+EJZ8W/2eH4TWIE9bSm8u4Q/FHP0c+qfw1QlPWX
QY5qobMMRn4s2LyBGaooGTQvJ++8TVgPEH9q02ObJ/yUlAo2J09sqM3iO82zetC0WaPyY9IdW5/7
6/5j5/iO8R7tmH8ukj2geIEJR/U0QWrdlgBqQPyZvyA6reZWoIkLSF2fgLlZkk8iJf8EyXwjOy5V
zBuzVYNdUhj2AqzclXwq3QY9cPeJHmdSY1iY+7NoUrMBmat7cs3tkFrbN0LK1S7NpSLqwgpR76x4
qEOYM81fs5DXbux0PrefSssKrpsBJhmn/h/zfXcdD+Y0EwrhkYnUWJ7RsxMkqAXTTcsVugJWkRaJ
J0koBJtfA1jzcW5r4TOQIty0BJW0ZIi2gf7+1ZhOFaDxrTkOVU0x09xGgIX6qVBWGNMe12JNnmqb
550NpLd7HMLCfhcv6CtgCSP3XmgpSzLVYB7PqelqxfTd/njPlM768wNKfxNZPunJDVV+BmyuO5dL
QluW8kEGdHno4YwKcIwLwSI+z/3TLWPSdJYA+pnc8L/x1QyxZRn/q0fRLoD5GM25XEdIwPqlJP2q
c2d2PIai4q3HgdCuNlz/rmH1qAMDHcSVpzq13XLHUqmj8zWrNbCfo2UwYSGcl+PAj++XKQi1lUl3
rvuTwcfS3yqWRpeyKZ+XqUTpJm7UoF2SF7kYJCdBL5IHJPxGjILvDMqIkXLjUYqDjdFRuGgqGNs3
InNyURxvXHsjP7LVZAz5ke2BwlhwJwJ3vGRiVxyIaNhBjxDYlQP8JQq9CTzMVfCEKXAMaPJ6m4Sm
5Vt2xwa2mtjg2T7JUfZl/rpslB/e8+LzAXD6KmO1QkqWjNOG97YwhwQ1MB5C5LAcHV5BqSgdig7B
qDPKkyp0KAaAmpGySONYHMdnZb2YvYg7jteHryx/ymlRLxqb7GfJkowX3xtypnlFrfKLEwftfnjk
OtldRsJVGRU9XIG/ilQ2shBZNwXdwOug7OiwQwb9TpJI1xTfCxbteYsLbdXrbArnDrX4T6J/Qdq7
YUcugwrvteNNGfbEvfaywwkX/9Uf7eXuwyUv96BMix0hzsTihE2bwzMAfhwQ0nfHdBoN30YGNzaR
O8R36g7UfCr9xADxl3TPe92FccomWoLH548idayu1XQioElolhGogLl5G19GYj5GC0jMQvS+drN/
wm3tS1Jm9u1ue3zYbYvEv0DGYnZNBST8fjMRYi9hR9Pv3OgEgrn4LLh5zaJicZUUuR2QFR/VioOC
d6+79QA1sEyB1AHwiHO7IBG6iy3TzJmZYjrJ0US28HYQF7SqZkWvP9pXrbjTrXFtCAfHTUdaxI/N
Mn6ask4FQMkx65f5DuE9XLtUcd4m6QD2cINg5Y/jkC9IdMO68tqwJJyWnxssRX1dNMIDZj/93aKN
7AA6GvodUlLIVux2cLasImB7dgO1ubKXTwGRsXjhH9W/JCMv575qvJUBlv7Kuazs+GYtTg+3W7tf
BUuY0FzKhlFQkD8jnlEz20CNyxCYvI5S07q4Pzpk9dV16VI5vymKnIHxxm2eF6N4czLRJ799gtIH
tEcYfDa0vn6X1a2LKn4hpzQXUguZu5jVJcSsgT+ZoqvI5P+0qUpqDH/o8sGojptcAzDFYhxH/zJN
803DljQ59GUvUzqVd5F2inBGNrALSH910wdQ2MVUZhedue/pz8QLDWMpUNbP+JkP6iSidfVKJRyR
zao7q+3dGPnO8DHiCvHvWlJpdBuapw6GGw/5cX+9C8TUHXk4JCJfOB4OeoRGjAnLyszdYmuwz1OX
UvL6/VTE3ANZfwAKc0JPC07QFkG+S4afPxoLv6AohSGLOuRIwYp6roLy3f6B0P668D6YYeqQoWoz
rvxWxny7rfX+imHTd9sicZE3sZvj+GX+iTWL3GERuFJdYWUAf6xTRriUFXXG3Kw7QoQPCq6rpAOd
6RZN1LkhSmEzbNjF14DYzxto3Y/HplD7wNj6mezAhVma02KfJSMEvwYvPVfw67joOBqHe2zLWEL7
IIlmHGDjglPihTP8e3UMwriJE03YRyesg+NVLdGzA20hEK5SjkCRrICsId8boF72lnXM9cbSMQns
SQlrXpMl1HI/ya2I0nwdLjLoA2aPC1j69sofB+ZnE6W7OCBm2+h6B6E+6Kcfv1xSJClsniC+X2bT
OZ7MHFzwsMmVo7t+1Pz2DSrmljQ5TJohMub4mtb5WCmHHZaMRvVfg4t852K6mx67bm0VtbOiO20b
QDolBnUDL5gKjROx7uOxNG5mZ2IPdXYikwKTwBCWL3ertsA5MvAr+NKzR+P0pBZpcwgnV6+9Qqaq
F+wrFQmes6pc1q1DAuy+DW3uyWWVlV976ziLQsbvkWEpw0EoNBCfHgHDcbMCE8ylmCIyA8Wh7BnC
/oXs2HrzFNceGcIdlPYDG89OXEUGyGYH8UfnqLaGMM6zWOzjeC6yQoZNIjqVfs0xGsonsueXyiR8
W2HiUkN9jH/oHI9GU6iNfWiS+WLye3wnHknjWOMRdtO47EklT06QVhgI1U9T/b5cdi2Pr9uVKGdg
hJZB7j2KXO7qtbQ97BM27mYEiJ5gRImBgzgozOXeamfs8IHv8Nrkw3DH/Kmo67vaBJGu5PrbEVxL
7oyWlN9azXl3JXQHh7Iht6RLbukkN93j8iyixOwiazjuvBep9rDsC+CyLailc5bKql12BG+5DdZ5
AALrLwO8Z06tzzfxTLbZEHarb8bUIKkMphKlgvO7JMLpv7rIAe7UO1jEcRL8Fi4wM4EZcUFNSCKN
jECe619ZD9/npg6FAGlMYVylFCVPrJOF9wpH4ODnd0Y3w+0PwMeqRZf3XvpseyDGutNGrk/09W7Q
G31zDyEBUXlzlYqdH5ps3LeCvgq8vIIFCP1S95ehvWuEWaK5EXhOd8VS3zr/SN6Qv0OEfUZ8JT2M
+eFhHK/G4lzrEd8KO63yZXRRxIqdx6MwHEk1ciJKePnXSFntiw9rFOynnkltkzSTALRd6mnyiF8Z
OEHymx4M1B6Dvu8vaLTPOLrcomG+kea2LFoHYycmOk5U4gTQ1Hw+IFB7bkiL4JNqW9qdoX4w25PS
hWeLRCylXt0DRbpkIJM2PvuZ5fRvGnkVU5VY4S8B1+xChVVCsBWd8A0SH0XqJNmWDbfXTY4Rfjl0
vR14JTV+BGlIiQNBodFA0k7GfzgY99J6HdnxabaPGF/2UArPp2yKIlCd2JMDXhIE6xqKPWg5hU6J
7OB333jzdSJUeQ5g8e8aEoNMqOdQ4fbYjNt6lDbPo54DGmg2/n07GdXdP9to1JE/Q7c8f1jZBiUk
nYV7S8utT7N6qkbZr2KbrULLavhDvIx6LRoDbGrSHXesf026+QXzeN+6JuVpFWlfB6a7UhLDO8FI
5vONgqAknTvp8AX/2NCvxy2eQfJQHIfXUL8j/71CHZWNakKUC2GdMSyOWIi47LbyYuHNyy0b66nr
hE13egDY8PtS1to9T8GmXZmOspFrOMIqygjNOIq+cbPXq/2cEgWiD3vMUCPSMx9WScxYYK19JFtz
lg1K16dRZdKX7MxFcEO723Hb4cRCKxIjskmd+5ocvxCoKM2HkgywpJiRBcVd1WSbSfYBQK54VxFD
gwknEvA//luRB2WFrgueKg0sBVs5sF0251HNhViE4/pNYTgxwqZcwerMTSi0KtTi1VxwswrdZGs0
siT8L4Ar4x2NPhR7gkYOM6W802wAT0k+yt3aiZiOxmDy09VZa1Am02lKo/ip5ePNbNt4gHtzYpYz
V44IRvmEw/AkBSJ/XJwkHUZLDWYyIki0IasRisUZGnRR3fwwXOkdrbsAl10h709YIEiXS6ldXADN
iIRLHkS+Mv6BnSxAc5RmmD+fHsB3wAQevyl0x/LW0VpcAOcG/iGDEW+lYF8rCMlc7Gs3NjC9Fz3c
VgPQIeAEOmaWtJf81cU2PEY6TInH5XJekBRO7D5H6Zn9N1PMwx66B+VOgAzVdmocZh3WjWH8yc4I
whOcf4vTEX4Dx0KOwyCXNgCkZS/apkNcBqsHA+J4VNClPoonXC1BJ2ZYP9hPgZZfPQlY9BScIbpt
kD248yARQCSqBzaA8bCz/Uu9M+56U8I5Ek3Ic32DfO8FOFf7UNgsoOFzQ4KzltNRbkZfYiLODQQv
/Dw1W5YcdqUiKF37uUApnb4w4bsdjg+qcZ4ZYvidSNtbjPRRrPGmpV4NF7KTANFvKcPY9SQHtgyP
/9B0HUS+MqTxoXCMCo+hEEMIvTt9C/kwxilzHC94Jkr8HM7KLI36kFmLS2j1xuDJLnsgizPMgnEy
qHZgjj+Q/gLKJ9emhys9nLxjNzX1oh8HYSoImGoWy7nfyxNcwWTk2krpNJ8H1bNRNLgpxmZUwyGa
V/aYGrHYIX6vbVOuzh6hQwZqIAdhRmJDD1El/dX+H9WlrAcLEj/exPQwkqfeJVxR9QHHbS1HgjLN
ZUGH2xAfi6c3FQdlZAu3J3uEKb5gnNxr4frrSvxlJ6ArT7kAH4EqD/oDb/5UlVe74yJUFQpavoHL
cbyhy+yrMLmXpIN5Nrtq4G0+CpJPaNGMQEOxcIg0oFoWI4aE091n+dQ01uKvPhz911zEO0J1L5+c
pgXfDbo0SsutZSKRcsxwliQSS2xibHs2AfkSIi+ujLH8TW999fVSuheBC7Ny1XZydZOfoGCgM/cR
1RO9X7vQUR8JuSu4mDbbu6ZjL7xypEEzw8lvk36kJ8GmZl6hNqJMNCDhnNa3GwWmo3hfGtO7e3MH
dqEFOiuOjCj0Vb1/L4N0JIGeRvcVLK88OhqGC3uuqKK9tKr1lBjDglq0I313x7+CicrmqkZi5U0V
gsVFsFlLGIE3H2ZaNDei/CKcUrqHPYtbpWEmVBfpQoeUy9g4lRAIaRNYOjcjywkxL4Wi/YziqgCL
bIwaiECo02LTuKqPD7Q078qN2Ci71WEoOLk8oCvOBjAx7jNoZMljmqWjal/f1oQY8C5vBQfmEb7Z
WaWy2JAqEt4giz53RdJimA8Ak/JRFPy62VubPJEF2SjBisFt7RsJ/kaAElD3QbArMQoJgHvlaEp3
ygNZdGifHP5rvvzPpCKvSDjSPasoMSpko8FKwC6aJ3D2nxvjkeQrm4fnlPqqzKdGu/I1sYGrSBXj
jNZv2LTvVZY0GKrFI8wS5R+6syH6V0rxH9IXfbTsiDdsK8TRvR4Fkf5kBHRL5jUjy4YpzWgwv+xv
cdo2cc0DEZW65iQmzsZB7V0X/JP/2zkqjPgAn/m6GMqMTSKt8SMqd35yoTqcZFB9+FJ8XmkChx9W
3bVtmz2KPG/30ASkMo5TQDkZfepBalQ20RNHLCRZSWVFTyqhAGQJCvolFLmjJdaxcc9SeUR6mRUP
eEcYLSR5hcgepMqdgObGtIgYL8qreSTuLHBCaQwCyxal2zQNjc9O0QPckTHj0GWLazilb1501vug
NG38pp/Sys+l/bgB6iPXlWxPm1C0nz5vshGGLWhHZeC5gyGtVaYoVWqYq036Az9IEqTCm9NHBmdm
H8pajy9AkXvp5ZKHw0bAueSuIsrFwG8rjvDr+uWTLW06+bVJipsxN/AaKeLZtN7Yy4kUtl0qPPhH
N4dFgzDtH95NKRh073QtdeGdrO3BH54emJwkiUgt8ciXFNgeVeetN7hjczg0BPL4HxXezB94CmoX
9phzElt7PsGXPun7pjK7xANtZZaeYZEZqOsxIs5qH3lZfqCeO7zKNrlIpp+3l98uLFRP3VxU0I86
cDShMiRbOlZHKGApPdAGNb/HeW5gHw5vB2/OKh5yZ+pDCrEu/XDMzqYf2CofSGhK/Kn0kVLldaIk
Vf9N0v1AOP01yXjArcP5N1xoTDM4r6zfM6P+hMwgZkd1Yz1HRC80Dbf3DmsXCHrMq4b9Nf3Qdshf
B3jXDaoDxEifX4acdytQKehpOWJsJiQ8KkJYu1G2MP7dtuRX1YrYEoXXoVtck2VNeOcxZLsB5qda
xUk/pJkSVjOs1YJPfPaesY/5Ge8TAjc4UlOKLJJRfCNQNWlZi/Lb99c6ffYLRSncjSrPWTVsrR6l
F4KBisY+Avp6phVer1en9/wZ8zKGsmfqAIz7SJqsPZdj+7uxSX+ZivByiJ/BQ9++wEK8Pv3mo4Pr
Tko42CkDdBb5/XJyjHqwdywdkJ3wj/OQNTs3vAMX8OkarIEk5wnZXVfhTGQEJYdxyIYGdbR6+XDB
j16sSaJ823TAB9Bv80siXXYOLCCIDpCCNam8ayTlx4CHRtnncplUG/Nz0HhP+fiK9VZaA67+5wf0
Mro1P9OgZpzgNbo7ecOxyKh/K05lfDbXkCYTW347NT0ynFDde75r4JFzsZzKMyD5b1Fehmky6FjH
miW8+6awlVmfU2YqDd+fA1y7TCn8rqodwAYJmdHNfV9a12IE2l68knyR9Jwns1SXqbOYsHI5xIud
3g5qeiNMNy7b1K5oVtm4tkcKHxKofvxJFWUmRh340vXiSVPcijsr8PePAAp4SpnOp8GlkxlrvUhE
TdNJlGSZd1Z1GQBVwbVI6iRw15o9mN+0xlbYKuoYQwBrhO5IF41CLL5I3FDQswHLleffWoAEIDO4
ItOHAToFPpY8skMpLI163olJdeIaElWNyS0CM7DW8/EzxBIpt0R121C6Af72y2Z0AKpXVpJarm42
gYroZPKZF5a8rmbn3UIVzddpQOEYDZavE0Rpl5eU2uf68m4ECaOvnilsGiRZy3nMQdM89U5YNsnw
hdtG1TpPFsWi1Lq521tBFSnF6IfaHm+BmVHJg+r73uJw6MT1sFKR04ilE+iOZj+/iAyJnL7SDApQ
GsgO7Ue5+p3zag4HHf9O0IiRMzKcOtPmWATV2pZY9Wo3lJVe4g35GD+usGgDQf8VzLpgLhm12pNo
Vg6QYmWFUxbDiMHPGxBRgDyWh6fDgR2m/24FB8+fefN48npBFv6qexa/RwpJoZX/yVkoWYV06Qci
Cdp8iV6dbehUFYl2JLBwLa14WVQhF6S1o4BK3Aow9a/ARMXc3Mukwl5nXf5oZAc3Wrjm3baFhS8a
cUc+g92onZFRspRJKJYRpi5500uTKOCFOczCHVWrbfG1jx6Sz+VWcwixMhI9hIJP42oN3T6PnbuG
HrnYj6pJZ1Z80/PSrrvn9+noH7sfFeHmLeiE63Ik8a0f/zwP+qv9zbgw3enRTj30TpP++GM0BRrx
TMs8gRSGXjNDXFHJvH7UCYpyusavMgmVuAa8hZRA1/pcsOvtJ7PN47W9lNGvzEvgNiVw03SRXBaR
cgfhP39cCrnFp9DkzD4iHkW4dcFpUWtraGsYLRaP+LZIy+32Fpuz96HsTMvLgo08Oth2j+8Fth/q
5qBWKUY/do4D9RktlioAVOdY+13EgpW50limWj2V3+GP10cHobisoOyvFjDj8T1ODatY2/XVCb2M
S6NW9V2IcC+mE7L7RwcRjeGM4Eyp05Gca0+A7KZ21u/C/hP+rA83EiF2c2cJLPVgE2AxuZ5hFM/j
Niaajtl01m9BBx5ZgQW4exEiAwzJQnP99cwPYO2yy5uZsn9KA6iJm9oMcu4CSUK7gcx5tDWJ2JsQ
ZJcKmw4005PFAkDdqCaHkdB6Pwx6jI8Ek7lmY4bJgR4PApMgY3WT8WLXMgFroiDh5+r9Cmrm05hH
sBBXdtTDCFNzN9jGIHbFT6H8o8xxyDV4TKTN6csBrG9IYFSJlZZJ5VMMiLwHlxFqtL+YHZjVBJzS
/fp4fqaFFSreFL+ruxPwUqlkPhn2kvcvf0TmB1AKX+/qJ8O+V18tpsC7MXfZKjWxG0rhWAUogKRC
dDGgQx8smi2lJuF+duksNbFakNMMfGaA5tO8lTRfpKi83c9vJpl+aj8xgcjmfbScCDy+YzUtCvb5
wxeyMoedgBPKogxC1DYzoqkrUopdqM1wpTJddG1MSgJCFC4JqmiH7RBG+F9QCVH/y5/g7eouWNBg
wn9sIKlhVJJ9AOBnn5I3pBEoxoiSsOo0w45znKweJ94rUOzxo9XivRdvQvIaJLgj7zC/kgFQ2D0Z
fomtY9zbtZfg0KPNzRWG20b5Y9gKmSXhxzkfnDkFR5jEnjLcaoR8g+XZn1DDjRwaZ1x6pSm/GU34
jl73sLvi8piPC5TwT7y+22RNl0J4rZXc4esZ64/WqHKfIbBo7suDZ+7ikslIlRj/OFXTAZGDyJMU
PbL5HwlBNmuBJbIkDrGM3ei/4wxOC+jXUomFEjWrjiIBOSmhGIuR9z43APSIigIWY7BIRDiVWM5X
sc4fTWisH1Jf23BWm9SQ5zDmWJJqNNebuNgfR0+ZmZaoZyxHmuuN2HWhwaa81fUDYjxV74bcuVJU
udep5e2LDGLdb9+hHoh/fHLPhQwohBx5aOw7OansZyoqM91JbOfyEqwDo34/luau/XoWkgLhKilk
aFZ3TrOANGPVLvDqlsJUp5PP8+TRLU1KgLZyQUxVHvo6glg+ENtNpkeOO7qEh0x4PYtbo5ny1u7M
MX2gY3BsMVIFwj51TYbPOtBwm4FrI97B3pXz77VAM7IsLvMlPFOIDlMJSWnaaVYxQ+Uz4BfwbbNd
bxxiPXToEfuV0ScmZOO3QOgp1hH0I7wFgnLM8CJHZM7/+s04OmlyyhjsNIJg8qtRVNHPFIU+ukdM
sGZRLrBCgEHPi4nfZ1GN+fL7WyJ/DxAElCeCYrQyVSAK+BCSxVn+mADy/CilN87cauf95mveitbK
QOFRQZ0yybLUrbhwYSFklkHbqiZBYyFOuHVP17svhAxpEU4zVQ+hOObq3N2rVW2N3hw+PbVc8y2+
oavgX3isxfJWl0c0OYeT8uNue6ryJhHqfMRlHRGt8W0Fd96e8SPilmMroglHzM180gmRgol5TEWP
31uDd2j8RPCEC3oscawYUQlH5OMKEIltXgNESgaMnTzRgTDj5H5l6JQHj0m83ml8HdP+LjUkGAJO
aISm0xfx+EvnL6jUUEguvCghw5mCntFjnpPYbGhhfaCshTqY47abenOHk4yIF/fOkkM0mSW0bXIx
stvBeqqnGHcKBZTxWzANoGed5EMmYs7crz6QMl/nK7ZbQZOWdGSWpPyyJhpMaV7STFBbQfSpzY2j
QRycy3MgUwNKGzTrU9Jfg39buA4hA0Hyj7xXxAuwzU5rI4sIGXmWd2HBniklmEBNDgOKYnObJf/A
dzhd0qUhpivYWHWoPeN8yVv1jAY76tQWTbOjeentVUwmt8WJyAJVhyOOF4ogBwYFQ6v9XE1vqCAW
LdB8cC/TZTX86wa/p+Ct4BCOrdqGqej1XiriYYRTvjlxy0OvmCcLfcdUCJ153YpvXXr3UnGLYCrB
LxFrHolgyXZqVT5Apnacyb9MCcTOVcHYTMHn4/sHXMfVzyYDkHKZUExm2zNBKkcBcBKjZ41ZhDai
COGbHvYEaoye+EbJdNbRIyqDSNfV5VH2B4swBoUvO0EnT4pD4aJACXZEKLNoF1gDNVBlBx++YMiF
U5R80XtfFDfk8Xxyhf76p1e+ywlmb4U3LwO/nLijucVPtQoSXMJFkVPa8jwDTPnoj5qd/5sMY822
DYzFsMaN8pss9inqm8MP5tEnP2U7FF5iKmNbhQU43hwQsazAcHKzAp/wV9g9T3zJkWc9at78fux3
TlyWjzlwVt1+Uz5Tt751JmSVIbz0wG0DNoYMejGH1C+Kud01DD4JPV5Vp/ZLPsPfssM3TCZew9E1
RqxI5rTBFOwclkhGK0Z76d8hNcUF19Pbey3iVqdDKseqUVRcoSD3GFM5+ookBs1/LDPTZe0Tc4aF
yyN8qYIYMX/JX4z0zAPYort/s2nSIlZf4I0mF5YiPHstKp7Mo1VoWHj6GgPECAKNP+/GaD0bH5Vu
507EOD+Xv98T+KfmAyib1qjp9Mgggn3ZP7KZelBx37B3xMsLT7azPYhejOc5aJxomRmWh2Ipgv49
Yd8yu2SFELOZIrLN4Yu/S9peFA/lCClKm5KjK1cBhyiiHnZXhBIR9y2lBfbs2LcrI83g9BB3jNeS
4yXqRWy4yTcB39C9MJ6cbCRoy62QKAYBAA326vu8bXF3wTQ6tnIYubXVcwp/UG55nCS2yKiPGrsb
XcilPKLaMzrFAwwhR0e4S70weft2f1Zz6g7cevLz3YTk+JgoD5hnOP+qy8CNp/HBa3IuXUz9fckg
1bP92ETMUyu/MuCHLexqkCxV9xqdRJU82dZ60QXiM5JWEY6UcYxVgANqfAGNKdwpCB4Z7jfz1tyi
foAjdTFMZIsK3ZrTO2yK5pibvEgVYqCFzEz5TuyJ2PaLsH05aRHkBoPio9rbp4fUYed0GDFjtPWD
E4u5U5kJNo5Hvv1IwHqUe2sfEuiij5AOwifxoVvLY4bWOl8SwbBz/qoaxRBkjgHfune5g4cAXtF0
nwfzku9zfhnRXoThfQ+Dr95Crm/uHgE6ZSFkQQdsZ347LzJG/kf9kE4MybOugZGHrZzW4uXHzsOp
UUkqz4tCx/2KNjGbjdVfoWiCGPDB9LnjLFtjmGV1pQ1TPYY6TopYg7Q09iBWCFHaVl+CDNgauIao
8E9wg0YiaewH6hblqhxh5/191BWb+9V1Vvkqq9kcPcu6FhcIgNS13hPH0FpUB4ec12aI2moUmKz0
J/tHBNR6LGPt0Ja/MiXzEPgvNA6c+jXCc1oJOqrwDcDwgYNLORrbuEOLxsumWy5Nf+GhmzOg6XEA
U2q2BTdzw9Bnmtrs19clob6KL+YXXSWzfK5OgEc9dWLQmlNt3n024YRKO6o6uGRaWpUV5F5fEYdP
SppAMHaoOJ2yr/2CmD55IK/ajdBw7wzZZfXf6Cf/BTWuLqEQ5C05aeK1q/61YR64Im5XbJtWfNVV
Bk8vjPlSZT00zonLCvKBTdFU8+Khd1bG6KbOmi1ZRwDMENEB09xnQ5SKQ6niunv4PwzUqFCv/Kk/
bmO5NM0DbAKhQZcG6A6benE1CGWEusjR2bB3FmLZ/7B9ueTFoidpUo3HQq8nwo4eQgFwkYHghAcJ
Osn7+HuJ4YZ6lpcJaBoUK4oXrifMJo1p67k7D71X35im9fXu5uEL8cjlhFiwtljQesyToPyVBugq
kcg5rHys4a1QMVyZ2aEo2z4/jSNOJNpS0YaG9OBCl1K0peYbbb/DlPYvoP4msMpXyiiFLIa6z+6u
fpiKsFaTrZCyG2NIxtlDyfWhu6+ofc7CsZCg2zoDYGIeOli7xDevnf4G7o+59PtjCdabgMp9Q45z
mXgByPpkvjtUtZl9u+kQBHYQrxT9mQUE/Vk5yFc8y7jUvNjCuknhmQazn704FnIsuaH+hnYusdHw
J1orOPAJgTcIFOS0GDOm1dtEnwwiGFdiiqV/4VAQdVhP1UHnOiODS2dsApFEGISYI18WlKqI4lC6
MCCy64rFYh7RnB9AeiKpOQaJ67xpiu3yQYEjstbtf+JMz/wYExaeQQVJi4XUVnMljQD6GYBf/5NU
KduGyQf1ob0M5d/0H7mfKYEx3B+fxk0bbrTDvSwGUjHWe7wquxcPr1fCQcfn2bAD6ni51jV9IoAC
xiCba7jDi0zg22++6CT4cLEXxh8AaFlBLT+vcCkDjNO2BDlOOOgcDP/76g/70JWB33+ENMwlnen4
1bBu5b7pWY60nPTkgyo/GLQoMr4AMvU337OdD0oGkO/U/T/lwFQzeQ9FVgtRm0eBco8SRf3uGqCZ
UFxMNp1ZGNdQXPA6JzCUHVj+B/J8iS5FHtpvCdP828ug5wyXCv9uGqsEWuUaCtkYPwcLYuSThZYo
MrYSm0m2yAlpdDNYjFjJHPjTPrcwcWptN33bZ+2ciV33tb1Dt1xzZBbacwBDC7xsgTsTYV1Pf+Xw
TmXAAOO7fsbwWias8hqNhUYOHHkRSMdTrIvGjBcyq6ZeGyERKbltRskH8mIojIjmyc2MjSQC/RZ+
ZpChT2dkJfDixBVEzpS51HEbVH/Yuf21DfCPaWm0PpWbxcO0fsqeN/pP8dnlYwAZTELcwPN8dsZX
asXF+nFy6d1N3Jsxe5upP4ViHkzFVnC2D/ripe+eJ8eUo1Zzzm/smfyOYv9s3rDBMWAZ87PKK0Xq
UFHszdh+KSN7B5NyrbeGPfhksRAItHkS8W/5uU9qhspJdvlua7Hv6+d1iXKZZ5R/3ZSebDpNplcy
xvsHyqg8abm/XaAb/sSyj4SBqpgcQZWkLZPOQ8OCkYA7TLuHj+sKHEunMi1lb08p9jH6GyBEAR03
itfvD+x+uRGPlT06Y84ieFN7NybxaIrgCtEhMOEVlC2GBv2F5Zwy5pGZ2iQ+QVNCd77iJQtfbdQn
G5Ao0HFT16yEJO70881sEp7BVvaV13D23HSWMLtrFkbYL7NWwUQ2RtSeOUz2UOYeStFsxnHLCvV+
kAiZl0OKaaDbr7sIBdoNGsjbeHBD+0rfKaB5G0zgbORnj7jtgr4CPGXWCAGNcjpt+ej3B3SFOEZZ
m6VQ0ggqFu0uOJh9R68GDBTeCgDwFhCFegPsgtFk12WxKQfdeT+9MzayqG2zoqeD5Mekqrr4LdCn
/1TBOWv8Gal3MRCHKBX4cctHKpOCJr5lQr4iy5vhMY0H9+6zh2bU5eazF+hWb0T0EnRcsRer7M7F
Ze33dnJv0QXRTiTM5r0GCRrY+rdUmp7v6HRYSLsx+6bVLMQEgCILCwX2U5aG41fzjrcIDln9vBHQ
4uCGgQzRSeij4F5SUyXecKm7kEsczdezLV1/BAQLChYxxwjo4XflrY1RTrry8qKDdkOcjJkycHl7
CnToNCLDXuxzcfylX5jCILlemXp77H0AwI2qArhuJhziuNRHNxOcTemOhJ+K8OCH03wEng212lko
Zbwl9uQ3Qz6rTSI9vz3qVAp5EOeNlIUruuzZX8IscPLs9H6eTEi8fz6ZYhrtJmMN3B4Hxs3Ws3UV
rIWapPE1RHZHoOcQWtmHXjd0y/TPSpEYcD7xi/O0M11SB84z1UjXlwf9imY6W3EOTB6KsTqSPvUH
e/UlBHzSpViy1swttudYwOipNdgZpAubTnffIJRCXAm+3jR9hexLtU7oGiPXlCB0xta6mTy0ddVk
WBVM3FjTpzwPuKpHdhfQ8HVJ31SDW72zz8zOv0pC+rqblVoSI0yJgjWKZdDGbxJ7u+xQ/F9CdVXD
rpHOGgArG4LyiS6tq0KUg9Q/NeyOb1t2mMgNbXYyLgJ55gCMqrFPOYclY8RHlTudpSqWY/TqBjpd
snHsErFTYeM8Qc/Q3GAQSuVOoQ4sRQSzegrKlSRUs5/x4W1ZULSMdPDx+ORS2R3eW03qMjF6HNzm
uPPjJZDfuTq6R7hNKpw6ZHUWPaQ9L9FqGI5LpPvqG9cw1amjGa3NAzSY8L0PS5BrZeqeu0UcrvaZ
/eXAOViVLra3JyxyEFskM2/T7TEmLBPEJRRw7iPVEl/D58TNVVFY6zD7gSlj1uzeyckf4/x3yp12
Kjse8dr0xi4v/OBSW6hNV5+K3lEJ2JLIRTHYvAsEze76BglSUIirEyEfJRNguQybtbNLtqDOZNZw
jlBGL5cQeaSjJ4LKWUhHjTfZPGpB2j0wEF++dgT6/xWZlthC5dcE5UNhD2I9CinQO1P8b1tEcow+
5rLKLaETn+nu/RiWDoHyrj4IoeTSKQZD51RyHHphDWGr6PUUROcM3FhZdmIrTluV++XWiI7rOu9p
kAzm9QhGJyTE5iiVeJ8yDNIIlyD/GUUattGXNcwR3I/lh+vhp4gLC8BHCijtuPR3ggrJ0FSAxKK8
6BWffkRiY4P0qflvAbxVrs7ioYo8NNHYDFoEjAt2X9swFVzeknN5dHc3A/FNabs55YLges59mrZ7
VfibzfmGX7V8oTVJSDXBy1X3tffnw0ZsoSTbHPP/UAxfvBF36KS3DydowK6/ttX5sVAh6irNYyE0
AGUif1UIVfsOQaTPgG+EMgOcEriW3jpEGaTyd278Y6A1Mwoo/CQ0O53NNNehk3p7Mrfxpl/w99+D
FUPdL7M/Zu4siwder2K638nqYbWRncAmlVKhPQZSaayl7PUjPk+2G9qw9A5YkWmj84hrFEGdE5T8
78clO/NiAm48DywLsxeufEPPOFGZz9LAgOXh32EDl0wV2dI770xSR73ceyTWBh4Wj6FXMsxfLReN
nCeq01BtBM0I7PHq/sH6t6wG/nYcxu9g6LUJybln89EyAHL29GSrhykfFgz51BUI53iPk3jL3tKa
alWliQohlRXwxgJrhy+n4PL6PN6nBbQcTlx0ykQLPBHOk6BY5ZuWqSgq+vRgQSXKH80sGFxHdxvD
wFuBjl0nZjRO2vwbW93H2i+jGBZZUgXrfB/aVUMSjQGxhW0A0Izbn04A23V2zJ8lPF4NaUyPKnr2
90ohk9YFpgFssl3MC4Z84jCqM55Zt5U5EVtc2vi/fwh/3IhpbD0kHA44AH6n/wv456BXX0gXpgzK
5wcSJbMsC7xRcKO0Yqju1/QVUQsDUQn2zTxlVAaVRhsKTnHx+tks7yjxNAwhG8PLyCdll6ajbggh
g67ol9/3pbsbN6de3Yi84yzdySPMg7q6Yk0uyoZ4ZAYnx4movFBzMvtSoqk8valFLru0j0c0jC1n
1efTKkcuLkPoNI1gjAe4kz7kfov6CvtWx25DM37v2r7ZsywlvNhKpCyI45chi38B04QqqZkpHNQK
NmuE5gFzo4ZYmDZJoNr2BmCUeySmdTkBXGJHZ/qEYoWxACqrkWsTVd6pChZVPyYZx0SrtGoJwTKk
ogURyOHFp4jJH5sCwBEX2dajTNneQDtqUwBv/ikoCCLt5UbprtlomNw2Kzb51zDhiSvxePhVZ8cp
dkpxlqP6wwDAOwsnQZMKqG43BX8JmUUzpYMVU5vW5aNbytnP+P7Ljv2OxYOd+ha+wWvTSnOOt3LO
YZ82uBuW1XwyFsLMAYUp8CqaFcBiSWwWRifr7EzX7y8bwH44qNJ3BiowHOyVRXEBirZI2X2eg2zo
87UfZ4y/8HF89bvV7tLmjXwIAZb5NGNLQswrCPlMA+bIQtlacUw1LgKy8UYDmXfV0wIfC6Z6kVMt
zzPLn2a2wTYtFaHGvWl7Mc9lc04XIj6TiUPAdLk0QZmYbhIxsErAiBsf7sd06migT1XIeLW450D4
RqMdu4THkXUq9QcMXt+yiyjaWuvxKouUu7IjeL3kJq3AebgiUfpCG2g+qhlqx4lME7qefH2bOsoU
AFY1jCBLH6RcOQmAX4IQUHOBtqyHYdkhNTsNQHAb2Fu72zWJQ95tZwgpdZi6GtRzVdc+fdd6pOSM
Llkbjm7yG7yZw41OZDRl4PB8YB9LW5JNP8npT5P5cSOUVkaiKmoHTuqkvIEHhvEgGnunaejebKOU
EODg5pnTBeqwqQWI3immBpXr6QmKbC22+Rt8bmnKd9c57VjK306eeAuzXVFNrz0X6GFqvWMrKRps
X2trvFQgOe8QkKrkz515hNbrUO1/Mzm1huwHaXKaNKGEabDv0nkB/GyZklHTW7jCGRQP0NQdi9KF
8WiEhGniiC3ef+AmT7rAZnx9vJ5vozx7sRlJ853IEpb9G5YuDEICGac/veanURsbeTQ3scM9oMkR
oau4R1+Kyog/EeaayCBQI10/9haQAQkdL8XTdJHcQInYxkW2iu769lpNsUlzl4RjkOJcx7LoFt+U
Sc/S+In2BEnkS93lW11DqXOyyJk+h0ASHseqrjCeE4rp4CsNwvfMOKeuCRDTpanmj0ftEPrumBRz
HYWqwKsYc2eEYz004WyS5gqfkAV3l3jM/ciFDkH002ZuJbnF2LLPHYAO93jZbo6xGhLZCGNsjHhh
3oVIaUmFgz9+MEJjcSq9vVRU2ZDMao90pGhHxvQlghcJWnD0f6skGEUBLAZ5X52+s3WM+0jQACE+
vnQV1SGQgbzA3/NrHsUjoxTHWccOfArb/DR83WBphgVm7JqvXwnUpKqp+c6FX8E1D3KIjGLHrtmp
Am/v1S0VUr/nJn7RfQRKQSMVi57vPQJ1diA0mjYujwMTt4bmTJ3xfPL2xLmrFsWsNoOO2ffgx52m
iA4pfOe7KgNj8r4UYf6Iww56omSK90/87j06PuUoZsbHXIkgwVAubG0sWx+ml8KznAVXDQH6MmmA
IGCj9eOPje3rBLbTIdV1qSQ6jr6NAJCrO2RIcfMKK6X7f15IBpdK5zXFx0sCjZTL1gYgoB6a6taT
zYH0ikxtWIEVyPCi3JrTxs4+iAGnes/GSAW0KfgIjTBmV1xqpiXx2++PbPeTpGs4MiQF+NFULbAi
sTJ9VOZE3CvdRruZljtP4N0CJ++Gu1tKMJXU9C+WPxU0+4IUxWcTdyjJGCrqtQNGs5LeQ8xYt0Xw
PNXE+ExMTMKc/rmkXSWbk6BBxSwbVAHIrOJjh3ZXFEgHV6sjy8Q0wJIsIej/PjD17gBL/gJEE8mU
evmWZfEuiCLiJQrFHnaAhF8oYGvOYyuAoVyEl3fTWPxuw0O4Xtxq4ZypWbrQyKdsXwEFgIXwmsMi
AsmHAFIw+LLI2oaQMPbRpVo0lR4d4Vp5YvkpwwUXNR0kkwSS4rCqzadI0cuHh38P2YFf0onOonWj
C7FNGyFgM/2j0NoBXcFs8RqZUuTPaMV18ocaU4xUFYTrPtdcSA2znjCUSy7CblxlVZpEwgCeuYaC
pLokhvoGAcggRp93ve4hB4S1TJhfcLShyv6dqXbLXdX1Js+dHVoipWg8YKhTwej4HgeDRbP9HHrQ
pOAr+b7WBHVtUMr87q63WNZMEEqmM3Kf8QRT9IlJFEtVuAWQn/iM9uHyj6Is+JXt8rNuZ+R5Al/u
BhRXd41+CEERCTkejA4BvldyQwbOL7O+9RNY+cXUSviY4IRhue0fMxB70Q+QiyrsWkwK+F6LgyuF
2BxVoYKRz3xrNtLr1P87fCKA5dZKLC91d8PyYiN4kJTCyP4emJ09ByznFaVTJeNMXxmpf/BYEmU1
HqKYvx394JqCm/8rG/2uU1XGLYQUdTcYA91O+ssaxYklGGMifG6Yvmfhb4jAhUoIsm+HRIyFi9Cq
zvNXqhc2dcAHY9V9p21NngphEq0LSy7Jw9B+wRGoL+JttlWWVqHw4st5PJ2H2RRdxSHDYPI5//rK
eucjtjeY+9uDZMDRm5M4iqQsaUjHDPTJhVy/PrbrPKM2q88n1+LBa4y8YQmXTLKiGHlzfDkXXHB5
IcaFeXVPKe+/KnQd9tpmDIM7FfGgkKgB6KImEPhfR9AKGelq19dtwj75qiyuYsI65aSqu/Z9+7fT
LyOYgVD4kkfUPA0dR4QPr6Z3LllyZiyAbTXItYD+gCacDW0JSioc8EVVdKTdSYWMT2rpWboz6j5T
QHq1YI4+ZhQRMZzYq1Mzu41w0nrXFXA0eyfpjwXzmy8vZ2vcgdsC4do+Eqmu3+T0k3OC/Os6vXDE
5lyWFTp+eanwIV4XIy15VCBVK35cBy6cixAiINAIQlEZrZCtTn2YvUUVfP9XOqh0/ayU2F9f4uWV
bOfqMlwQ1mL0g/eVt/IzOs0CKMkpbsnR0POtSsxYwyvJpvPPqKqTqUCeuhh6f0epwZkVoB3+CVqz
0JvNQelAd8SMcjc6X+dBVTi8BaM1XwGdqkQaq/9TYB5fMqcV3rsh4cbp5Rolb4nKjf1mF96lvuRY
Qb8C9nvA8PTBWVLjLCk4/PC24ff3bwJSN7iiZm6Bo9ocbHZenVPLvbf1WuESZcBN0DUAyb2p3UKb
nwnrwbmLTo8Nr/tfQkogtCl7sk0FRGBjeOzUDNflZ3671i/axWESEAuBZwS9AqYU0/qqkNIuBGTS
QbDfbdoGZgQI0ePey2uWGP7zIkad5H19D37KqGtsRp1p3lxzL2OxCvEmOfGMdI9QuCNxIPjDtSmQ
SazXKwb1CH2woOVWU3ob24uS2NaLAo9sdAu+lOiJNAQN3fMkUhKTMGYTF6J4E4UA9aDm+RcxJZsw
V6TGvljNV6hNkFRYXIbLXro23BPRjtuJfIlLKJSeMaEtbJHYsuRQuaSWhx8S27IhjHeZI6EC4tCI
gSQhh5mGTmc5iVoiTfKCSBGKtfMd0yCA/ulIGNPOHd0x1m0v4BnoG978Kh4kn/Ta13cb00E7Xcku
Xx/teus2J/mELzJmQVutlVKQ7NCjWqObXCDWyw8BDvVo1I4oDU4xAPsv1lDNXETPYOwWlIvpX3vf
3jQprgeHCQry4oK4glP9PBADeRwGNOwlYIWU6tpe1qlTy9mYw0kPgFu4icvO98mpeYRbUxfUE5G2
dLJ142Pneph7+CkZIn8ratl9lhl0z53B4tLrRaL88hwt7FOuw9BEzTXyltHX7a5/8aYxd3wZddEP
wnd6KgE3TUr0liG+xAAhlDmjHLyDqB0FVQO7ATO7LsOS3ZxC7YjHpYHVn6xXiSt/T9WIDoequyiY
FM7PNmb9UJUiUyE/XX7PxaRTOJEWwzNKZ4SRoZ+40yxOUCmg9CCCvySqQhQwgwLMYq5hBUnDH1/u
EHkB6SzjT62hbfC1ZLC9TDYWcYs9VGT4B+i+DWKsLpS8cK3fzwBeFQqK+OfZzjC+riwsi9mZY6qj
RANMpH4aFNkGxZfL70lvqFGIMkLJFtxpHbpd1ghDAfwPDU5vAH8cbtNX6ICrwOhz18E+uyRfLzxY
InOO620rE/Yc7XCbEVywyLLWllQ17IcYl+NYApqYMs4GP4Z3cox/zsBHc3cGsvFqPRDTF+hEKVF/
Gn3ktPBe7bgCB5rgCSxhXFYopRDvIB81obyHpo4KnpuO6EWEKlpkdKVt5Zi9y0CIt6yBBx5bDTXw
AswOEMlxr2t0nPTeMtPRYrXbYFxu8W+zOSNU966UsRqhpnCojuANZnqxNR7+ovDVsOPJVoxisaHj
ffVwodrRdtW3RzVeY4BHranuAJph5FbwNEoNikQC+j7iDITkgZHMpmPm7yRNTq1kUDQAdE4qdzIR
KtSsQVo3KOew/U5LPhbkUV4teDmdekY+cOPVW68faCXjm82WMJTDc0/GrBZfp//BdMuQi5oGYrqZ
R5IR6WTatES0fYUK1DG+IsH6zsR1lL8wvfJEh/hkugVSStlf2Vbt3MptJZE7Az44rzSgLu0YArCr
06Vb8ORL2LneapcLBJnpLx9eaWPPKYL5gMIVlaFSw0kyt7tr6OkhB1JszScH2lJ/X+8fZT3pCEhx
TCnWqqkoJkNH1PPgciUeO5upzluXbcu1THav2pZHdpHqJatVsDMXq6xHE+0S89DqwFbTGXZsiMKJ
Bt7E51SqhjspJ0jkPpBEcTYKOVAOIObnVlBLOqdlWRPcvAsuxw5ydSIxcjXVPGp3ORiyOClcH9q1
ucPO4mNGO5K3UjT3vAXOYreI/Xzs1MUOAoYFsSxF9RhFPm1RVrJnXuCeNfUR9zcQYjbIhHPgIj+1
YWrXbp8RfLBwS2SwIPlvgzEdVRYS6yvw2lCsUyd5AqMmKqXoIt/CTgkiVt+c27UC0ncJbS1viidq
IP1Yy1Q1IvBHDKb4o/Vf79cebc/0vMo8W5MvQg/jopA5s5btSk4tvMiCtwd2JJfLkdhgne9Mo/hq
eZs3aPxH2v8N45O+Vwj4YyNN6/JZNDq1DtibzapsoR0o8VYv/V8EvsZqVzjiT/b266/DCNKJb9uA
+XGgzJRzKRpsLQQd12FGkNhasYi2XstTms3izdEhaTw1LGdQM5ZszTuEKnRj2D9mlj85ilydAVAe
FQIDxTfAKiFagwTrKXRsJ2KUF3gg4En+s5aJMt4q1q/2LV1MA/chSC72pHkedJs66x4uhRn7UIuA
tUjUWIIcSkl/IfmvFLh4xKe0a0nvHq+uTkwuDNptbEY3zYFpBkjrdKHVmPOPXTy11SwfvqzZcxRU
CPdWI4MSpMy0U7MXemhIKf6cTb6hG+Yt/vIswpXM1nkZCiqS5U5hbt13XLQaDKc2vAq4E6mFsXCo
WTwuB8vuBqfkFUCSdfMBlvWrhhhSXREpbGxW2l3Z7qAOOIlTvJTCfJrzurtBU+Kbklf0qW0VqXy/
aJwmC4d/nPcPmcQOwi4CdY9evLz2nvYqsHeD6qQw3qAtPZ24LqP9jS/LtljoH+92l4byjcXPsWuK
b4BbFUZj3PFZaTnSiGzK5v43nyZkid7lFHMr+zjb3LS+033k/aOrjyR1q+ty3u5T+jkbli3Nquxy
y/04FA0049gSFvwaJAXvHPYv5dhPavvNJBUyPf/zsEU5JLmWlZkEs+HU+PJbrMTnu/2AJgUvyD36
hCR4UIQWBcvkaxEG2+I4AwYAaxJdEMEOH2vAsmfpt6n9HwIuk1wnEBfO0NIJZOdP5ArQrdNI8DYS
+iXwIxeokjvyfjeO7jppKq+kkDsC0nKvHRDdjXAoKkNiUjpRZA8wep/530oSKquVf4R35ZKpDgEN
qoFyaKPNKTXHLK2SpWcQQ1gl745yci4w5HO3h33VBJA/Lle5y0/D9VC2OXOnrLJffWi/+EZYnLas
xsYQRKZWOa1SnvYoSwYyboaCblGwJZOqrRdx0tjDG9JpNU2TBaXHiIyQrOjVpspP50VV7WN9EDAb
WxQFISmk2J00HJvT9Pte1iea/r1fPEZooZJXHUN3qj4lPy68kr1cWpkQNzr7gFlrxE0V/i3K4tSx
PdMr8h0QAtERUvRRJVhZL5i1SSBRG0oEhJU9SIUnSFCZTI1kEynLO4hiRwdHGk/ABLc9Nvc8zv57
HCoLK4NwqLQFCkQ6dQYikR37q64wzD8CvjfWJgjSgaZZwmdaAEmf1HubAb/qojPxTAxQ9NA0BvyL
Text4kAEXICBZwrqBDqgDfyDdx+DwLmD1OuTWf02BVkRCu8nELshSYZ+XVs73N6vJVh1gIOpAeQb
yzKpaJcq9zLM0WYERqrIt1hGfgyBLbvIcxDCl+7mjj7WUiOCgo4wUraEsmv1PPGY06459X+KW/GT
p2BB+K+nxkURMDWiwrnyucA2et8Z998rBxtLSjTMOMvcXmhKCSlp4axixnJedm8MXxJI/2Ohh2Oh
mrKOtLxigZMH6ENW/J1s7zqBhj8ZsMffLDX9jP93LvedZcY1OnVbw1IrdNm5fQIA8ZqFpmcbJArA
OnD5AMfnM33dd8ZoDweUC34YAG4IlR7vCkfy0kno2R3pt5thTCTWLB9d+5TwACgA0pYkYqynn1UG
ZowuIY3DrM5I37+PgLUt0Effe6aa6swNkyYtDSKDa9msTcSBe0vIyd7Fi8FXfg5E2udRV8YPsQVg
yEJRYD8fhh/Z0K/G3UAOsSTx29RGlIUxLIX4qJpPwP/kDyKge8pPflulAs75ByNsMxbVZK+F+1tN
2rA6MvToBOoaQ645sWA5qGpI3cdtn+bzopCq+x5NR5ddkR8i0h/z595agQyHRVSwTism0ldnueTk
zCNn+dvhbNVnHfMKY1+9PAtwvmx5XHYXJPGdDF8dT3awAymno2eWmNeukOnii4V8UExMAV8R61Ek
NAZIp+nxQzpjQ+nhgGcMBk7EgLsW4+LFSS9EJ4GB5p3PerDvxTS5KbXM+LqjREWY3IVegN/kE7tc
lN9YPmQcmC6P/IgSVfcJ3pt/3Q3VgrYYgNcWwu1SPnTD5KDL4Ci1zv9Vr9xcn/apx0VMmWEcm3BX
aK4WCX8CPAMiGBZEGUO4vDgKvGTCXSmcZgiPGm5FcZ0CPAEMa2GGkDAjNkoQiXZVobxyX/l+/mft
mJdqqiVCXh5RuvEzu3sxC0Biaqd2VNSZNEKIGX58HCAJk2zHsKbtDmSdTDtKU7EM1Ml7ZReG+Gus
om0lGy7HwhDLJtKKtfKsD+Z2ZMAgboRc959BQV8nrvqKuRTTni8+HDoqcqKhmhFOgOI/hz/sbnG6
YqLF6jUVQaztj4yySkV2GkukqNJFmonuzlJkXrN0UPV+84MpRyFavj+vnNU1u+zj60Bxl5a0705y
yLW1vtfZBvRumPN7L1wQ31etOoDX7Hz/5rpp/03+IXXkQEooxNF4POvq5c07UT8yNnJQ2MgTWgji
2ITwabK8PZPSPw3OQxRpeRuib5UtIXgHEd+0BHG/4ZkRT2dnjrl0PFIu1NnOcwfH7DhAO+YJvsRk
gsiyskxK3gi6lx0SRGcWq7g5CTIRQ6a2Kptf6jkeuw0GEDlx/tQ6YGlztvVinaj7ixSpqY1+8oTw
RRC/2W+FmE9fpAoFQRzlCuSc/WSk3/R9k4KrZbnuB1TXMjhhBQLGW+YIG115AfptEhnAUE4tvIBD
Dlb8/09QXqFbz74jGfXBIxmdxyFgQGTB2r3sJ0PjTSrwXd1a57mAxQ6H2j3NPIB2k89PPCk3DXoJ
kwvjC+zQhP8+TLDbgLFmhIqti9YNIXL/3fy4UomRc0QBgQal5ZM5yKM96nhnzwcamLsOeQsmj6tN
NfqrduXk8lsmOSlG78uIEDJNHz98T4R7KGrLW5Fw4Iy7hkqYs+HMeRjBECe5higJmjEY+VoD50VL
64Ok6oDPrO2ysJ4B1l0TqKPXZC+8XcSU+FJH81zwdEU0UqtOVOwZ0b9sV6OGodFUMrqxanNyRjZd
3vXFiXvXdfXLJkuTBZ0z94qFDAFv6lnKc4lO3jnDYpFledDSlYBgwPjPVjnsuQGt5D3Y6deg+zmb
mBqb8uE/C9ju9tTFXIIKhk+LH5LFnpxFIQtvlfBbBe+wo73vzRQa3ll/1goVvQRVc59DnUJUfiSS
B3zAWg3ugw+eMNEyuA6+dXAXFRbHNKMMi4TYqtZzbmfDEpEaiysI/+7xAyTJaK9/njA7HzN247aH
yEYdntVQPNGSjDh6yiSMjKdaZJuXSOh3FPui5rZYIO7U1QxqgtH0pgbpHMR8SoOZHbnEAHsk3vmk
8bXA3kcsvna3MZzsaN2iWoaimuf9w7NHis869IdsmXf6YMEIQIvd+4wlTe0uaI5Y1GvnHdBx+z46
Q7FiTLqUdIMzLYudeN3G7gXn9kXWGUlpjbpasZhfvRHp8NfyR4Z0eT+7FqxdLeeoXa6EV/DRKM55
tECBqMZ0i+xtnvSVj4+DZmuLEtscMRglUXWwQTn/v+4mEE8L1Ka3QGpth9H751BDqdcBc5KhCa+c
p+ZYen586g8hzR1zuwY1JkYUAd8smbc3N1lDzlVyX/hSM73nJeaxV64ynPTagwcafBxmYCObq+mm
2DTDrbZM0cp0u026c16ZyMoAOiO3VHwhr1V7csBaaanT09Hors4OlsB8X7cbQQXWU7tocEvFGcn4
UOY8L9WJPbQz0gKn/zw1eyR079Ce9tnSextTQPUXcTeYiJ4AkfTKQIbwrSObB7C3p5gTa+HsLeZy
czE/Fv9acaImQb7384IGNwvIOF8Cc8FRYb3CnDY41o2aOZW47+jETB/osYPnxDzZAD9mSaZTjPbY
nF2o0Y4iauEy7vC4dDKnRKxgnWl7EBBpir0evlyuAVIcnvpjwKNvxNSlKHin1yngfCAPuowY1rPz
CNtUvg6AsFhaloy3xavp60vhedu0pbPfcAUVBDGXvmUHjDR6AhlOXlqBSIbd4k8KRJ9wXAdtkCiU
uN31/xf5DVBT61lYw9oSMHUce0YppYfa4qkLc9i6c4aw0Z/GwTl+XvcOmb/uPetcqaokoL/KmyRo
XEg5eNU31qU1Zf8e4dGbgFl0CfBIsnWYovgpoMksRsFa3Ff6LROMkThmmbrthmAxtlVOnY1X0s0A
2t0z3oc3n6aZqf+L7B9ycip0u23bBffgHL2MSqYqL0NJXDZimIL98W6Ll2t8I6P43x7X1tVp3xGx
BzWlUAeTv//+Bkhv3ODHPztVEitmAgP+tR1PaBaAWwB9hRNPxS9N5y3yhKmNt4f7N8ouaGm6xKQ5
+OvNc+trtcE9/OdK127cTC/NYns6n3ZRAmW2zs6On6+W/CTmu5K1imynxXoOgagp0pN05PwfKGZx
P97crdR+SaReJL+y7YsIzIUvL2aqVuqGjwuzlRe08qgHhLkRGzdNR2NgZAacOlP6k/RHUkj+0MmJ
E5wgC3KOHUC+fbxSQkC3wI31vB0Fc3oUK76i5uttQ8Jyc2hxdJcJHDWlB/q5v178N08mc6Eb+ITi
J0pekEHISvy19E2cSWds56dMYPLq5+33/PyDUOEKMW9Rju/zb+dchjC5Nv5r0Ny0k1SBrXPuibCW
T/sTR9YzyzGYZkpaRyKeaIv/rCITI6xT+Wv9Q8IKTTN/024B6MqTeWkJQMJagfvE4YRcAXBBbBdC
fT4I4c2gAhjHrrBA+CmmswTFvBsM/MZ1Qb2eqC8ZJKGhyNUAXS81z3lTQ2m2e/DzDRSu+UrGm761
xvYUHYHVhEFqfshXSNXN9TgLWZMqDfLqe9gtvldB7aZWxyRA1YGzqbD6p2REJG0GzguP0Zv/IqIa
B25gYKjy3+qARwWr8BruI60lzTlecgel85mpwEe9LsL9rADw1CUH2pHaemJ0tx8/i0GipU4cLXDW
2pjuPVxTvn/Gok0coQG1xHKOYW8jBXsnK+0rktX+cYTgMaU2BgykJpEFQWay6kFg9jKpgHIc16Ta
uVVT1UbnfALsH+wwnwHc2pABViXHjoRXtTI75T7V0EQ34NCNiuPrJrTgsc6pgOP1mwWgNstOaxIL
8J8XP1+V88d1RkSONdORuC5ryDJ0+nF693j6MfJVNxYpmeuAhBF6VSNeTwhxao4Xp7uLoGzb4BMt
BdO7GtjH8oreEv+Iav9cJk06vCHdiZ1cX29Oj+g2e+xCxUDCIsrHa1teidmkYGGLjwxl1KQWb/NX
zKooWBMax/Jf8tJla9aBS/Cc3jwRArb1Q4Q9mgGz7vgubn1mCIlnfcwgKPV3tJ8mtIim476Fx3+b
P+cZp5hLGimxLyioH++Xw2KM7cJmym/P+Lf37hEIg1jP09S1rnALHDE1xrhkBh1G4WwuxcsF6/ZF
tKkdMrA0Is3hP7XMx4HRxz1o1MmnbTcMVZlDY4sxYLols7q64WxOYq1zJD5OjhRIbdmudXPHXsjY
KOhpphWye8QvMpwYGwOV/DOZn9aIXm4fFtf0hNhAwOmAUnvC8HOsHt01NgYva0Xn2jk7yace80fO
4ozHb2j1xXFDFBIUfE07Eb32lr40w5nZ281E5eI0v8l63ZRZWZGoBrE2MxPIu02cDGZl5m9cKQIZ
VHs6TFEcuLmttChb4Be1SrW/Mm6+RXq64OMTT5vd6TgIv77p82m19xPxONpaT5A4R8uwsiRNXRgt
tykpwIwFPEr75FSGXOKWWQGU76BVeyBsUvtaJGVQsvKuGTU89tosbAmedNnzwQWaLE1Mbm/Od1VO
XGskdze8Q+shhme8C4IhBoLfD1Wb5ceFlXlhlSwi6fQTRIMM8KQ0LJvETG7tT1F6Xk86143owhzy
JSQ8sgpLRpgsTtnXv24eO4EgUvrZxuMcs4gayuThqV1BaVBkT5+lwceJVl6wHJfLOBB+4vsVA2E/
nhcH4ez3HTJ9OWnHbt6mSLd+0eavXT51lPs31J9fnEfUdyf3iNbLZy17k02rERF9WDVexFpWFebD
BOLp7JXYM0BXdm1UZqAtyHD+s3QVGw7IlCVmYEID3v/75tLINB9XrQmaW6WvOmznk2k83YFzRHSZ
fkfjj+vqrp6ADhnskGg6Lf+W7JSBNanfalevml4geQ6crfVDLwb7I6gLV4pZvD9FXWg2m8zoMKy6
1SkWWNzmasdj+g/dOKdv8zOmmuWHjgOvLO4AZODUUSMpmZvqTxZliO3OuPqoJju3XYPm6YJ2MJB8
7x+M0vlM9IDFkYvGJPhh2puGwYT4xY3EnQWxdA6NwsVTn+sTJsVIa5VICBUsITVplJ6D7OgR79Wz
GvICzFsZuWrgbRNulZ6p8TbHZG3pVaP+qL/eeqZNTecrdduneo8skUDvSudZT1jP/fCK0tei9p73
h+s5kYN5yvx/1fOyP1u+0cnSE1TESgmsFEc6ril1HLF8z1rYOSuaYgLPdceKJw0VjgEX6CsRt4ul
rDTNvsjeTm1+V6Gorw9MJK+iMDt36NTvzZ4Ttc4bGv0s97ciRUYv10EbMMf5+GdCXB7dq0x1lqui
b9Kg38ZpglBYx44h9ViJiKidL/nzwqO71ggorKU7gOf3IZLrdVeLUEKY/56NuHFmo/UuG2uVtgaZ
6C3Mz0EMwK4s8pwrGs+ZyL1cEUT2MexjdeRlyt2y2rwmyxOqOtIu0epC7S+gTb5RCbfk1DVjhXFG
ZW14jQ0J/yK7ZTr9kgQQi0ToBwfVmE1ZSJmfKq1akEqg2wg/60+iW8d42LNzjAQekVUnvUTjcieh
vhbirZZgUcdyrSkuVqrGsxyDpC8HTw+FmFxTs7tKUHt440lAo5VjSzzNl06m5shpBcge1YFgINB5
KR8xIzlhi2rI3BiWbTYvytO0v9pTaJJlrQlOCPh2WxtU0aUeLhnh94bc5LO3wYBtF13RlN7HJFee
BpNXedDCNnppHoeqRzrvJ1kckGdSuUvvSuAcsH7Cmt4whXHgDuc+2AIstRA7hMjtFBfuUplVRX7f
hBDO1xsLMfNXZwrQtzgeAjEWiT3IlU8qYUaLblZmqhPfh9LRBQToDpaVSR6ChIfVQ5HmDubCHHUp
MIUbqIhiRQj2rMRGWBAg19cEnVpim8cpwtQxe7S8y2ez9pvY/7mPuaohiAp7r5wXzTdYcRXkL6Pd
MtfKUJILRpo5z1lnQQq3dwEbe/kDPyvZ2fPBgCJs+SAmIGWaN2LKrXWMzbPaNFREgew26NLA8hH1
7yfSPhftf7I4TQD3rOvYjtVO3KyonIlwShY3E5/0u2lwH0e39+ioKFgnm2+XCDvPrSPu46/Eu0T2
+wa2k+JrtfUf0xS9nvK3UN6S0GfImwyGLr+rUUkcFb/taRdmyf5Dp2/ecs3P5gfmfuC6c/b0hfRo
ghVyWl6LSMZ7NOrUY0AQfStgr+e/EwOLjsNyygfAoEcOIc0fJ/siqfDYU3Zef1dV1sPZmW+vQcQb
mGqlQPqwPXBKJ5bmD5mqO5F7BMwwYbfVh861yoljZ9fE/zwgjbx6ay2zrTDzO0T0PyX0Zwpr5oPl
tEwY/iLC3gXSoe5GYzDhY8+ILIU5AYRMPvWlTpFqA2TYst5qcZOXMOJvmfLSUKG/kdxv8QdxflIF
KzvBR5Dhe4EaMplWlngIy58tkLMMfohD0BO5psA6Q5HJF8f0KclrfiF5fB0V/ksp8Am6DA4cJ3oH
meSGIR73EQ32+ce+C4ECDvkP3HSPXqIwzedwoGRqNwGK2U6Vy7mvAXyjASsM5pK//ofofEHWln6D
jbVX6xEbvN1Y54FJhmIYD2XmB7MM/3e2szLfQoT7z9bzYbfNRkOmRWODqwN/nZXmIBZCa+iWZQsE
ptkSjILvOWh2etFdfijd06G9Q/EKHMJKXTUQqygco6WnWoeGzIL5Elv3AgsuYUHAQAoXdqGJ8BBf
EW76aXHyPpFMsWhfRKKHxkJFTPRA/gLlXIrMCFWwIopafoUTQntX9NOIGijj/iItpG7XVvqZjPvr
RH2Yq0I27P7Q/OjqQfxZtWQVzxLTtejEFzKctseVMSNciccaRgbDAOFapMKw8Mw46kciCcIQzinJ
KegkXjxCyBq5oLn1Ubj3IrnM1y5xU3pIvQEtI7VnFQFSU3bn9JV+ddsCEaCy3m+U7aoUwRTcTK2b
bR/eLNBTdMRFBNIf5WV3uc8MgPHwOtiI8yFtj1b5hsovGwYUXW230ViEWnRLolWVkZVvkKvWuDha
y7E3pn1veksEVCDuiQDmUix/Q9tkUrR361YoH4PTmi2R2tyHV2Q6upHUUfcmPctXrj5g5kFb4jYs
hWoaYDadEaPWOszoI74xe/xW/v/n19V58lZVvgEe3dl0+NAs0UQ5eDqHt9C0MvMyCalvxGHEN96X
VawhD12VrfcDzA+1WT1J/fkW8OVCZ9s0lWt3xWKM5zEJoVgnkivIUk+8P30kxlQU7w0RooIGcYyp
zXqLWajY3mRWgKMxi7ELntc7jM/sG0h+HD3QG/RJpIhXWw7by4VSZaRdWnS9Zvia+fTBvq495q++
NnlxgdAmd2LWJdKd+lG/Y+hDn2g5XGBPcmu97VFmqILFwE9NwwOu1N7126d4Sr7lIR+vQV0o3kWE
g21RDl78nWLWjp5IRglODxse6y6Tb9CCnuwmJfmxVkem+lbALbUXDrO2FbZ46MniDC/8MhTpKiEE
2WGraXCsc/48ATwP3h/v5b7GrGiKEN/DMMC6zoKti7Vz13BIZ9OnY+Hy1NepyF0QwhsNKzaGTeq6
nJKDTJxoPC92RvgrtCPIuhnMmkWL/NA4sI07iszkzR2faXZIVnVf2oAcqZyoQL26mbJbnWU6GueZ
csYhC4J9VpQTGCmGzDJ83GWrX9ihxDOgDYv7Mv4ua53Fyp6+mxiCbdk1yz6lCmxjffrCfsqFK7sT
9YXhA6qzwvUefuw1vqvSAtPtfx+V11SjpyjPcIrdFwVp0puCGihhsoQPLW8vzyLRgVcqBhJ33LI5
oQAIp6H3PyZkyG5A7I8G6FraLSX72Ih3jjjucQDhFKtDYxsJlJy3G7B1BWRlM47Gx9rX0QNA6I4S
qrB5nG3TeoC4IvoJHVmchiLGx8Mcn6OXIaUwH7h3GASwCnpeIwv28v6JdXIKCqnr0NyhKW9hZBiA
t1Go/OytXYoGNbLJZL4RtVkDaBC+NZtQVfGoTYl8nzBNTbDPCZxkaWXmHHxEJdIiWfUc0SLgPBzO
sgkNFmkbA/wo+DK8SFIm66YXM4Jmoxy8OZL3KIfYeMbuaVP4o5KtP2KWhbVgvvJil6OE7sAr6+Uv
tDoFeucmUtF07v0INEtAljEIZZWlVxD5IaMog23pp/p728S7iYCcWGwhT19kcs0YnzR3phq8/fNC
WVeDrktvlt05n/dNKFbFMvVI/8mLFWJs4yb6aMQ2vP9b/w/cIAv4I3RKz2VnH6/9yAMDqrxB3L12
klsWsmvaE13pRbIXWmzkhS5o+Ryon9MijN0A0OueJTRWkKlCw1u0my3dWP2uACx5LegSgixSzp6X
uz8XB+iRFVP1h8OZNXf9Wd1N0mo8vKqapPvKz8/jzca1Yoedfxw42NgV/hPm/qHnJT63h0VPfR1f
mIc/8fFKSOPAelW9nkUiGMR4Ob8ZpUDbiOhFW049DhlIxwgyhloCr4HXevi1AnwvxCYEEOpUn+J7
Nswxl+MMMCfcnxqgxhwoAQHvUweatmBHPCCdh7rNpMvHYDSWSAxaLDPz2EniwjpcgBsvpfyfbOTk
eL9zlyIS5TQHTANaRNYsXrzohvOozO+3V1Fvad+39oxYPSOBIL6X0rVMXOMExsKY751wWZwqp+NB
Up6mVPaa/aVBFu8EhFRcPVItkME8Zh76QFC6BfyY4CEQcYzdpFISoM1c7Pbm0LEL8lnitP9vBGc7
sPYojuCQ9Grv92OXm8AGkELEphrggUe6OyMHUxJUMTUewXiGP3JP/amc9x3K8ovl0EQayL7823dG
iNRG294aF0tt29UYlXndCT0yeEvC1BO/nNK3Q2VlwBTv3zwoGg6sbfPnDQUuKJyUnYmyf2gjHTzF
pgdUQ115loa26UKjUL1QxJvzkD0/T94DLFpbeGIuzVgIFZePnvzHDL6rlU3t5RbfPaLmwp+0v4EU
M6bevrKUMZM7Rr/WSHwTgK0Z39ixqe3BKtda7xlhIeAQ2t5PCPHhNxIefe54tpWiqv8u4oRU45/r
ASCIPYooz6ybGtR4TV8IrFNmJ7H3E76WnGoU5NI/35bTCYdPTy9l3lzBXdgs6ksMbWAK8jTxtVZd
xRCBBSGhS3pVE5r7LCNvyDC28RkaYz2ym22/CRFhtLv5rvs+FYdD+l7rXCi9PvbipV+TSdQ/bodg
l1zjjnpjwDAZsFVjeggVh7t5vfFynOdnMnvWPEeXvF48g3JGgFh77EU2EI+QSEC/BhcLRqfYNsop
ow+MWjpWFs1zIDtsuyfNMpIz9L1c32HYOqJe3dKLTSaIzsvE3tVS1oY3uyDwp8J9nvLlplZAcnl9
XkIk4fhtPZlo2r7SWqX1nSgN7BEjXKJWEVeWQAK0pBNZfxexfdIdwTTvWZjesTw82rlEpdKq9QRA
IEj9fwHHH/Fm//v0qxd948BMDfe82k8a01O3cACmZVIiPKwP3HgHk4/PpiMpc8vgdI+8Pvsx0l4u
pZNk7gqTlVDOzdqA+vV/6/6t/ftDIJOjcHE3ma7xKBa9se/+RK3q9qZcPPec57WB4HGy8J81xzfn
4UJ5F/h/9QEB5e+ALwKmsvEbDDne42SN9QF8ncz2vLlUSMk6xsy4xBMBQUQHN5iMT0ACv9Um8CzX
rTJDumq2lQ3yUMhUEv9zDZ2KEprLddrfaPJ8Q61TBJhnqp8ytULqRYd+Rb1O8tg0PE3YWV1jtj9t
GcgRx/zjZrc5BjzV8qulbT2zKUrzHR2HfP/kGDCR52MqZdCgk70FJvkppt1xfTRmqPfL6E/gZXL1
hzKhY7yPZ4qZaiX2h7bIMs7sZ1ox7cduWRY02VddRD+WhNv8YhhNUk5UuTxVKMq/iUmSADvbS/MO
6jsIIzX8FOjlUkCD5zHCNQzP/mGe27NswTk4sl3wg7D8KQeHSgLD8mrKRJzex9LpylJS5FTZIyHn
DM4UtfsF5zwpwRO7AtYJnY2m0Hgbt6OnInIGqpdAnGhXkcl6fD081cxeWNq01QwEs7prt4IZROaU
4RC5A7QLK13DFVC2JkSSUuo2nEcxvgjHoofIMkVf+a8yUoG/88trqrc6NxbInojsO+OdH3KRr5ie
993s6dEmeYmky1jh0SDskVrvC7jHMVzTaxgBtetkAVev67mUT9N83LEBjnYXlbl+95zjf2DWSklp
LK13JC+mMtCCGhRBwH4+N/LoGur19SaJ1R6uBV3bZ4cWoQlLk1zaO+XpOslKreP7ojOHErTsqFTF
XCPC09VWRj3kxkD5L5JNMSMnHte3j8d0mftlgcMiihw94GL0dOHX/iNzVdtNpEKmiyRKGOJWCqQ3
YhTrZJRtudsJAZvWiilyqZtGgmwwPr5F2NnPexy6QO2mZoOSy9j29O/5wRqqmoRkI04/O+fK0NsW
4CRhacfrqIfbUhy2872Iu73r/oM0gyQCLgb5QMjGgTblTFEXdD+lySYUBHemPPakQbNG6T43ysKD
q9wcZ8wMKQ5nL60e9l44HblejxN0+qp7NauQb5AFdnq/dh10qBP8z4TUIfI7hvLiIrTaXmdkZ1VV
l12ziKa4SfJaJ7ccedO4y9CfQ5mgtmN1w2B+PlpH85mRuFGT1pBf/Q/ilVXhq74M+T1UxBWqMo+v
Z1/+i0OL+RWwzwdHMpb1TXDa/57Gy+Hv5GTTBqHTpyc9c0s7II+IsLyjeVp4Y5bUipPwg6etLcNK
TQG/xe0E0AgezHY8NIjC38rwVHz4F9ltfXebZsg36fQs6pF2pPUJkQCUHLJfYCl/ZyN4zSJqNd8u
hqoD5Z2mOdfcZD2F3j3y9i0fPm/JgdirYFGF8vKuVcdylx/10itmffcw/xh8bn4EDiAWZ7vZT/d5
PLlyYB32UHlgGCw0hGT8h6o6QStXx/ra8nQqRd+p5n+gAMpL/V2o+9QkJytIy+IILI27DsXVql0i
bE+nO2/8CwP6iUjJMVcHSNmOytRuLHHnjPJ3WnJDVol2kPX7e9tJrf8F3Mbw0ydc97o28iDd7pDJ
XZ/MSXmKJu0WoVr0Y2HThWg9rK/3al+QHHjSTQNhbDcXFkzXRtTIcm+Ohx4pHlqEddkJZHKNI8TI
TF1eJ7acTxdQlu7vbEUIuOATgLFB9DdKhqZNLr1vwYNzdTYXlwOXQhlcg+RIjqcWOnxF6NsIdGg7
zwUdVKk3uWZg98DPzDVQVeKZYr4IVB5DFPz3dXIslAnYxG+QmhXIL99splOmXX1r4BA5nIIYIIWT
A1Ib4rnB6q1Z8596M9y1+Xajy9PQtsr3CAWx+exEPAh4lUZl8KTf+AM2AsdGecb9WO4SKcYkYUV6
oTV/vUD2ZwS24K9+L54NG5NWa1yoZ52Trrs+6Ef6lWYO70fdBQ3du1Yq76us4TdZv8P0gUj4ClR7
SayDlFCZuTrxWmjAz0tbi289KR2iVoeCW9pGblfykqjkkekPGldrLxTyWGkEbxHPbt+7FfaQuCah
J216BT/CjM1jdOG+6Cz2ufDJwMZgpnd2z3NihK5LgcXApu6fbbV2K1QYuxgR+aLAhg7WJmnQ6nGs
9vuTxWVwUYsa2COHc3FXF2oJYVd129KLKYbHmz4r+kmHtWoWpxpP3Bhp09AUf0mf50Lw1E0aSE+i
dSqFVKX3JNC8oUbEcDUjMeRbXnVFYkOGzsPV/9yON6Ul4H+BkVDnN4DYK/kHY2DJDRnUlqINdgfY
AcoOJWktAoUFsgjntNNX87jY+Z+nHoMQ1Smf1+WPzPiceXl4OW0j9OeF14zKkf/3nxyY1I1wOEEY
SZ8yfnkjIV6gA4XN1qy65oy/1MSqfsLZNSi6FkAiSd3heQ3bLZK4LSrxxNVQNHSh7eXdhPxrIJFz
16pYRGPs742kNLzJ7ZnF9zQy43ULW7qYa3Q2ggqzivdZj8aoTbyMerG0CPJDjfOpAU446Wl/hSxc
EQcG/H0k9NWGT9nppOFbWEuuZBlI66ezj09+Wmb4ENV+1vAVuNN92r6hmgjTqMxirRAZvnDIqI0y
2gP16K3+GAm5DC+Xh4ZN0Twaabmt8I8mDVM+/ts8ZlmFoPmTtPTC02GtyxVR7u4yBL2LN1cQQcaR
B9egDPqYgsPHvNgHhol9ZgdWr2Q94cm2xw5IMo9lduPbjBUtk4Y1/5ndVJgIDWuTKCxbHbVO1nvY
t934SyWxuw3FIGghN27/3NcRWxsjhDGXDoXfCDkxyZa8P2swU+cMbScVtfbhtguSsT+bF5PHw5NE
ubv2lNnSqJqB0Rf+VM2/o/br9SscXm2plFncxX7w6+XvpshiOx570ruIiwTgTZYzXKySj7X6Astl
q2CrGTZm2sOTFDO44cCaand/O57HEhNX1TEWTxT55DsXWR/ltTN8Ekm9J8kaC0Iug5QIN14hvsBM
mnIkgkIcfDG4htC9CXZwERoXNtNizzMzlLj4Av+BttOrp0qNwoer5HqOBbswky6nH9I7KhLlK8d4
+OldDi3LZJFCy8EaHzbmEhNnAOafuNS6ra7O1WGGjj/n15tlBEv7+ePCEexhLbi5lC7rUTXSqY5e
cW2j9pbFHZ1MHoXner2qB93sDZisqW/FNDHFs/m5eZiWvSEjfu0KPkaVSLJeo81kqgctjPBQeR5H
d3sQ0akPEoqhHaS62kdxGj6Xs4AvASDgXmLlCWwbTh/A/sJDI9Ysl7b64NsHdRkOUs+Ayfej0yA7
fQxohhUWn8px2RlDIKn3Wx5plCjAFR/Z/vGKv9ZAd5Yy3o+UwulCvZCvoqlUGS9JaB/dpAeY73HV
CAhrS8vY+M0abvlxhTkQBNN5CKmSp3qLmRdvQXuFZWqYlHa/WcK4t9sf5mYkhyhfSbafU5r4VjWq
dNLGQVgAco4p0upT1M5k0uOocqgSc0MXaXKyf34VOs5rwb+bD7UcoWa2zg4C/XTFLeE6MZRkqJcS
bJ/XULlsBUi+82uISX3tTnBTscSzD1Vl+LJs5L86ijLkyWlYVkVnTWdloQ86qBE70QbyppVSQeVZ
alp0DDHfNGwe8PvJ5pov4s+SDk/fcHYyn7ePggYzobcZHpK6WE9fCObUsMk1re9w4XWzLpzLxmux
0Jlr5TkK9K2v7vG+KII2WFYH/jKJOnWoIsRTHjoNc74hDetjSDtmjOL7FewWZgSORfy4sb36/NWm
XeyLdGCCw6/K3sA6Ot0OnSAgwVVjoGFIGBdNXfkXkCDCvBDucvmvMMWeS5YHZaJSJhWhf+7p4hC/
j647FQOvc9qzfdgE+5DTJ98MBMlyeTs2M8nvt950SRXZWby4nKI3BjUAqSrDRV1c8Ea1K1QUZN3l
PfVOC506MclDfT3L7H8LvearliVLcGMQ/LOB0WRkeWmuR9ZkBHGFYE0ighsoYvkb84NuzaVTn75a
hzbxXAWFLLF8ErwMADUKZTMqKAHWrkSzwJJp5XANy6vh8kfiFK3jBqmHNkrDzCIoguBRm8L0S8z6
C0IeYlRc1bqJR+pN06O+TP271xr82LXXmop0gu1fo55tu2Y0WWjrEtKYAhwfBT9Dmk0a6qw28w7t
kJeI9wUo5ddBBxDOQ4RFpro9gne3rZ9Ee12/cpfyvnUvJUR49g3DVcmVjRND8SIFDDKmBQDYY2s1
ey7Cwxs5VAceDpvrgamF7DjujzyWqU9t6GM1uefxK8H1vzzhdFoDMJo4TmToE5r/oIutypvSg8Ne
NRNQfI2+SsbAitgPGX83JD1x8Edp7D0OeLuwQ9xQaVG5zSamJuoAwqZvAnJM1hncbLR8uAPf5Ct6
xGNFRdG/84r6gdlnvki1+zMhgn1sGftay9/3VzBcI+d84Kcq1OXWW4ucq8GQVb8zktSh2S5v5GgX
PausZIXweVRWrV76Mzp5lyIEoZJctocjnqTH5TxWYUPhFWTAD+WW0JxxsaRMBMQ4aIp8te9GdzWR
2zJTI1nZ7yhRrVkZzFQVlk6Di4DLnFPCrB1zLeKbYzAZHGQRR95EehYAmdUEyLlNNlNqzPpxn0Wb
jCo/q1lY9l5OHuWGluNkCD4BBaMEbaYEYJ3iJyOhzhrzA7+IJ0iDop2Fwb3Wb7sGYm+BH2GWVbq2
MRbBK9jUPh+7Q/+Tg1ObuYw438MBOBGGh5noD/HhNfph00o9uqGmBYYkwvdG+J/Ht20DFIk9p4nR
uFc0eVEYkAvCzNZmSoquufd7bwyXw61SO71nx0SPETo5skdiPXE6P/6kBDtsx99Y3g+cGkZseCIR
yZEwebAuDr5U3+PqnJm0NCa8KeYz5a86XuTvv0R5V1d4NxUs/ZwiJpnO8GnQMeBeUYfLYjbqOUpY
gmuvvdC5FopCej6fofjAtPVGBM1AMr/5fapVP9HtuMXHPGOc3l7Y+OhYriROfIlyFec9hF6ULl4f
svuQ4SJaFpMPAMkg139QCw/nrjMvjW0WxRM1c/rCwAh1km5QcqaHuWQkIczmxbt1bDbC9VLFXM1I
dpSk2Y74Lahz3MKduhXP32E1B3C9u1HyyYHg6UWssyR5hWsNb6PtwWtpWJm5sQK9hTncnm4WPXVl
TgXBllPGOq9W6OWdUCDmWqtjq62n86lLmXeeUYVspNf1BC0Bl5cBEH71DyB21NjNAA1J3iRi3+hg
/TNH+EQ/eLopZlhcI6z662CfA1n79BlR5BEKOHZP35T8lX+NQEywxmN7f+jn3d0k4qCX9olE6c0p
ehjDu36n9nGwWZ+Ti3In25h3Vm2oPlOpmIhBj+Yxz4u4qSqssVdNxi1H0i/egdMfOcxbID8A+T4O
McYa0Yfh8o7DRnj8RdhTRBwNETz2vmzlMd7ILE0zYB8POhi1PvBwQ9AMERvPquT33rJ9r4mfSVIJ
egHlpH256jnwLBWe9TRb6lli7jyh4wkQDXkDna4+2DMgqzE8SY8PfQ/gCYqa1ecR8zTfH/ZCV8M1
Nh05n/CD1Vk2QovjtMyKUtx+18nflNeusrGkh8bzalN0ExWWll1h23I/v8kF5O6RMHyA+NiyyUhG
Wa2valEMbyczvtPXhJXdQMKGcesvnHEXUEr1rbp0KfQOfe411V4ZdvpMXeIZBLHHCgPHy2uXIkCU
4ruLxoPfeGmXuyZ/k46DxIUahxUaG/a78v4Mbf0x9dSr23K6XDj238AUDB/C7e6LMMJ94y8UX2jx
m1JQ4OHHc9rU1o0xYMXvjWll8+LzpW4b1Ywbylgt1RobgHB3ghJZ2OCSIvlXNdgZxuGloPBEaXFH
rE/7TEqXgUOOaUaW842aGm0RaNa9cCXj5PK3EjE+uTVWKqCocwCJwBBqFpZ0PlLvxvKpfdqPNqiA
LhObqzS1t52BMzWQtB2SGI2+CNayV6h0rqIXr+5k99lWt02WTLq/a9phEksv+Fb0iFiCv+A6v4I2
sfWXN+cuZuDpCF//fzXEK84VqMIoSKuZavbxmVhOSgpX8i45OboK731mB9HwLgb5q4MmnRoN/nXh
UgH0Xy06TN/ypOD4OzoyZJTZD08/K5mQs/7a3R1gXLIecF3oMP6fUz+dLnjWNLu/Nj9PV8VGv/Op
hmDjAPWh9zlvXKs7hGB2pRqdHb3DO3QPoT2g4bavEumLiyaGePBnjGaPNP5uzw0pq6EkFZ3TX49i
MrN9qbctHvKzaw0BwOwrT0cKMCaodmWcdoxuwe/HXAUAXuIVE3sxn38MV8rzWKBtW9KJteP0SelW
C8Yp2llrZWPR1drENupvRMlRlUaQhuxkF4AsqyLsGIlPexXhBYa2JzE/2zNRLKqnBze+hQ5JUKGc
DJxIcJlf6jE1alWDkHkOAdfWwpvt6btUdAumhzqh5V2w2/6RdkcJrKRvITgvGEGcCtX7X3+2QLRj
xBwX6kFDNfOT4vAXK6VVYwbRGerprcpmUpHawMcW9p8gvcRWzzKrFENXlxw3hlAjqs+bPVRAVL1Q
IvxpcGYJxLTcaDvyqOcNeBGWpvJi+lEqLqrhk1bWobrrW3gAfZV0V4Xq5Ahp+IENRpQTRHntL8ZM
YddU5CTAU0eqO8E67mwBAXrilsN/t9KbikeWCHD+rXQySwsTtiK1AAAbDt43rDaHtLfXrwD2JMjB
zs9Cn5XANU3Im1jtpE6O2lp7HLjrOQDXWmIBVMdNwiH2V/KgIP1F1RvoptJMTP0k0Aqt4xcKmQD/
9TbVon5Mz8jTZzdugIZ35WCHbvFhsPQU+jK4EV2J5YZahrfWoGO+jc9SxBCwAG0XH6nkKxdQzU3k
bmD5pmFbAl7FNGiaRJyhuvXdwqx6BSIzXU9C3IlHxflZfwwyhcOf0ZfAL2PtfSToHMYHGHBPvvwr
zTvck4/nLyKdU9J3K3rXsKlTS6Ex+kasQw92t4zC8HRilcfy07RhdZVFw/c6DkDM/u8ixoY3Nt2H
H8QdiRtiBeE0RROskqlm5tP/Y84pBI9d7BO/0kyYiujl60nXJ1B3k43aHo9agZkJxqWpyt3ICtUS
0dBCmlyo+2PER7Q/l4h3eh7IBUxysINVPNYS3jkStMnEsnXs51HpzQRHjhCOILO3OII9unbevaRS
Ukr597AW6TPtn1txVi4TENW7UcbUykuOdnqKlmSLFcecm1gX0JPCfvYfIuZlCAPivXBe4EEgiPHR
P2FkqkLhjq6xjgbaSuPx4pEGgzFFVohii5a3Q4Og1jZlYwf28s9+rrBzyDq9970NcbPv5PDgs4e6
ZvtRhSNSe7Nfa4rFBcRUyE8mLtJTbBplSnzPruOdfVs8KDDpLGaT+ncoA+HT+kOiRlBEl+Y0S1pe
+sZhsQNAAMBji1IcTLXu2NvWM+IadnCltTHKwVSPHv7OLVIb0PaVsgOuexT7TN+NFmRiydN94z4D
5f5BvraZzblKHsiiNvgHO6Q9OZoFqGEjjRlMJf/Wqo08j+3NHJINwF1d1OzXf9pLafdZh8JjnB3X
exjvgDYghzkG0rVDSac986b6WMI+M9TnmFh+rOKHORlCTFpJG5+BZuEcsYSBiNz8KAk8GsdeEeWc
gORjAf8GtP/8UNIlGF/vnkTYqmuRpY9gcGQGkK2zM+Nt2L+X+IYMvFGrdiC9U79YIgDT9bfyfKEK
ay8EcTCA9bueD/0CNi3/GGSUl03s2V640T+PRS7LOYfuNo9HNYbwvkEkB8prycI9eqXji54CUYMo
ncd7NIYf+fediTyALDpJhOfHqFKF5qaRUYMPNYu0BHZMsHw9Lc/7gVIuAn4wIdG3W5R33r3CVffx
YhEQTRhZweMgKr8XHvgxGenW50cGZ3lIIRxlovV2tk09bol19O8r7llFShn8ae7INIZz96YTyKA+
W4uRFQsr8Xl9a1g5XQrbVNwk7+GfC9ro3MZBSNiuseoRAnBofpO+EZsCGRZuLYzFzFzhhIDs8TeN
wFxccErhMB+EMejqHG28Zc/QHOBD0ug+5gyrBC+F3QUNTDLau7oIsewxoqRkIt/+TloY9FwNyvdo
Kc+n6wLKCW+NlcWTAhTuxNGQsBJJuiudXwz/f0zimMGd6GXaC0vBY398PfB7RkyIHGpOYaVRm57+
y9w7o751C6wXbdg+pwXcyuTNe+lw3CBbpRW+U4u9Lz56ncGuk0nKO1lIdznPUlDwU0Bfq+nrVro8
yndA1eiHAVNLfCIA8+2YWlraGC8/Ev9PV4ejk83UJPFCI66Tnaadt9pnAKw3kiZhNfMj/KKxIJBn
QHsHSkeTJgunoq+pmzYXuuBYqBf8X9ElSNMcdlMr5ke9y7yRll6rIJjxJjDRTY1T2XXa8057C7FZ
ZCcFyMvJExrVi4PYQpVGU+8mOH4NT4p+zsOJPpFHdi044r3rA4959QfQYyfHdmffEXd4fpsTovlz
2KOTo9eyvBt/Pp1vO2CCZl/sT5FSYyPCE4EDkVCRqxSzN2Ka8J++ZCEKY5CtlhoR1V2CmlKSGpE3
kP2826//yYmbESA2i7IwsRIfpN65fsp1SlModYUAPVkLnOM67cqNpiw68nv46piHiXtc4sTBnD7n
B07GEAnydfQVPiQH3QBsw3m82jrY4zYbPqtNAcu80g/2ukOrSY4UoQG2+mb3QRZmod5XWm5gu13e
gyCLbtMSs3nKFOCwGS9sM/YzD9p5atRo0bTtkcE27mXZa81UqKiqju6atxmzMEJVNiAqfXF+4mDM
eoUxiEo08jmllkJuGS2cSTsV47tNAxvtNzWTs7nKzk+4RZgFAe21wPQWz3qrzzIXyTGDqfMk+IIo
lhM6pugIWpv5GJrRKMzhYBFVDX7Ya4+g6QXO0ObJifKqvBrVVIxGKQhk3Ha9s6qAjtgZ1lwjZXlG
M4b42gjd1za7iUkVsdyfPchbmuGw7aOKI4E094CMDjuLmhmH3A5zhZ4QcOKJQ7ebIRtvUA0BLrO6
rm/DVx6PRJA1FkLLQVxHYQTnTrVJ75TKdVEhirtQ8njfKWtIJVZ/L4eWY1mYFhO4+qTvtE3sKc95
8mQOAEzjQ+l3zKp2QlxQu2LrpcYwlLH5P8op2APWUKzAu2lBAcIXh8xZIHeV3vLpeuhZVgS3UBqi
ga1cWl+OJI9MiIKx9DHgGzkOfG/xL05QyotBPcYSbgAkt4Oi5fp0v3H6Jb2EgoA3Jb5MOi/CoDWs
tlG6qYUXAKYEWKrODuIYdjYN6j6n9/1+SBk6LrPChAmoVK/WWGel/WtRe+jE48lOedvFCYzdeo1n
xhwSq2qOCV5dWy+hTf80yufTA4A5gNvBHXJe0DExJWv+1Wbx1ZxzVv6FkWTFJDnjnCBIPpKY5uBw
Oig5q9kZo21U12K8AnYMC6fnVpF19jo1vcM8gDRok8MQ18fj4TCTN4h7DA6JcGsNS32OkdBa678k
BKRhOd8+pSvfkqxK+CX4J9r6ePDVLXk4cOroDohP6P8VCDqfSqLeC39MTM8AQQjkoHqyh5bDsMgN
t2jtozkEGbBeQBGF9NetlkJjA4LFe9jBQ9TXD5ubuoiOSonbWlzUGABraMvgKKBVypEW8Z81UyAv
mjBoSopcUEVyEpAJkDIBgZhUodYHjcUOVaoderaC9NVLjv/QVo+sZEQB9DYZat03efsNMYILaRQy
65stXFrpbGKpB8ASjwmfH2Ik713qXQ/A0hjSZflgAu3GZv83IvyNRqWUA499WdiMV/MX+48lFRO2
BSMH6JOpvpVeRzfxu8xJp82aV1b9YAxLiewVnJO7ddP5P2a3kAz/AcCcOkFMkUZdHLtp/OgeC45l
6lM+kA2qrJqJwd7g/UJm4s8Dwmg8vUVpRVROaw0VrUM2YizIO/x0n28iHAev/kQT18q135nxaq/5
pk82l56SPP8Fwi49j+HEAnWzJtObzykqjOsKOlN9jFTO7XW8SkezkeY4LGPdRy6MHVKj5/rsn6Tf
6CHDE06cft/FtKUXBaf+UMX8T1TevJHttBfRVQLQxErSjU+Jhq056deKo5o504ZPI52nbZhBMKvS
yNxJgZgc0iDnMMRhV2DX08wLMuu1Di1q21fEzhWENWCGMrcZLC0E2ziHzBfQo5xVjruJsUZlkpzi
UyNG2GHAi0Q5J9TQA8frDI0am8l0x9az1GUTwZOSnThPLvG7bEvDN2hy35K1qc4ewDuIhJe0UeAr
O6/Rnuv7tSMGFXeHEqY0YOx57hIS1SqrKfYoqkPP6eGp8vYKlMQiyfqhHYfOM1RJp8HbqOgkPwHi
IpGI3iDdJDncZSaWUp3ehKTpRBk4hr8Ba/Ws/AsQtNMopknwotCxKazmGW87FFGX//WIF5LXeaQe
4Bw/zgXJ9vgpq38oQJc7JAnbLbxIFSBzPHf4DdOTy0G7yCBYMpQNYoWpwDGudnXmBXLJJuJQ4LKL
/2m2e3wZPsDPpUj6c0Yi6VywNS6RlwmlLVBMi8zqDjpQLMSZRAPVyBRZCyek9Ebh4B2wCuR5NCI5
vyfjc/xuUfPY6q7gV68bQFCZs5QM04qT6hnBQjXXx57g5IaCHrCURSKRgP0yNFuTNAokmKlKLTZz
4w9EkbUIuQCCXaDeLmZy2VGbxH4UYd03m9YsIrbULfCW3Qy8895quMeLdG1bnA3UtcGv9xPp+iXO
D8FoMDtZ6d7aINFd/KHDZXjGJ2Mu+OBvww/2MdARzcSii3eoWQ51U2K2GVaW1IgNzJE6Q9btrWl9
XsbvhWWM/x1eaT55oVfeNjdbONBBc4sRXZ4AvnMLqKthQqGqLNAEK4EWhvg8XVkHg3XOERHAHIge
SYXb71V214QmfXL/tCjaArsv0QryFhBusfdrR+RpcDp2acJc/HIAfU274LTD/0pYpNeZlw+TqIyA
EfdQGCsjfX9hb7n9JqIXUxNkmopfMeJ1ssRiUZP/pSrevXP2vfeqmagh7JI2sbCc3dRyVbOsbBC7
XB77Tl55LlZ8gBxycrUnadSsn4vg5PRPSsxvvdkuYQXjz3M1MejHSeM6pjMZlPeyEXozy7M6cyXZ
LHkM7387pk4r+mnSORVdr/bAAsHKDYS5rZr0VCo+8q1a4k9IbRZICv998PYkAfeT/hWpXn64cCrB
Wt1GfQQKeubYcMsObLflp+1QKNzItwieo6BL/L/757Dq9SZZEjEQeOq9GV/TaZHydpI1cE2cwYmo
EhZYUUB1S+9BN1evCAnmnp02OskoLheM3820w8OqnkLRtnsAFfokik/VCqrMbWNnqw4XQC9cnzME
he0lQ+fMEvXdgbjLLATslH0B3PZ7hkcLdrKr94btFiWJfwLsqGxQ0DFAAAhRCw0iNR+ePMZey4wA
Q3B7QCbVdVSQ4m3OdMWKhX0vlYlbnde9BsLWXcI1dMIKmvG3p8P+9NSKxm2FCQqnwn9TgJ9bbuIp
4jtRSXMMTUQkFv2fydKhLC2lL8OXLGv1c4X/Hgr65yFvcFW8gFU6+tWIl5ZCKYWUggYWzXWTscD+
p1U5DGvcJAISzmfMJSXTFiYsBuEYolAOBp06LWwPpVbCZYAArWJQzXO2VyCAU5iqQxDLK0wOAxcF
9Ql4AIJ6yx4aez7FFBbVkYzNNqEqoIMpo625QYyeTi9xnOqs+YROo1ivKlN3QWPvJVlyIJbZd4X+
NmGwIY9Hgw2pNt/I0D1k5GR/caRcCSx0sIh/tIaZlGpY5to8Q4z79JaLYI/Z7L4ketrFlQDYMaUW
7isO+oAHTEhcZP4BCmxHLR7NePcm+TDfxyPbaLpzBUMkkd20bY+sxaMtK1SPk2nQ1dUG1QUPdzsv
y1Wr2veCplk/l5V8iga2iLQrEtE3tQW1XVJ09gTa1+9YXTjIglQY2rrjtpZvK2OoyrQD6u3SkG8Q
a6mZFY8R6d9TkAF6fSJprlGRpeqIlJvr0k/2nU9gwzm5UNVEKY20/QYYnCBpbYY6BGUqttQ03UVR
JKH9CH06ParZGwkqRsZ0CfnQNnD1xyza4E4lXr+WjSbWf0q8ex5g4YiZLl8g6rv1iFIph9L9x1GB
DKxSkHFjFXm7zQiKebYW7cR0Ty96G7K+Td8y4uyUe4g0bZw7H5V5JzvXjX5sNYnI27rj+MgcNoH8
27TpQw4s6Du+LWoVF6KMU6q8B4n4MZyk1qTdROZWRYCV1L4Gbkumkza89TOjEs2N/o/oLJ5jviid
RGgswcuMjErtHtoOctyZK8wc266qy5xsfHwG8GmNepS4zQw1wq8QKXFLQJgYtoyKsdjuGl1Twc0W
L5Jh5PZnmMo7uPAS3AlgwxglbLvid8MjzFMUPHq2bLTgbnlJC4Wz0cNxolvFfaYcfh1LlPsBx/7t
7xCHLNXFAiUjiJkcrYacEiYb5zPFZq5dtzIEMUGrqe1JfCBgFabvHMpFtF4InVrHrtpa2lzci372
2R+hQ3iT6dEHkpM+ht08e2gyPPfbmgPogzywRrZugZEUAEhXiPGDue6POIC4nqYhCh4LDRRluQ5g
eX1m+BXBj+dgcB3dGSvIZvDAh3JNAAB5L9TVwyUNF+SKXY3E6ytbVvNqIZl0ERwM/lztBq1+sxiQ
Lcahy8OR/YoucCRk9SDKQICOKrLYN7WpzcQ6HKWIEbxnF2HeVnKyolui0xSI91Mzmz0Bj0YnWOfm
9jfr7e6jv/0nsb8lUKyLys9gxrJIVTMJGLJk2SXKZsUhIbpRV8RisXZ7ccaPoVMYq5v5xT5wm2a5
ijW1yfjLQzYDPNiBpVKxZG+LglbO/KolV3yxiAe1D7T5rjPQhtfRpX/04xnVQ8Rm87Dmiy38fYB3
6rtLM6pRSYp9LWrQuoc0bYzFf10kCOUgsBUQaHUD6jeS2W0S7F4tQDxSyueQ5rUApr/3XSJctpcS
IGVtofjnPoDAJoeSB1WSJ6mzsq0wCsHtD9lay/DZmWd4djfhyLslEHzSxiF17+CGtZMAcRLAgRwS
x3+A+RwPnWwdO6cNbwHvDS0SPOvF27qRpEz09mPW2qTZA2AhiVg6smQzqIyEFt2n31EjKpSy+jjH
V/2rvWMWN4mvmgtPmTLKYb7kqd6rJVxxKQJ4xwweZQ2a8R6r33bJHJsI6c9eMsz60FZevdFo4bdh
fXfDylnQwJqAEDui7A5JbHin8+Lre3nz6pnNDR9N1gITEMc9w3bVxug60Ia1/JtBUnZNGtjncR2f
d/TkrzDVko6BB7CIqUtRR7l07aXR+RFO8cDPZu5FldLegvGg9TM7YGjlYOvTy5Fgvl4r0UrprM3s
927Sm7hSBUxhrXhL2U5qmEnT8q4ejPeJjZaegg6GjYRB5w/b1yrvC6Ix1+K1H9q3GNJ2HiFfVMeE
wq0Dp3QvCxDf9q2F2O+ma5KXd0RC8FJwiIirnzKvCEFKzlSN4nbk3kVAd1AwOBR4oJ6iZaCT4ma3
1cuUQ/MVO/AGvnbL2IUe5aPdHsXvsi2kQNpy6Sudsp3acHuZ2EwV6+KWSaVn5YJTS7OQI1UKejrK
QrBqLJSNx6daltNgHfAxs6IvpA6FgOU0+aJIwIoDTNFar27KIh5tdyzI80nhsthL5i4MSK4r3Oa8
boXz6ZpT6rTILjJn0xhv4XjyAUjrEz4jS9wD9ycn9K9H9Hf53qEgAzJj0jf7D98jFhQ2KmIyBrGM
89l+lLNDc8GG7YaMM84tVvFo98N/zGxxGgPeCTM71zZ/6e0/vkkvv5EX237XbfNdOwSkrrrF4NV2
8jY7ZceP9uGKUAKxNkXRNjkzN5ultHSPdwhpp5xiXTySAw5N/zUyTDj1eR8JfsJJNClGGZOfzGnQ
e2bEz8vJyCn4u2OcJWan+D81A5SM+2f7FP8pmhgkaxbCc6Bh0SSQLYTOLnhRD4pahKHOJj/mysMv
cIN2bFLwVPqlOFeq8DxOWtv8Pd6y9Ey65/g0c07BDdz2MCHTRg7BSrGYhPkM1Fx6g5LjoRe4Qmxv
r1ge2W+e+w2NNUPIRszEqbvVqcyVxFV7hK9BrODvc9f/3Zh09dY66yFJNsn2IuRekAWvAZKsZb+b
gV4oYoANMzPhmb18vFCCmMGNmmPc+tfBInk1exRR4rrasQgFjeaoofSGSmSoZd5+SyQBtJDgxRcb
KJtb+im6IlxgoqRRWugS2/VCcUNqYqQWKADd/Cml5pz6b5qTsvKh8EZV1Igh64Zo5k68XXeJFVkN
CGjLrfyk55e1LN1I6rJukkuw9+usGpg9XnGh2aEpf87Knfg71Fedx8xRiI1+wUFpjfJ/ViiyHfLh
OGlyFbbtUJD0nlIDtANKaQIYvjDpqwBldvZLjaGkYWuabVBcYzJAPtrt+7KU/WOGQErUW+2iP3Pt
2hrUivuQg4p6JLutW7Wh1VZyJF5/NtWANCu3tKr1/NvTZdidFjEXSBx18q9nk6iv5FYPgKUqQaJd
dVNspUuJ+Q6p7wGgKsauUDlOebFKHk51NPk8Ng/myIOmlLjGslyZsflKB07wMNEsGk1bUeR6oQTD
U0HkUhKX/ZzOr09hzY/jxtb+NWeEtx6SiJatkEf+76tsVmUkC/QniNhK49DFFtWIxRzwZiWX8Bgv
TNkCuTB0I/a7UZPXaMsyE4R593K3NOYgv8yccFnGsZ4OZI+rWakovI30CymoHtBb920ttzNhSdib
L3ekb4+7eYsPrcJQYfZhC49lw6K433I4JC+KtZZGQDY1JqPB2+c/unHh1QCUdfA7l0MU1vhaG2eC
eQ8Bb/ZUgkiiPjkWM9RsJWHSM8wi8WEMqXOJm/rszECzaONjOEqdUdMuHYQBE7ljJTTZ5v0ekaSv
yXqGMhLgeUv6sm6cF19MI2oMnzIy33UgDwuwR2j7OlqoE4ofkM7MWAHnmOd6/KUEvKXs1wYrNc2q
Ts1sDh4sN077PNWHCgXawtiT4jW7plOC078tXe9HRQUFou5H+4u4tSsJShSsAMFSzswyMWY2EKbK
mgT/Cq1W9CC7rA/iTeRQrTCEd9/r1Px4KOWtrfI0g017m7Tl7eQTGCYUAJ9ZrgXVeDloojp8VYqj
qpBMh8N5kr/yC6P/DBUW3JAiTX5QxZsmFr20kNkaDbf3fkj4R0dQdBiXSaBgFhdd2TOW4OpVUo+8
8TR3SiUkqQjWp9uAMi6pFLptY40sVdw5qgd0tOchatLKjq/IOrUW0zg+dm7aiBSJz7smU81rIs2U
m1M7u3PUExNxhEdgUFqpmsnDvlLUcECb7CYgHaRwpnyB/LRIQv3y7H17uHFPY8ftGlaVjmiYwSiz
09Gcgt7MTFd8cA3Vng0X2d0Nhmg0tLtQSZ4ohxcpn3Mq51NANup1lXR0bEhCE1vwmbRqle2hTBui
CrstJtIU/3Ol65KXFfTnHm8iElzz2vReD9HNm0EXovWtZHFZaDf9OXKAP/7tBQ3mozQoVIwHaVAc
BTnwdV9UbTDq+6eKRqozjofqlxqPuwycU7m8L23xnWVWN/ZBOxoOCQmormXC4lkdu5VcqfEfJT19
lPHdHh0Hnzf8rN7I8IwBcuJFCziWYxi/j5G7TQxyNqjnb+GsGUb04aHDVEmixWKQzorpi0dcX8Ld
NZH7SnYHRWbcyveOHs9Q70TYZ9MpQo7qjLUVpppCTL34Gs5ZV4dU0sIip15AQOahnjWJwrRmDNot
Lq4e6MiOO/WvEaE+xsrtdpM/+vymZ4+hKfSqjZzmZvDYzud5NcqY7V4td8GTZHJ4PfA1uAiYrqcs
QdkSc5jiQef8+eCO/2kbXLQy6RsJZ5VCmvY57tC93K/JNvy0TijQCnYgKNBQRZ6TP9U43ahA1Bgc
GXEPJy479tsrN4MC+rczNW0cXnhwHZCMKWMGk/0lFv5BqtRX+AnDqOcNPWi0CPYmoMY/AgIASf5c
pNfVP3s0H3QfSOr57zPL5P7AtA4UnEIpxsxWLAZHS+70/5D155DCpb4Pe6863tE4KPBB2G+13DUC
dZbb1yQDh77sO4FqqeewxhCe2G+NVGy5x2Ibm+UKbhQssUlpjpEnGfrrCZcCizn3UZHHiumfIk5s
b0zGly+poAGDOuJakZBO40MjPyRoFU9l1SiGajawFnvc4XGcuAq9QDsPYw3N5zm0m59TNGydw/8A
I0uXmcXItN+q08XtkkX4bWZs5TGCQ9OpLlw0zmpypCHBlnBadf0hoqJJXkyQJePEaACrDs4fdDCj
AROIGGorQrFWYPuz68jHBqBYMoqX00wGEwghCiwMFlrrPy0sxMOJzQ5qYOj6O8OYmL2mTOIeH0u3
qNhWstPYjaH6p3d1hblG1mcW0ErAPbgdnEaI02rVUtikmSl6kKBY6j/PMNlH8U8EwM16Skg/Q5I1
YxRjfukIm7oZYuij8Nps4LPm7eG8SlqBpBRgnIpevRGo5/PX++sntLODjSVQDDBsaGkB9T+sPVPj
U/37L89aXnIxHKTrc6XPeWPbPyo/7Gvp+mK6pLNXCDukZODVXx6vQvaeBch1xbakv4RjPMbVgX2h
qfLGNbz/QwF0YZYRXsS+eC5snuQG/6qLOVjSdapi1UHcfEy4zA5lfjJkGRg+zYhdqCDy1tgGizO4
fsTlZPi772lcoSV2JLlElw57cIlPQwzDxjQxQjqzAXUDKjT4b9V8yYwe1TvEUnsFvP3lCeb1OicY
r4q9nnSHCffxgaPF7re0slICWXy3wgoXfgYPsqoExdP9QXRcTiMXJJsL5lEJTeyGklZrvym2gstK
29IvDsttq8Rl7rHpH5OsyyKBqJSjbTE8EtTNTW1u8G2VSml/hKxEd4W0MEmXbNOSvdjIC5Fp19zU
8vaUiKxQxuoseFLGA5vtKuMpUfbryoW48G+Uk0G+CXwoImhesBGBMBh6XtKIuCVV4zBcZ9j2OMm4
8qtuAbirqwJxuzUnFlNSvTnQw93MmPYl4ZeF+AOoi3PHdS3zsRncGzJtL56ro+4BaWozbXDZcMYG
yuzQ7x0OsMv7RFi5Sa0h1cst5tg9rzdjMNauuNlwqMqm38zrK1JTEP6J3GE9MGr7AZcS2+DWO021
fDwsfedoc1vCt2ahHo9FaI/BuiQTlc4YEQ3TQywuGz15qGzWmPTczZQY30w+V+Rq58gQkkinajal
KgZCAAyis/l0lI7Kk5FA76uW/eY3CS+lf85w7xLplr2VLuFnYaMirdI0hTYtQ5UGiZLr6VWyxSn6
VFsahUeyjkco169tlREUuiaWje4olf5P2c1pDLHNlSxqAVPefe3gTnEQM9zq/swDhAMX2c/3qKRG
3fiKD53jiH42OkocOlsK27UPuUGUieejNbbzRD/fmJ0VF+V0Hvk3YlxCbVIq+6GkZx4Gmu6MFilx
j98R0ZK4fekF6KlYF26Jf017I/h3q8/MYjtrhWGKODI0suLIy9a2OZheu/+t20UobEBF3XXE38LW
sZ1hG2NeNCMIZluhjLdYB589HOiV0DL6B78LJm7bQhYJ+edoL1J9m4EfG0iqSeZj0Kk+ccDrJRjs
DzQ2Q1cxEAoAWrauQGJyaVt4Q9DEUSxRSCuP6gNWC/qTis8yelveo/j4VZvVJVIdsLq0+eD7U4QT
NWEyIt/ISzy/ysqZhUDGYBRRkTuojhXj6SNTprji4ZM5hEcGLYN5tR1+U1a+kKjtPt26XmRYmGBp
3gmE+vytwCiq28b4FiNWdGxeWvYadRtqoxsS9Gh4uFfTXSjuZ85GzzxGqcuvF3gdKhdczlHkNYaH
zORLS3NIJwW2VkBoMTOVorbAO6eSVpvzKLTMxrb1Q38mtYDz+fr4sQlifgA00RLLRI8OLbJjMqd2
x3H5S75bs3S0sn/ysMgb/l/CUkhc0YUYMCC0PgJ1VUuLLuB7XzWxgtuI1L6TmlUhsKOr57YFspmI
ZuDw5eSbcZ46h61fjQnA5H1paVomuxC4TgjBqlE27QDgyvzCBwonEezysVD9w26scbHtlNkwHoRk
olLpHSWfh7gPoVf9siGr3FMM95RYfJrzJMsEFlFNRUTGGjPQGG42br9TuRa/zAmPvFfOOFClX+GB
mQBILMhdH/zY1JL8zz+V/bJhSGkFat4r92A7NDaiTVA9rZl7euHVec6wCawlQX9TwWb1Ivh4EuB4
bH0dKzfa6bmRMIED/UVW5nGmIc3zjfFf8fMWAQ4D/rG5Lvfe+UWBcznycTxa6A11oT6DqXj8NL0g
Y6pAZKnSG0TI2Z5BlrEhB0Z6Pd7EKDsnalY9FWP0n6PAfOukcsigWtbIwAjSrEKroIDJ2mLLyFcZ
NOBENO2Gxb9dBBT0U5iM3XWuaNI43mDN9sLbz6vRP7l5jVUW4PLBbCSXOf/Lu98sJEdsa+jx0joI
a4QM0rjx/jGDZYc41vur0ViXcAxNXGXfRwcYZkRPR/GmGkRI4MQzwbK36tZx4yWrAwuHaegtaFhC
9z8Rl26lXgbVNHICWEbT3MqK5ct/YP7imtY8BBpmXmoaxRLvo9dyAQuIN+058dAjBsgsOUO4+cFj
CYw+dYK5XnhR7glVFqjRiGks4NEQEvVg34BM8giit8zC/Vlk0Dji6dkMgjy/noYXAENPDotrWWkT
a2vCbr2i5s1D0BDoUicJ91Tm63oERIPqMBSW2KJfSo/N9wf2KUXLzZDIsq6oTjcGqEyMdIq5pFZo
Brce6rFP0XIQpw+9dSIEWHJijHA1CWweRwloAqBJ2rzjIOwbInthQAbCPLJsiQquSxtXx0w9OEMe
O64sODFT8UUH7pp8y1Axgst68+44Kg+k9yQLzxYcF5r2WWcJ5TQwCprDvy9ZHzKhEGXSdoBg6ImE
uDK/l8o85kRWNwifENwBflzy2ug6N8Bgj4sD8ytQbIUdS+H2lpd4O+gGbpUkMgUpBr2kv8LYQeNT
Imn6OkyJDV/e/4bAE35yLp8v6Y0G/ud9vxXPC9kLHkeOQTY7Tf7pCEvhVUvcfR+iUduYfzUCK4SF
rX/GRL5GfvsSJrrsozrwczkispMfq3W1Qg0DNyHqE1XSRUpBq/CHJr1Nu3rKbTHD/mmYc6UUg5PB
9YsrApyQcD/d95O+AflgsbH27VeQc7GqhwXarXM2z8Ua/6Jj4cv+gStyVC/Ao65+QHgjPHODzIhJ
Inh7ZhAhrsVU9fl338NN4REv6+5JKLO/o6gq5F3i2kwbS0O5Ty8IOjn+d21Qt7Kiz+pN7qDQ3X4a
F3ih1X+5ygEzdYXYZi3T1RZQNH4fqesYqoRIS11WsR5S4/fVgs2zovPeq7YqF8+pDTqRaLrzdMMb
VAJokI0OuXfr/h2K7xz4jRqUnCuFJxrovjf51iqndI9oUAPtZgq6uMPvPtUh4e0Im30zuOjaCrc6
az7dYN8nPQN/Df2H4G5lGPiY/AlMuBVbqNmD4FGBR3bNLIURud+c7cUmBycFDbxw2pLNwHzp0NMz
c/h3gjqin5GwdqKMhYKp+Jr32b4p1FhEfRXiUR3wHY2BWbRPPId3g7Y3QAqqs5qwGYyYODupy/Rv
Tkzyy6QNbfbcKQMNrBFDh7dstZR+PfbMb/XSrOYk6yiBragHO2Xg6JcmOBXT2oqfdRe9u5Lq5HwS
AqSKaYJvfA3/mW6lT0vJMoFPKRtJvdwvZ8Zw2avUJ0cOrnr9UINMGWW0KWmmpW8d7F5CXQyOUJL1
Z+MPyhqout/yOYT4LFTuFae+8i18Hd+d28xGv+zqOy0m4j+WwsbgBa/EvxKfCZSOBuRqsrN2psDB
xlu5fGCPB8fp/OJYynmsx+ksKZYGRGjqf13os/Schzs1mF5sG4FhLuGSvgxGB8f1ykJi1bpzzozQ
6cHiZ3HIuXkp2DTD7L6x70xp49qFQ+a/lVZEZ6Yc8r/chvxmn8KgIalQF7wXJfWvygQhI5Qxz4dT
FykXQ1CluOcIBZCktp/k39NR7jpW6WhU9BqqZaZD/cxn6Vy6PBA+bSP2D3QX0gGY0uyfsApw9Ljq
2mPW4OOtBwhPHFV9O5PvsUdIdZidw5oZ4mZ84yDJoH+IgMkyrIS6qky3Lc4TtAQ9ggm88hEOhOfE
y8hAUnmRiSfaAzVm5QPXXRcIn1KivtSdcXpVMmPE85lastA+ITP/PLPW2vjDzxDDIjrPiEcWuehB
/ck+rRfqkbZQSYy9aqJxGb+8fEUZ9yhn4/u2oYaj4Go1mTJvw1AYpLxGm8T0Df0RhYxKB4zDG43i
L7XuC4/nRQ4Ww4Ba0nnwSCYpF13z5MvoLNglEccZR78rphxPPXnSro2ZGmF8vXdfmAuUKXzc73tb
GQBrLvfoBgKYEB+/uqZt/s+kCZ9EZrxjilomxltxuMgUHq/f2WdWGsKYdUO20T7VOuyOz8bYVa6D
F930MukJicG45vHT1s+19xVL8cnBTnBSymM6qLt0MPjLbWS/AY+IRDmf1nldxJXafYcbuCe5CgLG
e4N+37R2mIHj7ysNzk6zqJSd7ZgJ8whotNF/hfxe+aB3W782Xe2o1Eqtc2GfG9cuhe5m5Rp0VCyG
la19NbF4f4Kk8VIOtQbv2zi+/AMkOJ2azjBQA7BFvyx0rqkBhZutsW4Jk0dkCR6XWTLpwzbcda38
11WmBQLqU/aOUmDJs/0k/GggK9wYvDFyykYpU1Cpw0Da1f+nBoD+qNpZyZ4BZUYiiRGriNdgj0wB
Roy/UuNTcd0HXZ9lsNK7j3kVx7UFr9gDpVNXO0GF0wIOdQFEW3C1a23PGCxl9yd/hhE44fzFitDS
dmuBOHLAFgx40e7Jf6a0B4krssjcGQ1yq5Q4jSkO1xF99thWCMwJWNUSLFYOkUc2wlu9RKa/81Hy
wjWpHWYzrJojcGoeATYG27DOeryoakyVE+xzi+wpAl3mq0sw1zVTXMT4umSwTyIZ8FuZJCzKHbs2
lAsZwANPTwu2F0PNKmyXQTutzGnEfpmZoHUgAnn5ujAZ2P5yI7T0cKl3u5GvtYcudoWwjW+RCIZh
eglEXIC6Gxpycbn6Bfh8Op5Eo3navYi3WcfgFwzf8kxm94uzCB35BH/ptb7PLt85Jo7vA2tlo04P
+ExoufKrK4z+7NZ2C8musj5BtOIaB9lcnV1GCSyfmQ3kiJPDU4FBfALJD2GH0woXEiJsxEij5X0H
aUfOVfrGkO0EvQwxo+nFVbE7ccN+ibw+ozQOAVs9JWsviVrsQcVHDMhtP0H0d3o09cw4WexK1ilQ
uxEDAAncqU7W85l7Vifbjb6HJ6QiLe3I7RlgYTOmJ4MmbA4CgXzn6RQPmZ+lU5pln5obUJXvT9SI
UFBOp3AbUkvlpxyC+aXUYzUNZ+wTKqbwLxq+ud0sdMjEiufOIYNyEtdHgA7MXpFb7WS7Yp3kidG7
37IkydzUniCqu54eEFjUwAFUjH3gw1ryQZzotuGiDyuEsK48peBCXVpFCovYih9mL08Vm15DoaXC
0eczhjRBlEMgY6swwTp8mv1++XC4pirZ596hYsx1Zuh8YE9kpNvIxw20mhrMb/4LZRtLo20igFwl
/74NKInEQ+z0Yfwd8np6uQgmk4BDOjhGLp8HzWRXxfFB0eTV8JQf0hcC2jKbfJm7OAeftXRuGjMo
U4ffiOORV3HA3+KCRmFijLw1O1Gcznlb0qc0nC6WKAgZGG+EJU2ukV9hqMlNdQFYh21nv/tsy+Ov
Bz1iGqRMVCJot+5t0MqQgnAHcxsWAlW/b4a9Q8GvsXQpQO4poq2gjOu1m/o22ewv11eqCPRT//7F
4ZLo4HQ/B6b5s/PX8BCc5x0HZkR9aucak8XZShdoU/7A1QIDb8SZ1RXGc4tVbxupTX+s2mg73r5C
tcN9WCPE65NATGZfiwvMcWG077brVDuIl1qQK6Uppy5UbL6oDt9gLL2vNmV+UFiLJqfsCEnrHiFs
IOb7Oc0ZhX+p26q4HcyvPbhVPV+xDdeZKCm+CS6IOAruZboKA1qpGbatw9o2u/N4tfY6i9w35Hxf
pLbtdAcg8CWRCL29HJ+jjZHa61iwZoI80pvISnedCzW/Y/HR2ioUxLKZhh0UUOmQIZAwHUfNTgJt
Ha3WFjepPDDMNipey6Slc+lTp/yhklf387zw4bWLikNgNfX+NFZ/xNMEQosSbP751KFhxh69whYi
Jj8KFNLWXksrgg8+IskRAQ35dFAVz9NjLhi04fT5fJvGEnCubnYQl9+53Rgw+fXOp5HhhZdrEy+X
QV1T8HByEcexsNWRQYADBY0pCmHzXLnin4G1D+mPcOTBg2ddAVIOJHkHHQOnN3fXXxdZpaYI0vck
K9B5unBIh25hfxa8xXXLgJgYBNEoD08AFFapq7BbFZkCWlXeOK4TgECtp1Wel0X+1dQzpfEQ8qHt
Fa59ZYZXnSVbIkx/0ltZAs2TVPfa+9szhkVItxZlgX8zNfa6T147pRbQ4QqxjBlflAWYAInbjwfO
gP/NaIKMs5+x9e3OBgQEGPyUy/ItRGF6kYWDnUHdj8G2Vrr/oN1VFw+jGyz+Hc+CPCwiMwdwqzJF
B0edGnUrSjuqEWFYj3UKv8hcsTKLAjYdWbPjHlHU2Dfq7JFAQzOeCyNL8NM5mpXAypVy116DUyce
BkoFQLwv8Lkm6vaGKrIXeRdlqfmNEm07zzLmynrSw9PtJT6m4H0DO8QayDm7lxVoR7GxT7HxaPHr
iQg7ErfB00XJx/NfZPW1ocGAOwdn8iVP+tdm+Is/vLd0ppCsWaKe7bbOUJlC2AIaXXNeEJRZGc6R
6uTQuPfBLEGfeCPIjOyB1/nt5/pJeIuhEJ0cSgRSshllMc1Y0/6OJca7/I7edf7rlpeGGZ/Anz8D
yJVc9DcRR7pwwYM1cVHUkXtJIsKlxxH3Qn27ZZdIFNllziCYSLXeH5xGEgqNqnUrdKlJH9qRA9Jd
XttTqAkDAOcmsCFqqj7vOpWqpslE9KPPiUqtmjxGwDCkuExKvluFWi4/X2UM6BfdRJFv6lfONnJs
MN/Wt5sBEz91NG/3cYYQh/pP9VuexXn77cCim7vjrTUdF0IxLHQ0HvjXPMsAiUC9BBf8bvfAol+D
DGjk8mTcdk1Sn0BMI3/sbS3oJgSYnGCSo03r52UXRd1pu7JAKGruAHKPnTDaMPiKU1FBoSFZaT0q
BovauZfMi6RII98koPCgBmhZXGj24g1hIPHm7tzzi56rCeDc4ULUYkL8ifcFf4BItDqHvgc8q5Ql
s8xIKeMWmxUnk/COmohBupS95unvy8nBZbkAAVZ8DzcEoRpFG+SA7+2mIeRtTi0nAfTue65N4k/+
sQRu0Pw4fGYOhcpIDXcxAfjGImOAz2Z1zHTJP5o3vwo8lSo7gDcKrvfLU3F3EQM0xhfhRhI/IFvn
VR0y3HDnxFfz5R9nzJgXVRo4xEsjP3yWBWjM40/K7GvQvkenDG5G6tjIU7znt8mPFspfl2VNkJNQ
qr/sKwFAmvGlfFxbT1DOsJFpVMG6pSbT1XAaPXkQBsvFo05QML3XH5HO4xaKQc+m+ut36XfWd6Ke
cmLGmXXxX3q3DxDA05uj9kzOW6tWOC3rnXu4/5n6InMNeBAuOQu1KiFukYvT/ev7HnwrRLCBvxKK
saify8ePsiNdXvCKZLexVBegtrDUO4WMwq3/ZMmGA+TfBYwjuh1jRL4r6jaMIRxpUsEf84twTarD
dZZjsJ75vQw1c1F8NiYpDqOjDNYJ/KLkVktyeB7NrRaBNRu6uXBYkfAxAHK1mVBQ43zZknezLCRW
xILzhX0Y+4YSsT4nukqmetZtGayKa3532IjLbvbMR7omKJQuTD3RqzLRbRiE7A0u4SngrcQeSiB6
lRMS66e9Igi74oDtOGxMJsFwHyosrHgoi3+eWa+nm8pV1d8xcwMEtmfkPIgzwRSqVxSa8EYwVewH
3eqDBs7emRXOzXwLY6HpHuKd/s5PTn1U+OnPj9MtFo0rSi1ImQagPyopazC+MGv3VL8M0N+EoMOv
/JuUNRgkNqknalfM3JSdCU0MMMsk8woZ/LadxY2lhphsH36YRZAePOqCnmeodo4/SIZyLelJ0c1A
hJq72oMAIHmtqhtkCXGgQ7ECaUQY5II18Ps3QX6OERbldJuFZPxgYokHfAI7RXKJhOAyjrcaf3Am
xdDz93EDtB8bfwIFi5RF3iBOUo/42SbnVCk9CyLrYFx9drCOCsCQuEDqPY608WFlsc82HVmuWF8S
y07cRi5x15dAO0Zg++sjdxObGud8HAnUJNExpiWe+nUq/wcsXVZE+dpXvdJbTYBAS76DCJJQ/3IS
VgwAF1g9lsvq+NwCHg+wcjM0S/I/nPrALpd2HfKyO2l9i20f4YwdOwdtyzEx+Qqk5F7hv9tAO1wr
Jxbcyb+EGXcdzgPotkhnovjs6pSIqbyPSCapxrglZ3U2lcmgli6F7MSCUouN446PBijYyeO4kH5A
paurHTfVTHrWKXzuTlh+rDC4yLJ4s+zrKRSH4Qb7BxQv2ylDaWZycjIbZRwmb6ewBDtJKWHP6e62
M1AS2rPcea3t2HhavuC+r0PvGQ1IMGEIM7eBGnxaGcuks9vCGH6IuIIirbCA1wdhRoXNZKE2tqDk
KxODEEUHxN22lewDN50umpnsLWk16OvG28Yw1fG6uJnWEvlU+INbEOVQeaTOkhGzgBugfLgImkTw
tRBVjQlXQFHqRrqGLn30Uwu2A2ee2ZKieCNcp/OGSeXM++tT9uFS6b1412mqUIS5zG80Z3ToLxzO
uNB4zHU3sRl1IWxnDx72BriS6IM3wdcCEAGcdavLEXSKJ56DRvAd36maYMq/gGQ7K893nRgV6sLt
V3U1zGrEhRWD6rD6Qub3PqNxZT+mLygI+h7kdGBMOrUXs7fPomPMJDQkaSCDmLWsvJ1wFz8ReIQq
KGPvcq/VSroydld6BSsHF23S+kjECww2B5NxCpvKF0PBtJ6vjuhWIulwXdH4P1ni2whLmwlyuJBO
ZjNSzI2gYKNqnjp8PHYLmCMyaItrdqH4F6T5/oAIpy0p/N3uYQrayWd4QxwPA95BQgIheka0UqSp
PAN025PZ+nvF+pvksvyl8jYCzQcAwWtJpRDqZdrPbGuMN+/dsFPL9opPe3ODUV/xjkpYuYonIcpg
iBnkT609Qi0OHQEv8E8Mwz8PSOCxzFGFWuN2a0ZqjG5YqQyFEgUj/wMuHBhqjFGojaf8FsmLiRw/
mG3Am/Z7OfGmKK+M7oh4/qFpIgiRHRuYW6Fdtbxd52FE/RZiKee1GWFDvq0aalBx835hO9j9wGSV
dRCrribQJ3zrbE90txX4AkP9CyVg1do5/I/Cb/8HBLFg3fxrhOJbuTjHHb//N5KcspLsvPMmJHzz
fgGVkHlxR1VaNG1Wrfp/Mx2vVBMWXkwyrzTaUOEu1O0HWrfvOwW+rfqsDJwlJaXJDVan0lzt6fNI
TQVaMk0ezSkYDoY/6JxgXS9J2Jd8dGPASdxFGW6u1yv7jjZSVz1sVNqa0tU7CBYS4IkxFoIlBBSt
2MtVO11LNxVUSiMo37akIHZMuFr4lm0EDndNE2Bpea3eiR6FhPqnrP1VqCu/TlHv+Y8rBw0HWA2Y
mHvgQe02qaOeeAtsdw1nhfbkf7v+hhQ8SfRExvI16MdWdO0EwWfOm2kWZcylHi/03XzpC0j1PLbv
bhK2JwkzJ0CefXoJtuHxnrP05ZObp2gx0ojkDqfe9vzd1cywJ4DxVBpG2PWfLCBZiUKi0yew2WSf
Gm2kpZahO4/olpFEOyT/3WpPjN6sKf2vyMGZqo2PYmP0FQW1KWuVZ+jYkq73mTMFBhT56qkpCgT/
jvT0+P+ya01msIKxGi177ICat8hK7T60afAx4OwE+8KC1SXIzH/B4VK1wLlQY9vfkVH7BNTnDCjX
MzMBaeIo2oExJhNTwQloZ2Ge33U1i3PnXd8pnmTv0i97bqwh7DZLl4v78HkezjUrwNjHyKNPdxBn
eEdTPYkkq3OGZ62+O2PAj94VXqJKPUQZ/zxk4WkAxQk/cVFFFNuqvz2rhG6FjR3kDgoLX+RS9hoJ
9GB/Wk505LIZVY7IkBEUB1L84fjeQAVxZpbdG3ciuTkTgiDU1L94koCmkpEoLRhWq9efhJQ6zBg0
z6AyOJmhR7yPw67fyI1HmBRYHbjVfPhQQYJRXbsCCnqZQnQ7rSbFwdswcyrJ0bWSzCfaRNmZ7MGJ
kmJYDtvYgo7RxcoFIeJlfjzc/jcb/4J/NtmJGcD+lEXq9DAgpEzA+txjSXNiUGyeSSxhKHTj7+gZ
dqZwfCDDC7AyoBI40SXabGh+1qQTWgmDI/iAaDcr4SOMieKS34FrbmfHUbVdrNd+CV6bMYlSoD3D
mx142er0wLJNCitgPYadhCwlaup6DiWYFEIo+PIsgz18VyUYXgLp0g3VLDFtmvYZAjOT/hgPJakd
Y+fDv6GP1k78CiH3qnpIndo9XQqp+q6lIiqjonwx3GB6Wb7SK5VRH0QJX3BrJH8wF65Ck8scuWpT
ZQjd6hoYZEqa14KD+RHWQR/FLHweui1FzVAf5m6K40bv1T0J8UicTOujoWzmYnx1BZ1TsBvuyFrP
ds/sMmyPDmdiMfo5SVKs7o0Oxa5yL/oZllf6cEw2LifBY6C9yUbU/ncUX3kckLs8apSNnCOmtB04
EHQYzDyYuqIohsEt5h2CCERS6vEn+f22PTwWyFozOAJjHnj1sfq+OMfoVxpHJtRSPZfA+rYCeKki
CmW0YG7HSojQNPKeRo838bxNyAQJuGA6WSbYZGYA73/sBfFI22/liOEb1NqTeBr8xwqnOtdUpVrO
ZBcI5BuUH1GDuB9L1HoRpLgKsQy4yshThpG1x6rUoN9iwsI7KSYo651ZL/3FTrVk0D/O2Mwumcnd
Ys/FH1eCPzp1OrVoQJEcXeR7m3HoddNNFeRZHL1rIYnz8tReY1g5ii6jYbD6uN19ElDyky5Ia37n
vKUJWPPaMNpbV3G1E6CMnSK07SH3a1JmONlX9pBURd1EX+Ly2mUt96O68hZHmbWK2Wb/g4xUbK1l
TJR2RCNmQSvAZY/3y4tknckT85iap3WhTvsYvuNcErJh1Aa3gtsG4T1qwgDmsRNBrEgSi6K9pbtQ
r0knnF+fiFIX3NzG84Q6l3R9KsfTf8Jl3LB722MwXjzLXgjlCoEO73EOY/QyijGgwNp06QbfUobF
9LFNbKcNjDAow5SgzGLFmibMkhoKELA4JnJjhJLwIpAQFD2yNu1Sdl1MC+4+Tm52oCtDJsH4Gydh
i9fZI3RaYcPuuQP8K69cY+mAwcC7NqaGyPbAWlsffQCsEGV0LMMwWK9m76rSM+qVdvSHXC2Gkpk8
A/4uxLVJglj0uSYRvg8be+wp1Ia2499XVwy4C1y2DTtPhC+s/6jcVlyhqeXqR3G+I4dvmCC1GREQ
+hoD7reIQRVmYCSNmt23GtPCwJFoywrSl9fTx9TImBFJszsWF5ROurWr/ymFgt78JlcLZUYrQmFr
5Z3pIQLjSNle9TOjOOGKyHu2HNYTnnECZAz4SoRfDgXe2Uk4O5DGAud/0YDv0TZ1DE8hotK6jtvP
lK/ONfKlDyt1R6R0I9frdCHxZMjNrCasQBZCn9Uety2evLscMSLqijMPmj0RxHSOgNRsTpr7g0QB
+Rv0m/fP4yjD8xZ5Sayyg5oW97r9o0Pxz1DXt+LwxTQL2oNk+GLawPWV9weECRt2t5J976HzFm4l
k8hZsp1QRvvMSoUOYS+CYt7LuYJlhR1PukpI7xpMDqW68LrnJpNmfQumNJP4C77hldEx662nC9xP
r0th4vJ8ytNV5P7VQrq+VAJlep9CSbzbZLZctflkPEnTucl9vugCEJ1EszZIpYlOguv3SAacZLMo
U6orwEa+g7kx8daGSPJXPA72URS6s0Xpf/87P0vcx4kmCNyY8sAYzDoSD6QI5zhSEyRJlRwizyOA
UbeUH/C8Jmznb5jyWftphPBAKjGwhKtmLWLpFjsGEjXq9d2qrZJrBa7YASyZjipdY4Ob9npfvbVF
avVasLY8//vDhlsJH5geM4+DWTI3NwPV/w4gOa+4h3/avU+fNSuDtK8fcHW785kXgEsiFLKLL+Sf
J6DlLAUPYTSSjyR7J88dQNMB9gJ3JH9HRMitSNvYua8K2XNvsbTbVpwFY+xRZ4I555HuX3GAL/6O
Qx52bn2xvlyFumeRI5KfS3sRQyJIYh8XtSbbS/jmUl/TQJ4uVO6X1u4REX8ILq+hMR9Yt0Bs+jDr
xnQGCadWO5mXr4E/QZ7voqEtPBjWKXQGvB8Gc+JW+BTA9L51ILxtOF4v9EMQFn4f39iiLP1N4byo
rHGRVWx0CX3+olfeXQBiEmKKE5vJOszUGoLEKXFcYvGuupRBhkINglqVIM0Od2ONHFbHA5UQCa7N
MLZeZ2Jf2ZMH0Sj6VsupEm9l2UkG/OscjiJwiSNqkmrndWU8Lj1PJotDxvWHQdcN7ZroayAdQhzo
rSa7yVL4WZqx9gZ4d3i+fy8xFRNXsJjPwQ+WIg1bYVySRRCY4c50hyHoYwohlrt8YLuFO+JImFfd
a5h5gYwAKcpmlwP/xRvWEObjm/NSCc4L/b6enh/Lbi5o9UtqkZN2aYZUHJzvb9Nw5CipM4Pnh0JI
0/Jz4F38I1MYIbpQ4MFJnqUYvKxLM0PozOuEotQ3LlKNTHF5vy1H++iPJZUrXk+Sesi/J5mxciBH
GVLe4R7DBSPzfpIsTbnldrZ2kIThPMS95hwzccAeC/xuBTVMMwasxHfiFeJmpmNzn+SLd7Ylb20Q
6SVcx1ymjqIpWH2AQpXj9c7xeHQjK8OD0644oeofJUfDPwFD8415TU0P91xBFwqfFYREp+Mf+3O6
MNbyBFHg8trdAvFtHdM/ibvdjEOGZ+aQIR1v5wrgvVCl3ja/WEY7B/qdLdA+bkQb2lbHy/ksy/nC
0yCJ4oZRakw6XBKKwtT9MJVc2nlULI+HW8PTzWIAoe7jXjrOY/E4tab0xnGN3eLAqGBUsQ5ZbMjf
Q/nECKlarb/LPuLoF1yIxrIQUx37Y/+KiEMiwIGyPSZhXRbrFOESGnua9dNbcudHMK+PVuGinzIh
an1+EiPZVrU1LZARNO0WpLjiD7OWqkVNbH+V9Zqf78nnjK862lSwxnO3ixUsO51Gxbv8Zm6rtDLJ
tnCQvNXe1YqYl4SZwBWQVPr7cELH6ec5xyOeR8sGop4ly0d9E1IIKW/MtvAKxbcw1WEmoY+c8som
L0BNcWHklp7VJLbZP0WUeqHKnGEkHbZWKANBxLnqkdpjz5iwCsWDkLlUK1Y2S0T+VuHzWcwwX283
4ndeIRdV37DYx+ol/wGGMMtt3F6alq6nVIGjPVmAeskzbsmJlqNey9/EbO4K9ib1QJX8asTTL8C7
35pFgbMtBfrr0AXUeAced0ggGPYHPB6aLwk1ROhAC5xxgYrVpNmQy+/r3zSjLI1Rr4/bhBmDBY4v
knzardNNZCgyrojzBuHT8L48f8d7ZiBNg/OubooAIfbPAxQCJM0svQM6QTXi92GQ47UIYQ1qxDvi
C7MyFpAE7j8nYOE4I3J/bCZEWJRu57QqeW9Aei+sJv8uHPhT24ctTuwALyeEVrcBs/2+MLrDO4nv
/eg7rOUlx6Bii9FUSb35BY6pApB8m10YirIOaXIeVBhDMgMSCriuE2gajyQp/grP6ym23A0AL1vB
rKq3qmPyymoOZbedeyez09NzopLYkfV7455rAgoNUnpnpM3SNJkiYiGGBeo+K7Jw5xalPtZm9+7A
4tsHO+s0Y8EUph4PEKqUqhxTR04XtB/5vpz7yQLcyBMEQ/eslfcdw4URO+2aJGouuSFxFUdUvvzI
Zxo2Gk/w4DuwGv3g8q22eGVoFFtzwCp5Go8JYW4dtyodU+4adOvzZiWUKcVnFpYyYQNIP4UI9N+r
Zz44j7e3T8g+ZFva7QOqu2OJwkmqv4vNIVME6wJNMXxiGCWnjviUcOuxPXEA3/ncWIJsx3r9Bf6g
P0xs1eL329GKFWvKGHRS466kI2niB1IiVXB96RmeThAOlk0AEKHmrE6Ym1cbLi3+fMo2q7QFM44U
NMpqLqF4bjHp/xdoOOG4bhvQBrH78v9Shjv+s8bm5owCD8YSWZmMKxndnXxssDG/Qgp73S7peemd
n8WGJUA/pC8TQiTUCgQG1MPZmr/XZ4GfoRBLmOqEMS1yUZkOfLnLCHynO1J1aIeJh+XjJFBwnWWE
bWr9C4db/5IJKzyjNSIhyt9Cr3M4wEf+goCEI6t9nPXQFaVZWjNW2PchcOQO7/KplznwglvRG/VN
QSe3FDRXklA4EZs+6h8qctjlVTnPTcMtrzBzns3eJ3BpxLcYEPCNnvslDNaiMcCwW+AHqJ+AiET9
FYUCZ1FWMZLTL7Yxg36cuzEtVBF6hU8BHARNuekOPz0Y/mUeOlG7apqHVNvVKCbGnm/Y+4ffHUL0
5E0t85+J8BPx29i/Y3fbIDpxQnHSVaPHOtE5EDOMB/0XrZA0s6AhuNkwspH9XvyInNevj0QlpiAy
fHsgn/OcsmuAgnLGWx9PMG/M2vtb3hZVbj2copolKjzElfSpZ3ioK3I1K2KJ2eERHNrgrH5H21Zc
c1dey8B4N8EP7a0EKQMMJLLjx6QNz93im9Dh469BS+ug/MsKjM+XJffHFdBOiA5oFhVewEc3tlUK
XWO6ol3B6lDwN/F8xWG0jmxXskebJI91wNviM4gDch6EW6BAFBvIN9v6X/dZekTOGXzn1wVjqSVl
giGuCWfkUoOhFSLsl5xjzgpxay1lCHiMYhFfoPKafpBXaAws+Xuivzj/u+8A4+dgh2NNihn1aNVE
ZHBTMVdXMYMgRzsVT+1Fk74fkVDBqHhg9llM6SKsh5SY8/zpFNuO2OSReA1nmVvxr2rSvsEGknu2
4rWn0YCN5YP5UzjEQCzfeX/EhCs1Djyf+S9m19NK/YNWq4d0cfDF9p+EQGVKBuBnkakmz1uH6Cgn
svgs3xX3y/2oxwmar5blml/h5+JrMbXGq2qtO48qmRGYk5rXPB5gIymFYkrTtPPW+C/qX/Hwcgu6
szJi785ZRGGNJAKAhgOjdyziYm7kb1m4MS4V6Yp99laskCW7dY7CB5l6mGLhiKZh5FBoKkcE/Fh9
qHP7g/kNLo88lfzzLmqiNOvUk5vYLGAeY+GwsQmkdsxldyIhb2mnIFFAhTCOJkyvCVevaEHHxYUI
RFtUEh4CPYnxp3JA7m0zTkUm+LtznLHmsQv83nn1cr7YcGDpuRjbJp5PricEi264uoRpCwnTZR1k
EHuJIzy6v7qhhmcn/9M2dozwLuNBOUl1lkuvJO/jjInObnxmz2Tx+KMcPYsg3YgBCQT84wEpKRpE
Ip2ovZMYGUyl9PY8k2Ndb4xrKDBe1/96FUzMrSwKO5lqV0IOUeIUk70682QnwMufuJD6rPQhVsWn
zVSWHrlAY2bytlZRDr9pwtxJZd2q4mgTfVpGFQMp3qj7g3wafmuypGhfOsWNA9n117vY+WFEc7i2
cMFrdLfjYJSJZ8u+UF1MH/4LfSQB9AygF8FR+QrDSd8AbiqEFrAgFQfZJt6LKcxZf2Y3QhRvG/uS
buSfo89hvnUk9zkUxJAwhBKZwM9L1ESwo+zV2Vor+PYor+k7xl1uvKZZtBZ12rKkZozjDR8diSkY
TRcbeNhXVHiPAZgUOX8e3QUbDr2YlIjGSEe10XBZLQZi+P8zwEYKHD9Fk/CVz6z1PrAuifVvpGW1
nI7XgLU4cdV3tUGxwv82Yv+rp02C9diyaDi3LEqyCwo4086ZbKR3Cw7LcY79W/O6aNNGS4Vy5p5S
wk/tS71R4xrlu60Bg4c5X/dU3knb3TrrPk9jsyIXYSInbkTA0JfwnLDRBPnJtiHCWJbKJYK0FOLf
1asSyQaTNv8tfXgj3PsbF8sMlmXe8u45UcV/OEvmoKZAqBL9QhbNd64yxIltnVGeriovFm78M51e
D0BuaNBewqS7ntyesB0352QFzKDpYE1nsLpINGbYEdEM4XlDKYlEV4OrGZYZdGp9nASLdTigz7cn
nwvf4vT447j/Jw0Z9mkr7PWlABaxFz4gyZgJjVcuap8fFFPkT7XwpISRXp1hrzMLKObr3sV1ROrb
tojeUaRFpmrqusegu/EM7Q2RKb/6h6DZO1nWBD7bUGNPpXEKKEc8j3psRSbItTOlcnsgot9Km5S0
B1OQYgTg0dpPhKpyb63maI/bjzyJy6NeRGVVamkE0+lWMJPdyJNoMwoIYSZrBzjNoF4sewKuJZnY
82daE9Ac4YSBe8jcUMyObR+q9TQ9IgufwPCHq2B1NAR8ZifuvGBpSljxVyIpIOerrEWEDHxJbuG4
CleWBauJGhePAZ096PnF759PuLfxEzmf8G1BwLF32nwCt6XJ3WpqNshDHOfdZQUC81DBRxkCj2i7
op99DrOEPSEZrtctVERJ449qamWDnE/kK1GUC7K+kMTdBfO4oESExnsRPdMIaKrKkVvDFlA3heFU
N6FHBRRHx8IYyQuJRkJM8ua3IYx3iZ+T0HEGg6cvSIHSIcv7Ti8fB8nZEJvAaEAqSzbEneR9zcAM
1gldqrVCSetgZR8zQWvVhoFIqNC7siWpWVMh2h8mHJucRWATvpBIRXCSyKOccfJKz2K0io/tZHb1
pZeK9ItbtCxJ+t0PGuMudDMzgKAOgKxfZ7ZEuwXsm1VXDUs3Ni3Wp3dc+FIhCOSBkyVTQM975cFi
5gz5U8vZNxEZInYYDqRUOWb+/nvKUAgpnIqFrwmyjoIJtSqU9NWeXJX8kw2bg/oJ2Mqge7qOmtsG
PEhL49UjtpBC7A005t1qmJZKCo9TwV6W+VejKjGkS8s4bRDwzKXp9oDxknGSuy/vMEKYi8molv4w
zA0njRrm4BrA4BHuBo3v/dtTVO8DhmolpOrVP+plZ/FZLCznilZQhZPRoWoWucuCZPfhu6EkaHol
KgECzx5hyGPSBfJHr0pdosFeIPQeYNsUxfT/hteI9rpYmwITwXUZKiL4T/9KjFCMWCg6xZBn92E0
Sec6w9tj3HEagmM89KegLLEbk4jkjHfs7fqeAZtHKBJJ5DyKzuZH5WkdPBU4RhjVcsd46ug1+Evr
cVXF8CkfS9+AMapmq6V9t2O+MLT1wX5C6HinX4rgrhMI86eJPxG4jotRPZPAl2bkt3lIRHLy54ea
qEYtCHE8wVqJBJ2iNGKqMYLUNQ8n0tZSwNE3qszcBfXIXs4O4RQpAUwO0C7+lxu+5b1cDP+DJTlF
GBiZ5YaYWJdNhadsdeIqV6rzy2iSfD6WJgKzv37mGNIzvTswg3P/thV9UziZrF6xHW2NTSujwg/n
31YuWGDZbUDUQlFcnwfIRA6S91A+/f30Q7KOOJKYNPT5OJFTZXMRo9j7mIprov/yxOWyLEMz9Mvy
YtUhrg8U7g9pcGrxBUrSZv7wK3s02EoyVLaZZ+lRVTcxse5jLQUMOrwjhDC7Qdglf8pyCk6oQSJb
hoffBGdRRHleaYeC7PTbrY150TvrXtzl2lSkHm9T0qLNWrifFkDp+ecrLQ6o3yKqAUyto53YlQNx
VzrMwxoBmrT3NYySpBysXFyiQPWkm/3mjCYbNzAsL2Cm4rpgIuzvOOIfba64dFAGjnRJnFNf0SDv
6+e2NX8JUfp6UuT8laHzAie3rNygLXruRWr+hXlx6znegLNUxEDCXgwVPhk22LlHHJX9KC6OM1J+
JSfEs/j4LwKj382521pBxs1rjUpSjUUKqYR4Lqen4X/BIeUrEaLOwKE57vdx21rggRGMtSa54A1r
0UkebpAxipnp70SVHa2agiWnhBj4XtnsmSaU+Khv/GFizbTOVmIlbUdkvtwdTyYhntutP79u16Da
vVHprWWthiwg+HArLrsTx2Lo5pOXhYld/fumAFgTu8LT/6EcdLKQ0A64xLan8Lo4xhGo0uKbiEA0
HyWzmPX/WQV4/YleCqxx3K5BZM4Cop4lfru0V2LWWpJsWwHOs2c3ahe5cjUFXxsqh3BOcDH+6Nov
1JYAMGCm3N8KfIXFLgQwc3gEDtBs+7zdUDWzWpx2Mdpa1oQnujCE+l1lqbOIA5Ci35VdHJPLaSXT
PZbLIv1tnp1tYnjeF3RiIdlWiWdvSGVysZRB/z12Y2RDz2MNCdGLE7O/ewCDe9xdarxCG5I09ct/
v2OsNAznT1Ehx6kOv1ymDWFhDFpLTXSAYc/twgpSSok/Lch7xIyZmIMuiPmgyqxNnnVtisPyjDrX
7s8up4wldJHCyzta633NI5672mzNtsVrqv/WXEzlO89EJ3xshazozgtQkOrVAzdf8jywJB/zhw+O
1zQhE4zgJ4v71GMemgcf+opYE2mBkbymgyCBaoP9Nik8DjFBpTPbqW9+2CeDPa99aUSNGfBnBoYj
OELnKg+eMHF6xEQ+Ua64Hq7QoNor76hEUB8h3OykiX1zIgGj1xk3E0ZIeJI+EQSS+ybZ4lm9X2mn
eUSkStqSIl8qqke83scNvewBIbiEjr0ZQeQrTP/AN1kgPM01Fki16+np5tzcY0VADi2fVaC4jymN
RTM0l/IjsdX/1v5VeHbo3Q0KgKIj/OkddxvlIMR8WUjLCdxGTw8QoH6Pys50kEXg6B7O8DrKY1PM
2bgq+UBLJr70tj1JUjx2UbsuOuqNa2pCi1A9VYvNzxit6lO0yzY7mN7jOdd4RVRWEPEdQo/EuEc9
3h0IFhV2lcvaiz/u102BfOD9Hrh8RpP5ytRoYqy4owK4ODPgfOnjnw8c5yacVAqLf6+f1ZCussM6
m3ANz8I9fQeHX1PuuT86VsB8iB8oRWReiCu8hyRFTcF08nFUJDhxeZ//bHPJ19krPykkTpzm3v24
g9QwaSF0gx5x7q6Kn/89CyguLcmeKOCpCMDIH6SJkJRcQ4KBccEYsOYn6Lemx4SFI3EC1aynv4hY
6mE/BWKWchdpQ/3M6ocOaCJIxJx1aivyz1B/buHyWMFRUee8aEWXLvTuvK9eA4yaY23hfQZcrnNp
TxsWrxZzxYvwVvVXWL+SaiVlCvmxR1GKXT2o+peawPbHv4RmDRmVbGVjTW2tx5d/2McpfbUxbI88
PnzbY3PBFHgLver4ixu0nQ2xIPIrOnklWKYE5iCQRAgGV+EjlJbcr1EjVpzKNPYGY3y/sviAHaEJ
peTCiiPU89VynEGeXQ2+zoKmQ+UmC9eOD6SePlTmBEIcW0/z+bg5zTSnZOFtBZUALbfggJlWjloR
LViv35I6oh8pVBiz87PhrZDqIY134TWiQs/tlWXk4OojSAIkSGIhj9k6U7/vw14ap0IS5FrCvx3d
CGdcKvzYp+cto4ZxCNP7OlZG3NR9piv5fFKYLkdVnVLAQ2HKQ35xvQU0cGqvVlT3U7GzO/7MaLVG
V4gTdbOC/ZebqBJH0Tt2QRvKGIMtpTcEI46gtL18kYWOOcZRdwtau1VVO4bkTkYkHlPZWxVuPo/q
aeVGUbLMjQv4kKTTAyYLtqxvZs5K/iw5lxMX22c/98UUd13kA3HRNsP543cLvKgEC84WfsxF6piX
Bi2bFu7FweQ/ILDuxrhV6vBisyhaU6o6I6taMpajvJeYP7intQhurEU883VsE2I7sWBO+aN4dgrK
GGIeo1yJ69wNxvGHoKPDDXyVHQvPMtsaYoLlcdlNIj+yTKDWk82uW3rMTREuIWaOKrY6UxgPhCpj
B4G4fM4InWDOnmQ4HumGpeJ3MW3QZQAWRbdu6T1VzyNupi3vrpjXvioASOlROoZIuIwn9mddwQkF
lMbHxwcfCnJgUZIy7rORRADjrLt0uVmuNQl+8up0gsTlEeP3zjykeuvkxFzJ8H+yZB5xxk/h4Td1
IJXrozrrufcUY8yg15EnBcRxdTQWztsoLvsLwmmHeDaqUslTPS1+ePejU7eZZ2AGLUc9edlqgKeD
HMgxgQ649JJ+5Lf9Fekkut/uWbVCprYSl3aDoRePfq2ik/W7oS2TVS8CvcOOryVqcsjbwNHRtJm7
nn3QwiLu9YB/dF0XTsKKVWM4PSZZzLxT8xKiQbjcaJf0Noi+N/iV72xfYHyvsh5gpoiDDP4/gF/l
yShBbcYruw3bScTA/EbSvD8zSSY5PVHItuYNk+ZlM9GkF9DIm6gT9vuKm4j/NAcOIrptwe9wpz8/
f6U5d9o/4kNRFN6KaoaJ2sszavMNLDObFuRAUFwVnWVFbMLmoumXiyJhDIYKPVW6EUIgy0pGMGkN
NsLDEimsW/i0zXNu06IayXYuCY5HccHSmR8VtGK45ud0LgYZqXdXU58JdTV06oRe6TQni0lU1/Q6
YJHvzZk5KCOWx2Lnowl5mBXVF7VOoo94uKAVfoCGiq9pIdmsgiYO/NRX6JUlaGAglBhGjVHRhjwr
lzOrn7J3lVWAcq/pA2cPkwKQb/5A86i1DXn2t4FJREZ4yREisgfXqvwnCyxyHUFzuCHCSQOuKZdO
84unu1W0SP0tEVTie0sSwdBj2kKqyp2tnsEH9mzcrwMiJgVTWkTExQ6Nezr8HgiSMMFmKqpWH8jv
IOjO6bR4FwZIcms+3ymPGjr3xrF5kV19SZ3rvwIA/tNkuW4xZFmLiJX9K8M0kjxHr7veHs9QGs46
1LmIat9YcEZxE9qrq+tlfEK26lpA2MnHNSCRMHaahDY0RkOuzw0S1QmVSq0GgQktRJbePlf7gx4a
zxt1yo13d+vHsNo8Tx+jy5Jq1aX17vm5ZoRhA/+YcvC/gx/BXjRWhUGS3ZkxcJUoeizR4FVFqM26
47Ez1vwqh/c+W4jPYGqnsyhk7BhnVBr0pDw0DmAPLf1X6vZn+7x/ri0IbD8vXTnaEq4GHXhp9yTD
5RXbngWRo09uuE5yWOvzNXjw2U8gEJeQRfxYsiKMTnlN/LbPVj55qsQlZtAf7UO2mLJ9EG6relxO
JS8Tycn3Nu2F/tAFlKwJTMc9ulbQjNqmpslRERkEFlxoqewf4pAB4KZW5976lhm2GjxJ6KvMSBpB
GepNvEJLSKxNnhg2tHqTGskEH+mZaMz2Oz3PeyKILYZ0wS/jHRdm5EuhfKqG/HJYZU3lWLf6Tj1p
u7+0axQaOmjrnWlh+hBDkvyj2wykHhYVRXMTusrHH6ni1/so0ZUH1Gj2sT4kOTn13KxMSflWlp3k
MnPV8lm6+KWyiqb1WvoBSKzS9Wg+LqFwCfHNAgBxtHPD/brPy0QjLcjdu1RtWbrECiHYf7YnAHWl
Kh4t2AdIu7EoP8j1srUjZgbncTMOwoNKZoBmkGvSnUzq9GXZfHowfGj5zVzt/cTOnqerngAeOIJK
oe2C66kMitZjhbjUz8yNjEhpF/ZXhn+8VmIXzQGlXcZXPrLoNImR8hpxVabE+IScxIyjyfLQeToy
JdCw6/mmDlDEfzJPyE9w8fmuBzgzMndMMmKa6MF+ww97XwWsOV5y0gbOvPnToqr4Dlw012y381MC
hE93uPn/yiH58Q8SDCLkFgmZ2R3YrGwTN32un7c7d5sjQX122xsqbDOSusHCu/akSaLHLoTz3+tc
HhPuNdj5/s4usEhMxXUndYXNMoufMukNKGjKs1a288f2Nm6bgMzAq7ZZ9ZUcbX4jAb4pBfZvOyGM
yaG76+k5LzM7C1syTeGYV0AZ5qYMfjdFpkpoHpew8jNd9OR6lH99x2SGAaeuwpvzw6WnhroPgT0s
5g/YW9xZcrb/WBDVpRMBjhmAbcybatIEXBXssWHq6Kt9o01FW9oSprpvOoj2JoQe4IMgGDiCKezO
E6ZpAJMFD/74VqXgg0EinjV2MdgHHJVgcDKJvGljiWZ2eIEYsgfpMqOSanaUzqAYTVU+sALCJnMy
g9E6TcZruqdLJM/LPLXIZhE3VzYJWYVorFLyaQW6h4Ztuu1iVM9Z0SWC4QHN5Zm/w3NqLR1iRHgy
kEZaXSoC1PJfEChR49VOiTh+CFZPIKOvCNeboUm7byFQGsXfcIss45G+d6/lnMG5cGm/nGrRvKmf
l+CtwGJ6k6yYXfNu73aiA3PXEXEjPKTV4oyzHIZqGUNPQ/xWO4L3Tkw1YFzOhRTU0Gwe3RYYITnw
zclJKlkmJYt8lS1dU7bepft+pNDbi4IK4vJUtD6PEfVWKWRR9ro3qi0qj/3hq4AfmVmV/fwyRc8N
g1uOpblDg5bJHuHEv0/jGzhGhK709+AsV/9eu/TyRedKudscRReVy3678HJKU0roZa0Gynnny/xq
vtRNbKgT+dgomrlcsxAsR+2BwabpLQKNbdh3O7h4B/mW/+Zs77b3b6QJxKbq07ZtCOnADskPquQz
15m22mmbfmkoZpanWdDf129XZtiU4yS2CfgXg4drlT6KV76QonOFRxy/l2nlG+mSY4AVbRwkKMfm
ecS9yq4Z5H+XKnaCxrz8oddMjLRzlqxAbSmKtqFlauXaRH8z16gw6PettrSFC4i55ROF3UJdqdmR
Ck4pbXhMyDK/A2umQU6YUHh4qedGwvUEXbq05qOyHHsnFjf1C0OxUW3USqbUNgIkh0I8KC6JKi7A
BgDPvZYJ53lUiK7rtGawrfpcAmyDgTSXzBJY5Gm1/I9OSH+1o93w0N35kwhy73wpC1GTGcUJcqbO
9bkT6Y0FyhcTIuzr92JontzaoM+W8VvvICvjOtk32TOdjiOrUmdM98PiPfaTQ7wXbQxTjJp+6Jt3
f653sJ8d9yGjLXJHqMgL51rtGy/cnGgO4FhGvdBe/2VQPQxn2YgBLQguIItYPDszRMuQF1tkE5K5
KcdbFSNQwmkNAD6q6DI5/Wr6hkfW8ajO1jQ8f1wuNZWUE+n4QtzjrLDRgLeKtvqm3kr3VPmy+DB7
4DiSWDJCnuiHQP0nF0nwjXQbDDDVsvjK5N/pTxTK3ShAFnV1WLUl7jIDF0NAhHh/0y/tjYQ3YX97
RPatiUT8VXt60b1dlfOjOPLMVzN4hf6UOQu6iIMkF817kxu5yezR0+QuQYxQDJMlSX7TdPEwCMoh
fP3rk1eQ8xW8kksSDiLrbtiCtKYAGCRPw47rIcZMR+9yBnA+8qPjcDHKpM585GNG9CuZPI74kE7z
I+hqReX31tW0CWVUoIwlDbfBJkcSMLlP1o/9V4xccpZZLDisekc+Yqt4+Qnh21H2uGcr55gm3wyl
Mo/Rz77Rl8pPS7EdPEMNcxuMKMCiaCptSMKZSs8D9q1zQWvSf6KErRYSJc3cbkQD5EAW2KCMEOkQ
0A+HnXF14eT6L9fMJ3EJSvwPYSTIKiQw10gtpN/yXLrSz8FUP7lFaYgoptHQnSpCKSJugdOQQora
WnjFldwYgIr8VV7lFq4/p85CRvRpcY6w/LTkFGKL56JSlsnRV0EdLR+nRn4IVNcHX55Wn/0hcphq
n4cOz+ul3wmdwzKkfjwyhZ8wZ6T1cC6SyNidbG92PSHo3bJfyinjxMYz4VSUGzvEPceeFb1IYQ5o
3y0gaftiD/NXyiJrdg038zR35D3ZFq79NAL6+Yj8oqY9PSgFZZsAupWczHX9W9xj7NuIPqF+HDMJ
1ptiT7av9p7FUuhoXGoDs22+cOguz+Z+Ux8InqOnMiApuB4hoWJkYuxAWc+u+w1TqA06hACOgcur
tOnBHgYCZdXN6l5lQvO9lfJSvw0rQnL0gTr9CDaFdxvaSrscqn+TPJjaMoTTw6TM3QUQ/iAWlNEj
ht0Kt4+LoWr1GwXycTTLnf/wzFVMADQR7/NLtGKCl7qNmrh47+1Gxyum3UAXHabuHhX/PKAWkr12
ulMOacpgtmHVT0d6HGj55jM/Q7hcQRba5lCSMwUgca6gpS89fdSkRcZOfY54IEk5AYCTWNG3KiNg
ghFqTBHDUQLJ4pufCuIRCvc+zaa3fCTDd6II1X6PtfzgsB9pLeO5buu12FbFdkhfG7MaR735vGET
3IhOurHZBKtMdkBFKE2eeI4jaazTbNmuA2WsS6Gev2gvpRg3i2KeMEIdfYYmRnvaq/zFDsPxKZDJ
WzeFiMRxuY1Af27O/htCgU/rHNDrU/9Nb0XyqtOSSQoWoCuCc9PiziE2Sh/Jjm6tZ82/fh7H/OkN
AnZ2LPi7+G5Ych6kZI+dOPN99K/vGWSuhfM7k/HCW7SJ8zu7dxI+Ez0rjL7KmO2m7JnMuH0lssTd
AKYIQmtZNLDf2UMgRox0maqEf5IgpjnqXGeVV7Vu9bH8P7p7kUkN8y+rbRIzyQiRiw65WlhREOo3
bJgJk8BwT9jQfB51ZeJlG6vKHNvoStIYUfUMmfUybis0Q5HyKTwAqkRM0Jo5ApoLDA3B/+K4RSiP
jq1QUZAoMdKQ79C7twY8CaQuUfQ078zjZ4TVNMzlyyjylrlG2ncEvw/uVR8pwvgPJgDtI+u3KjNT
x51ME7qiGAkZhlRqN393SCu9aox25fugCVp1QdkI+Pvl9MUEszn9dzUDSppypKLvKcTGTyhgC0+x
rt/iTA8yi7e8WRIOPlMSt8PRSsqaVp2/FoYbiall1zgnhB/Q2dusDYHFJV0TmSTeBv1Nz+r3Oc4g
z+FalDywbOOuXxRERNv9SEwkNEycFOFReqU3FL4n5fm+CrXEWGr54rsi2SNpqvqF0pRd3Hk55FFH
PMQXLcPcmiQ6d2HiQFmKys1OXjoQ8HqrP6hAnQLXLcqI9hzi3RRdgdn6Yox39ak6RZ1JH2rnpBSv
YVQ6er2M7PEl041PYSYD8sAXS2oRsPyK5zzJEI9BcKfxIHzDoj6hNnqCPlj6SErFnK2bMvEiVw2d
NZD+Vl93qJY2dD4qCFih0EW871azU2fu3UI2YnA3ThVq1F1hYj/P2loqYPcpKbrtkpppSWGYJnBm
OwSneL1X0/tvWMvt5MJd3Uh9ZJXHlxexiO8ZwcUw/ZvLG6Izb+/ejzMsDfbE8lNbM2xyzPMM0LQY
SuDxC4xnZImEGe+VEJT/Ns2OGrEyWuG/eBiQJnNpv7ckJk4ashM03ntXAd3ueeM/3PqS87puG6Mz
q2iP2Kq+RbQGM/mfkBjvEU5/UPfE7pmojBesvEZop8AT/wUJhZYiFf8fJvtloezFLTH21rgjYZu4
X2aqiZbCvZYxusujZWo4q9Dtvv0UeIRoYjysEqsSyRiS3qWS7560JLzPfVler/UPwqE9tfO1y85Y
ZqSflNFLLx4k6k2qPTwz/+sWOqviWHTLLtjWnHPZUTbXQbDwGDuhaLs1E9hUjmzKl5vGpkhEgOgW
qa20S2i/ebNX8zkUER9DW5X0TXjPXjHCJzGylK2e76XYVdVno3BT2CJvdWFOXTe0k/Lf0zr9P23L
UXli36Yz+E3wSBaQVNKsXLYR8IaY03yYB0lZ05gWpZCz4i7oGitITKZud0FZBeDzz4vvpWzyyWxO
xeI7US9V/3yxjQheVfGGyqPTuitmomuGziVo22yfJjGKgkExYyhsgbHfydPXvuieDy+D2AOC2MfU
i57+FnXH+U+1mHdgqR7WtFv2Uem0iVC/yGG1ThfN2sbGXCRIzh2UT1UQa8DdWBW7jBw78EIwukv1
+dx8jj0mHjcTuOKDyjmvASR885wFkAKQlX/G7je2+POPzn6IxkCpr7fXe4EXcxV7BaIWQKeF5CDD
ZUiQiYqmE+TNmSNwcnBFFmXNNgPDFjcgvyGmPLYhnEE6vfuOsJUkOsinXFXKKlYKAIa5M/J6aY36
f9WvwFfqsUinaIffWf6vDF+82utUzMHF5NNaE87Elwlymkt5z2k18pVMDubFBKGvmk3e4KJiHGpK
EEB027BTm5VAd5jyiMrosRmdnPiDjoHtC8geWKCTfqsObvEkx4NQTgFDVtrqP2SRLgQEYYBX7v4w
fCp1/Ih0rBoPUma956xo83RSXN5IHfH3s3Kw4LSBETVqaSCJ5XWD6bmzEIFNX7ipbqoqaYwI8+WW
N4pDMLCS7KPKWf7KALHOyxavhrVvvCKnmzGSWlulsvajo7oyMpqdrS/NMeYP4DXi2yySZ0WVaK98
W543Dbul+pY/26NPZrAwzMF3nnWBx4zciLtjvZu8Ot+vubnPkJLdW2Bwlh+cNiHHY7EEgabSuft0
hmrm7LFCdu1BAmOl63iOcO69PUcqPycVcUVgadYfT3giYvuUvNhKMmS1RNVYkXIBh4A1N9DbbWYY
wJeovolw09Rm85HYLZY/BNu47riHU7TcHTeNgh2CWTpb9xamfINewS8RdjemtmB1l1pCEP/gK9wK
XoDJuHnxJQLunXvPJwsok5mMwMaaLDZcik1PW+hyWHiBjrdG/gfWZwhVZG9jatXKdA7mk6qodOl/
pS+T1ELdVt4prppRgboFghFLCqfkeKMveDwGjOVixVU0/Tt2YWq0ycQX48UrKjFNwvjSF1ZQ4P4f
jc2NeVS3mObUv9L6AROa816B7bA1XlYjTW4UT/aEKf4NUT1ssluufO4PY/+TXGAIuZgHlDZxgfEM
MZoMMl9A5dDleHDf5GX+pv7ddePJDJzS0CxD3BeTkZ3vUl2Eu+Xe54M/vyCG3XKhQiP0yFwIu+s2
qDtZH2hppsz/Az67m7UnCEXBiBWI/eUzmJ9WSHp0QOf3+7fgL9taWiHufUJ2JbCx1d1hBYGWNoNa
qb7U+nnQ1Zu8/7rtRDgEs2G7+QRuDCrx3ktNCaRfuC3j9wviRsGhyqWEzKdeynyr3ZzEeqzIHstP
zBfAtK6p+gpt1egzCno7k/qed4/k4nmgMpvQQW5Wbnpe35ZSNranFHegiELka/EyW2au6uvnvLU+
BOfrr0hzuFvVXI9Xr2EvPjJp4SHDvqc27bMOeQ3FpZbJBJ4M1wOI9KIdc5nEzJ2LtXXv0Atw/TAw
9vqYKbM/tvAerQykFeV7XRDs3theGF2dljU0AUjxZ9zFF8udB0mXBiXmoObDYdWK1NKyDuIIWwk4
5cOP9siOSgcRTO7Df3m+5md5PW24C2NDi1ES4q3PYgtIfpKhyUFLsYykGczGJJOnmaWYgBi1dpDT
Rqlejg9Ej1T7qz9jwc2q/PO73CVkBJakXwpIrpJfYI0ULOGUBW4YPAMS8B/yZ3dYI5WolkIrQyhr
Lat8VmSD04RWk0jJdRCgwkJtH33EZsAb563JzNcBH6odAq4GrKjIoCesYGZN4EKriLXXuw/7T/dl
WWB5ychrZOuvJTcwz33fda934pmeVjFUj6CWzmeQ3us7G5K8L17q6nwmiCwWgEmJIFnYE1PFvgUR
mfPzKxS5eCG784tGKZHoNhQaRR16fUbDVkThWobM77L9cstWCmpNb/VYP4cSd9BttiBzscRqMe70
wOgBw3bpbMaMuMjRjlLicasQESXRS0hxnHy7+CCgp80BTc99d8VbeEUAAFicptX4wZVvfphbaDgN
O8vOdDzITu2XZuF2lCM3fBcMAj0R+1fum9JcJVSUzX2FtQpdWfoetiQQM6k21ASGEzZKrkgpOvP2
IWQ6InOiIIfOGgK5CC8qqjieomZKvQMKivNpDaCaEDMrMUSe37OQSURWFOHbnjGYirVFgkvSaBlv
xDFMu+xAOURVJLGOD8wY6gK2knXhJt9yN9lzqJQgnwL4RHgxSEdYGkV3xt3ooKFCweDPC2QFxfVo
0LeM9/qOvj1VRz0cUx7PaduoVj481MwINIf8YSG1aHNdEu7p+RXdr6NP2T8qWFLeo7JLi7colNlC
qVaZr658ZMv95Dql3oY948UnVLG0MKapYEZC2grJBFs4y0z/JI9x0AwioUfOdBKlipt4d/iKY/SP
A6Zpn++T9IEtFcVzbLrWDw9u4ZPWSE+R0Jn2tHzTuhvjhrL2lPIvFjUpk2Ndi4IRpw9T4FTwXtlz
KsQencFcg8X/xpKZDoY+74ZD2c3MK5ygNC4h6dIIcTm92LcLqUz2IIp0IvRUPPjOR+O09WJeyfbB
8Fab8gg+atVktvF/XhKzvDF3DbuahFtIOk+YKgkeTOa+0f6UNgsmn7+4UdNu618qVUD+7bMdFb7/
TAVyVyxGKQrRudkLF+GRTjE3ZxHV0KpNwpHNqV+sdQ+cU/4AT0vMDxPMlwvQnKaHizdlx9PpXLNB
9ySemPlRxyonVR9gNAs2kTyeZ3H7xJrrvceBlJsmwCFVZgjVV2euF6AfxoJFlnRhKPy1nQxkUcKb
fdw6D2hColKW+jEKM8Jh1wVMrTIqmYv/Pcv70eeIQ88ehEmXsdN2+ND7GxmUklQYhJskLEJX+XwQ
oP1rtDzjVrr996qLcOp6N3bgsvYMvVaTJPJnfy2eb0QMbbxb5mNl5fYZ7dE4Tpj7/3Fa3YQdWUe5
tKekBSxb8cOe5gQvB2TwtCkPUav4HNMFq85aknQbHsa8ogCGuT2HSu+idpgxoiKQz8QNrMSzroXg
+8T6qNdCGkXbxKRoTcCabBWsmGuK5vEK9edP7x8/0QFsLSEGjw5otHuw9c3zcz9n+RlQK9lLO3em
4RF3oyHJQPDLfhwL7MAMWWPb12pCRZSnIEvS0VDpHv4IEW4Ks2fIEzIsojI2tTTDMfiOyEaApZxL
yYQPr+JatSnH8MXnk+cHk3WhVqseZb7f4hQVyQ2rozaIG2WCfFpIkhUY1QeswxlPWHCwKEiG7ERg
EJI0E21dU9608l3tQL/S9JTfbRck1PxGr+hwG7Suvd0jFl2VgIHoyOERCylO8kyDjmznSCrxqo+N
SgaEmW7MQh754om2f13wsezzkhEEI8HZLivkr/TO2ggr/1c0SGzpe/Qq/Z0XUHOAnBO7JBVddf/x
8GOYvZS4d4nTpFfJtYKg5T5ITvNTDe/cMXfKzupu8WucCWj8MIZ3ZLKKURyAQSk8qqovnei9eo9c
dE/esar1N2qeP0FuuHiGoBuPtcL7KIXvxf/yf4gVxEZxdvCZ9JSil6J1ycvUTYd9VZgoMP47XwTh
8iL4rqa20h75HN5z3YXOOZZhMDipUEy/3DlhOOuHKorn61+riylqwSGEk8evWtok1Irp2ftGYno6
cFquB7JGno5re8k/W+vkyOiQuoMGEwbFMw/lzsOe78A440bw+vzuFDTBxBrgFWhWllDMfZUQFoxn
mFl0MghMjSIXyMbaAk9YV5FJkJNI/UEqABJSEz/KpsSV629rRihjPQEdn6vtgC+8UfaglphKOiH9
WksWKXQHzBgYFuxy6SBzMNRYxnaGb5EOcnf94LZI4vdADuetcgKAoPII8C6dLdhaKg1JwtaPyGmI
XQgDi9SoXj6kL+TMyoBtNf70i/YT/nC9j5+E/tyk4zYkVHCxTGHmtP0DnJZHc670SX58ZQnajSgN
pyZwLnqwsrpxRKFA+BP0AKubEWbx1ARG3XSXVuMGb096LNekJ0/Wd1jT8PgAwlXQj4gtZ7baspDx
L74NMzSkAiwNO9Nl6m0jq+fLhPtU/R2cDh98t70SOegIfVgHIEQAA+6QxkoizTDGzodAEg0h0Yh7
8f97uu10EWdCqB0N/WDBoUPNWH50KrvT544o/r51h2s3zflHxBk/YD/pKycEoH0fQEvYdcENwlNA
Ebw6AlDHJjff43m2VurwKDBuWlTRIMU1JFFoNORolvpBPYPP67Eu7XNXzPdjNItou7lwkf8HF6zC
GFZwnhiZZDtvufYuAVNuKM+CWyrfUR1YveiTPANq5S2zzAj5cSUeAtkgQW46f8jpQk6lIJSd0Y2b
3MTjsHcLDXylU0iQmCJAm1J/1J3tnndrytHQHPo7/w6cPSFSKBpF/rgGrAmDtFXTxU/sP4TyR1G2
Enl2gc7lau4CU2TuE70asFA82/goRXX1R37riC53AE8LolDjNf7JgY4K8h4pKEPTEykcqPRNSzs8
rHq02+ViriqRypKNXLNLg6hn2eF0RRgyF4e4hqudiWJMohQKj+P97wDREjORhHwTwCdq7BPEm+7f
WSDtxKyLSlgfJdAQl92o1B4A/n/Oetjckf9+IXfbRCneMhQpE3scg3JiT3/fgitvWpZHyrJunfI3
pOgA2aDXsbgYRNhvy4P2XGjyEbYRst1YurP4UeXWeQoq6lN2quS/RRP15BXpIN9VN/cTsyJBSxw/
9mCpzwkLKnuSNxAyWqoAI23dKYN98DYYO/EHKOi08malGyJrYArKjQxmCcKTJGf32j0Ukdm7wLfO
9grlgJ+mVUF4p1sxIiRFxHcnNkyjL9bPVDNiCki+JpqFAzh2EImSn4kdJkUfPEYPtgASYwt0T4mx
m4mqrlb51dhlSV1amE4R1EZ+ZjAKgayzmBOSkIazuNvf786yE89lNoeWvStxqlCl9wemqU92yIH4
QNWzo8LYqXkGDYl8VIh+tzqGQHgIPeanokRZFhhxUro0q4Uf9hHNInwHgD8bxe+IJUz2b2YubVeB
9IqrOEgcAlff1NwuasEl7T0aEmHUBYn0leAFkSpOeQm5cs7ZumCL1DvGbcQm23blNS17sPjFUGAV
CMNJajBVoGDb4bh0PxH4QxLDCpQtR4TCUm/33A3YXXOpdCYm3r3AUeIhCSNZIgNRk6EDmBiAHX4Z
mH0r+jlOosMqMVEgbDqYLTi5gtxejyCNEIjzsGM34MoL/c1uA1z/lL5QRCsE3E3UlIIcqBe5ABpj
OpCZqGdYHraDm+ewMeD/t6QI2KsbGVaX1Bar39vMrNhVTMzHV+Mmi+Dl4quneqHzqZcSoHcDSEGE
oXhjxi+Cy8u8L/cvPsXD7q79ie5cxg5mef+7USyTK/NtrPMzoiRTfIiUnUiCamp93r1lgFjXTFXm
dq0k01oX29WJ98sKEeM9WFWAVNmsYiDDHNmb9YuuaZwcA/x5IW+owamdqFOLGs0dp8lXz2ofsnEP
QOZLt2Fs3/c/3Ex1vDpAM01JOtRFfPnGfYJzUTUvdF8oiLV8w1qTlqGrPPIUlq3RfoQGOflt+iYY
b3tIQuFGPd94cHjMm9TJEtWNFX/czMg6YCWuNfrlh4R3dbzne1HXn/rp6ejmIKZKlDcJzA/xPsTh
pktFiVZp3zSx/KqkkM2H/aEMZNB1ktKhVLFHhZgE9W1kh44ciuPZSQUw9GieID+yOI6Ozke3tjy9
WFLLfZAJSucDQxokm7CboDNp9BLCeSyG3eA/uFfjZIDXyk4N4U/rpGf7YiSjKYWChJVpc4dnmXHj
eQXijhKNaEhI7oHXBZoFtsFA8yDCAcJyBU+3AZWsVo2nv5SvLUXljR8awa21EYfEvfWrkG+F61KN
5vtLbrdIaTOSMxIfgv8YDuNb9OXfAHYqM8bUsQluVLXrK2oCgWWYSdh60jYBwTRXADWTR/AZvz9z
NyZbyGL7VnH+144KSqJhQ8knF5GowxXepZFTeQ0HA/QcLV4HCwPjOeDzKcQ19Cs5sBKaHDQePOQE
3VBHmuHOwl0PpaREqRuMMnjDavleKH5WA4SCA6JGCDfQVw/OqizG266TIipKJXhTRWtI1uuSOrUA
yUcN6/VtLgNkJrq0UaueXh4PjmjIoWVmEmMtpCxxFzo1iV8OrHErtNuhfmy15HXPLVENCf/4pXQw
mSbY5uuDRsKmLYqW2GgpjNHUz22PuB5tQR6+GF1LYvQ0oIgihgGamlxdXDLGHJbYfvb8HNbz0IYA
Xg3rkoHppXKIVH4oD9N/bfGzKijqr/PUgcep+ctB2u1rluUjPh3PktrbgFrQzR2cv8PNF0FzWSLI
UjwQ28f/sQ+SJJ+Vemvdd5BY+3VpdvcaSYv2ZeUHDUzzKHbB+hooX4AztAA0QlnFZyHGVAktUDnW
hlYRblXEe9tPyG9tW5i71vd7uVHH94EPt3+mOkxt60oESx68UEFMUttLD8FSHFJtZ+Age3Wbgfgf
OG+vpdyOv16LveoJ2jc1O+9lCHW2AYriDZVDEmx/cYnVYGzpEpkIFUG64gqn0Tim38a6hoQ873vA
JCoNId/ak3rxd0q6/WUtbKJSNDU66sSu9zOEqGBRjjspJI+i2NN/A1aOUdIo3yC7AdIOENn+Z5ka
rHQVXJyTyIeHYaEBTGoCjMrU9/A2Gr/6Lue7skz+jRXiy7KwcqkT5mLZXeMg04lZmrm4eWxnsIVl
LHDeN+PaA42wCK1GM9DQiZQXWRKxZVyGyFXnJXonaADft+kmoA6DNxNfWIVsp8WOvOCBkTJzFwnv
s48XAG2JaJJfvEXlWDOVKu1oojx6cya3EmORPE3FK0/uL+rA4JcA2IpiupDCtJdT3Uj+9BRInGBp
Q8idoX/Q/ARggjyP1zfQyqlRoHAgMAuaZbOkgOA7uFVQbyagzY2I1okwQGIMo8OI/u1C9QILdYP1
hjw3QD99aPbTWtzXKd1mf8D1lUA6eIMQnSpKJLIvJvtVAJVu1cXR1Xei1sJ2cbOn3LJrRjWwFbrL
pKfFpg8RmHN9UctR1qKNqyRJUVNRhdCOdbPQ7Q22joUMykAlL2tLQhNY4BLgdiqhxMVI0fFk/4Qy
hN2bQ8HVoKnyBO2OrmdE8/tQ0yqi5Qb0WGjEiKN+T//EOrQ4KMYwNBqmfrAOemdGQCUjDbcYaydi
QqdQ0ks4sE6RWkeTHoAIBBYpzbQwK1EGG6qpPEvz+0+d3AbsZMKcSWW2nyLG8v40SeTPAgzED4cS
UXiu2Jdlsn0ovxN0bo1xUh++mbGxnsiLXfs4BLfly9+ILBYZQDY9rm4Oeaup2mPSOppqjY9TFCw7
TQsxfnwOZlnpKLRQPKSAC4biscqOXHU6R/n/WvQj7RTDEXyTe3qeBl2FpWRPln2DxaUEUtZFrUCL
SVLSOD8Um+v6lxFFT+jrFcJUX7A/DBmkpbCx/LR+J7J8uCafyh4Pq5X7C8ns73blwzLA8YsoSTzH
ocdVKky89co/mPCY82C2yl2ne6xdpjYHarkAnsX/cSuCmJmCyC5ZLsHCiQEkDngSitMk5GW0qKzC
KPNoXo8vzE6JqgNkGkfYLhwgP4Ts30sI/iTSkM8DMNtZs5VrbKWEBk1IypsMRjrUQQqxEF4P6xlP
YRsL109Kawv9fw91JojT1JsrS4G5PfKaGK4Ck3Dy2bPpmGlhxBEJfnLMSOJn9WzqL5zc433A3jts
Sl7XP0yzO0N7+RJCtCma+fl9On9SZ2AeiTzlRNmOqaFBsY7UUZCEZ21UEnla412XCXO0gW97cc8R
Sh04knkCfas/1hhP2c90ruEKxtqy7Qg4ZEpuiDMGx4h8fEME3Kw6rc00mp9NMFd0M39fcAzlGZ0N
tSPRGtE7R1JBOUjgYfd1ABRCEuZmGYPBoaVGTOxUo5f61cl2k+NS3e9hFL1LpqWKjvN1gLo6heGP
kPD9QzbFxOSqdd8Dd4+slm48KUohG3rqJ6jlSL/jBIlD94zc16gtqFOS8/nz/S4jGNR4mBJXZVg6
2yFv4j/tK7Kre4fp9q4jKsYNKU3UXB4cjc+tqbCDGXEYPfsvD4abzaHCCgHDm4igKJJi5utUkq7m
S/E/kuDrYU9WU5iiJ4koAhr1NhpvOLNGy0PkFhFMaAQI0uMCt87dqk9Utfzn9cEjARGpKikOM51P
ECRG1sIazRE6mfMHlMw7B8dtWWDkr8xkEQe/9HSJcZ0VGB57xp5SdRrW2+Lf0KItNZ8QfA+/V2sR
y/ldA98d0RCTp3BWbRLj1kGfq1k8fC9A0CZOplIqryHk32LL1lR8AAP1yXttXJC3lniZQpU3ExCO
8aO/r5erTdmw8XDHb1OAVFlyhMZxlIweJcMztmA5mulmUVQASy6X0JQ/lVzUa5I0RAZ/a2ZuJjeR
mGnkG4CVLo7FIlqksqyRuJlxRS3a8qzrmZ5bLONhMzNMxR0uqvaafN3LSo9eifpdjPbS1XlRdtE+
HLVjGdYmiTBJWSSgufCkaxfpxBpmKGHfqQ75UuAHo4lrjNf8z++LmQbT6BFNBNMzr4w1OCr0v+hg
rl/mg5OsSeHqof0QoRNcKnKhzYtpo3ztGNpSgvOAOb3fdeXFf9r4M6lv4co3mnfDDtV6P6RKYK8C
m8o4GA0p6MZN6jOOm964v0ttGP6vGPTGrA77dFdeiAgMN/AARqeFDvv81nfTYB0E4qQeD7HK/FoD
Dzn82jmg2uKln8FyBL6ABSw+qSQIa1GxVom4INpqRhp4kXWcQU96SS4KYLOX7sHiq5F/5QygpJpg
1FLZgRXWxObr9iDNUUyjLaI1B6yhWO8+P8dIO0ICVZLR07/TXtOnntSipFT16VpBR2M2yFLaen1X
06z9G7MqyGTUUyDY2/ytLLa5xscgsg937YGDIzuwyW3eEe+Z/blda19BNpp5y2Wjl0azLkVTKyKj
l6/W7R4FWUFCd2lI6v5vB792uYgkTh4EAvfYZGXg0c3Zm3Atmub0xg/54fcHzcg+CaWV67tYUFQm
ifpU1GTHU14rDMtV9sAwVx7CtIJoP7znoEmPPhH5KgIGv/7o4JO2Ni7QW/YAt25NhjkM58DJQ7Ix
YuBBC5NW99chOj8Hj7bZo0HdqiBCX2GZo8cdHEzKNJ5qrc0SIze91yeJL7lmyx9dIcgvpDqNQ71a
getBbleUGJzNiXSDG8ASYk7fVqunY8bAEhNvyPAOtwnT+YRXgAWRz8m9BSj6NuDUOIdi3OFTzOlK
U/K18wwLj7E5/7PER2yRpPWMtjPfdOk2LQRlYhDMP8AMLR9lX1BHZ9183T1gQFSY5dkX2heZR1tt
Dtq82Wkec+uXNKFShXB8nZxetirIUzTFFwQL2WN0xpKEtbv9AOeBuopRjVwUAuqJ6sw/21Pnwgpp
er4K/6SaLHNdpOo+K0nKzN1/VQ3xzBih1F569N0Z+WLtOYrkMk6CHThICnIQc4SQUsREGRRGr+r3
6GId397BVzhBzE52jzKWH2FCIY869jsc3aU7kUuII8VbE0Skh2U6R56cjvMk4W/al/DItbFI/6/X
IGGkNWu8uilZvUnU5gEkED3VoXNVDFKyi/4+Oe/896gmYq+alJ+R+sMhFM1uVoly6UEj5L8VmG9V
ZvCwFqkPiX2XdyF0kQbgcT1FOSge3cEgawx70i0GqakvOHMkziogcSBbqlMV2h7QiWIFkQ9TM0tr
y6asVAX4pc0MtI3XForYKhxpUc2jq9k+AMprLMksej4aVXq19UWbqhEBw2iBnOJJq5bSuHb9FUOz
Pwip14wMFQNeNOUWEd2Q3vbuxKlJf7rKyJtiQX7wUfuS3coYLyKQSP0jY01c7bs1aghnAhaPqBbo
3xj+meC1foRs/mUImZj76Pt3Afrmh4uaw5dzuIdFyi1kDzrnBtHZA5q6eO7coXHOT3YFqBpOYO/r
sQ6+fkiKw7xCD89MDYu+r9eKpfZ/txrkr4GEO40xlfBE6T71HnaRBLea3j5zcphvP3kZJnam+OKw
noYFvKFjCH2VuH2azesBdA3vKbVT4qNgyf9wb0MpbrU6IXOXUKYJ2+jAaILNhFwm0htmHhrzrtNN
PFnV49tF3HE8bgSlKgcLn41nxv17zRXJEiBO7psE7NkF5h3+CCdLXWy042IS/OcWL0bcbD8xQvh4
LkYe9XMsJtVqL4EEqR15X0FomRFBHwRz2/glefw1GoEdydtEWyCzfQ+Fz0Gromm1niEk/xvJt1TD
mONdrmk1YifMnVdX8j4ykgIt9q6zQjnQmPCT591emTBDqgq/KcwaAqLmNheHoxCCvuwgv7NO2o6T
akzYV7IVpFcj3CWoQTjDXpvzry52MutyHq2I2vsvxsNHZouTab2JV5SrrenN4X/OKMXxTngrC5iC
zA2dEeWn9mQo9I7nybtaNOQBhkWBjzFt8IQIy/FvXppMgIeg13DMyuWhUwBTowV6cH3XlvvQrVKG
ySUqp99PEK+l/6RUW8+xjqlmWnkZe90Y2EYxwmHN9FENgkDN08BotyoRD1og9LpKjvcxVrnVfDRS
GUzSvC0jaThasyS8euJLhhquzKmEhLmA6R8xvqEtn0es/oTEeooLDWYbaQeEZmv/9vIeHXpb9Jc1
u5aIzLC85rn4FLDE7nLBGAKEVar0KsnXMUwVuXCJNLTOkNRinFaV/aTxyedatBkFSrll8vYU2ziF
pUkiSVmg4+Jc9W9CsLn4h5fVChs5EFCwhDZGWcEZQMyvDr4u1dXWrJRYKNg7PlR3p5WrJ7Kg4kat
a9ebFzaMkvDfk3tBYMn+xkmnGcU236B6kCq1FcHsdzXkurCxuBbIJ3S/WnYs7xSvLyby2oykqN24
4Ou3Zw8k8RBPVB4hNVNhOQB57BDAh+cQtrIYZzo2gicc2qFA8CjmIiXCFaqMeAnlAzooypZyM47s
sq9nrug6sdA0pVKyYvj77OiBk/bbzRHNnXmmo+ZpqUMoPpuzBj1jcdNmymSCXTbdtBXc5F8zkSjy
TSm9vnRDIbACjSypl+wc4CSnVv9piAesBiLrzLxwhzcx42kIHFIaOcHzsSPa5tai1bgxN076/3+z
9owklBHhDeWAEpWUP54yrMta63Rnol1lfJR/n3O3OgwTXTaqpIH0EOtWWafZKkmh+LtBbzOE6N5U
DWItxT+qdZP2iZHsm7ff/Y1qGTJ3TIQzr0ykWZD+PieDnHM9QRqAejUQi37nLT0P8HLKFPMCIldd
YHgEd9Rwv9FWXWaO9jsIBki/hOkxfnrOREe3zUaecDHOuRMgJZvfxdToncXzZx7ntpTyUbyaICcf
0xKINJCHT8DvAI1tFqVoVk9e0XKkYJV3rCv1fj96ZmFzO5qYGELc5Rw6m8Ki6m3VmUANzCAG2sRW
UF7mOEFLU5NWn14+MDm36s+QOBaea3BkJD7L/Brpq62zzbgWlPgi2k1dyB5goRvbbZWC0SxbEOh/
85cL0rcHhbMKqPtL/t1qsezBzyHvoqB/k0A4NgdY7Ma4ZcdXOHPqy0Um/kmZafnWG/l+bwYO4W/h
SvN4xSFFhPr0GPPKXXWtlTJOYHGogv1w3w0hiYqDXW8dxZ1Uke1VlFHHOo/dLSLimQzWUIG/o8kN
aPtcjRNLOtKKjcGAFxMQ8jotnOFr0GUmplltGld33N7idtuvqDGDYDiL3v9cqvSKPagJc8HX/7d2
E6ZMxb0wsX0zQQ3ol/MTUJbgX1Uhb53s5QJMl7qh3v1fmiElLb27ExsxUbnnkrq8JC3hSWTvmene
3gSUlL3z+bnDMZvcxveIc68nn4EQkwGUYjVPdlVtP9SP3baQijv4lpIgSJV+uOOIC5C6QIQ=

`protect end_protected
