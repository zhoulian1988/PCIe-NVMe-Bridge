`protect begin_protected
`protect version=1
`protect encrypt_agent="FMSH Encrypt Tool"
`protect encrypt_agent_info="FMSH Encrypt Version 1.0"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2017_05", key_method="rsa"
`protect key_block
OF9jK6FaHrF3+0KczNfRRevBO2u7mNjeaGESwqNzuDb71Mj/Wbo3RHVd7V7nPejF9clixjfq+wtB
o1g+yeyReumA5favmBnVUTraoQiF+2+02KodjkZ5FAotVKhXr2vabOjbC7V8Y3C5u8pYaQF1BKq2
gvdczgRD9JhjLl6sI3TpPj4oyN8A2+QJwH7UvWfPYbVdwTY/fiqpyUYmWMLvBes+PDI0xPPM07BN
/WmAnuOFzrRScL6E5NXxEUiyAgUhPPMm9KUQ16V624sCRU6+FEFaupc+7/wL+UjkYWTZx3tDh2ZH
H17NuH1iPQt5Emmun+bBM2WB8sxZ8X2x7cJuZw==

`protect data_method="aes256-cbc"
`protect encoding=(enctype="base64", line_length=76, bytes=214080)
`protect data_block
4uEfULHnBNuj9+6Njl7KX1OBWCqnAwubPyZ5zmPV+nJdysSaJdiKqanUyJGX/moPrLC8NgxGqk9l
BVXfPhPDfzH3OUA2nqpwV8Ub1hcZYpBaMrOVXsftmaODWCm0VP+4z2pPEMdZzotWgFEJ77GkQ1ur
Sa75+FRySrtBW31fQuBCf6P2HQZJGUcBxi8BwqLfW9aA2f6tY9e+Yu/leEEIbqhgELUy5jnUEqxe
1gXQeFe66Bpk3nlUhKITLbTxMOb5M+74aMVfiV1qJjV+semxKw2sko/EuSaj6888M2gpbfO9NC9A
w7FjSrN9Nifww2JAn2rqm4rFzaHd7USaiAVLEdsuAxEV7U4VTsOmUTlvn3p24U49uSqik5kai7RL
iTCAqqOcgb6eA9RJyUqktuu6NnY8kcj6PBX4Gn3GP2unS92UoZYqEU+FDPkxYrw4BOUW0xJaHz12
e1VUDd225jhTR7nPaRpetc+xymJE+m/A5Afu+vF5w8lfVFh21EPB4Se71LihLF+asJnvYoWpT/IX
mboLfCBeFuU3v4UOjERnrEvcmfDSKT2zkzbIS6+Guo3dLhvGUJ/wjJnOCzus4Zz/qTVLWy++dHro
HBBM2zdKenXk7mJ+phiAeXkfn8Wfmrg4eeh8Ux5Ng8bHd3rz6pYQUGTXEaJLdDEqY/bYLub6NIZa
tgL1VMwzl602v++6T3kRjZKY+Y1hNd/MwIsly2jUSXn1kqw0Eq/+6kupc9nItIQYnYQOi5631WPF
6ZmhXbx0R/bVKeKWJEV23LeHT4TRWo4Kug/4KqMwC2JpAg2kYjJ7Rcssx60DBe1k0G1xKQxEXfy4
6RJCBESWL+BTbXBouA/WmvUo4qNLi8Yv3EuzzbXlb7vPlAYRG5lEHLYMjAM1kHp3DSgAztg5tp9f
v3hybF+U5/HcXxGsc/0VeiRrEuzHLXwzuxT7AS1Age3MUig2iG2JwMpFsWzJQIbrKp2WHuN9CIAv
mibhVDZcqQ8NH/sgbuOUpVEjdsv8XY1+TAs78UFrVysW66uUaKva8ssIpAo+Dx6sT2tEwH5M6mM8
0TCoWv75tgHEJgYB1p+mTjZv6ikkeX9qb+sZLzCR8CwHTj2EDzX+N7DLBJQYyJTrJfzXPiAZdPnJ
zRGNVW0kVyiyLsq8G6515zhQi/CMuwCc+WVV8YV/byb2OaAX3PLthJgZRRC1lhF+sMRMrzpzPpau
okA1NDaGGWXsZZuTP8JKo3dqGUes9WwvT5MC+X6PMbK7oPz8seOqWYewTbjLxClrE0rw9Ijj6lNd
/OK3O0UmHgz4zDqLo2lN5t8SwFx7JB1WiUQ13UKHy8HKRjs7aZU2IKASHMEIVhqbkVhIff8c3pNh
1VfyX+XH70oVSIHUkg41snhZpkAaB6VuvQhvGC8x01yPQSFTcXN63mfvCSC6TH2Bw8XGQs5VHGuD
W8NvruciiLuw7JyUkmEU9qXndyDXeshQqkFEOSMSwp2OeDt4mmf3ET/jH5kOVPZyah957HgUy/Tk
iJX5b5xu6a3jM2/zf+6J+pz2Ye66iI20agpUcGMMPdcHUkcI78sPx3lxBTkq9OSMeZIQYGJuG3Ft
vmUeZ9Mw8YcngQgfMwAyKgrYAmITIB3sOJLG2vQK6T9pDoNndKZKuRtwgGBowEdIpHx34Xxql1Io
uUfFIjiyC/eM1OtS+OXCcMoARzRmNPmJ9PCqgWDV3x3z56KJ2cVfwRsAMR7RB7zew1BYNyMxLT16
dnJ3vzCrncx7dQK2oe4/7zCfXvoMdo25I1anf7IjU6WPOybBVuH1FvdbmAXhXqI1PAS/KJWinpu5
84pvLSi9O/tIeIB/EBK8v57QCBtr695FFdKxwUVer1C0HvPek3rO1iBBLTijST94mFW0YwZlkW7f
8TTLhgWn/9DeLIiexu6/2+PQldr74s/wQcqqiWJtOVXyutDNBtHTTgByfeIkJGNQ/wste4Lh9myI
TQ3asrv5tyoWJLyizv0MatKbOYbNI4lOrji7/azumaabjxdesk8JrwQkaae7R9+ZeISIekKWM5UA
OqcrNntbvfTmVTuIj68LH9wcXwj/7PfFKVJcE7BaWpjN3J/8qSwCUIQkqUjumBdxUoZ1F1kJATI1
lF6I30/1iGfUcbG1GqHQeiVnlHtW6pfFQjrlG9Hta0g3gSNbIrknCAzEV5uYTFtaJqJS25ccEC7W
6ymzlCpuJMat1RIngx3ehgnLaiY3F/wNdRl+FY4Wn67kY1IOVH8m+A5RcT2cjz3cFUqmMYEH8APK
BIJzljPTnADXCqL5EwoqKSHyzmcT6If6o7XdoZiJguS6mmTt/33zNHzp+GYbWY3bJBxudUKnAYvQ
Zq9uamhILf1w9lg9LirUOTd9LBpXvvPsE95XcqCOE5uyLBdy88Rn/R0usbwZxFIVrM5/4FdMFrgc
P4cf+t21cPsk9F+ktM00bjmwLp+6evcVlKT/da+nr9FJ5+xKAjSFnq7Qb7EV5hoLDze2LjafRcS4
BcRSEyUeqAbFkwyAPl7fZfts46J6Eda3NuSVjtqLG0Ji0oUcMS43Y4lOHH211bGKiMUrFnt7V0eq
K7xF45UVk/KFRmvvqGPhWXsY6jQmrf6tyOFw1EbbsaDxF1yAx4Pqx280a39tbohQGwA7vOGBnrF6
FqMqhBoN76+4nJ+V6J+0F/WMirLGSub/sRIYDEp4fsZsEcvfbpPw8B/nnT0hSNZ9bndnOFfIoXiW
j7kA4DrrApX8U2k6r80Tj1KL5LzMbexWwyhFO1+kF4AcuZfGhMkdsdFEqB5mZNplIQcafPBIVckT
V2q9YhAhlPpFN/LwMGUmmbtx9qSniQMzHvi9rmBkaaRHcwTfDlrTstka+AiWXCmH/7JCcQuCw0kK
GFdJayXOmUcrIjYY19KPEOas0qychCPEQz680EN2PFBJgoTJvK1Eu2VenoP2xJtKw/7o/D9KC+Qy
eyWjBP6Rkc+2zaiWo1/pSt/ivjqnuTLw555GTmrfuk0DTX4cdPbBZWvUIQ5IDt59/iVztdSXUpLh
gQID5sM1iifT/dMlUxVV1OCHo4RgQit9n0gAN0T+LQPyE3jVnfk9TB+mdtuiCQIRFs76twwACpTm
WrS7SrXlTBPaX8D859kqhIFW2tu8ApUzixBEvcM7dBnvhlHWvx+5BVGkFBq9+3e60gYhSk7onSis
y5HOvYwRH/MwNZfFeDbHhbtNhx+d+VHYw0Xy4q65x3xdh9NhYRjLEGbsMC9J7rXwdk6jq/h4O3+m
qPLKRx0CylUH7FPSlQ+DVBgNjvuEMqIT2zrup//gJmcd4D6u4NzWjp+v/mg06yv1dpACBiUAiv1y
rGjfLM7UcuFpQiULCLLoilOQzdInrsTK/u+V8BRIrlTWraiURY3vWAewRjl/eGEdf0UDM3elGj26
QmO0P8Doin1NYhxyHwiy+jlmLI3P6tNGYg2aG0Bw+vtsHQr/8CwHA54z6FdPzu9lK3xvaGgV+kP4
dfSddbPi5i8oGWVV/H4wCyeU2nPbK6VGGULUhR1WXvSzwu8qqv/jta7vr6vutHmCjmODR6+At6a9
dHUTARQV/YXpsXeuY5NANM5mVMtR2sasQwygfWHX9XWJZESBIC0t6TAkOkurTY1UMaMnY/b6sGGi
al+7OG5HHGSWABguC5fy8fL5TPU92CaEtpxfug2DBIKLd5GKOenvcQ0DQIjeFZ636IWClFIwGPns
hBrXn26nPFlhXJZ2fpbIUU4g0NTc1PIAffFX8ohxwfy/N4Yxqi/jfIuyidmIfvQuSPFl5qGiTlke
vWEw1t1q3A29aRL5Xa0OKXQLIBDUCdbEir3U3Ne83FqYqy1QuQl2YReTSeLTF5QhApAyCZahp6/6
3+bDZ6m6l8NRoF66E+WHgHwtIluRaMenIDiU/hhMVnUm/Wr0+EsYWdQJFnV2SchqpXjmuS+L6c8w
HAXKVK/7d7TEXyfXyapATBT+TzPSz382KywlDcICUriaHfhobA9DlHNpC2UBLhiuGz7SAb0/BhK0
UTKWBEjjas7RG8bI2605iezicfq/q/ECNVknBXmCzJHkWnQX2IYDSUDiEInppP5noJfWHbacHsyG
uA0fr6kQSZ4076AsPpc1rFJrmIhHGxhLhPA3XY/s2zVh71CS3f3sYqicOk0S8Jd2OBnXdlQYdBCo
L2bm9hI8JkxbdlzS8wiAbio2yCDJSM4nuzG84Ygq6Tbkfumy8FK+UDt5DY0NKROwtIqd9UgLkRo/
0I3LqwNoOil4fbgmvw+j8nnlYlDyESyftJ3jrna1s9dn93n4dKchw/eGS4WKOkKoiMH9iySbEcFL
YHjBQPOm0W27N3Rx03xcQPLoIPPs76SwP0fFo+UHnLWWjbg7HNeMk+Rzmm+4URqMsZIe3UyJr7iL
MHbU/cr3S7vPZwCHe001Lahk1IlUHx752M79lSRjZS0QsbofrrsC+HlAqrCU/ijE3Wz12bIHKGpE
GkjrdrZ460ICL41lH++aJT/z8JPf3xmO+wSnyDroxJ2FVg9uiRg/7vcXG/Nol+XeOGCU9GM+tcM8
bNplNX7XoSfIcN2oFGCbqozFLai5d4iFIdD7f8iivxt8kIiZ+GK/HPv4i4dQ+xD5JsBqFA0jafzl
Gr8bR7/mPlGEh7lDIYVNNZZ6XO4qdGBobHi3MIsBsE8/Mq5uXaLkoLWCTo30oq20/vzp+jPjI9R8
8labRp7t42jT3l5SV1wGNTu8LyaAiKtancz2ItTI149QlzZfUCziFRBR5C63zDhJxHv52oBMGCKS
ncijjXEEeGApEEfIsRA9C8cTuUES68xs8NSgcsZStr5hFNpfaM2CkpVyAew7ceHuwuj8Yr1ISdwF
EmPjBG2YPOpgua7Oilp5pTl2A4fwZ8l8s30N7+50IfXXpf895D2Kh6wFgUyumPFbgvSc3uDFQm1O
0Xx4tBCs7vbsM36YjrcqewlXZcRUkUw6FBqEiExvtRzF/LArHZv31isD8pBI7Giu/Ci+JsPuN+Lr
2mETbUwcqM3HVoQWlzC9Y9bUaahg1yYVeV2X3AP4hzsz5U3lpKryQfPihXtvchQXEhe7qURYzLNW
BVaVnZeOv/pXpmdQptbn5HFr1Qat0le/3+6Su2ImQFWSCEUFx85q0ImHAf11O3rYZTlbxtV14CVq
uLnyTW4FNzgU1E74Q3CAJ6fJ13A07xGOQFLno8arv5EVSX9FSXZByxxTQ0XfwmT++KwfhuJouliZ
Ry2jSBulRyKU8FMBFZ5Pr+Vn1WMxKThbGsXOh4Y5pEFdWsC2F7QXCGZLJdeGclWXBTJzwi3wJ2T7
aTNNr+V1zkaKHaJfoTxvneksQb/lpFNDk8IYRhQ6zRXrTlWsSFb0xJpp/Czem2judWjdfWrUpcWc
TwvB+xGCbomLLu/mfXr1bV7C4lTOWkXv76HUmmoZdaf7y6aIJOcBmxBm0NhlBO2FdygDGHOrRolU
QwQC0SJGg1ha+yb1dmAVJv4i+zEXKzs7gTOpNPk+JPBnM9Ffe8qFtkPpKEnINZh9vk/9Fs+AgGWp
ux5ChoNoGqdFrjBy4t8EXipXh7dnhNXssZWm9GviyVFv+RC369HjZ+XIQIkGF0B7OfwBaVzDECfI
QIF8TQMiY4zw3xcrMO9rn4NA52Yo2qecq7xJuooVfuJBqU3ubX85VILG+oE1QWft4oxP0jpa6kEQ
NPkcNXra7mrl+zx7vhD7mmh9SeCD4PdJfTF1rYDI5EXuPjX21IJJtoFuqks6zpOcaf3Key1HE4Uv
amMjpVtGW1Wk6Gi6YY3miDKiVTl8kCQun8HoBs+J1C3oCpA/TU4AF4Py8dnqjad8QncTfPMVQor6
XQjwFsdqT6lYcsX/uYMcz8078DYmHoTklDK7TxW3aoAOTGa0B1YxgxStBytJ8549pwsYvtv4LEhs
envhiYaojiJUaZycwMfjc5L/w4vQWMikGKSCzpBAMydOWogznLdtJvS9DR7RovOnLinQ3Exb1SlQ
ivwJTly8FG134hVqCs6KwsvtqAYhfYZ5yfkJFIv7guPQ1M1CdE/nn5aVOHwEtiPZ9/w2i03IYYT+
btmrWNXAjo1BgnWGau9m1qyTR7t+L6VfcPnOQdYQq0wQqng0saT7649FAsHPdX87O6C4GSNa7DBD
K4f+BzvpMu1JCRqUttmhHAxydklpAXy2029jqUXM0XwTJ5YCSuqWYiPIrcePjlPiVr1bWG4FzvrO
C5WvF0+oEBpzEJiKOddq6J4SMhHKLV3PUMWQXIKZy3M/IbwHMkaFUjAt+my3mIwNkNDyoGPpe2v6
oJ+aiMECaRe5lDhmZHJUvgYBxW3abpDOlZ/+iZKTXKKhblSUpqdusXHTm3WCy/saggr3z+VajZn5
5pHSn1AbSPnYb8RLn7i6IrTcU2ZZCQ4KrL+40szSSC1TYdqLCz+a6rRl0LbEztosxMJibiWDQz2C
40/n8Gw1F3a0d29bOExNv6IAh5iTdzm4gpR5pGoOy+NXqhsastWd7wfLWu3qhdPM9yccIuFLVXb4
x7t4gn63oyUkQIUgkfDystC70zZXB8vcrnKJiktvfA9bSJ0i+qaDGgxAb25X+S1BKmUpxLcB7Pbv
GzgeYVJI1C7SOelV7KLlH/GCv8zjlJdDB7q5WLGl27Lr9/YoHxrOx4Rj2TVR0oTyHMGsIdw49TBx
9X4ZHFQMtYttehcCEEI3uTKYNcbwKerRuYM2TnD71xko2IW2RSf09XocRXZWNmhIEXKiX2u3J8oS
NO1mQeN7VzNUbl7rXGhyoZT2D1Ib7ptY3+3GdtzR3wGp0dPKFCsGa0Z5ghpNNbvM4Pol6OsEU3Yq
3/J8FRRRYChcwQ7+ROsgrtbQUo0kB5S+uSbGZfDKTuX6uT4nvfkK6LmeVVyUofp2edQiw7/5CYTN
jpEt01QAnabm7iu1FNyGu5oxdqm09Ju2nNRw0yHqX10a1pux9qlyqiaEJlL9VaiIWk8vKX7NZG82
8SIOnyMAEiPuBp7AGJuD+8Pzc8ZeMEfUAKQMy9Zx6ZmGn7tue0tcMDCtE4lEXhGxMmnUNmbChsOr
6er+P0WGnfOTvaKIfyQGjh4pYUlFXi0O0K/I4OXFqublJlG1if2rmv7bJSThiBZlWTV+yOvqbxyG
Ok9CJJHrVNo/Q5yz+/cDl/5GKviwL6qyr5+mv/EhqR7gH/68an9uliIc5UqgRYV6GR4GaTvEQRej
M9a4Gk/i8cUhdrHx4HCglIVlfcW4FvxsXbO11dwJWkj5jKCgMSUEcb+rcS2FZmawibQIGBM/bS+X
TZKPbcIGECfLS44/ci6UwoP82Ebehj00SiqCn7iUF/kX13gJOyIJKm3LbPOK39tgHk1rkQaEi5l6
HI4n4dINd/WXM90s7vQawRJ+HnGDGfLl/KH4h2zcABFrjJGb2dEV0P8ZuPOYRY6k1XovhzVazn/w
gF2fmzgGjT27yggqy1/9uR0TVmr3LbsVc2VdgkiFwVbDQceqEMwmxDrx3NLVKygz9I4y0vgN1F/U
D1uIl+WnpcHdbsSa+RbeIhD4GlF2uWK9ORnv7hfyeB/huJWhWUgZx7y7j1PwKLpl8AyGPzs4A0Jz
RfB3HNKz5isKCzsQP2AFHl1AlyxY2bAlw/s/4JQhGgWCx3vrxN+d49aXgy4841yABcLFrdrPND3x
cp2kYatqxehpNt/4/f3E+4R0pANqhhZf820zzHWrCzTDe1kgTwXD9o28Yxb/Suc6oDqdWo8OcRDz
UL0VRQq34Qe42RFgkNaOfusSLF+gOM7JUnq5bxduAnsBE/SIrINJ5apnZp236eOcUvjtIVOjXmaZ
WiQ/gtKnR+TUBXICLAPz/OfBn5xBvYuSs+8GVoa/IjyyL2GVnboFyTIkXL1oTM+KJ7+m65qm/pqh
hcE7ZNT5IXvqPhnH/gnRB2dutgs0iUbfaFnaAIazsvl/tBaXx2UHa6CH+mE0DEnz3Mv2yYlC6s8e
CUvA8kP/2SV+4ENC7Zzrr4QfyjkjMANa0Omgn5HZmGbgZafnG6aqkHcf8D2VsnwyMy+f26LScqNI
EBaJgqY1SAiHzlUa3dVazaWdpvXuCUGF/T1NdVLbSovLTj34DQE95tf5lypiEWlTb1XroAvg4zMH
o0Z+vGKDnlUkSqdtSGM4y3ybqU4PmBP12KSPzzWdzqHmBvXN+jYvZvkJovDXMw+89TKmYb7KqDxt
Cn/NCbvmmYlc2XvlZWFGf1yhqUEUT0yN45Cns+6//+u77N3f6F01fY3tcj4AUqJb0DoQRqXAFQ6k
k8EtZihqRKXkdtyK20UdNyCnDftZFsQ/i16N55TQew8znsAjzxcb1JYikeiWwcrSCFrO8QhQLGrX
i9D+J0nz8UKUrXoKIphbOO8gV5VObkj8qUfDr64YhZxhKCT3tBfLy4KuhMjIF2eUZCTf5JbRnDNC
VNkGvdpLNJRaBL8L5fDn8rU3dtW6Bnk7qs9sVllS1ZA3urVMYsrCqcBafZcOeT+fvn04d6y2Vv1H
v7WlJ/LKHp1SLcC+Ygq4yOCj33DvuKGsDvJAkCxISGVY1qo8an9GI79IaEghCohWXl02wjqWkd3C
QhGhNhXox30ebVBIfRihAKqmTx6/qbxV+QdpXKWzdJ4JaiLojo3MdumNvMkUy4OUguktaOZuq6BH
GutiUjhf7TpE9hbc7ybKU1BVclqrMT4LZC0fmXIn20FLk68PS39mXbU5EMZqsogjw/1KOe6C/Nf8
zxELHYgZfdbaqtnUoZZqOZISGeSNYg7TwquS7pAD/EB9lC8wjaaGp/h3NDS6IZGX0qcdhCKyN8ha
NYxGvR2cIWc/kmQO3HSLrKFJ2D7revCkDJtfBuE17XxLyoe66JUq3993DmeqFAnW/jsi6ahe41jc
KAr9g1Csx03xN6/Q2SApMzoxFCaD+rV6yCLFWyMEaLUXUoa4VlBZ/7RLMHg7Q2VSATemYBU4Y3uW
eRklDmd6qjwSI69bSvwwABC4+V57//7QNgH9ILOSw36e3icUIZXRpudjb9rCeO2Y1eM/Iiuwrgoq
hHaj/BMy/XZqZ47sBIx/J0/eq/ITKD+/Lsn1OZZXZ1oiTtEkif3ALotdlBt5TpKgSXkQ1nSNOBDL
T1FLIt/5DofrvJs8+ifZnAdtglkCS26055f3hhRytQkZgSzHkf3ixY7hZlWCcNdYW4jQNwZELLUB
Y4oRXh/OQycrad5kGU5YDyVAvd/OQaaTm0HNv/wdaV/7tBPcAOT+2w5oIpQtFGFTkT/MpwK9XRlU
0ZIrKbiJxAnaohcf3h6JqNKdQh9+KF8hhePqF0XM9NWBNpYmrEBMnCA7bURtHEUt+ahe6qTBbn++
pJt6lL+CjVqPd5266O7HIrLf3q5W+HUQNovMBU6dDQYKr6Cztt5Tnj/98kcjySMJvkpz14WSDzao
kk09JO9qQqYrZKBK0yxKtDkH4JMuHpynamJ3hQp3th3uFW9GQJWhHnC58p5aZyB24mTRyNOD2SmE
J2ILNPRa/sy4QtR7sUy/Ay6HEBQkAJ4ZJko7crC7KFPzuOolbQAoOQuyE8gJSIOBNk/hVtzDmMT5
qhDab73U3P1y8zGKt7mqW/wSPOTRVULl9TLqSasYkJBaBO2Bdhgl01niyo3HK6P5lwQh/tafZFl2
TnxoOtyb5/XvdGCMo+TY4iHK7lNjJ8+3VeuVX1iNJ67pQTe3mzx+T1gk57HE7E6f0eBvLiWAwjJX
5rv6A9kd8hypJ/yIu5LYxJtFwg9dd338vhP8RWtBn12UFOu58C0Xi0yWwRsx3+ZJTw3sHhFGnK4c
/zna2OLGWr0ohcwZZrsGBPfxUesqorvWiWK7sZjPOGc4waWfsmcj0MxhpbC4bxOlmCvOR5mfwDdn
T40Ou0DPY4+uC8pDrdSCWeqYSJ/wJI8Jp/+q37jvp0/ISDIkXn4lj2mE/tYDHRJJvvkMZ5aiDNi0
FhVSh2qpW4WGvykhQSp6TvJP+Uj1GSJzH/hs91mxc2Nr6mXYBcN6M+UVd5JQ2sqlaHgjNn6OBKhs
gSfvInA7+XAHQTA8PIHt080dMy65wF8NF+TrbAq/rMRClIbUFHScoIPNjdEbvk+zRo2qfGiXb2nL
JR+XMPlVOfzzR6OW0dLFM7FLrrcVXAYL1rA1s2SOSJB4ZEZtOV1MHXJOkLa7sVld3/3Sl95D90o9
dYc4qa8rH81pFTXmYx1XpCV5WYW5arI91F1POMvyzJHIOz7SGgYjsoTBP4KxgvKWR6nZ+mmTd8K8
1tp/XD3b8h+u5rSEwk1RieldinE6q07tQ0C7J5w29Pw6cjI9CwAW8vjmTWp84aL4s6gYxg5eM1BQ
+CRozGZuR5LqJewCTOwp48BHs7ff1xVyHRhyWZ4BVPymX/r4Lqjw4n/jp+bPHH9fVOLAm547oADB
p5DxO4fsHz9BN7j1RCNZ9jvYXBZqOR09yon0zT7SZnBqLH3iWhzhUnjLRD549UZg6qyeRlV1aKH7
hWXsfIFoOq7oWvK+PRRA5onUhFIkwJv7QHNo4LloouKOVSa3kpsihunxmm2YgO4v1vysDmZjl2Uz
3/6AIJgyUJKtd3NaYzukagg1nbZ1U/VJvsEctTsIf+/WnG2m2a2MYN4TUzk16ES6zQiMIDd4kR9T
7Hxi5Eawxiz4lhLMRZKLfl2I7ouOZ3ExnxLZX084eFo/udLV3E4/6JIsm8A4h8prV2eoU7Z7uFBm
epYOQI2MFnwfU005UKXXvCi6erMFY9duJtgioyymP7dQcQg7bnaUOAgkOb1nvfcrEUFo8/eDln9s
uANRFIlbCjEM/FuFI8xNvjAzCfM3NPJoXA3s69p3ckKz/mM8W8dSrkqF/pzvk8XM53zzLxQf2oek
66l1uxOL7krdzHKH0ndTqUjmG4yKmkxviJhFxdfLWIzMA5D1dkVGZ90BVV3muefPQlSMIUg+6a7S
YPYVnc2Dzbm0kR+dUVYcHpDSU32CjuMg9iS1z/2MTJtvayPI0rfy61ipTPzcWSsVly0bvTmoS44w
tPosCk0F0P/56x8PRVju8oJ1WxE1C6qdAixK7EYiRU5vaKf7CM8i9uUZzn3O98x5r/kgkBTHkcX4
aUCwPgk2jKFGqPiy3RkWYaafldgOY6QUbw05mLCBn7V2ITc/HhX4F24KKA2eWRdOUboIf/KhG2hh
IGEQet/DneuQ/lEo4iqVjaFJL0SjuQUU5hfF84PM95dhc58GHbdFGPIbwSvVhRUtmH8lJyKl6kMr
0ZaWTDbggVkt1TOmv2+HpKyEr2V2Te7Xa7+0hPRuKnUPUUY4Iylv1/i0kz7jznPAdZA2z4nN28OJ
JniZX8LuBt9EzcQxrzzSd7P6hD2I0fB+7RkEFRWfooq0xQzH7gcPsf2gxWaiwln7hQy5IrJxgXwU
lgrhIZadBe7j4kOcTv+fACEH7bNzK5AHohX/PkIw6PS7chb3hZLLys/GwhswD8Gh8EKTJxzM7vTW
Ytp9y6kCXj2TqIWBF6KpVHvaqJsEfmbd8P0OxEDV04L4gsUcoHr/jU9BHTMAB0mgknfVqIBxAsqC
2nJNIxTjN6u3ggptHFOWN+yWMzQj1U9ZWojX9hLfWZrDFnDn2hUVcTJ1iWDL3P7245V8QeYXemMk
2Q8Sq2/CaArUvp1M5SvctSOL/e8UQRmuHDGsYlG1/GeLoACMKJ/ghuNpPQuHXh0yLZpxPikk2xFY
Q9ycBOtzkN7ppcwdEfGFqtpjo3roOBCwBMWlhU2uhHA5gziuK3R5llkSG8hneQSwO46+fRwMEZPe
scGVm3DaYfvNfDbd14e9vM8tAuWbiMlTklHyHikMKRYlE67dmVLpqK8ZxRirFfqsI7z+iwIaKphX
v5BoFy4LcEM4RgQG/F+XJf46A6oV5ZX53fCcr3sSWKYXQKT1hH/27/iumkECWAWY9yiK24RcaHE9
lwNyqNcdP6bP/h9cgzwg6ho5632PKRCqCm4KneucaL+bhNcN9gAeND7aQJaTCV1oAg3HU9EwquzL
MQG+RQ4JSmnrkEcnUyP2NTP1s8eefVtEoSwC0UuQSV1Qdb++y3V8tgZxP55B4wcbQ5VoX/Q+u9NQ
fJOwVW2PR1xX0LUhbsI09Nb/GkWK4dk/MWvUIURZp8gxPCFmEO0p6YC6UkWlAGXK0bJyHnWFsZg+
75Zg0FIVe1myMch0u223fdxlH5uy0Fvw/LqziGnQgn8p3L1lEsjes9ipjbnKmEUVby6Ai4JzJ6Or
iiv6kGXEC8EfHRFiMbB1/i7eaWyy286sJq+lZuP9BRc7fapsHTthos50mGbwEgS4K6KRJ2nAtP7D
G1+eYE68can8KKz0NUyQCxsHDqsY5PiPTfYlj203TWv8RC3r6ggMNCewsiSSSgS3rcIRVEviaLKG
4eZoQ9LoayxnIX11fB5LMOy+ZSevZ8KX3Katg70P0BILWr7QoOiE9Jsm7NHgZujnt6KqQSZNPFFe
ElkDxJ4zw6h0yV1vcoFVmw1Fmg640cEXg9H5CiZqGxR3zE3ChakD27NRaTDmPRQgP1y2uPyf78q0
g1p/wzoLtuPACIwT89Ky/phYQVp4JnoqYQa/k9+9jC3LF0Go+AZsSrZeuJ3fStVvQgD95hYqN49a
5Ev/QewUQv+TYJ4zX0y2FsrNN2gLTxBdGE3L1LN3cNMIDhy22sOqBX5Qp/awnG+DdeFeIvHuzJ57
ZrS+bRqGHBYC0P1gC32QLJ59l8gAErdR09c7U0TJSqCu4vq2TPYdv2UACvii/EyAASf8imhvarnJ
ROX/M0a7PuaUEtFG+mm8kblHfHIAdzd+kqfB/M2N1qVCou1PyXpvL6BOfLi91J2TkKJwrFEP6Jlh
MExd5FWPhQprgO5daA+hm2H2qyh3IUOU+WhzMY+FJFzXquWZ4CGOdyZr1cJvy7V6UlT9jsEsMqDt
fCivklJoqQQR4m338EJGIB6foromCtP1dl0IJYXutdkez1rCxlAjUCFscjhhNQLB5En5+waYyTdm
jt1UKfI4Pkaw4vFIVjQtxTUWQwIkzVrSzCoAhAeuHV6o7RTT/kt45ktdJIU7xTuR/VfCUnrwUgaU
t6IVP8ICBcoRtyHm+1M+NPkfjLaflRdj8fDEzGuRZCvQ3Eq1Xp68RJMvPj02W1I3b/+XOd1wEwmW
PkES8/W9QE5UYRXFb4nWH0KcOlzfOwsCekLlhAJY3i7mo4aViGKbDYkKu/3dmxMa689nTwO+8ZLe
3tY0DWcHBf6tk8NIzmfBnInPhgqhvWiz/3TP3rB8U0SOrm6oAFO+CtCKttZV/SUp1NcngmnxCs24
9UYebDwAKedBK4l3KlYCjJomBxxOb4j0+SBTGOvDRlFu1VKo/FuNjQvBk/SKRm+1XhxbPYv2t1Mx
IyEU3J0+nGLPfRcsh1TaQjs0dRZl2Gxifa1mQE4vq1cKSwd6LPbwzUl3sdkXnUVdwenDfwjO/gDH
aSCgyBSNK5YuP483bhN0N1mwmUcf8aIVUimzzspxIWvx3amOC2AKCfyceOsDN9+gY5QYTVI+Pjl3
z6bZAbiyQ8iDgiWYeOGAralOUAFBccE7ggyQSvpOKdmgWVXE9kKWt7Y3BtAVUauGpS17NL7Focur
nt/XvsvgYVOxFsoh+cBeQ9HM3kgAplpQUgmOkubKQ7DzUvGtlaP+z01748xeNOeu703hrWST6Tfp
0yLu+tQ6f4DkJxEKJjicierwbMdd+xD4KQamUXy2729KLYt6XkZ9eIM215FRBWwMYzMB+VYB6uHn
J2fsRFMbwlTnCCcRPWGjog6yLcNVN8te3fW6dfPUa6DX2gyfLuvFZXesn1HLkjS71fEX/8YTrK+D
vLeTbFF/sNSpiWUuH0ZXrQ0r0xg01DALxgN6UAwTmJQKz6JaEkN7uWWq77Qt4I5iaQPK9NK2Xv+L
vgTY99OU/Rt0l5bY4gDBxsv1MdIkH+SruO/JQwYnPfAmDeak/T0g4y7UAj4QtL9Hpsu6QrXnr+M5
/bJ2JcNaySi6t/CTJ+vsMhklOoGqhlDEsnKkOL37aZ1obQvikbVe0vgD28OS+cbDpChZT0nzB0cG
ANgxG31eKxOgLsGjxFVJxhRThOWxUewdnovHWWUPpXCpqTDOzkyDitxkRxiRRl8cqGPULNH1LIa5
8ZAmITY4KfwFjl8fpBCX9KWp2+6r1Jtyu778TKIp1gGi3foxhg9fmjYvwW1wCFdOyrqnnCtiFfoE
r25Yh3Cq6g7Da42p/pKzWaODx1sRDvMRShYjxk/YO6FN/xo6ZuQDIaSkbciy3kReCzHaeLVG+wj2
cwDRD6Yopa01YsOYssrsRl6hMtpFK3PI+UsMJtcZYvdyQ0VKOq5FkBdXwx82iazfd9/bQhtqcmNn
4VQuS68WFySs/8w/qNAeZnZt+Qyf5WUOG5yYsQ4byRrhAlcCzEimEwjRMErGaH3uQz5WjbNKOPoS
vZrtqZcEH64ZzligfgCompe2nE1hPL4h5EOAJJYVIreQW66N+RFYkKMXe/Lfh5GG1IRqQpyofOVN
coB3CvdVAXDAxcQYjBEOx4IDB/m+gaOlVroGc/FWr2VSLhwtwzWihaJx+2LdRF4XNMT8Rpe0BHDS
bQntuZ5o5b7VJ3I6vVTDDH5++cBu7W2RIG6mdbk4BuKPXcmw6XLfQetak6s1vbQMKlqh6UgH88TP
E4inl0UuN3Pc8CHIc+YwIXMF/ssaLfpicSH6iXGLWSuZoQfqGD1u/zyVq9f7hzsuJtdA1WFAxZXw
REOm3lZ8lqOySsdPhuRBdVjX/HBjczE+u6xPobU6z6Ls70pQKVz80oeO+ynSXBuFwZ5ECbIn9U3M
idx+c2UbYASJMOjhvdW5Q17Sevhs8OHfPtU91zUJByyRo/DjVvQiD9nf5DwntexLj97YyinZDp1Q
ZE7ByZgKv1IRUIW1UkfIeV43x+AFLIg+4xn/JaX6C0a5xrLk+Dcj9EHMF/JnfnjISN12Xk/vcwij
pr9F8VMsPg81hSYh4V5M1s2Uii7Iha+eeZBVOm9w4EkHiBXsCiEgRLCVKzr7GiGu3QUHupuKIfoE
gadL+5s81ddETcDkgsJScBfHey/rdgDn6y0cbcnBVoeeRDQEomznabehKNxyG/07eyZWS4Gsf5/J
whN5uXm1bm0rziv/D6dw5+Fa59FYHhRQGYor3T8rUbLxclgiqE9RhDZN8mBK7esgF8dMebe46520
ndIbtheR+dekQlGd/foNbX59dec/UKd/D5qohbkEqoTysXa00mBIhe0Vc6tGMVifuyGdisb5Mlie
9z0MT8EqBzvlsFuT3HXIBRNkPBhdWWwsuOUgW2C1Mjlztz0kA+nWo3g4YScetCj3qmAsRn+Z3ANA
ylGQHfAs5qyAR/RmHUqrSilXZ3JTa10TpAH56hK0pCRG06nvvzLats5l6W/Arp/zahoYKEgw5YFk
xsqsB5BjRlwjyk+jbO1Gfxe1KFHuIykQ9l9Irg2CZIgFSyxZiJ8I3UhjcrhrtfmTtOuKWs5BlUfF
57FgnUqt7rN6us0Z7L0XsD9SLNKRpZb2hJaLC+M9uiSUKWaIvG9V71aliD01s3nFbtNxGZO/wBEy
k2QPOD4pjeLBuWQXmCyRpdIDKbMjocpHv0rMsTHjHH3uj0pt1BsnMRd+5/7qA+PG6j5/aIyzFZ33
y7VKySPIEu5Wio3h1aYSmRxUfeGS59kou7uvOUsLc5oc/U4++hUwFxAFiZQy0s3VhFKGbGJvKoYY
XCnXeHqZA7L74ksP966Csm/hgyJ3m65sM7xSwDps75cfw5AM1b7CFtbnLKtmRFi99DgejZiNn6/m
oUcASFS7iijusdmYCQy34VUKDlSHAVygnU9Exmzqf5eAMj2lqluXsOxK/5TbfBJUjf3D33pg6NXV
nHa1225Ep2ztkO5T91jtganptxtDpS9U0JNHJ0/tH7ebsrSIqqw0/2vwxaz2uddulQDeukIxG5oL
auFlp9iTW5C5kCsoFHr5FwBNNO83n0AQH7zzzfJCiDEWOdP8rbvWgy+lQOH5NPZhk5NzA1FOW8IX
IWrzV4iWpIh9A6vhFh/gFkgg+uv9zlxuk3oq3aiBrDj/prDfKgWmyFnwEu84+wwZ4Qh0O3o2QF12
85D4AL5VRWWdzMMa1cHxiZqza0usZegyep0pIhSPYLnkwr+0gbM+ts+OsaxJpRNbfVvbA6jHCtDv
BqtvDuo+R2gabC3O+qb81Mo+uXwqMdR7T4JB9tOvouc9IRMyvoowlqnUmno/I90YvDNH14JnE6uI
4o/W7PrgqcaR118ldNlxn26XrbYfr7bpCvQhWEasYXvbfroPy6CRYY/f7eBy5GVw9cIpxH4XRHgW
12TrvZ9giHxhWAmSlHBCW9F+YY+mLWBciynib7Qf4PnNELxDdMiqQ9q8LVb6miL0UAmTZIp0PRVG
R6bN+qKvidTIRiouabbeb8DjTrjt/XYHlNJZzbpFAr4zKVmSIrCDyu/T8iynaOj2qAsPQi6r/3tb
Ly1c3XvIjcz7z12NaiR14RCC+OV5L0N9ImmCPtbw/4ga8WOCcc8xFQAESzb6uYTAslNWhwnz+Pyu
8NTb9AXdJxPJu5uii45YVR9NffFv4geJMnuTXRtoaw0EFhyxJ5WNx2xCQUGgVm1W87mGo5gygzG+
psu+nppa/Y1EO+tuN7IC6vTLLsVsLxavjKl808XQx9iaMQ3dVnns7OlENbhCR9qXY6aTdoVuZQ12
W4EdE7hHk17GJKyhkcDniuHQ99tR8pluTgUGiiCC4yqakm38+Bf9Az2rMyCKT29Fg1elv42AJvqX
VQ3IMYanYAqocJr3tHaKCRocyZSQjRAEVnipf92ACNAOde4xAcACx9FPzGVQawtBXAuhJ6GIiO46
8pMPkjw2zAwYDotOyu/kqFE3a7Zp1K72K80rro8ARfiq7fiWJPL3g22a9o3+BlC4i7lUbKRIpbLy
e5a9Fy/txTU0GRafq+5ENA2nw8lwAeFpqZrD1Tx0SyNk65Xx3c6x+xSwgn7sYhptt37GJEfRcUl5
UKzQjH5EcvIBLMvUteCdblWlRUb1baaQzTaSXPHEmpwgQPlbaLYHpWEDlAv5TnnaQELRvrLbbXFN
UhCbAyQO5qnYXj6uG9ueDM6aqgB/nQ68rNFqPWHcOyg28cSZVfA2rNWHxG9jmu3q4oDQ3uUXZhEg
xfmRhn1wZ00nElGgoroNs24cgAfmezmQpp0qiZehT/EdBOy4s98KtNeA4E7dHJGARegiS67b0rlo
DhGq4scDQUwyoNAZhVG9YCF4opBggisZy412e2W6oGCyGCutaurKvoIxVshj8VVEFJnSBm5ZGKkg
vrA/dhDZAHZhU5hG5hXf25cG5EdRATlRF6eel1+jKikYRitAuAzTinYBUHK7rUKbd4eR+5t+T5r9
BwxXBiF9fEh0qzCIT3DJLPMsWJHFi2djztKirMy3PDXQb7q5vtE+9xz83peFE4ouNUmt1FyAwVOE
CEviCTk/zsashPPNcKI8cdAXSo4Gel1ZhQXKhEr29c4VcX7xqghcRGfw7sdnSXuPZq7sfPCgjLqE
JddY0zkHoQ8joznQNqAtqS3s85aKvfSBLoSjcjusWm0lKVKu7oxaA5T0adV2uWllC7EP1FWqd4I8
t7n76ZKeIbBI+bFz5dj5CYxZREODNb17m8AAQ0WLg/leOxG6Za9XO2En/nsZvfxlL2LcvVCYNHPZ
NmP21hIp7dx0uw00+ImIjo5vsXCApm5arO+2m2/V4Eq5ql11Sq0VLN5NGdZ2Qw4nhDqLf3mKBKrM
OrPWEljKW9a9E5t2yss4cLF0AciIp9tZlLWqi+YuDGA+w0cash1sS0WFDkaP2Iu3x2uaNI0gFJd9
Ljm0lqMjCJN9VaSn0FvxzXMmHYi1kizLq6uh7hDAgrAMapm+lx2Eih/TMpxoNoExnIWuqk4uZSoc
9tf7cvlJRDnae6JWarP3zfARPyCbW1HyEXYRBCKGhLEHmeSbiLbsqNgXVoXgLfOcdJCzAn7GWb9v
H8jMf3Ay1DE4pCmMiwcKwMDB1VRmnhCNmD6q0LWgw+nzlVc/oLry5pKbboOdZ+SMu6qZY5UDlpEj
iFEY4NzuMx219tVyf5kcX9yCeGXQcDjeSMFVAasKHp2tcsOmdKhUW3/yQY89t5JwJvukEHqFPNkn
HrAGCI4GJbNAtK7FURa1JlK2qLKYM2OBg0tnEMcKEwVPbrxkLlMoAcbHgwUWxWxBuPksl+tTmkS7
Tr8QF2o7uIuiyxq3WFx1eVtrbgNbGzKLdnR4lpFrdO5dvS2LedefxqsLDwom4LUjCLHlOTwoUdyj
3S8lSlBM5N4pYC+F9KT4lWIYo5DVaVLFvZcnVClN4U/Y+2Q673c/NdVHjk4BpmEZVWg2mxX1Q0Hl
dtJgXg15m+vYsQ9QDCtMrl0Q9dmPud+dKD/cVTuY0Tyre8AWZeT6hKsghVUIz6QnF7OvzAcxKONx
SAEnfQ31ofGIMJIu/3tIOaV0PHkw6e6B6OcdVd0QSdmlKRaRLlC3+eoxf1+Ek87h5rjRvefQ2+PW
9bZD+y4CG1vFI587TVmB1XmuhPj2lkRJyuJ+y72BBp8DDqVeFh59UttxbhF6B68hFjxg+Q4iXGs8
sKIkiu5XJDD2PYeWoWwkxue1PprQ0LK1hVYGP3ccbYTp8jtum6vvufDsz52ueHeetaxEn5LSZy/F
x3xW39DF2q0XSjfYRvSKokFXsqUW9f18GGaq4hCNUaMB4WsfXiZ164bJbFYlUjCcHewLNXxy8u3Z
6EhcMRJTtxwW+uQq2Kmd6xN6xMwhYZqwoO3VGgrIAq+RsXkCJwiAyk+qQbAJgfenxx/eCXiGxarM
wG25Ab2UMMmkGvSeWI6VJTAl07xyONXBI7GYQ6atoAbIWD+wOZXJ3AV3+C/celMB4DsJrt/fT8Dw
bCiEoq1nff66zCm/GpeBKIrE8TpdbNkHjJdQPnod8dXDTGIE8b/m3qUf6A/JoXwot4rFGAVRi8OB
GU52vOo+v9uttX/XCNA5wV1u8+Zu2+iex2Sx7WdDYPwvSN5GlTgkBSrX0HXg7g+KyrcqlYS6Xtcp
Nzczs39cHHKLDD59hDpNOji0lAhCKxNccqGF1oBFGBxRkVcZbv0VAf+3ypOUlS3ZNmUMHaTMXzqC
LPLw9Gem0tEIXntdDGeMM7HEd5S4h6uW4T0ZpzO390eHpzBawZQHIIf1nki0DFS24z0ll7MnVmSu
XdDn9ECO8M5Rzj5LfY5jZ+6hRnUJb/CWdEi0T0CKOiBfyvKjwkXq5iHFqiT4y7Fo2a52MbTQ1Ru0
ybV7hWEP1OO/+CiANbtHYWg/lfE5hUVbhs2ZQMBDrOJF7yTLYVAGp15hOIFlbjn+FH98nZZtM8wk
kjkbu746kEAPhoquxA+qfBrkd9QaPbcCWMQIqKngViFtu8csw4cWY7Ay5vgeq6a27xmbIU5VCnbT
hSqBKF/tjnNMLZktGzOhlpq1oFKfVE8d/9E1TZhRuYSlI1NBipAKdZxurwKuL6PUPS1oSSGZHTmF
JM0HYN4OmrR3ARpFchf6h/XqOKuM3+qx3CJJxinJrcyzfpTaMOotCXLhTyfn50EePGYORbvZ8/21
tr5JIb2TBE6pw1R4tzVejTr+Fms6UpbHDFtbUIxRpjnZzuYXu63KqHLCx6KZ+osPpWI6Z+iC3ziC
9ttrQH337yVhT/eT5fCDiKzeuOI9J0C+x8wLcSmZGokIksbdQMupeTgFlb9eFibKno6FPbJZSoJG
iec2Cr4LRFqVkMw/Lk04y1QfAj0Zb4wgKOGkSwXLiUU4YaUhFKfK1sfkoDUZI+Ua3CxAtDy1wJBN
EMT+JdAlHXDfHC2zNzixSH5rAVGM8a9Ex4U09UCr7labpMTNNFZ3WAJpYq8AmAK08WVe4dF/3ORM
tGdLo9CfUD8iOPOQ3jG0MVjL1rbV+MzSuU95yF81yj1Gm0UF3w+qgR3hBdUqhCOXuHg+qJoVp9CA
WKhukPPAjpBmgAnIZHHwwRT6YHDawYLMaJoUpDYTHNh/+XVWw6BsGq/h45ZC2cWDh5aH0Y/52B9I
LyEx7vP9ZNtB9x0j1aqlFP1mqu69nTKg9Xq31QGlc3Q1K6yZfr1gBJt8vfGXSNwG0iGeVeAPBJhw
lO6aUC3JP20Jc+RTgZuAl6SaF2udZ6ozQhD+b1QMUh0Iy0nmbek3muMekiHBHFndF0MBqbgzNTgr
6Wxsk1BsfTDmw65iEd/QJmJ8RLtbKlGnzKN93ZvxXjJwHhga/Xa1NFQqZUD6GbIh8/bAFqqTFXef
3Xine1I8bNUk8gXxKS53gjAqrwv8ZQIjXSXb1LTm0B/gFqOSSbTbs/4dGV+5OFJVTseWKrT9G53M
I69q2RE0xJ76p3oHyvY0Kdi+kUJTCXYHFg9ObPuYQ/UAP/kdZsUL0Z8sgMVny5pBQv5Y+1UsX5LL
lLthmPSHw4lzfOelX4wQHsIr/xiizAi+rv3o5NuYpm3dAwB38qb+Gaxp74JBmaTR4Me7YxfeMcTb
mq7M1k2GXiXq8LvdW/XWLb1hIPfatQo4m7bT7er2f8BLClH9ims/UtCJ/2CmXehRF7ORvI/pTrRK
Ord+Nb9JeG5pSmDVwViFiu5ARnAu9V9MI9g5c7ZjPJgiCrLDNmQWGknbxuVX44XacjHxC6YOosFK
sJR/iF3M0yfYRERUXCBLP3cioQ9DWd1S/kX0wF5o5OeiMdJ962nmFmu31aVoqj/kHSS4WZyuIm+F
ef6snN0vItU9NkeWExcsFvqfQnMuwcsxQ9A9IT34egenEDgHoDfx7ZNo7ggAShjuwCWggsQz56hI
nQUo1fUQ0ec9kvjKFdRvXjK8YbnxBFr+6TLkXRrKqVyInQyi3SmZvkX04JAsE4oF/DhzX4loinvj
nUoli3YWzhWYnWaiUdSJz5fGzNc3+Vwky8kiZ5IXYP5vohGo8KPhAzeEV25aEHyelb4QGyDAB33i
bf4VAEI1ArwdCd43I0jfJ/0qo49ClSgJNOAfkEFc09iFN/YpyRNOmWzsH1/oGx75NLQfuVYOoA8g
RIzjkiUfyrvvZMv8hEYq5wAPMVFXtdmgtQ7Nqml2R/M01GtbbBECfezbwAJ63evfxNhVmv4N/YTG
NQPPoyrRKo/Gehq7OwQgxF7pgsVAVNu1GZbUHHixq4ksjCMVIDU5Y87nHSr5iwm/atyvucRumORF
fIqKvAj5aO2ST6aWQEssLnsmd5oHfW8bVv0aUnR7hVdjfi5WxjW6e7ul/WNszMIYXLIyuG4ysbHx
rR0JL8idKRco1NxYKQAwmhsbfnlfqkFMJGwLnzn20W5tA/qkaB/XWRgev56pB2k6VDi6waFphJmN
R2NA9Onpt7xnK/hD9jQz3TX7BbwN9PsHh1/qL3urMzV00NF63hCgXB2Vw5ffjhP3GslWnYx76ISm
VHUEIEIMH2vcOMjf7S+KudmX168Lk4TutuwZHAuiqtDqU2FhC97AARdAek+/wEAyXwjFLAhGXSpj
hZ7WJNAh/fFkDDlcCo/1ETPjAGhO0OWxw8Bpd0GcAWPzPgs3GFn/e0svHnv9F+hunRWRm0LGSdbT
b7hR/d00EiBRNHUpZ2WHUwG2nhEVGevQaLmKrIJ6kNEsJpZtA3WtYh5xj8fHrcDtfc2lZv5m53iy
8Z1HL624w9z80ayPeRN/AmnLg4HTiTlTJ2cf2nC6BkAyB5O7c66uuCNK+6EBSMkyZv72u3zUiBC2
ZuLgomv1xEz8TWcx9poPPdbww7KLlR3mUfxMLI/7fWt8Vmo5buKpQZFZyrK0d12/T6JOHQVkzeFL
RspKQEoXrGBoWiVB6YwhUVhnKqFtuWroq/YSIs7n6TjCGUALrR0W+yZSWF1g/G6BTNA5/GOauK4I
k7wtSeem6K/oho+TrFFzUD1ongj4+43UFSV0oFcJE1arL9X1yDMHCU7Cj49ywFyDhGfjgRIwuBh0
vGx8EyF2aIdaOqmv+zTHFShVDnWXZndrgzFljGZ1lgFlYGC9ZcWus+YMOG0nz3pQ7or+0tV9NY1g
ABAD0383uXVt6DkA35omNhHgdDptSavgCP19E/C8WRyySFCBHNRzLC6Gzu7ni2iMW5abbC1sxv3t
jMOcxWdQOzTND8m18z0mk2r1YuJoAhw0h0rYre5gXFGnlemo8E33yxRcrRT93ts/Ul2VW7z0qQ86
ZeivJylSnaFuFQK0G3awSPBPLe8RBJgOKgRqU/smX7t4PknWd2gh/JNiADwkw4/hQBj55S+ltsjn
3Dwr+lmBhKCXgbswoImQGAJ5+RjKoOSpbGNGkhwfEAnKm2Pak7SAISJdkoB2J/ou88hDHjvpV74h
hLjBAV/sY2XvlZaomn6aQPgkzga4JAm/fHndSIww5pyju4hu42GAlcI5b0J1FWZs+tzxcdCuWCQL
Sq21obMAjTGFXZ+AwAhuR3Q0u3UVTpeGwBteMfiB6GuI0H00/lu+ENxwhEgQyVACqYugwGVgZ5Qv
jn4yIitncwvScUqiGoeYBqAZEMnu8gs9T29GTc1YmbQs2wELSpxpfwplnluDN4xfRJVDiNPg6xng
4ia5xN6ylOECrfvqtIN9N1WebN1DkEn8AQFgqyWCW2P22q8KKC2M1PHvKubM7Hj5S8XsJWd+DqIN
EBiAYT0RomOeJ9y2kDA0NOObY5OGCEyKlwqjrDXOg9LCRuDR65eViOPFXWIEsHxdc5yYdDpH64Yi
MQZ0e/FOgmwL3AG1S2JlRvzT8SFBg56mcCRBWNA06X9JERI0LiVJwbkT2UxXYnknzoi6PlQ/tevd
z4LRhUJMLw0DOx+9pmU1LopXIwMh3bKFbnOe8UaRh64F4bvWXTUW0Ytgqamx6oyFceBacEDIegXA
Ft+xcWevoGoDlDbOkiS9aA4mAFbMkxvauOrjpCXZnjQEdEii5e6PzZKo/chacFSnkNfwW4YLNELV
g+X8bBsCmMq0HhRIWHeqbr5++W8Ngk3H/a9bFXXFdTObChkFV9B31dlb1xGm+3WZWC5pAADX0ipn
Y4/JJ4J/CucZC3vz/ZshR93nK2XK8mmLltYMBTWf0kJIREEcf2YZqReaxKxf3VqSAE0POVwij0n5
bV/BTwCXrkAeYWiE/UmXh/WfYMk8Z8sGAw8AM99ptkC+zgS0Gks9Wr/c8iTj5WrorPl3NEHK9W+v
bwHdyXNQow1M4//4qxXxH6ng6i+/wTuNNqvZGWTg/o5zqwh3G+qV1nXH7RVb7OD3YHXIu94WhETf
SD+WHTzQAkA5zE8CEQkE6ZqnipXlZzRCy78p+A0/b4YjoVJQ+RREo407ANVcaOZp0CnfDfMS55U6
SiTamyMLqmV6PiLfCguZge1YsoxfdD732WyeaVaTNu9nhkYu50PG5GJMoKbyFLZsQ76NrqgVERmJ
ZX/BRHvecSc5+xAQuCmb1Vm/S8q0Hz/WToNlHtvCS7X7cnxYOR6KlogWQwklEGutfkCKcA0CWTQd
KvZxjpYhMjiib5FmpZRqGvREbitgZmizi5pcis42Z15ZXfCVqk+ZijXL5zt3MeNXIEv78M6BMDbr
jPHL7h5wctLXot5xhDHxLWqVRljvRURjCZaifS6WF3xJJONrCHcDF0k3Yv2ptlUPwxVwGcG5lEVK
hSuN1MpLeMYsl5Ea7/JJHKlimUZ1ruCu0SCp9gCrAi52VxpZjy6HkJsyhpsbLSFAFPFZs2RmAE/+
7ZRjKF07CJZCA9ja73s6h/ci63+Pxiy/Hj2xXYB80DpFeOyr7kSGOMpY1w+gzoLOhRlZQjoXuuLs
C5cEU5HAj7TOWI5i+5+YzIkoNxFNzZRp7NB8hdekD4RQ35AMpFXffDtX7l1wyL5ewDIgrHP45uzg
7YqEeD/D+KEtABu2OUdfm/eKkGwP/cg1Ej/v3gWqzLdGA69a73IfYp+gMX+b22YVMP9lWTTGTe4X
WYuKUtce0j4orSpu7YAIKv8XOCBCAMmSfGwqL5srvsgG6kKOlz9VMbac+erd7Kz3Iz3tIOFJ7fTS
IJn2poidFYF1x6O/6qJUwITtBFWFTGo38qkIjZOUIkCyG92HgfAajotYDGOfdAiNn/fO3AeN1P2h
Q/C36PoLmRrW6TfZNLnWBoFSXkbl3aYgsZQz6NGqgzP5oNLBH+c+yzNci3D9fI7I5i8ogLvVd12Y
7dKAVALfcKxu1SjKeCdE26u3SlCqPzI3wSr1SPZ2QRu1ino5O04IFv/0aiifLDu4GxMhX/ITYjyH
96byY5lH00vR18DWM7M9/kJ/2NyxjmlaVYvacMGyTmkq7InRiFPmB0zc2M6QYS6A+6HEgRtG1Y9O
iPIvq3Q8A1iwOV5UZDJi4Opopn/pgNrxLLTYJ+4EEmlNLwjv8IEV3VT1aBfnSKHyXpXs6zcAupsV
9BCjbqFxV/xFb8L2pwhMfyZPLUuGbDTMXBDpyH5WJosVPEOkEEGPFI+PijaD659bXy3O2fRUqv6P
LpGoiq71cX0ZZWeyMUAOKH4CNilCTkGViDbR7QwqN8TMFWux4v5joAQ2RMjvMsRYaaK9mG1z36CD
Eb73Ti9otsWPBV7c3QRYzQwrp+mPUSbPhZOJHgudWp1TXruXfmFOhUZz1xrUrtGROa7txJMaIZjG
NIRDd0CvH0PQaiii2EOAS8Ct6E8oBLHi0gpOum5fuuoyRi8jx+QTI5VxJKcX8Ryw5yh/UtdFLK5b
VGGewYZf0/IB06lxbggKTlQj9Pc45NjYGbqZAg7x9TY5TZai8kwNW50dHqF1SQGuwIaLpWq+pq9R
3f6jBjL/TLY0XER7vraNK3tZirzrGFtE3g7DAslX9+oFJrjeDJva1+/xr/jSiVpA33hVuEVz+kcd
lU0Mp1vCoTC9byJZOh1sM5icJsQXq6JxS6qIcha+wzcLdrclmKh3Q0Sy0SDOws4dnyp45UM7Wb9T
6eGU0Vm1BZAJfJkpDlLcrfgfcyBGjWocIbeEgrzV7GJ11Mm021JQqnXHpOtHbpH17A1IjSPOFL3/
hv1LqdFhEQFAOegbXnaE1UG0EjSQPy7QQoxo4EpZg8ygO+oPYbmK/h2JV7KlgXeVvuOSR75ddmT+
d8Gb1NbGuQSltDgxonasJavaG1453XqVgGVAPQhRLn94wFjVi//hJxsIpRmiYpAyoy8SUx0tApA+
2amd5Mhkvj13JJ8SO/f8Xtde07829UkRYdDCu5YofcLkG727c4z5houAnAivaJu5JrrjZFLri2UB
swuohYYjgKOe8xYWpBuJxYfMGLiVFwyCEydHTvRG/+rlS6b5aPFYwgCFaDyJAzuypFIfXC/tGWve
JCE4mVbpgQOhpuZycoSnBbuA/mOK5GPUCX3xxrwa7CXNqzNEGCrXuHW9OmsiyaE+TOD4EuSFInPw
al1qXtKuV0YSNVoSLruowod5sxezY05pFfFKCCAF2oL9ccz838e8oWmNvALhGFzSspIUT/jwma6r
VK8Ds8Lg3mOx4mlPpoRRzmBciub/9tI9iVe3A8HDUctaClWPDyknPyen6wM19LdKgChPGDO1A2G5
CDrgH8inS9KsZ3Qymby2Vye4W6pP2shvwybjD1M4k7xRCPD3M0F9IcUoJ8kqafXylml/8EgghGWZ
0+oDxAc18nkisD2Gy6zN3OuF0Na0oB786+sxN3npjKNtnHBcYAjK9Kj4SiySaG7t68ixZ9OjU04T
TepWa6f51w2mqmqW+e3P26G9eCZojH4//5fWmMWLXGMz7+zuMB4xDaNJgpksjH/obvW0UVouTGup
byU4sv4XeACo95vc+EDqfbXXxFRObLcLUFXwQ3LDvGOdpgdSXRDb55BI+knps8QaygEt9a4YxzpC
btReLu8Z3TAG8c5PnNBhPGLsAtnWaNWsPl2rju8vaTku9N28hDAVtIm6EH8Y15t1hwAuYTHo1NAK
Kj6rDeOOy3dO6kBAc1xKY5k6bz/qeQaYkPVyREsWFi1DcPcNyqbr7Mw/GHAxF7Nd+fbsQkX6Opfd
Xid/uTXIxRIQRS/JajtswALzjmcHOeCZAqlYT24ugIHDDrEz3NfhmBmIFJ7fACAo5+ULFNlE0LCM
+TB2LCPNY7pW5zn+kkR+RfcT1StolhcL9EUkROhkjNMgVgvgtREj9tDZD1T+VVvZwbR7zXv8DGpA
vwZa5CLknlta9WX5JyrEKYDd+RjyTBES6ykXEMoS9rfllZ+iiuA57N7wCo9XEp7PetLGQsijLM2o
Bi7NW2KCU8z6lwcMo1DcKhbGADIRx3O6AOZITqVAZKdvVnxJkAOfLGMQElw+e8+Q6Ppeh2rD4Dmf
oaanWVbWXNLKWqLVfRYCu+tUcnf8/8B5up4mC2blRc5RoUhK+6eMWmQhGSQIjyjXr84nCO6/km71
+A8IzM60C/Rn0KoTgo1r5++UEPIFn6gyA5IdGx4qJfcNs5RpGhDDAaFYFyL5FbGl4XdcdIu9vsSm
Qz/y05QHswH9nm5MDvsk5qxewfuNrOXm0OA5hfo0K6cywutPDn/T/vFS5FST636YrtxpvN2d6JSP
iRAj2MmqAhDAGfIrOnH9rqQHTeaEy5XfOTl4LVb3dUJxee+/WOO7QoC99/Noh1g9t6Z69Bru4Ob/
nniJqBjCYnvukNcMHm0qutQsAl/x/u1y+LfwGJD7U/l8PN27DPJSwjp4FeAboB2RA1IWZTq68aPW
ZGv58GQZ3Ia9flGEbEInsYy95NA/fuvsGpJOarEoulp09+Al3yIJlLKmnbwFPJkGmhWRooYGAUrG
vBfe+7wKRP2uFd5L67nyu7sl8/gK3zcD9ZIecG5neymcHtd0oFVN5XHtujjFT/ZVxwFsYH3OsgOb
/BihGX+IttJLVHlwrAbWjq6YVbq/F8ziu3gz7A8j7POZAKfXSEJ4cXYv312vuPi9c53ZWllld/LR
aTCK+pdRC2je4h9T8TIqt1GhJqOjnlCx4+LaiB9EskzZarF1MHzKAxTywm0s0BoWRtOKEDbGY1BQ
uOZpMGu7FMYHmfDbPNrmkxdRgtUNOXUx1wNs4lnvrCOzD5+46uGGmF2v16uEsWETM+gnZiNJXK6p
sCtQSU4GtVi/Gh8eHbBWxDgNK07NEToNJgniBRaXOvoOy1HqbG9gdFEek11yxlvu6yJQ18xNxJcj
UqjPZvf8n6td4mwtEJXpDycnju4zVCPTz9mHZm+e1cHAhVY3nmI9wJS7M2euOUc/lyHpiYo78OwS
/Y99xfA7tEtvtwqImfsutjgx2VYN/vTQt/1Lkb1Hc/fvPIQmOl+ypPbtp6Ua69kJfd77vIRx09Fy
dj+B4VpA44Rv+qbDWkrlUtHCc3Yvd8AOcMd/1hGbJKCBa9XakD72QsLd7+TdSPZjyX573W/4twqd
fjBIYqdC6vhvtcpZzlFBvwFnERgphTs2ooPFC4qWa68Oc+iuKBfISSprwUZmkN+2SL+KBhi9baI4
LMlQOZPeybd5w1laVJTSirXdn/3o1D2gIjUZjkQxEHHJiIZNRoZ4uu+/gs3sWjqk29aeR4CkygD2
rDBtvWuc+pafNnKMx+ILhi1hbRx7apuofOg4wE9azJaroKFcqyut4M2hJREiJPwDdXxP7a0Qd9Rs
hXDQi3tRrhC/vpVUkRjQ602g77qM8leQ+VRZF7OHH7v/Lyx8eMtnvIebovl/IGEchBCZPt2nal3T
kPFG3KAAVXThEabaHMCCkniWYSGoeH6cB4hRfBxHpqxz/YFtQRmSFKyy+UQ7r9E9fWKGgam68Tlb
8kNqDEeyR+edaKhrZMvLszDzf0yjZKFn+FjNkev27Q+kGvTW1dWXxCD23Yvyp+dhIi8aqRX2glv2
dNuBrBH9MR2atlQohAMiurIIU14EWjL87TTy0eB/OUOMZJVSzjeI4K0+i4iDVxJ4QgZ4VF5g2LIu
iUmYelRfK1LWmTcnzxeosWmseJSRrHR3hbpwUSIr3NcjWG+hMS8OXdr4GnBK8xpdrBFE1u86mBin
27NkK8edEd/ibV3jVQtC3437q9b3BPsE/MqijTnrsYfvdQPxyTmdWsGHtwiS3hc0DtYfaIk32/O1
4flfnFq7615YSuZZpOLqxVw0p7fo286OHKoB7lncegOzdk1Cd8CwPuctsUNzzHFxRCPFquzsoCGj
Jz9bMRWNb6Xl6EgnVgvExSCacRPRBNGOW42yKzZUNf1a85sf0f3ZfRVy7+IiTgFahrKUMdeA7D9a
FeC3LH7x07OUvXJ14X4wV+1QagC2tglifc9JAjL2UQVF+9V3XIjrUlSe+6cedWHIcGFy9p/NQPo+
jG4LD5FSrm/Re+zIpC2nin+CppwbrVxnpr/J9dBZn1LfaUsUogBwjyhJyY5sOM13LIC1qcY3V1Sf
GrzI+tHXE4/eKCGXs2Lt7O2iEMHMMGsa7xGH5nWJEKp8FteAA3FgxvgNj9QaErWCWV/wbjAjLgjF
Za9ESc6rZ1IGdD4sC0gVksPAnJ+0Nusld5SKipnTVVRO0YCNtKgLwAACGKs6EAHhfGllQU9IdlR8
gFuE1bKSUxCBmC/HjVSN2UFonISw8sop8fwYXSUiZlH6rN9osk0D1+1Jjx/s7bwucDqYNJeQzHk3
9VUlDGSc/T9vhw6BnivSZDyc1nEXAgUlBewF/VaLGg1PsYKhCuzRJPuFkGH1vB23sR7CuYm/PjKX
SymZcj7TLqJB+QOEs/m6YK2jejEuDvr1iO3j9NbAoonvtjHpJT1xfZf0mzbVd/wECJVzA5crBdse
kpG4gzevF9AjBtS0SFy99xLQmMLGwOBNAYvwsdVHDDRWG23shoqzN06hGP8fWJFphhTzttull1bB
m5By9e+nafJxVZAFk2+LW+eRChPfkaydtHu2QO/Sr+QUNPC7TmvHEW+x+aGC1sWQ4GU04Fko30Rp
+dknevWSdqevT8vKJEAeCe9CCER9EsBFX/mFkvfXeYlTNruW9KAHJVMfFSCjGtunm2AB4nofiC2p
nWaxjfgX9PZ+qzYPE2dNvzwK34SjO+XoFkX3ZGaUCDZVsdHs9uIbkQHfKEyDZCJ4HSRgNgM6nn1/
KbiP3b215rRiNFzacj0P79OJf9BypHdcrXjOv69J41wYcH6+EPSM6PX8zYs7p/HRcdsVBgKRdJnE
uQKO4x+0IURJjajkpydEA++nmmXS1tP46YYa1+P3M8hl4LOOSsRLBGBPqEkEo+gaa75CYyJSQhGU
DdA41SlOdjsOG25PXXm/j1pazaj1DP3j/z8jRMd4oI2L23B+8KSwPR2UYVf1mutd/JrrusOJElcc
IMHLsXEbYon8xSp4qKwnONQer/Qtr+e0HsyHkU0EZZM6EsbQWiWgO+t4+bJPE+S0DiNojwxd0jc4
l0nJRQuUopk3JZ1S15HfS3laT4q9j4+KHHW1lQqz50bJ9QOjFHdb+kucnZC9+BICaTfvNMIPG6n8
P3jk4y6/3ajR0N+K+OI9lYjdMzk/n2IhXunURq/Vuqk6g7qqBOpxDVyT93ccgXB0zh0A1Rzm0vQ4
zyodkRof7rwfUgAme7F9ySb7UDBjCtWFRGgpsQ4PzQVob4b9RZUxrqdy58oAVfXfhvT9mv3xx3vd
j+R3kexgwqz2cdLgAXP+VPYEVrInZ3QP55BXM7EMLslQoOm2clJh0eF0ysvOy1BpS7JQ82SSun94
smwMPTizwOYocG2IX3+qspCwL1jbPznqeLWt+b6PCpMIKLc9dShV25m5VbJ16PfFiORFUO9mTgj7
jjHidtLJqdXV3jwXWkDp6OUGsrLUxNJFJzUfLIqIHCOMsbs9WqXGjOMl20q6Lo5NsS9zfd9gQDkM
faQBty+GyvcxAu45CnOjZY2DqD4N6k7Uv8Nv5HGJRpSXwu+Mx+qktX0n/hJubMoLGpMs8qrMbwSI
GK6NoF/E6r/19A97BgX9UN16Uw99phJSyTEmKX5NbDyVcSHSGd65IhNaYojvjkV4s8wkd9Xpb8uU
YFgQOkgUUJrqrDnC9P4yhAudfJf9IV7GSH4ItLANj6qv4Ck89Q1hw0bSM9zIfyXQvzlcFcyhgmJz
VHR42eiQSy8wNE8CLwcskPPlf8B3d+Owkw+2c6ksHenjQpbx1Lj53QhzhrDwLMsxzWbRE1kqaVGY
zjUgKNVksWIgESeYs7ld+EYosxZzst7r83hH685/37/rGlIliFFFOtt8zrjItbsZLawXe94jwmQz
dOEvF8Ev4+W5HIUUFl3F50B2S+1bXUiHMWZ9tgczcAJJFGLX6t549sAqom5Yto6eS/j50uqqq53C
M9IUsiHSMqXPTmGy1tzsq91gABAzb71uCMNMC4C4iTxYYj1ioP6xWcP9hNHBlwCrCnSRTKaSoeDs
H0blpth4umPUuGDFErUdqAtz6LkvHnClE4kv6yAarH5k4C3W1H4h0tTlkKgly6G6snBY80n7TLLa
GTLlG7xIcEkGdtrnf9RWxTnnPWb/bNtdl6q4BIOoiudNUadqdXIO5K9GNc0bpmeu52GI+SZsxS7y
PfzS9Vw+wLNN7yem7FE7NINv4Hi2fuzu4ZHVZDq4ZH+SwL8vHXTF8YCW4CXddlQxFYPnHs9qzLYD
LLxcppWD0Rhf0t4scTlnH5nOsHybI65scluKwg4unJfPZyf0Zy5Tdo1vnbStoOB6ory1G9Bo3fXo
H5XLVv4J5vM+mIzBX6gsBY0YHYdymE272qnQEwXP67TVAn7jIJdU7kG1Cc8AvaNT1bN5V2S0npps
qoF4oBAmkrIPbUwRoXbfWSOCbIfX31q38SDpg9yIkIUwfPL16ECcrb1J7d1rnp2cl2pONBNiklb2
6nAgEMbiu2HvloqSDISf3b0J3VDGCBvxSvrRWUJSG1oBDCavQWvOND+FonO1ShZjmfn2uP39EFyb
jW7lQ5Rr4vxrkc+h9miHAeNSm04C6X7N2LE6evBdBnUXpYoIZTUFs7oM6zyFBxHUTOPLf8SSw32e
f96mtSeNzmX2h5UbbWUqJ3OkVKixzJWlOMRcyLnxFgbj8LuzkQOXe/GtJh/BiQDHyADpbTsSkU1c
Ozxa4w62IOlkN4kF1+knjhm3Hlcz2MWTcyRm7q0XGQMqq0rue2miWMwHLO11Oi4DQa1rLOJ17FsX
3oyfFSbfjbndm2xPu6htmVv8JxtuD9ko04Hi8Nx7tJjiIKG5uiGxF5OCz1QRRfW52VzQectCNb4I
H2SbyYBg/FK4rox3TIKcCpYWh0VOCsNwU1nRBW0r5onUhUyLIbkGVv3NhRuXxTHKXtRBqXQZAU0U
mn94yZpLbG22d9b7EPR564tsS0iTciol7c5qu0VXz8Z6qflPuk6KhvdpNwHkSUNwmNKMxUoqPhbv
ae0qfdplc7zlQwQRWbftGGTrfReiqIMNB0JwOWTwaPId3mNXi1B5E1nShSE4ZrGU2MgxZgkBEdoO
64aGdMjRaEI14g8vu9JWConGD+ERSdDKqhyq26VGYF+BsK7Dw4ekxNS2zxbcczAtL1ncsSb2GlTh
NLFKsBYRQ97IAdWgiVT7EAAuVLLpQI8GztKxPL8EBWp9y0yO6VSlfxFyB9RfaLUTPy3QbRa9rPRY
N6BiOF+xlv7lgoLmLIJf3LSIwLNNjMsLBv7w3n1QMZ1MC/Km/gUbUTNX9ViwL2ExY1g+YoxaGoMv
XtA933NlC5Ko/3yIYn8S6vwxgdFNqUPcVsFxBcxx33V43IeWBwFcXlwr7JXFrkVyTBaBVNCowcp4
Fspe6jW2ca+noYoYx9Rf32wdogL6aFDtb3NpYKKgV8ewrPAOhV3tUNS1lK0IzAUynAZ7YJ3mzttP
crWFi45/B9k/6J7yGNs3VVhmjPr3BZ/d6edg4LvCmVxS8wNbnpUOTHUBDv6AODGIypbbaZBjVjLm
SjKF5H/aYK25UFnSQWuvDv7RthI0kz3aw6KR89A03GN/z1bxV0OrSmqdGzwOFmZav/U0c9INEkNy
E9rXHekZsoE1W481YGgWUW1wPfxtvYjEn7Y6lWY8/XrZ1JVU6fAkNDwKN3prMvI91ihzsMR5v/iY
PyMIZ/e1hlR+zQUYd7CYhe7oQeVBi06l8tVTwlBnjXuzMYyJGjDuMVOi33Zd7EgjxSQxCrjQG3LP
UOdiPllOrhTPqQ7gLtzmXPdiG5xyAingO4LwmaJ9EMYinXRRAjiAfDFhr4V3cUX39PUn09y526aL
RoEVFVeZNYbAeoI4njkqEKzgbjHCD1ua/vGXD5ZfFu9cGtajnpdVg4Pbp2wSKTCTZQFd4odyOIQs
7lKtQnuXh4XhHb1qKCj1KmjmHtjEZ57BPFw/LgoD+tH0+8mMCJF+PTdRAe7pyQl/ZeRaI6psxPxA
gUO21CH0I3yEi96SNbAhrIDamC66V3HH4Usd+xGru93Q45jJLTgo2VsGfxIKoh39RC3oHE4hUD+2
meehuqz5OjH4a7vT/lyJ30OcUqevd4haFKRmbEZ0Y7UoFFC9uC94cPHMRxSv9uYoxSr6A9m4jnHX
NbCm1Tn00mulbaU+s2AeHj7cn40zhozo5fxX+2XabIfJIMWDIj7U3L3m9fI2S/AurRpOg8P2bnJ2
ZS4R6uEQ3CR3LA3o5DcumdSt+XRTQ4O4H8HFtx7rQkjVOq5TmIPOCMQqssH4V5XySRTENpnw0NO8
+swxXqaZeaiCjTMkUFs2Ip5MYMG5vC5xeU0kqbkDUc29aABmAYaJTsRhgqQ0U7rlpPPqkjzwwFn3
4GstfxP3rmWCQbCFpCp05QhSE0YySXgusld3b6g1pLUaWZgXKv4FRjwDb2kIEmfyiBI1v9Fv/qBh
5W+WgE5Zyw6WrTLVC+G9CK0nQLjo1ZPZTMHkfdtth+K02unD83cY7IvDq3FcaTiw/QNknAo43YXO
2766LPT0Rxz/qC/5jig5+FVkzV4827guP1jRC9Ht/WfIIT1q0rh/xsmS+Dtxm0UR4+XPNY0MsHSP
FVHcvFle55V9Ddbil9Hd2bcIyU3aRL9hN0iPHQnHzH4NeTq9LTdnpdJ/iGjove3+a0rOEgcwdObl
Ll3Z9vHiNnhk7sB9YkixbLpiD1VdUwy9yGuMC+1SczoFKjNZ+AVdYnyZiXCjTFtDN8rke35rC4Zi
kAcLNdNnzhNevXddbbGrq1pmWZtLM/xFxTsdz9EIhrXIBrLaA6e1qLyquqFTfE6yp4j65alv6EFM
phRF6LhfVQPPiQKmkCBiYqxWQm/G8x+nrzcvnL9+EBoX1HSFEwizX0lD7Sx2qQtXW9D6aRVJUwZQ
crCARX2aLTlpL/S4OS4refCpPX8UixDy+xvlyIDll5S+LBR6lh67pD9b/2KEe22oXeHZJoiLSdLq
/5Bx5UVxQCRccBJ1+A90VZoKJKusvy5jM7Hc4sQRQA6Wj45SzKTXY367J24Zg/yQfGq4UZo9gSsm
BrDTyhFHl54z20gJgUIRKYVAZj/BCC/4bGDStlyKVDvmCjcNwK95u00M11sPvS8RyXFQzDXHXzUd
6YPT+NxfGS0CuOnWaPDPsKo5CWFdnE+4vUNs5FC8FGYzvwHzQWKZ63v5r9zcOt4JmYJSbUmcpDUp
w1iZ2Qr9GqlUCTQF8a9roj+Tj35Ucd959A0sVPT/FQVl+q8zyELbB8zQXe6Vu7WB4oXE0Xg3JCpS
hl8n8iteABLU7mBdujEAOXQ+Bd34G3+H/dgrUCuXUl3wDa9fDslJoe30wbPpIu8IHG5jkRZaTETq
0BAMegSz+wbFUtmv+aWO9ZCSp26RExi/zWTR+6s0AbHcrLs4QHMhdhuEqHT2hORbsQiCzzd9UMBU
gSIXK0wPR/XoIIfJhJb0LBAJV7gvTfSGY7KmlQwkoOkJ9A3nJogWjGf8ytFKqlxuRSkCtuWf4BDV
EfrqbId0uQ+8zaoddCa54bmbqWkqJ2fb8HD8WJ7BNb3Z0YDiKuO2K+ci5uy+wx18uZ2lJy+8/Xli
GP7ucmJBvwWB1Q7jLxaCgHpaJeOZgWL/oO2v9clUcvc3f8iAViMXjNpTWb5bhghUPMOgzN3LsQJ5
2IM+ZYZvbwKha74BPM2VRxaE5yBzV5cBrVuNENuT7x3UUr/qIcLF7SRDM32H/GFs4I7B0innf8VV
klzgAkAaRzbVyPt5nwz9mYd9PPOU13/OlJh8J3LJyCKkIg3fUS5jjzhvcbujrO0qf8IMJXnwkKwQ
98agILQvuiYHvFtx3r79jle6faM7C/igFjEYLpFrWbaMGTQgJKbODqjN7MlT0/a5DP+PlMZ2vNcy
NRkRl7d4+RoAF+RbGxttgNPJkWotsrdidAkMbfDYSgvmhiBoL9ckQoMHQKM/6c/6CA0H0yHiW4EE
95qVhKS4hw1NjGx/hIA2wGG3YsFE1PfBaJ6q5DBOsq1Od2P24hl/zQoxVfo4Vi/FBcAxb3MpDZJE
6MYvp1ZryfVVDly3wfODT2LV2I087bvqG1v+FKUtgIwUufBX8UOBr8g7KOdMgXpWQ8RnepbOvEXU
Z4sFR2AkoaonoXTvMDvFBfxZupJJnzLbXuV2V79GYunk3HEretJNjqjUv5wEDujYk7D42lRc9Cw6
h8NY4G0aGi+dVv8Y6KEkjZWZv27AVW9DnAdQ+DFwGr77ylC4Mcu3KVJs+jbPoUSU+JkUfAouYnjd
SztqXIfP0Zvkd89G4WFJGSrtui+wtxvLHprUny+4LUOiLHCd8HvQ7qgurmLz9ctC3R85VWF8PWYp
H54WTApP5PAXWJR4iD8SxSeEdGEFgRCcml6dFkNPxxsUj4n8E9NRpboU4pYXYkU4Z4vMwcVSbseh
NlzqF6FCzA8Ibw8Os1G7HyLZig2A62UQZdv0usbeXoWbB7ppkJ7rf5JxjNkkzAx9DXf8R/hJkncD
DEfyfv077qVD/P0sWRmQXiS5h6FUkaNOPPnbA1Qhki5c5pbCr7hSCjaaf1KR80HKk6R9Wa6SjUSx
RlE1rfrxQub9VgSUZO04AA/aFWGgPdEW99GRrGRvgvYQY8C0AZpXyNWJyxE6hn0xp9rz42TeUbRC
LRF0MYdO4DDvXyDOV+oAF0f1iFZJOOd6w1dvJn9ffYiY4heS/+Tb0oVXdsLqSkkU7zdLvL1l58HE
6ZrDxC27clDEVb04iS6a5r/sH1omtyZJB6KFY29NwX+QYDkWNoqq17eXMKXOtXDtXx7ZvgLGf9EE
xHoks/DNcuuZGJyBLTFRkxHYq3cLXQGlVGXhDSItT1q1XB76W9xiZKsLmS6ynKKoDqvfrlFvmzZ9
YB5X2Gqg0fPTFyYQabr5y+ZnDkaXCiilBlBHN7Sid0P3HcRjrMFCXk1Se1drUyVtagYdE0lbVPtC
adNoBjA4AguCyWCphcCGaEFoFY5OROSi4WenGTk1y4lADXj6nlFEuFIEyWO5a8EDaC0o3VSjaD95
l0TL+jH5yX65W4GvYupvc/kEVfv2cCkHeXv5TfHnmK55nfSC1YoZFIr5UCmKS3QwGiQ9fLScUkxe
xRYol1ltuSd328sRNn3TC5YaIOsdlQ3isZxesexWfW33AopabgyH13W2yZPgm818buxjj0C4ag1T
8C0ebSQ8CqZ0s8h+/KuaKngEZbmzMNWslQVCfmjO2SY4x0a/Ikv828J7Z9PVrtth3wrjnuLWcwry
6LpzDwNs12kyQFFuf4jKjJb5UCAvU9euD/5ifsj6vzCXxQXnzX53+TS0LNaExmdnQRw6hcS86ZGa
/3NTcyfDEtgwg4t83dIxOF1lbLLM5uA3Y+aQ4NsoOTSdG2hR4/kbmcuNNi1aKVFIPLo2uGylSvei
S9FpEb0cQ2TcbhqHjdbFSL0+tBrEL3P7FhiTLqB2lLufx1ydSehpRlTBftKyphrOiEecju8txy9s
766+FRIiZfd1NJgatBCEXAX1Xf5mG2LtnlvtUxF4EFnzvrWJNFntUJ6DEGjyrKwH6l7VBKd6ZA1n
MvGMRbqO//5h9ceZ+KDFE9SVh+BFh27bweKLjZXR/iZlCmkEIZhO7yTGpjaLpLvJrXXPhICvFSE5
GYKPDPiixXGE3HcSOTQV1SVphU4/SjWm2zV+Ibi+EX+VcGbXzf7ZIkGrK2yRf21qYpyaRt1uJ6DM
w+s2+xxg/o5qRNnyROqmQKDcGvXYcRcDW9TAsp1weGwYp5k1RKQ4GtF+ZZ43GUcAIpcpgCQ9Cceg
4E+7RH2rmUN2c55f5/DyD9ICJ7QW9YqFADKtplwgNIPO+txg50iYtzjf5VfXCUvj6yJ4socZj9XT
sdiLrZiiSJaMWtEfmHkkCSXvEbscxKBFXV8auKY3gzZMpeMtt1FbLCYBCdufMfS5iNZq1EATN7x/
pBQ5M99Yvg8w92PeOrtuFwz9UoFsoU6UBjJzRAwUSYYcgaVKfjNBrYBJkTaVcXjX6+w+mUr4UXQL
NaVCOom/LCg4+tgV3Tt5bpvAopgZS7wKn+t5Spd/xJ6RoeURIDfBct+fTc0n3uPK/TiGNI7tLWQB
P7JCvCBB5/YFD2zczQBFUrbTI5bU5TlPDOu/zgmncFB8nTyVvMBsAygCnhJcnot0mmyyCU6Ytnu+
Bo6eSgouzT692Rv7uty31eyA7sfWEZ716tbSNaZayigjQtAWM/KrMvbBtlO6aowPjhjHuHIlSyWn
UOidEMwCyvY9pOAkIF3VSQDxQBNtXS/iGqlcpUqepCz4b0Db0pT0tTjBjP7VKAQvRGeyX+HtmYJ0
aATsCNZ0VqFEdLOWV9Hy38/VQaJnV1C/fiknGFQfOy/spUodNPb1hNKuCj828cMH2VWEwarZrhlp
aQZ7aSX1MsIANkOLKQnwzS+NmijxkglN0h0KrwEGpodJbLZbDKscT+aqX+uJqw8rX8Tts6Q628tz
IHYJ+dilOqQWoXS2vrk2S5gnnPv7Ki9AF3GmJYcNgEamHiSiTJJLCu2PRAftPzOxPgDqHgZki0Yq
JOamTu5ETky9WWgZsiJCWSaOAsGCgFngseGT6nRoVj8NLcYpNsIIJoXg1zCD1KqppQ9Oz9ldJWnZ
0YhJ13xAo6yoqAt6Wx0gyiaNAAaPLWmGHSlgjmTL+etLptM/WnFxFkv6D/iG3k+XogvITyl8dpQX
FNquTzLlYXNi7rersy2jI8WLiCNTYIshGjyjHzwaF7DbPbJ1uiFmWOoGWlZvUfZ2l0l11pXpJmwI
VB5ATQayI18/0LJbtH35Hqq53necZjeJTWGox3zDfinfSaMm9jM10iJ9bp0Uh42l3UXD8UvmCm9x
TksOg+fuodMM4KPyRzXyCJDEG/VumBNOl6fsJlVENW0Waao5xO2xeXTPa7XujypBFyMLQr1majWk
LZVL3liHZwIXgSDQzTRK+ljw3uIQL1R0Ido/Vw0r1GsVbIqMR8G721vXC8sDEHosvctoSGp8HEZK
CXF8BMd3Lig0+QR3nKUyEu9mBQToXiIuRsghsBRay3GJV+VE1umQdR12pOeuOIc+1Kpi8meh1DE2
dcNvXJ0GOtIozgEN5zeK4TIgr65aI1QES1Kk5qoH08GUTU52cTIXvHVRRavrJpZ/f92/iiNeJYpI
VKTPvifL/O5WAj9WqgjwqmjgjECA3CYTFTzpK2TqDrbE3qtmIyaSTgYJz6W3cuP9mnAFSu5LGdex
D64nJAPwJXkrsb6oqH7FpIvs5S2A6xWhWVlhV9kL6Zmo8+pr8T19QYgiDx5Uq4CXmGNIUNzgW9Gs
xW0/wRW2s5XFcBycQN95rjtsI30LErEC1+fiw3VSRVkSAl7KQWpQg7Y3VvL6oYi2AgBzRXYipRWf
Gsr7NC8+s00boyY5O+BGQ+FrBVrujRfEXVSF/CeGBoB9N6ocwJaS1xPILjxG9W1xJJ978QnXR7tr
zQbhki1xANp35/aTzHCR6oEF6EIOthR8IdAKS//n6yNkmTYlBe+1anIWeiQQMEwgHV4yCkDL0TmP
gpBwnYvJIqj6D78iVIkIToeJ0CU9n8tFSgOvjHQ4IK3ihYdSRed0AjC45OlZCudiHBnVnlFhKN7J
cg6nHzCVx3khGj8lymLCl3tnX+gipe92KNF/xqwr5XG8kJuW02zK3RZ8s2S3DCNLEjtxgpuWxtB8
LgmmyZSuWhf9u0bhon5zM2/e/SJEVFA/gCH9/tZjv2WiqEVQ0Kxvm3ePSv3UfZU/p57SE5RYpc3X
yDrER199w8YnAJSDB5CUSn6tY5Kjw0NkXx4pM8bdGuUOHchUmBO/UKknQOXEL+avhfW+/Sc0tVp2
6HW80JX8s3Mrlt7TuP7/bsLLioEstQnLB86uKXzZkW3vpabyUzZfi0vPeIOZI2ifYHxeqrnEm/DJ
Bix2r2jLy7wHW1lK6i0TJKxgy6gelwuEuwP81OLtH42pax8w1O74vcyc29CB1K01wvnioUOcWZJE
14y8kyZddOU4eHW/9erQwLnjGBSlENrm/Y89tE7Bi7aX+vdv4YqZfrxKxFwQqOr9RCx+vwPu5ygw
byUS4kNHwcHSfY1hEmqfMbFIdoJOWr/KvSbdWMzUnVS/qtxbtjgz08T5gdQ5o2RfeFi40B0xZRmK
LPV1wwpvGv0CTa+/DxLNdolGYW6lakzb7JGcJjF1qJ1yFcL2SkO3dTZkDyZJyj1C09IG/ZwBstOf
xG87wzLmZbm7p7ZDja3//Nzg6x/A3SywJw/O8QPXx+m9NDh+YovmU6uqYHkjnC34SlljoN8H/uzJ
LaOCAm2Bm+6qMAoYWGIp7Srp/t8jme3gmBbUbSGrmNn2m6ZLsAGA2YdGwP1Q/GEA2bEMxCFe2I7d
INVSydnnCyuTB+lyC6jzYq2ud4KphbQA+KEcUaY7Vw0aILc1VeGBsY2AVA2oUztoH5YFwb7W6bT3
SLZ/neIUhkou9HTge2IIUislp5OdcHguVUPTJ9uhsHMfUivpjo0bb21DBN8sK/gkqLZ9gLn/ZlEw
tjWMR92zU3e46+C25hmp4N+uUT5/FkrFRY8PpMnMIg8YJJYWWy2wmmo9YzRaOXuUdWo6qEFaCr0g
RIq6G4is6eluCRu5aB73+thRsecIAqj1IU8Nz5gRYLUOAEFVLyL5Kp934ecHn/y77wfeYTNZqB5d
viBsTARMhgf747Vz+v2bPbj8iTxSjewcl/pY+BtOwPzFoxftlvbyOL2+hHuWUuM/nQlHxu3j7aCE
i600ZVKmLGZAVva1rlJ29D8gJfqnL3AmJlFE1XQDzxqolbAGWJz50Uyxg2/sKC9DsnoX6t9CTbnN
sn3xOokEx5SBfjUWuN8tIVEMngEXMXi/dF/1vE+0sqMQbQo1DQ/QuZQGl/9EtzC4cIYMaktQJrU9
vT1N41X3n7Gy9TFBMH9F7e9WcFCtH9v2G+3o5iUGPUlxIxR2T5xYFEwhWPDsZjMqpy9nZSRfyri4
c8voz3kGcRxJv2Ma8DOoyt4PepRtwOjy+aLivIRhb2ps7aXBbdHCwvS75cwqUhmewvBtYL7HBwML
E/4hzu8ui2/kYWzTPNr9C4y9J64xtntgDjn+AL6G4E1E+Fv9oHheo8Vh4gW/qTxbV77Lm9LWtHR6
9dgwCBmbJMjj8zsYc+DUG12lftBO+oy6hRAeeHwTqKI/EiD8zEGvgwUXdF5weGFXFk1hmDljvO5c
dkHOa7nDnxpMOpORb3rXD2YDzrfWL9A38z2A/dBIexPdnSZgvo9TkN4E3CgdipKDZgoy8/Z0M+6N
oiUutxwxZJimtKx/3Q87bawfEYBQlSYjI3bv5V0rmadQqTU/HvvG5q9w/VI5xyOYWx4bjBpUbMQp
l+HWwUvv+auzw61JmkAc0F8RiwSF05gLc94M8IxCYBhtMkInd8gHJNOlV/vuEfpYa+1wusZ9RjZa
8H7WOYOS8SKsGmwa4at/3foAjsID+wH9WeHCu/PDSK0Qa0qBZ2n7b4TGbDh/l25QrWun+FseGBRE
4n2YKPOp1S1GJ0y67gyiqdUfLdUt/w5YDCSRCNGpBII90g1jmlxhDnn1I16phOKuocCp3qrhFNkx
s0g6ez0zlKmzgBJkqPWWLoVPgOVKLxAXfFRk7GYcQ5kYBHzs/vXF3zlu4L4fMBhzKzkVbw+gUUyc
reeltnhEh0Mhy3w3ak3HsxWzYwbCXAalrkS9iMo4yT9+2txJwkzgumzjEpOb/XjWBDpN8X/0w9Jq
7JqeVtJQeo7aUwp7n4D5oQgKZmEYOiJ2YnsFSvXqmIe1F4lYRrRYBpEti/mxDIDbANXKR6aqpxVL
LLlgH6ftq0n7eH+V8SNKCpW32EF7dj4+gWjnWajfUeTobhzRKRRrR11E5UuYIBF23KZhTlz9PK8c
6pnw8J1WqMZ9E/BIRwdhWllYMYsFjCpSEmTvNBaZ025t3/aZKbG0ftFd/BVKxJ80sxESqUAAWJvb
Pe0WKDiByfdluJVIzQhlgW+uh3CMqIv8FnAw6hn0fp2Kv/6SrvryhR5Ra7WQA8dHFjOyeL8Zqpd2
Z2sTIVO0CzlvHvX/vhlwxVvQ2IwUdxBLjJ8Gl0afbvMjflF+PQyalB2bu1A6jdqBEFpu6EehjIjG
hD0gpviRbJ+0eqH6jOGybieneW+HB+hIukHr2G/0/xLIvJpj8WlcoGkoeXUNFyeJooygMN3ehHGJ
OXoOlccxTBIZh0noKKrXKg6jmlt/0OdB7PS6YdtJ2PcAl2ftbCM18TO+dm/ccMOsygjwyqPI6NTG
KJR1FyvfskepVfrb/4Kg6YVZ7oSlTRAp6Rq5GoHgt27bjVPG5XY5WFMokg091cvsae1/4U7fbObz
JA10Lm1NIY3V8PJ7BG3Zw3uV5lZs86fp2E2u2evEzFUSznnNFERCY6PRI4rbfis7/pDYx4RshKwI
acDrg9RRj73W5WHf03IzHQCmlVgx8sYLpJ1E3aK94ctMaKzphRwhYYEzpKX53VYkRSgrJyuy8/cG
uu9uEzTrlZCOFSb58SZAUievTNcz9R2MAmq+r0uLLQKzNNGaROGQa5sWSAQuXCjLtf70N50/KaIN
07tVROtno4nS2OfhnkylWDcyr8MbVDtLkvrLRGbSo/REdHGQXfjWz7Y0u+WzR7FSa6YvnLL8xV/5
oqDwimU/iZS0ps0i2PEdYumTQlTNvVKCvx+9uc3wshExxjXmK7tplHc1dVw71nHdCh1V/rrwDTIe
JSkL1cf884oI12P69ujp6gaxb+H1+RQzC9QZ8pckkGeVrW+BYO+Cg2NgCr3O5P9QW5L1hjswee/w
iT/jBAt4ihV0+sVeYUf8sNyoNtOlu/QQgkvzdT1u3l+d8mgm4kGTa1uoJzz3D1C6SsYXk9A3GHIR
BEdgv3sNOeiIM6el0OseE71Yd/MmWScVx8SyJb0uurQmSLZPPoMnatFlV4z8KJpwqGN1chsJn8Ni
FwHKJuYQpl+qohGd7IJ+TsxcZ9TYatFrWFuwkH+JFknwgU8DzkNDRljI8ln9naCxOZZmBtv6WZjI
sHAODLAsJ2kVym2iWdiXIUHfQmuzKDdM0+aPitf9/Di+/I1lDEMalXhml+jkCegTuH6iWkl5o5Ov
xA8sSHeDf631fsrL/HjjDZCxzZcfOSN8QcTfhCPmrsBJ6upb8d2LzRJfmInFvAxyk/I6seSFEobE
NeDc6ftzIdnPxAVEwnR3Il2I4I83hNaVKYrr6Hw030uCBLePDAVaxp/5txFAqTAnrU/cotH4AvEz
zNvDX9YoIiELzE6E+njgTdb8uLgsIy8Ji+djyGotBhafEOHkYC4cL9IWtXrcAfay21hp3PzjQo0N
TxXX6XjmuFEfUksahWQZ5Q9Q2Mvz8U75/xLCM5a/8/rgO75FsjeHoDEy4J5/QlY6d2J/yUpGdQ7g
VKdEhmm73tL68T8JrE064U1Wr26CakN3SLwnDtAXaTiYpJPJVxfq6ledNhOeKjeoCuJpaaVpnneM
IfK1b0mD36EHff21h4kk2fD0lOhg8YVtGBzTfHQt3sf86U/3NnQfA3Ta28wGHbIRVENq4iuhIA+6
nI2TJ9Az6qdyUSieYWHrOpBkq/uzls8EvzTkw2yRXedX4QV2GdmW5ge4cLOgif1isuCPXvUeSMTL
JICffdvtTGWgBWywmj8WetAjEjX79kK39Ig6pUvz/dwz8W1Y/z6OYx0lzOhVcxvD9KVMK7GpPHx9
iD0P6jOQpRRp1fFfzOFIKwBUN9Tp3tghZjeu7hLccdXX1BdJiAT8hUdUvgs9cjImAT3zlq7jg+qU
1dxfdLNHRT3/H1vFPmYHzvbGEZaCp9tUMZng/GiCP/u8SrCCNRx83ZCP8i5EgO0PcxcI2H3i3jQQ
WxLaWEDBV8fgu35TFkKaD3qifw2XacsVhjWuaDHBV8VtvSJZ1kSYpOQi+kU7HQtVrLnX/yY37kTv
u0Vjv+K+lDowgR1VZ0iMC1tsQLBtNFWsu00qVTApns/Nu0rQmTWLv8XPXkBjM8orDhO6E7oA4o27
IXsvDV129s0D57E2JfCtzduPpNYRxea2wf/4RAICZLTT6bO11EGLvBX5hZoVXKjkFFoGZjmw0/ms
J6Rh0GPnTChXCht56UPqTg8LbwlPwHYTEyqL1nKRBPt5S3tsaqlT//L13zoGDA8DEfBQXemIH/yq
YENoAgJEtICOeN2xMmYAm1YznrdZEohQESUAjFgtNiQbcZWj7hH/Rw2V9fo9QlfeAq6DYEUu01Jb
+qa0J7MOGQAFgQ+eJRVium+WmBNB7b6MKdZ1+m1Qtf/gEYGvBTF1j21uL9xLNfds1l8+yAxUN4gG
ohtuQS++uVtN1HYuE9ubEhPAd1NKh8I850BsGr/A9lz5sNb+UUiFnZILNP36lKMDnZatLR+ygA34
Z8HNDfn8Imbo3c3DzDgoNd1qy3JDjo7PS+Bd/NVLGD/qGhKh1JbNjcbtbVZU6/NmqPOvDLG7sWrX
pOtP7L/VkgPtJgu0hDKXCNAlsiZPiXDSTir8SbicCT2iF+SIIDyUrZi3maPgC2cakOvG8TbgvQZo
LXEg2W0ejXg5HFShQxd0VxNfsiXX/NcUxJpFzR4PpqzkZuuGNuDL1MgCkfBACKOUFz8rF65w9qqX
pUYB9A6qibwPUAyQqi00jm8ViG2txMJuJylsMtC/tno8M9IuP2FpJ+OzylqfUfKz6FEUd6sGujbS
YEP0ytKk75Ut4XuFrVLzFQ/caz6XlXKZsZaPdVMM6u2qfcx4XSuR+4RLdNP7p/nxEiZhPnR2tHrY
y7XdlWaavSAPpMSs4lKPDV16+DD3CDjp99Ds6NFRrVU/b6n3iOCkxzzi7SOdcPqbqphdMPLslCqk
6Ptdq3gmPMMWPLjXjAgiLfY0W+lg8h7fKXsW2oeZxABxgfXqrHLTP6duopyICR2g1v6b2WUZ9j99
fDpFPv84FlbPbG9ZMNmB2/28OUYgXEqLCaeDP6tV0RV7Ovu6avrQLcY5Mpu0T2AxVgug8eeeEyFL
+ElKSdmGKBMmgotY4zE5s512C73L/+3QGNnujK3IC0v3cGpEqQiZ/I4KdMk5/EmsGpaJg5ymQo65
SEnOswS48z3miWVx+GPY4IupfaVYd7JNpLkiDvajycnfqxqn4b3etx0AJKWkzjXGWPFiffGug7Uo
VUs488Wz51vRkL/b/wwou76aQPitw+N5sVv1FvgRm+Y6gLViaqGJ3d1BVKsyGdytjiWUvu056hbE
JnhbVxOWeanY+DzHqzV2OXbvz00SDIo+tfBvy+7juXzYmqNH1AIXvPcFpjqoHONJkIY75PkiHMcy
wnv6Zqjp3kP6C4nwxsP/M2ZT71XcfkDftdTTQbW13seYJ1sMgnDh51mctXsN2InBexcJVFPhqzbJ
mTzTICwzbc+Z0QoUaKiAIvhNQ1irxX6BuoCvsZG1NQ0jzCjxU+SOGJ3AysqhzPi17aFwEoSwgt9m
QfXqtcXCHq6u0V8Of1eyP9gqm2ZlGz7VMQM3Cj7XJ5C8RTr/atx1dui8AAHdeNdeUSZEY+yzDs8E
Z/0E9yeGTN/6Gf6wkTFY7tmuUgg5NVyecRaUILoFXrG6SGUrj04LsspWHCd6kFmpnaapmCMK1hV+
9YDx5z9oCilIdZbHcpQ+nvQqMtUT6SgL1LyXopnlN0oBFmyCcCFghJPlqjehC9RemY9ABT/KRiyT
vyFD0EB0bbPYCxT233BaoICsQW8Cmm+p7q7BpUyDYN9/X8rzYUWhzC0CYDtG5N4B/zifLc/QnA6P
xUxH1kGlz4EcZa454kTQcLGdY++AohOKu8nl6BTAf9XLGNBqquaWX53Vc2bOtN+XyJDQoRtyu9hj
+roIMtxDAv3ZndQ0JzAPkZhLdVZdDfvv24//AYlCUfBq13XxRtv2HR57BU6Ko5r37RaI/YIzKTtb
ub5aTAwTApDTpFd2JPmj7/q3PwanHOMlddgKDVtqQREl7ds51eRphMKBAdoxMOAXZT+OK5Ygqzlv
NFdZDvpEO4nyOUeQGZx4z1eszEAnWQF3WCWoYaFHc1HXN4cX33H/o5tlClCxtD7pPPMUSfNvUtkh
DajY8NbzInLG5UVj+Iyy9qj/Mm2bjzkjE3qga3YHMgIznY+J3UpXdg/u1XSi0JEyyB+Wo9CzOzOV
NJwVT9Q7EKwu31zWy/05dbyOnbsYxqXswMnEdioKnaX01dme5Dtm6wn41rf+5wtlBU+ItFF3F+/+
KHWUi0ngtAFLuL7/RCtF+1pEro0dP2p/7wl/KhWzeLVFr7HwfvLvNLWYo5QLonEjfBax+DLNhca9
zYljSZs5BTYiSKgoH7Ru5+OL4r3Bj3VlDkNDpOMZ2h13o+eQLJdS/voibxi7Ww9unjdSn5oqIbIP
p9tekOypffbjckHoJ5mEVNi2jRjA3gLXd51cgGtIGPwVFKh2jZFG1VWOFEHhE54ma8OceH3Zh8jv
bf9eCmB1fubDAvGNOfUGlFNeTvxAenW+grAfWv7pz+K2pYmgEC0rWE4KmhRW003MGdzisHS4FBKK
0a0geHLuo60JAZgdPubirfkx4UzfsV48hSQ8PUYNmDafn+Y0pbHzmRan6PHOZEumKMz50g/sUwkq
C4FtSxFBIRNEE59EGPcCshP8YPIgRjVs4xKzGEqS5EywDbdK9DfOlmzlfcXz52oYv723W1LCKydz
WFxuB3LudbNMp9LPg0FexsKbmqn4W0Li4iXSLkW2phzoGqYXBrWaGlBSkxnx9yZ3OMP8S46guhr8
d4to3CCtkcZGbgQaLmqrPj/UmWx8u+GVaLWPrDcQM2Hb6Xu9/05cxCje8jajjSW5idnwi9zvAC2l
k8wZ/p0v9CLG/TtBMwfasKOpnpL0hM78oh+1AYikkFEA4ixjVorjLyUOOCFA6I+tZRUC+40cX8Je
giWJSWxFQ8AIpcnt1ibNIPWIhaQkYWGc+kuT7NYNXwNfrrhlX81i3kycRCLbY2f6+oLldGRFqP1Y
Qw6qU3SEoaOpz3Z+ExGfGBnmbWbbB+5Ostbb2v0iE8xDQflFz1nXD/Ui/3NSQAtxUI9m5wMvXxn6
3jNVxvsr6EFqmea7tDHBZLXEwm/YK7co2owfkV2fn1ZI3c2G5KY+XJiPkB5Qj8CdQMT/jG86ZI0b
V3LzHj9pWIhWKPekCaoEhbBwfUeUpFc9ghwkKjb3LJWJqRMD+bgRobyJCtYXPLOcka1hj5ddWA4s
pUQ7Qrzbki3l1pOW2RsLnYvXx5tNTdTgsrAbkLMiK3RpJDolvZuyLperxyedzY7pUdBoo9uQvObF
9PKcCoXYv+M3MOrx7/y7/gscaER8fFFXBEznJ+SqoVWBifS7AHkSuN7+hjV/LXesn/WJqBq7RUUF
MZlaZn59JkrxzrGd1JJlUHX38kB+pfJKcM+guSulMbxAR9+IR/ufrhm6mAQ651MmEpouFscKB86T
cP4VsGCZ57qpVMvjqmcR3+Zf3smmXkvWp0lkyLeZpYmJI0yh21PMMlSQeO/BMdGFo1gRF5k4MLS+
OfBcCXnRr3g69YD9Au5+/BoOZ2TMvgW39zOQFbS4d/Nyzyp/fPcV//NlXZ0Xz17C6d8sy4hlhYyG
IGLLEqnpHkSwGCpxuwfiJ6wgd/Iw8omtA9iUDNsh1BPJBM0Yt4CiNTac2K55o6D8skHJV1S8QIlE
fcHea31Wir+eif9VUaLIU/V0C9BnsOBas3zfKz392E5yyUhO35qYQ9CECCk3+cw/NlhAKYom22c2
7fnZ2YaZxaQqXL5knkRhXZs9rlqYl31y90o1aGIblzS/rDCuhAO/QIdantiXM6EXYsyIpwBYnnV1
TT1wBITT63tbMRqlK8GjdldxMh4GYmIL74yOpZyltG4N0BfdTaWTGMqCCIE1ezEfn6iW1YAVhntH
H9trZ11klf1JwDojEJIxQfFf7Hq7TA0mkImPWazuGPZRVyKKTw1DtbGiNCW3aN2J1sfL14Ky822V
htiWoVlcImN/lSLS0K6vqiSRqwVF9GamIa6gFRU5Ue9nUwJlObiSfYc8NZr9qw+hMiqmBrjKQx2u
TQzVDh73qIv/unlJHdiKeMSk5D98Cqv22wcsORxbEK/eL1yckvQJ0EFQysnaF/NBprFpPS0slW2B
eVO1z8LRgI9JWfOYeF5raLOdCOeoacwWFNtbTsSkKh7xfWHxgLqsrJKggZQnMAf09g38/5XE+v0J
hYrseGwXkUUkpIi9tJPloXdv3zhZq9vZiCLonsZcwFYs1Ye/nUOOMYEgZku11up55K3Xz/wVBfpW
x5jXRwQ0PhQnJsnM0NZSOCUFwqvMgF4R9h/w2q+TCoIbAblJYGItrW6Vsxo+oTT4B2pEMAIcRTXy
cghkwH65WybvVuypsh4AWEh1bGRNv2aytPbIBa0xb/H7be/rd724D0eUQTBaPst132xpc/cADxRL
QZOuwwDOX5dVF48yQXkGEewu0RiVOaC4+OCVCdceRkafzeLplQjZLzRsby+lb1Y9pJ+JaOn7ZQdW
BW1EwMJbJizrwzG/okhAJnaW41dIiZ6gw/Jbo/GoNjyZ+RTMnNcoN0McbEjHlG2EyAS16+gcxUj8
kp4KXNGi4EqgiYLuKK+OW8dVkQK5CB0BPGmI2+1SG8udZ9fETotcAw99pr0kx2zYq/tG4U5D01vi
GqZAKqFdS0Ed7ryit7dB64iibkmn9fkdkvvjKr1YWdm6ppTsBm1Xbk6nLGHjVMEeH0XgyyRXbmkJ
ePDJiE4Py1xNvsAkELtHC8S2wFnebUFr8AnQQbBeNn6eGv/FEvdnKfpXXJdyLvnhc1yw+hwFe4RO
PiMEa1qFkHvCcCwHAhrQ7xbJyGM5sKzCBLhbQRK96v5LqgpCo57zTPxtSsOAExjZ1hRbfTXNBlIk
BRcK2iMIyOgxAaNy9nRv1UXbK5UkE0xvIqRNNFGGVIl+TMUXv9O5IAkpIppOP0DwQ7VhR6p5O/sp
uZe5xi306uc0aRr1LAhrZ0g0GxhYWq8NHlcNl5gZGYgWymVS97OdO94AtCf4aode5HGztdv+KHDP
YKL4sjQnAdIqJbZDWL+bT5+Hs+LgnBd3j9Pc2KHafJay22y2Lkv/86y0rUd+z7G/2NMVQQylxdCK
sZjPYaQsioCNmtMlY+leT0nndjtnF26xc6rGQx1kaAwpCr96f/7Cw+aCoWGHST05kw9mv58yVHWs
PRO3GYBwwVCnnLOjFj0lj44TpOANfVps3zhPFW7enIUyzZ8JSIjAa8imoy18YTbcpwe2z+e8NMLu
zEyNL7fCKdbiQayN++PPVesfovI0mjje97spyi+4jcgB7+xn8pPzVJgSNOO9MV35tEhrfpQOxcCB
cGqn5sH8ia/YleJlUeIfX5umhAkxfUiYrATNzut+dmpcRFgh1+zD/ov8XE9WT4ZvzzTWPe+F0pq/
fq1MfiSGshPMnPu7LSJuyRv6osYXp0JNCrU4powi/fLslmtBmr9KozSB3DT7nOiQnnW/CVnyQtGr
A/5snvELWV6WfDqzdxO8GPd7G4I47imaDQ/9syA7ou3+y//0sZjzmNi2fRmQBf4Fo8elcwwHdsP6
TF2JHSMlhkPbuvSiCJmJP4AFuU6YrzBNQaDQwdR734ArkaEgZsqegIhz/zrTZE7+m1OrOie+kSBp
tO77aeBCfBbMhPw37H0iKMNVgCQJMBi2hvAODNjL9EX+UrYrNphkcmLDEZytOM3pIp3dFa1bmps+
Z6Y5oGZPdIanRof55HTjIQdPLEOPile6tQwkUFn0oXe2YY9mNgDidCNUhd6QpmgUhjZjkPHZAyN9
IW85zm1mcsKLxbQZ7QgSN2e4deHdpxMX7QBqXhTGhGeuEzmF3LICJ8RkkqDR27LZOJGamXEqZDer
0+S2F7RkO9vVs8apJuxV1I9fAKA0mmFj1CVTdV81/lgy8sMQr/eJ6b5DnQSp1/x9p0II+zq3ZjC3
V1tdh0erZzzmhkPKTpgWQw9uDRE6AddoDdBbjiJ9ZWd8ZJxXc4AxYHsTTBmvfu+M+wflIhVjzBvf
Iab4ENx8mN/l1QzsrPW3C9jMMgLMwfVQXqsxX5Nz1t2OxT2SK/ezRZx6kg//YVR6+xuoOuD8G/ok
VbGtqMPBZNC/QFlSIQuLu1YG5zRbzU1cori0kQlLOdqaAQsV67gLSyFIcsSXsQdCsixlaeLhaMCQ
Ezk30ud5a85F1oBFSX9jkvm2GxNUv5keh/p8irgoggMIzfmmF0ABAHXTBHzojt8mDKXtNLUH6hfg
pA9nl1emBeswLyVmzhTBz4X2HvkOtfrNjvoAsQT+ucUNtRYZdRsspKskMiBTx/YiK7MOq2ePtQgX
McAAayLZM5uXbQXzJrnfX3i1oOxDb5yS1zbdo2PyFWZubuBh+DJbFnMSDUjO7SbiUPTUKt8BSFIU
NejgKjWrQOUa5EAKfMjrwCwPwzDy/1emw7W4RWI8usOtL/9O+EVNpCZdMzfpgEPB7fOcWyyOuM+B
n0G4lW+8cXJd6kbXKZWk8UHpJv/dehXJ7KyovP3knY2MDqX4XtPwD/KTYBIKylELw/w7hIyV55bY
IbjnIpVVsAuCyvbdIv5yZZsXnj+RA8mKMmiCK+hWdieCDlU4z5Mw6/l05PdLo5WcBqh1o0j0d35g
BdV7Vy8wKkoFp8AMSyAwLwWb7lSGVFumQdvl7OMw9iN+L/oacsJY/Or1HP5uqUCy1z13junoaHV0
KA2NvTkYXX0M+xqzqRg78Yh6KQKGUEA+FAVMaZDKZsS2Gc8UHLOusjncN2sMGoa4qCuqOJEQCKf2
JGe800rmoG9v6ig3wpQ8TS1NHPS0WikLWe9lrpwsGcs7sIs8t3F3neDMvDrsHPNcYr4TeqUDXpT0
XasK9x9DZzXdalMvUexXe83sppXjA/6RLGJy9CnYOgYWMYrNXps0dhLRANl5gaZQLW0m2NjC9TTo
BMn9katFBAwxH1B/P+Aj5cf19t7AfawTtf+Va3+zhthAqhhPb2gXi8UnUKPlJjUp/ckPXSVRwtEK
cap+I7EfRajHyLcurKf60pRlNKde8wNCrc8K81YkzPeNguB9BuzZ9AprJaZrEx/wanaXXWK7S5MD
iqhXyXXmBKGwhSS+NUm0nKUytkkWF5135NnI1itUcyGM2BYj6udKPTz5ttCxKRz//JgKqpCGd6w1
/TXhJtIm/ZFMkbPpzAMQyPjlEuOvlToIWMvYAAjmeD/Ku2DJZULPz/Yk4G7PB0TV2JoFNfHDHFLC
PIB8r52yYAeutwnCUnuUoyJt2Y4sO75PVX30OPlNWxNWun0Y1ecKXxh/skegBlo0gbD6lHqdNxT8
qwKhui0SXB7/9sAyZJ4I5pp2Alpxw4+1efIu3oQBxlXh5Gf8lYyxC8Fx0byGe69O4Lcq+BKYC02M
LxySOnppia02r3pki1UA8Xhb4yf3x3txXwEHzfmz0NMm7PUe9LxeeLP/2d0Qu23N6Iwg0NB0xBVh
YLBjdZ5VqooYjISVrv67M8hsJpLWzTNW7vxmSY1zVi+9zFCAXsnybPmuTnjCG5t8gIpvwVZ6ZyeU
RKwk3dI6rrtMDSu12j5YE+Y9KoLXe1SjrWugw95lGy7uPf1Eo6tAHp1a9pW8eiG+aTDOWGc5gmMc
g0F1shbOy19uQNMf0hyC85REfJGceADwQ0GMQIQs25tDVgJOhEuWRJTzOfh5YjMuMLhH/0dwEkT1
n3iIxL/iGFkPbku4BA7bWzbvXxF5DvbxXkvf+O8w94kQ9zLnN4WQB3A8p7jbRF35AQZkaLqEYCn1
bi7/T5hiPkf9IA6hCOAHig1wYJauVEXst1ZxIVM0UEXSL4x6px6hb7bvyWteEXyno8yMFpFULcBm
yWe5HRxCavDzxJM9iXrg8a2y+oBqFExLuzGe3LnDSda05pEJnIX85CKRkVj/L3E2gmmVv1z9YTeL
NYUZjqc5eizhg8m98SwNAbqbxrLXS0ZF6W8KHLYdd4FBpp41x9uydLjAHIklP4kN7drrOV3ciilS
iThm85KbyCJRtErATAj0/2zhQcDG1fWpdjxiCoGFAHElquzDvEUV1i5dbG/2MzK7AMC0qk0x/4FV
c1Wto7+GapwqpTF3UY7Ezbfyo1blgrxDB62lrSh0pUihGQNFUJl/mPTiJ4eaiC/Oa/5gCqkfX3xx
L5rHNj+fm464yYWpHWajoJP0khDJ2ZEqh4CI562JqRjV7ryaripRd0rfLcOfdBigMeJ/0vaa45Gf
Ed1iIRGBxUDdeHGuTP2E2asaQSoTsX0xcmO20WPFioHqYONUQ9MiAbvv58n7C4fwYr7lNJsNGrMO
mVeKpbn+dInBNd/PVxNfa5ujYKE5rd6qOmNI8mXUp1juXThsITjfkyaHGvLUxQL5/Dh8TEttvq4t
LESHt+aNFObJZoYmVfgi5q+8vYX5kJhKO1J9PnYDcgveprk8Tqk4oinztlQitf3NbsXQl8V0D98j
oTcNYOA3a4aiDrHlB56E6lnLBVe4KKxVPzefW2Y4PVJVqWuP3I7drqypHxi4tHx7ETIWiAneQlTq
aZo2e0xl9iSuse9FlHw0N632JIPY1KCPXTdAVr5oibZWzaVu+RPfLdc8EGAN0M2VZ5h3gj+K5u+Y
1bGzCKLxF4gzXpxWOedb70GVQjVW7byLuR0b/zWxMY2BPY5oRpT33wZiihyOgLb7y4Sy4Ioi1Gqw
DkZWZ1d5BL1cq0GjarfIoMwjmxFmb3ncmTnqroxCFeR9uCCaLbPGSrbc1mlaHhd6ol1Mva0HJdoF
rONnIqcDD/I+t0q0iAlm8IV1Ie4W3/nCFmNhMOAxGaxEwgeNqpokmjZ/0i6ZDmor9gJqwwiR815G
tAv6W+xaARn1aQo5z/kvaIbuO/JIEut/hW70/7wsFW8lgWiNB79Noto159s5WmMjzcgvvHb/IPAE
qZ3vPt00SbjSvcIEpOtKhlMESVdl7cb2wSXjgMcNQH2vPO6RNPXuM0NW4KcWEQWXke3t+OotYvRj
DTwlhZ+3dfJsgETVqGrpcLgx7XsXFldUCBWJ3hS8SgGN7wKPi2j58ImcBTmCjAJf7UruSQQ+7QbZ
Ec6NvmNmWn9zAkkwpG+PO1Jw0Onw+sMgnH+tcnLTBwyuLmmSYaVTU/obueEcZynMTj5PvNoNihpd
dgZ+c+g8KhxzEOCpJ0B6GgLnR/Zxd6T8Y8KnGNT3MRR3411TU1fP3xyz22NENHVqtKzSyqkUNomu
D0Sq1+nV9u+3d6UiaiA77FL5NDb0XrYXJDEnu1lJ7caQ/WiXlOaedWyD/WgtoqEQClKT5TlQgIch
NNK6+qULUZrVYTGkllSvShoHaZoQZqSFE0Bih1xo1eoht96FOaxG0blcM8vfNpeqVfYrpzyj8RA3
o2ShhPcFncP7VLdaemWfhBPR76JTDbXjqrC0ZO7VjtQnp3gS9kGmPeOzMCrJfpTzmH6ZjTYv1DPo
/Cpc8zbnlKhasS8ukvcusJjR5Cs3Q4iCDSKjPmADXT24be2+2HrYBUYsveeDbttQeJhw0ZIHxC9/
2PTYj2eHUTQwvcX0eOYtplCANCw582vvfbOmieRVH5I/W7AeWKfqeWjOrG8iZpSOlzklz+TW3Jfw
z/AUhvhHLvQSqNyIhqctPOgzcZymcfBOF1x27U17uyApLVgcMbcPsNlAHn9nuLndZN5m4LEioSTC
5FFV40S2T1gRh7JFWmQ3MtKiYv09PdL3wxEAxXaE+SR3oieaVCUA70q+1MYlc9KebcyP8LuqTfxy
xUCecMdYoWILn54xfa8aONhBI8k4qeUffGx+IfqqCHQ749gFT7A8KPv1Frbc4BumwQ0D/HAMAv3/
4eqQiR5Pasqqqy9TxpuMr3XOqclXMOm6govVIGEvrcIcGAue9BRmbReAXRaCMK4vnAucRLxsTjzq
4v8m0Um9uvAMeyW8imkyQT2ANGa4jvrsZI9726jeOg6riZHUFI5l2tORW1bFDFvOa4pjhMa0/D4y
MJTOqaVq3YkipyJoKsj2jv12mIWHQJbXgkHbPI2V0q9lTByPyyHfxVBxasm259Jldu3lZf6J76iT
JGBa99zpWW5O/8KCIqQ8PYwv3gNKXodV10/YiPMHvVNeUPBPnbVTTYGysa/N5R+IwdVJTcOdgjhk
92H7DJC/mjKZChZHm53NsZzGVsingiDlcVidsgfJq9JaCTFT1SbU/p4c0vwkU5cAqLaLCaAPTO41
Q2cMcZFmacteQ00+HbY2KaPQztQCSnSinn/kv2Zj+jGPvnrSwwOA7V82j15bc/CitBke9TpYETGQ
LVjC+nExcF046IQbfZqvs1mXxgHNDMcwfs9wBbgc3zDPWrgBihVXHM9BPDbX1unjj6xfaGHM5qfX
+d17U/2wfXOuhGRVOr7ZVz1jdzV6Gb+A1IyINuxD/f6suI3QqJTrtk9UqsoUYrFdeqCjD/jq+M2a
nMpmsZ6dht2cjXiJK4Uf1kiUBow5ANM78oxzX7LcXws8+/I1CbPcP9HA2N6OTsRetkn1oqF0D/Jv
nklEvp5gIjTv66xiQzpkV6+FZ5bfQZiyRxuJQJr+tMs1oPYvWbioTwrsR5Fm9BCt0+iiBuByg96K
bsoupKrcKJygZOXOFXlB6jIXs9b5upBmCNwcERmjWRX+OqHKAguHSvlvPQXCCzQhVCatZbJgA+8Z
gWos5okwRiySOUo1tW6zWTpLskpNu8wmGhokflEiaVUND6uWKSr4T/f+NvYY7/+4keSuITEyFMbv
Z8NcfPwqxzx29O0CPzPnfpbNKUuZMAoUI46PFC8g0SJN4WE5e9n70sC6hRZwJQRYVuh1hxupwQOo
IsoTOfE8jbvFuMwIX0Y+jcLhrHpq2ou/IEzDZygD9gvN0FzRHu+lhL4EBkaRPOWno9H+4NZ8eGmE
gs7T3rXl6bjcDbrLZm6/FkQlmu2Q/kzNCXT3iz2pn4DwcnHj/UeK0pabkRiBXiJzBs+FWtckdKlq
i2ql8XvUeMIcXQKQlt3ylGGJ+AsxmVDSM/7zBa7i2DQJNK0RBeKN18SoMbuJxUchSk8joBApF1MD
ZgiKYCcqcCD0UCpWyJplOaaqNl+EJ+YsDiGAjHUDTiODq84k5GbOH+3RPHRGkb2jyFJS0iyrDLGc
XlXradgYJ/Bs528/+lf2TTkl7zmxqQIVc7kkNqU0IGQlv1FrxKcqy6SQIDQh/HbFtlmJ9mhhn5Qr
wTcvuTTD/DUYkG6OQS/h2EbxigJPu5E3i8qg112GUDzUPCWNEhjX6TOnwcqob0MqdMEI9gB4sEnM
S3IWWywiTV1yXSECTddvjwhEa118TqZOfxKY/gijmEX97JZSpa+eC3xpKNgVFpmCKnYvWUMbvkEF
cuIQ7ewRqQhF7KzVoLhzR1A/8cAPKza+YHDafsm+/c7P1owlUIHMRyAudx6pNfQWlLPjZBVVtPWC
Roqj8qR6fsjhoaeNGCY6nNO5HbJK65U2pTPrXV16dI7ELLljf8TreVZaOBGoIE28F9skPoGaToi9
8hC/JEsNhpmdNa4thevlmmG6nDJIFE3hG2obBinDOhxw/Qknr7TgFRKWP0MuYoE8XUng4YrGe/d7
814Ty87wEl+0abH02OhsoPziUM0k/VRkaZDwAF6zr8XlK7Dp8pclxdgS1Gk8F6a1lysjLvb+Qz3f
MKtT13Sya9x0q1PpATMd4GHXlNu7CLdM6ANPydlsD5ioN4eeH61tZkrkTw5c3cWRrg2sSdQvw4IK
v0EBP/xB/9LEjxSthrIJwEff3G9/GLMWrL91guaFaqfsm3GYSa9kCV0Qx76ZOur2NhO5TjZPry+Z
NJveEoBpR0X276UuHjGvfPoveJRMGvTebHdfHb82h6kdmxajZtKy4tNtEN7HH2bXPO8XyjtDBojV
9HwqP3KQ9Ry+AwLl/EiDzMQ+YJRmn37mdmSh/FgB2O4iyQ6Vo/gD2WnZCKIETyvrLcX10q+/jfnh
rJzyK0u9iJ/p8REIeI+qT6vL0HaZQNaL/NMnYpEagac15ruI9Z9RK+GzQeHZ0iD+wTF7XJzxLZAu
WlJj7LYN1ooQ1BjEfdGnHXSUeHLpbDdzcKuzAh98Z5uxdHcZwI7oMMVEzUZJ3iFyd0CsuIEUL/xw
qtF4BMYmCK9wAYudZ2jaiyzr04Njy2lzMZ0/NIHDF1DC8wT/QpUG4pbO/5C6eTg/a2Evbh39vQjl
VrrH1WkIx4z1zKYJXKkFF/NbD4gvCTiVbct/NGMojd2oDVGIaDv+A9nshj/YplI9nMthTGaXL62n
HJyWtmJEcXQH+0m4vB8iCqLxUrXnDEufcZhSbdu/HZRs38DFTX8i79ueF+Qlx1asumzWE916r0aU
PYi47JyqQiLB1tGSjDHcZn8TZjGZ9kITNJqKXi2wfQooIIto97QnthWcCkwxD9u0cb+OeC1Etzt+
qmrh+w2c+1TTV0pf0udk0HPvG9utgRfPX4Nrc4vQiIDtKKI8AyvviR6uMzPcj23a+c+UOy0G/cFe
CSk8802f7a+MQ8r91IIY327o2QVxmA6eJVoUFU0Q2qHowj5HnHQ2/4UmHwyLCN5npGBYPXBY9c53
iKdGFrs4Yp537LwMK2gXk4ztkV9jZgE9SsZSaCPXhZGvaoZb5ONN04kNphBLxltZQlF19rLDC38H
MuFtbDy3szSfPwmj8HckrvMdzZmhIvYSiN6GcUH21dwlTFXj75OmIpjvw0OtJEl2aJT99fS4E5hx
WmVgh9E5ZBBfY9Zeocs4rB8kQlxZvK9ZIS8B/wwmmKdBtsRkz5dFXCKk6QyqTHmU5Jrh2vj4lvzp
BnAQtq56617n0mhhSKWAhHnbr2Qwmhdh2GZPPTMsjD69uZZ5bvCCe/d7PpBsWmBA/7gXxWAVGZNt
SdbWGlNhHs3pUhU+xlT/y23v/F72YqPyxWIXIA5FEU8duQELN3/V4HzLNcVOKfhMC1I5P5ZvfT9C
eEnxZvwMKqcZNtPsJrwhLaYvteA7LFGCFVBFXQ/qNvlo0pLdoAQtS1UIRMt7N3TN8SNpJ4KO5Se7
PgzWBALpBwNAjA8RRPn8+3UgKX9+ivEU4jKmCkF12pA0fMhWHpIDvA8ewNV8TNm/ujVi7xBdXEP8
hcEKJJdhSHvm6mNGGc/RwD5GgQRdXJrbuLJfQvXApqWD7o0p1PZTr68/YlCSvYzqR58oihYIkTU6
djemAx9B/TSZgeMUYQbD+IiIP84DQLQcgA7ruu5lvYHzJCC0fbnEPmHxmfyXmNRnMPxZEiLK/l6c
NXs141FrXWWUpFx3W6fDFyBK1ekIJ0fxWglB18OycCyTXD4fnCZV/jwlHNcU4lSG5SBA4pjGPfS4
IiDk89Hpi62LHUsoLtACSYEfhD8eEe/DLX11hpi4JptrjCSc/XAdrR76Ibe0EJjpw6n4C4SyJYZ2
sFhkUjPhaEX4kYx799YNnZJhK/sRio+HBnh11Gr++V83SdYidV0TiLWz6RFs3yTUTxA6UCjBUQkt
nl3FuUUS5AEsLVKuMEG2sWSsPxhQ4We3hfdMO0I6kgDhdF9tWh3IxVUivLxC+JupdAPaCB+loM5P
HcjNjpl9zjNcyGSuD0gqMK+LgWAFi+VbYz/mchJR665V9m+orYlNrG6IuSjVCZ3Tg66VWebkmW6H
FartrcdsU/lxQE68gqNv96ysZCZcuMAdyYxKnKTHVNHmhpqo7lf0PPKFqv8Vd+9K1zD6JWuUkrMq
tiRE9rnEl8rqgCkZaICU7+oe8bO9BgpcXyLtn5t46tmStONoOOY0rkOSzvN2bNm6pwHt+vtab82S
RuVWDj4ZJvUyuihj/xFYAWdqaG/u8EU4JTNb7gOFaUHOEMQzkVxwCE0gF8DfxmOiTToSns2k1ghW
2eD8G/OSuuLot4SmycRX2c+ZSogSASQ9uOVW05nFQF4djpRkM8h3SMKNNjMFXY6hpKbnq4LhKDGO
CEziLTpvPHP+m8JQ7vgASkIUgS07MD3nZA24LjsEgQMdFvm9hCwjHvxFFCfdYKnZ8ZhRYRiZbTZM
+pOVglmVPRkV75ADCXY6ef1V0VdzcFVPs0OJ8aYX6HdepB0797j6DKqcmanD3gkiKPer3yqhNYd4
hyNGFPTE4ee3BJGEoa+YL8Ixa/JC1W8CrmjeRkjAfx6PAz87dU09tok5EKp5z323G/1gYwGzUMGK
kw9x5SuJU0ld/131YmEr+FXECcZqMZOMHZ1/30leOtiYPRAWfF1b9QN01mCDWAtoT7SLMjrZIb01
cYDRe1ymmrx8pd5oy3HWZnsb/ofhxj99TqUxQArS/hvq0zT0Tkpdigzgo+aKKWeQ4Y1L2NiEzw9N
HT2814FYIOTK0i7x9qmR4jbqX5ibPHRUIJnemvbcfvBAe/oWEfDW8LZx1w0ZHatzb7C77INf1Sjg
Hfrivs3RPRkaMOAGwkNvD46OY7/h6cRgP2IWFjw2nUwflwY467wHU5dvvLGdMlXPr5W/rbMHvlhR
g+LqcvgbTiiYFbnwJb9HSjII6ZF45jq6YKxjbkFyN5Fq2xrODm5kQ/9y0Ovrr6HEAv9dKJD5Tf5M
JfNIRtsFiDCcW/M/CttlXr8PFEeDDBuxS4GU+740fPTzDSTNX7+FmG4AJDORxoPj1DYN9E6aHUJx
QHbGIzNJO2gHobrkRLNp/cO9+BQmhZmhS+or/A7N5W0ti5Wko7i4qvuq3ZCmpnnkwC+yBcn5n54j
HZyDMwGh9RIpPPV5oWudiKgHAI61IJL2fwYS3j3J1iz0qkRXfNLUcak/BxTrhCQelOV/bBnc1X4n
mW0kvjNEDl3K49OdoBioScqA9Mq5TNSdNvKPusUVuSujHQZuuDGo3yxyAzriZYAScuztdZUcD/gH
4drcir4KJjuncZa1OGb7yogzwGngjJuIBlUCfYUD7Ec7J+3akJz4pfxa5WU2ZglkgPWGBzzXLw0y
5EObGApe5ZXFHKpt5Lavb7QFWs5tBDa+mSYEfNr2f3c3D49gyMQ21wzxCjg8H1PD4W55kGTUGAwU
qusJhqxEz4xqbnSYUUSQhA/7fCUdPEFe6haY7wsoI3dZLE3urUdh3wGy0JIbdJDJ3EXnPaTWzeYn
S8KFLWVS0ga80WycnUcPFHTBOONx7KDkmyW2QDLkL8rwkBhct0GgjFVqDGVSO8Qur1x0R+Iz160b
iLB2Vk4y2fRnttGR41zYrl3yGa+BqtGJBb1Z2MiTuJ7xJbexQm+r6gCukklnWrnOrbZrJ0eMB/fm
94sjB3qCq6tNaTotpEfuVl0Q8mb8SGjpL0XBS2E08n1hQ4QL5RG96StdfUsRKBBuYg4l7bo5yytt
5Z1y+yfSdzjQ5SkcNoEh1Gv4J8sRSA8nLjnvyWs6IvaiTxjY7ZVDZ06GelDry3p8ycRWc6TmdFho
Jilak6sOK7vDOgGaxhq13ciEXv8A8TevgwqrMlpPsVJB70fh8gHG3Pnr+pIKnT+URL25t4RnaQqg
cdINjZvQDA4b8Bod2aFxb6xSzmFawNu6xEsbpT9Y7L3D5HtVFx2+a7AQiwWBLeGbHSYYCZBwcNcY
gwtcDZ0z1KBSAB3PBpqnUw68RYOuI0qN9oIGwHuq2u9WTCzQta7A1FHXPcSJaBImyD6z9amZe8Ms
0PK6w0DJtwikoKuoaVKFbxQdd3Hj1AqLPilzbe6cFCj8HvGqpH8iYgljChEdGMnALBUhkL9iGNj5
aLubn4mhBSs0ay/y4qnaxhcY4oTpLDjt0hS1snbVza2kwfESsJeNjnYm0GG2QNOnHrrS853YsEQ/
15o7l/DwMeCOV3ZTHPm/2P3PlY//fHEkuLis9Y7P1ZhXvYd34LRPXZpJfKbhzyIGL5TmyTDLwJPx
Nb5SHDxVRZ3Ma4pIyxl3HWcxgXAdHIB4TFRMsEcGoej6xn7p0fKidSRY0ELjJQwPFyoxQ8fdoDDU
mq9zKMg2YIcyjwzHMMDby+mUAPqGiQ1/pEeqbBk3B6lXDwIBhSoIgBfDjPajQDEyRFPHrg+5DklX
DcVg7C1amEz6xTgj3g/3lSA3Q6xhQDLRvPQ6uY9NlXZuliwtZTJ9bOfIwR8tF3Nj2nshm4HQedAy
Wzhv7UHYre8vr9oqyUvZRL7nJGG20q8HNU5qursiwlksq/Tunmd66O+yxyTOSljGbomzhMshLqA3
L8bfHutoRkZetvBU2NMG4JkACDxSASksK5h9rxnHc7Y4zysga/foZfSy50TmaMB/haLezvNIDeqB
mspQaKbsVXqdo3u3wvfuSrmuTWqq6sTJgGhsSpzd45o+EaJxgttnq+lfEFV0qEVOGC3ftnsD/Uzo
WRGyp+5G5/dai88iiZrt8e0jrfXXify/PZ86SrHCasX13SvX+NawIKXWzZRM/pyVgUEC3WwnHEk6
pG5gqepZgwghSYor0g1UJUa64K6jD7+9akHKfj8gsbGfGbpX+GSb7DEyQS3cpY4CH0b2UlxfCvf7
XwBgmnyc0S7SaKZDwftR6nsJJFNJ9jVbUqRvf/6rdsoWVA6tYb6I52/Uc8E0We8q3PjbnauBFt82
AHaGkL7SWtddUkpkPrxejvdzm058cXD0Ce2SPLJz3nTO9j35H9kjb9tgqd7hm/bjbDlZ8dHIBnkC
VS7lnKj6dCVnk8YPiizWPulboAGhkCxEh1E9Eg5pYv1eKpoappDK9fVcUtfrGpufLJgZA81IKDWr
4yzk9VeMmXaJgrTiT9v+rHm3fhmCE4UZkVmsEWvL4Twa09OhyL6z1F7BelB8Y7q6p5oV0iRNFf6m
81QPSpkj0ERz+2ak1yDea4rJaHC3DBmu/ih9O2yAQRTW0lHQqh6uNllbI7fX7aOpavud50NwDoDo
YG1FK2PM6K4W0a5haBQupNm/q55Cs1b0OxUrfW/YFDSA1ndL/KIDKL3yyC+uHD3SK2URYf+zGxM4
mhuLdtgOyFVfzSH6zBkAEoQDpxcePnntvP2BqDx611poJhX18JUsiyMxjHi96BipFxL1XFuq3JqY
ZMdXpxboM8HDCMibDbweBLlNbYth8kDm/U/YXQbaniEev+JMarbYg5qeD0mHbB2wI+bvbLMHanaH
rIJcNFAEEjbWtbzX4GtwzgV8jJ6fBGVQcnVyepAVOiCON5XPS/uGUSkiKmO3/jdPM2wWurqu4PnC
DI2kroLXTUX4Uhg3daFeuDsQ87Y8vVgbiBezxu2SXDkR7pvcpbTmHEswWngm3FvLbrYRLF3JCYVe
GD7+Z7GWRK8rErehviMHmgaVHCmVI9Ivd+t+THhbxRB1rh/GgjdkatLcgSqYtZPorq5TGPrpt1x6
SXybC5q0h6dmXU636IlAsRHgnKESjEn1qI263K9o7HbqiKUHK1B1j4rkAE1e6GmT9QvACI88Z3ig
bZOq+remgduxCWMUlsz8rtjYDDrHZjtgN5m7AOIV9CxnYcalPSM+MLlQyfrZP8H834G6aaVREAE+
9F0DOvamjMyKJB5STZ+Vp3xT9IoWNMqp6haw7KJC3EDuKWqKhfmdKz9ENXx22VJO9A2s8Go2JLM0
U8GdcbFHCuAQyhRxvr00ibQjxY4Tgb2ETmFQT1pX7tT9NiU3u5BrpDrYCfEz49NiWwWsM4cknp55
PyRCf+kwfzpDP+zxSxFh3VD/d/AZscU/Nox9ymThk4d8Dgps7cPYObPQuNkfLPqKjTkFtVilA9mg
qt1UvPPXsRcC8/6J63sr0v7Srj5UKgLEwdpTuvuFXcGlvSUlc/eVJhDVP7fhj0PoKyyL80sUjMqc
rBHFbOOI2H/ZyepbPjNsK9iObLRxnsAU8X1hHZ+kLr4vKg8f6JjkLTaXij6ELaBah/qgQ8FXbRbY
jPQOQC3DWJUOU7GVtwu48PqKA9QuajWisAux9E9k+WCe7kmZO3kg4s7D1Z15KXL4XJ65LXaO1CiJ
pIHQhnNZY0hkMLeyv/BZkvEXUksZVldOxssAJ4JQUEZaxrm0NrQ3naymQa8CA5G6MJPn+7qTxkDu
DLyDC4BnFiYCXk6DdgCz6iWzuDGd72cvnj6/BeyVYK8DJKuy2Hhbi60jqigg1A7uvbWmtAuHi3Vg
yI/RhDfbWWk3n5WdX4aHzR1K7H2kybElvYVRIyrZsQrqaSvWrbReTY7OxJc5LerUTGqUTmZ1LnYw
ofEcBytkTdpQIm66siJV6OuiOu5fVVkcPbJvwmJ79LwrWzGPh1V1P8lrQh45e6/7qkRjkh9i6ZX+
Wka3gF8wfl2Exr28xC/0HpDdVASxqHcEBWipbQRgGCH892kITfKGzVbEkE85lQEdWPCmmUmIa0VF
o/9ZvR+94xjXMXcb47XNwZvEMPY4D8Tk0q7Px2BDveAtvwqNgGnJ9t1pKF/HamOcqSZszWE+0bQ6
kyAFx4o9fFa3UwYZpNWjkYJY94rhO/D8zePFIYD9ZODvbBRUEUX4BKH4l9YEbT76B6OJ+HsB4Hj5
H4wtbAMRzyLhCJxxNKBTBY9tVZvrBpHmpSYc0Ezc0wSGnUv2tWcX4miGDP+oLjHPUboOQI4x9XxY
A4k1R53GVxPHBp1yJ8RUQsUmThhhLlv7RfMm9Zh+Qzi+K4U1pmdSbkI25nte+I5CnVuQVfpKt9YV
FlGz32p6QeD+86a5CYsmrWW5wyJ+mSewZL309k8zDaQrTLZZJnvFaZCOJP0qyuGKY72Nkjqr7/32
ZkwQrIYP6qa4TPPkRG2lLGxa83EFNVogDnblNgUjK/g9yUGZ2ZcId/J2zU3esiizd5VqJKRjrNhO
wK9Z5KwWI+SyQ9GmvLFlKxZF/aPDqyt+36e2u9EDe0KjzOftzrTr8YmKptn/2v2OZJVtxT+xMkJh
4VWnfEMTFSW/fUAyDH2vNwbpHi97Lhc25JD4BntPeyUH4MtQKeIGchXFVNeJBpP/cTvHROh8G38X
C5wua8yl2BAvQU42dWUDZYg1Q8Smgmx6dM9VPH1kAiovX8F86mv7vt0KdpbILei1PTUWYQX0pKXG
k4phnS/ydNJqVFSjqcWawGUIpxvno5no8KN12Io94XhCEmrPaggCJcH07oUOHz+TRZM7NHsuQqfx
o0cMPSZOFX/P7t21zeYcAty02cXpHci9uehf/ncZ/B72V8q66iltySYhMNHAhreq6xPh4Sehjc95
gKFlceW2DcWjMAUb2VURoZTs4tztr2FqyV8ne+m6C4XhXmSH67GppODbY9jfmEJb00qY0YLicgjQ
JzCJMqT5QjLDQNHJooK2QA0ux8cKX+HJGVNdJV7Px1b5UUwHB9fkPYJ4EW/CIwisbpyclXRwu+bH
bT+szAkzH7XGqdpwl6UmWx3eny/fC7FdSLJ3GvazvDnW1bR32mhfDuAcia+lv87HK/Eq8ZGHDO1r
JjCDN/v4PNniOHD/ZglwpPFrXrsZVdF7aiOWXuZaWfTvl4Ptx0fXweyXddZJd67KCgs6fq68VF3m
tAYFtwHeItsbqERSQDwMC/BIlHNk7pQJfp2zm70Irve+e7Qt+Vv8l3522Q6tVks6rq+okMtPEtfu
nCI3lcih78MnKK1Ub109TllGWc/G0xWGLDNyuPA9ollgo+1b4fun7pRkKcgv9VhYGl7u9XdbxNtu
49XAoitr5lnjTJTbbEfMXLtR6iK/ULuZ18b/kFhAl14gFlPRQutt4IsZljMIlCzDakQzVG84mnNe
019e9OwYRRsX5Sr+/zVinTRPDhNnx39pEbomj2k3F3gZ6hP+0l4uciJP002IwzierwR0BuSrP9bZ
WohjDAc3lBHaf9Vu5I2PfYnP+8eYgsoVwUvc+HzTvFv+WUuGifnEl1wROVjTb6J3kzCqiekoDjxH
8VdM7RY6s+bXkcWVCvdUrVugfugzT9eEuahl3u2fNhQrOz1dFVcJlYO3kVaNt/7oNvlxSvHCYYwA
YaSiZk7ZD9itRllkXsMfXj2Ye299XcJpNStqPXkPHwsSpPV8Zxye1isrSHbQ7Plt4PAIauXYBvd1
+2JR0aUZyFAy/PNSMUqoSYEI6VSNo1E4sckINPxU5Eh85MQ4D4PYQvkayA8f/amYWS0KjCtL70mP
snz0vMRETM7fZuaakRohhvlQVdruOZHr72iy3lTW1lYhwk9W25eMNW4YgW1/7DhaHQhkqJ+rAaEo
F8zeOLU6DAAaoNqXW1DjpyDdxnry3jVWCy5WF6GTgrG0UXpOGotzhSnaMQkBGc/LkYYTYfw4+jXq
CzJ6kVLyG9nrj8H0X2KaCtWzSZhUgjTvMTxKUmDAtVWSHonp53oMdoFvMyZnKcBHWKr9oEJJ2O5W
EAkU41HyvjqSj/YC0aVipBhdiOnvp7IQ659DgATzS6Tlr+AH3v5mnHOS4+pArm5NXG0qHI6AaAxG
oQR0Mgi3UxWmuQWhBUG1uPBnOM21VwXJINXmXHkz/PMwI7AnrVqzo2rcY/goCEhSPBTohThy+tau
FSaeUK9a2vbSRQJ4m2ML/arGmVWmxmDT+8ZhBbyyj31gEKyENFDc8Pm4oMsIQtGEIuxbmp/5ZIMW
hcEHbn/Tv34zMHetkTJJCnDqfCVxfRMokxbiPUzikHSwkveZPGO8wP0uuclFeTf13UeaAlqdk5oT
VAgeN0H2NnAlKKyrMOc2UmmtgqvA4F7YImrHio+Mu0KKs+SFSiz1fvQR8nDoAqTdkU/hPH0nd8Vh
STtKXZAwpLEgAOq8WQ8kq80ie6iftEyymjrekU9h8NaHCMmqiV897uoGwwE6QjaW9kOD91c19tSo
ZeT5sTmLXId5dE+CnL0bckXM0dxyR9pWHMPTOKmlyyXhwkznBXccDV7BuzZXjZ302oqdXSCdHHiJ
H1ESJBSflJDuPMMRL2UFgtIxQshvyxicZAa9MPRQhmlRW8U9QWZLW9fNWOHmljYYQ05aJw5hV1Pw
FYIHR8miE4NRr1sWFCiXm/ek+cuse7xkhf7T2Puujn6iO4Tiiq6xL3xOm1dBMybmMrKAg7m8EJMf
mBG9omeW8mfg+EMlRz8y3hxCIgJCHwzGQLc0W3XrRBHGFhTdnh5YtySx8jxedJPPdllMQZXpg6iQ
qIWgDsdhKHw2ZLsHPjFOytcJyMKEnbHu3IGA2Mvgh+73WsgoT2QCyK9g7dokUTpqWhpTiq5Et2TC
fvdhb84xH40HE7cAgMKAe32ZC1CxtYLMu2AkY3AXWLZIT4GfXsE/YgvKdlRHNgOr0iNz7Tuwfe6T
7uihFTsQA9w+Retib0lyHd/HWaMSdMUMEupmKmlre979Ilw08ngadAi+Ok/Ft8tzajHKEcczvSsm
FRHB1JYBvuGwW1+zxuy2zjw9GmKSJqZhXZGwI2n47FS3NrKsLg4BZ5rkMzWe8iC7cJ0vcIhtI6h4
EIrhPN+si9/CwDvlMxm6mwDABqZ/bkB5ofR7xmDirQRl3YcQ3Jkfa93x3eRvMUQN5mzM0DIR29tv
ZiCjYKN7KRIdk/orcB3n/R0pzhR4yeV2DItA4ygd/3vENsCzP499V01VT/pRRedEYGy68LEm+4qP
EkXSPUsmG9yzCK33GG5uediKh/o5QLCUiFFrC2Aklm5fYP6UO9oRnpMwv99Vza9DCgOoWsxqhuvF
tIjg7owhwfofnThy0cHuKIUdH3SeHDNAxUKdC+bCPgO/ibveeP7q0Uclx5hSZD/tjXIel6oJ0+l9
2gFc3BgQfoAH//w0ApyEL+QcjKuPja19VI9zaLsAT3sUJ2AuSWCVpkzfP6UhJrmaaV3945q8DM8P
VCbrCuCe6/Lh8rNWiWAavJa+2u0Blen3YDuJN6jYeexrYUrX36oPDsrCgKeMj8DSgsEfQPr+Pcq/
yUlWR4E5NsffanANZrbfvb7LDi8jEPruLY6ENC9Mj5b/ZqL0nMHpI83v3tQyoebaLqSg9UuT1dHu
yUrb/4CmAWgEPIo2Br78nycj35BOmu7CHdh7+n+HEAychYcP4ea8Z9BpptqgD0EP3k+T36tOcxEa
pvJGMK2dKBtPd+5b913yx6G9htELw91jgFH5yE77yduhvQgEbLmDbgY+tvDho3maMrNFYABBdYGE
TZAnK0IGBSZmR/4qj489xjaG+HkP3fSQtiHAjXwz/YE9QbbsGLU6tzNNYaZtJF/odU3EkqfsDIOj
15Y7Xc7xIxgWb1gvsb6+vfcsR+plxgrVpxUj3Zw1ckRwC4awfZnMuEpaSbEz7CsH2Jkt6Yk2gqUO
3aho9ZS/bfp5jHADXulAF5DDgNNfosi9xF5NuVhtShRjLgc9qo96l7YXQpnBoiNnC3beoAjwewVZ
2NOH8vSz/nEdlku2/kpPn5zcU3NuXTXEveIJ425s7ESNFTtQLFjo+0wMNk0jjp2H5BlWF5lRHe+c
OoudqT29pgzv04DIZ9xIsm9VNX3B/Hg/rFV1QqrIFF66Fx6T3h/f1L9L/kuXNgfqCevO6FEt0uOw
3MDUVXSiBi/C6YZ2Euxas9yAtjEslGewUxVgw+WvEq7RbALc/sVnrGTlyNc/JWoaBsgYYMcHUBRo
xJHuehmtlgtqXAaRWDnVdhEushzAMZlzEPF63kBV0MvJtOsR+rBxlCm+mgOJPSvlKBIMieiJB6Eq
D/ZQSRc5azKWg+Za0346s9UEjn9oNqPcW8CnsPHnnRYNp2fRgbDcVs1Q2lMTaJHmAd16DAAY0XEx
Z+3tTLmMuXyOyvwEp0kl0gGgoYVrO9/8HbNSQkxr11c1pQVcM93Fj+JPKsg7JDXlvXRN6BMnoPfR
yF/muW0hCL3VLSWqNcv0g5jw8W7oOhzdGKJHLXPf6b/B3OLpsflU5/Qg4KRETomQvIPAAaxsjf1O
lo58Tx0Dv/iKih/NRrx8htpFYFoq3Wo4z4QggcTc0qAbRLJJl9yKUCSyLEIkul7mYVgKBfer3NmF
20rqXgzOyl0dtjKyIPIrvf2tCfDwbiR7nLnjkH2vHpqAu5E+0R9+AGBavIxqDRqEQU8TazfDH/uH
UqFHRPcF+IDG1j/0iIN8p+42nKsfEy/QRNDJCXDdg79+BwbjVjQP4TfMPFrua6xCQjBFFpNBaVUn
C6eoDxFwO2BEoCECUzHXnSm+wEMyXw8qr8e7oRRtSkM2G5vqP2fwzuzv4KGbeAx+Km+/mFlI80j/
MssbwNeUSu26MixBGta3q6qm5eh1Wp8OsJRTioaKA8i/nsqMODfpyizoBkowikRLgQo+3X9DL2mM
SRPli+Ntnzh+fY/yXjqZEq/2swcb+k64HQMK0qGUD3Qn/UGVQIG6/vMJme1Doc8Jobhfau62Yv0Q
n6oUKBX9mKNn2cybcZuoU4H95J0krj8LitYCaty8mGkN8pwLeLYK5NZqbUVg7iuiSKckH4HjrcBi
dkxD/NKS+ulKyVK0k6fxd407lN+Pz2qF+3XL1yfOHU+rGP4bmqMqQe1Hm98TAE84x8/CW+3xkfcG
mjfQod/GVaR9JoZeQHl11+vITP65FazzpcOmCICbf0dpZImn0nVQuAuae2KAhIC4ivOxWkPIBSkv
M5pzBLTolz2GN/IG9ZxTlK8EJ4OnO5xcNLtX4FyHj5vGsgJc92Tub5DWUWvK4GWb3aBDjFaSfkGZ
m4chD8DIVpKu4fBYBWhtqpphAsBQdTujpua8ftrdCYxGQKarAaT3MKwucz6W14BqlAOoiaasOxHI
4FE9Jm32DTfpg0s8pOCirnHGmtn6PTk30TDRA6U1jbL1DQzQzz+EBZtX02dYTXuqP7gzz5WlOMhF
z6YikYlb86CmQZID9SdZOkuMK+hDclW8DHSCQWR/G2mLG3NJMU/tRzknVwfFaV8s8B0sHrtumwck
9rh/U8E0+cv7ENqaWbUBiob+qw2X8vbXrVxv1fzZh1NXvmclTGv+lztqT5/LobA8R96fDr7Zx2w7
4p7T22ozSVFh8ebKuXt3Sb0KB+lpmJP+sH7C2QmJfeGOwBysDYfSqgAo0vx5+j8YFAb3QEHONULD
yZWcsETajN9X6eX+xJfS0qfIXeH7AbcffYsnyBFtew/AOGl1uY8y4Nn20EQIZF8vaQLsVGrTUglR
77zZ2Yyi9qoLgCKS1yICQCswN/bQg0+s9xmpbX+O7vW/sWevuyqqEfK/ioaEIplKKqAqDT+gxdvL
keJUVBqAuOhSFEFulVU6DN+62jBQ+dwud/KVLj/WA87TTMWmKd/I4GpBgznhuD62TWxgQ0stwWdn
p89tG2xOXLvJIqVKa+/iAA0YES777lBq6p8rIwRs6y+e+SrN/Usrn4fdAJK1+iwd0cRXyG2k3E+w
oDJHvnOVEOmxFELOtKczc62rUtse1J80g/4oP+DJ6Txe9Wieb8LC5dJin0/SvkaifPjMSw4RJZrj
SJi3EdP1d//0l8zC12/V2nTTPAs5CzhzABX6GMgqINocOWp1jUPMNbTy+XDtmV6KkIa885I8T7um
JFzIXE8t+mm/Rnu6IUSkmC+H6iiaw9aU0FSZY57GurLJvWXrX0whd4Ciww6ZITcLuNo9yPCZSXmX
Ph3WlA7DvIj985qqdmp8PthzrsdXUDXL2UOAsHRRqLl//2i4zY9AMx7UzZj1vcmF2afCL57NLHqK
jksiigIecFRAMuX7++ldjch4td8ZAJhgRIwnYh6M1JBOTeiEc9GGVAxocVzB5S1KK1NOn3FSAr4k
Zf1mtxr0T/iteesjPLDt5PmykVVdidiHDho6T7Bxt1R9V2nom8ZGTvwMQBrQoCqtWoa+fwnFVs/a
ZH7oPHkmfvmmqATnjeESD13/cct2YCHqNl5EdsSRq2gcpirq/48vdUEXS88jfzbxOOmJuRkONXke
6zk6S+l7oj1ja36wG+FPzstrbllR8iu7czRSxeLcx0e67En+fgRIoJiX6is4bFC2aJ7NjluZ8FIk
NTzH3rchPsIcCl4QNcCkv6cMO/qqjCWl2CiCLdDNxkX/vVt3Qphagy9MbDg27hWMxOCBNZWLBV70
Y6LxiyWt5fih6vNwfzhQ43QNRmEyO7mDWulWsmbmfp+Oa3aYaafebishhbbQWCkBf9pNgCNRWcKL
kXQ6ZWyYfie7FwcrvEw+SWShR6KCDjzPeBA9guvo/VQpvTs0EHGoXRYXnETKxDTIQWADWWYTQcxB
QiLOxPK9EUmWceceGKLKAE4ZTgIBWm8JYAashuyPfrkWNNdia8wIQsgH9xJ9oLiGHxL4FoTckz4G
hNoHRi/aICpLys8oKMNIIFEWERpgzkdBcD0wS+mS9h7LZRwqmvg7WetzEuGbe+LeRjX5ef3gysnz
Ky60vT0lOjpLbb8asuvHyqnNqLA6Vi4nk2J3ZUNt/+Z/24fy0UwLzEWeZHzYIadfPGBYGZt6SBbF
sQUSAEEYawPu+wws+8w2TQ6EuGVDVE+B71vLj92bzjQoM5jIz8N+/7Qesv11/A5wc/b0Sg9Ywnv7
vy5oPjiKwL39E6bTqxCEJ+NSIxwC/q6XvA2hHmSNxw50LOo15G3WnJbWChgPtnxwNgSyYqi5uQ6P
lWiUpOXQNIDtmpXpKP5jDoPWrtuuwnrVEzA7r4nE6ZngjN1mTUvv4RhxeNdlgr6OgnS1ceweXXaH
XVTJqECD9iVfVP16gkvCBOoOzmHOntIjgxLYoRTQ+inq/MkbVcsA57Fs1c7QnlFiRhfsFzTZQF6B
AmdtwO8KlU8bv3lP63mG8Jm8qYzBvwS6IwyDd2scLGjRYNCxO/2SAyutiz3mCn9uhVrz2k+0XRSA
I19dZsrMHu1iuKA87xTiPpJmMzTYqsWeGMQY4XUon5hhMHWv1prmGb20/XBxRNrc09WPxPjTpvLK
KqThA2uwUEv1axKkG0VLB3J29gS7MTruRs0RZ/3ZqNcaLx6d/hGpAFgItJ5mcMi0z++GKBXvQtGL
ChVTPKeG4PH1Gjy6mW7EwGpOnZjwlO1ZpBcq75lHvJ0Mi49Fz1Fyhbb3k25iWdHn+6bydiUlE8cW
6n4eQrd7BY1y2XslpsyG3PBeABbueBGNf7cR7FV2gCt7eLDObrjfP5afC+Q7VmWROLcBL6nfIlko
5LlAar1rw+0s75ob0YcUWbdIl0QZUetldpgRsofDISOIh/Byn3PD+RI9HJrcKMIbp/waZVTt3kAf
y5zl0tFrn4sya8G2z+jA1fdSI4lU9piDJ8jl6hULEIbJTnLz+U8IqFIrPLiXofJJA9XGT4eQ0mZ5
bqewc9ABeW+n5jWyDoz0bZ1I7s1LBQM9tTqg2EnwzIW9n1jAmdtcioV8YTRIJW2NJc7W62/MH2St
tmSzJrhqocryh5GJmEa5K3nHDiaiPAoHXGP/5v7uhqiJAGECV0Dt8+VK9ynkJRScK41bXFuG8ccJ
AOcjPwEOKpgmb5i8j8CLxAvkp7Spi1cs9D5s9LNLoEcLc1BDfbediJa5MQQmtv2i2B2bq+CkwBht
zKeTlPpxCRuvzxAbpGLlcbsI81tZPJAVxRyB1Z1onShZzc5gi4MTJTZgf+XC+gWhvVkPgy5Mi23R
yzca0DQ/O/t2rjo1RsxtTIz14Dd9yw8zzHav847rTK6bclSGPrZl57XPFRW+3/Ti4PawyeWWPRQ7
rkreRf/xP77Vhfw9s7eB8T35/oam80gjDAWt7umNnjfIAfLHF0dCktPsl/sXKL/5+N7b6VlLNXya
9YFx2D7g5kfVq+DpZw0+oQKy4Mri+EqYFlpOmXxbm+Z7DVUSEKB5Y3wEexdP9qojxrP8pfH2AqKL
CmdjwzOT1lcRnaRK1scvvGdI0OVl2sG/4Kjqb52Kt9xZx7Nf4TnXt/EGFKGMVXGquc4EibrDSNXR
6ufu7O6bOMkR/CW6DR4xpv23yds6gH9zsRJXyohhyGDOvwO/3PyEDf8RPR17le9wv9t5ib6Vz42i
TZ+JtgAeecEekbnAQywOdxHTfkVkqTWRbkYg3eu/VICQDiWfNL5b7nCnW4ByjyV2EAyPoNSzZB5B
6rVjxO+kyV4uoIHtxonBzm8jXxY0b4PrVl4CaoZmyv3KcmiTwU5dAMuBDe+G58OxCzqspGkmzysu
TL7ogNvYCmCTxslAe55rMVyaz1VF5/Zu3W+09Kj0hHOmYT9nll0n0g7FbwnKUwHp/Vbh6XcSR1Gv
FQ96UAcplcdKlIjwxWm2Ry330pF6Z7Bxvu4aaJD7IJNVd7y58tgm3I4LE2ya1+f8Ofzao0mEH0iS
sqF4bkDOZiQoiJkBezD7Arkbch5HUlW28EDnmEhWHPiaqaKFPpmGg1eNf0dn87uYsZI4ljKOLjn5
zDzoBLJrrSXpRzRW3pmWvO+AagDmx38TxFi+WscsCfG5Bs7i6DlytaYyOpthdQMN9Q2x3X8CtJYu
a48x7Vd//jrn5ARa2SryOPrDTvaKRARTZercLtyg5nsoizWEY5oLw93fnUZcmZtXJEImATTAdxC8
t7S0wnkkEqzOR8vG22y9kluoSvknHxe2Wu1cgD+aqRjSK/oATOQ5ztRsCSjyso4fW5w/UNeBjlEk
iifgx38PtLB9znR5XuJbyHkJZ1+PqU2GS7iRRxG9NCVL0XJbyI+JkWXei3+tc+9Vjfobvl4Q/n3x
0FV8XC11V8KzIoAA76HD85DTv3BKyuFUsr28/awoTljCndA+OdqDhvee8EkvJlXWdd00DFEckHeY
oUh4yNh2r+6AfkvKEtJE7Rp1/p0hstnTFPQUaAclWPsMFYZsX5Y/ZxjbKYtqRSFPKkaGMwTRR1dM
I6qmgEU9zyVBvHUzudAGd+kZa86vvpOcTljTaBgG7jaBQwUkF3hIeoLe+90DFzzctuIwQVGC9U1j
Pgjb8PQ9PpTeBHIk7SZugbM0DEBu9rzAjBUrLFKmIWvVUB+HpwMdoa86dIBzMj2w+Hj3TkxGXbPA
1fvTu0lDYCkTTTpoy2JIo4sDybTIokpFqWhjiIdAC0iwlOKIkQFtIsaT576l8+k89l9m469j7VIQ
BUDhRkCr4Yhqh+UzGxqGddF96VqpfsSyD4JQb6rTK/88MKjJyIWtj1H7Dd/L9j6Twowjk5oJ22Je
+rVgMvvahGhhluzUtEuBWGJX4dMjxAMuPaLTMwtcNP8C1xY3yg/7Ww8AOOeXPbrDVNpbRMvZuIoC
aX8TAtAP2Pv5ii3VjzUJP88WGv/SrJpc17cDBb4b1I+rbolMxPH48h+CRP8K22Rb6PBpvtyy3KkM
hH0yWLrBo+GyPjwO4nyJRZmc56wldJ1C6belkZ6F95ZwCxQfXOn+ryGPvUAY/uIgC/7lMq3SaX4Y
O2Aj1JXj5T2xR5It4HXaF+FfI6JtLD644YAMQx5dYbkUg9EUwNbOnnW6JUvXD6qcHbPEYvFsn0yp
e88QSZOj7QOAit+uHEquomUsnK9a3vjc4+YXv2dWiHiZZ7I8tD22RLj4P5kA9a5yZP6pHyK940O+
a4Eg/KW+ORpU1zyaR1yCo6J1NV+XWkwNn9C7A7DCklOkuwcSsh0rfmsvBKMl6+7smcwHDA+nIu/U
WIWvTqxjjls81bjRkcQmF+vj4xZUGTXgcWjunNGCMJIcXt49rU81gr4VKJr1jEVVns19ZGoAeVE9
FGPwbaSsTacNMnsczioIxRqBpYsKyUXpw2FetxRWMU+eIpIhWgrbPrU5lCZ90hvmYgZs3DqF7bKb
g4vS0IqGYaGLOpPet3L4ldAXsZNRYpVINjUS/TqF5dBT4IOOlSwWxKtQJ0ERKhwbdXeWW2LaltA0
+wGMBimJUc+IR6C9X036OaHwpXGiNh/C3+NtGsN6oiDYlrzi8CHXT5DYGoMFos7zdPN2hi/gUSGV
nCCzFnHFF9RqOoRs7RHAIEvZk48xYEpx2sn3YDhtqVKT9gEEhtYgNvx5PRIGz6DVxAxhuZbjTkaw
2QKM3AR3V/n3NbpHoRgbFshHHQOECvS+K6Hcb8+6jh1SxMwXMTbrFjK8JYRIMRtLyWIS9JH/0fMm
zWMdnRPBoVws19vO6UKZhJ+Q4iSvqwMCe1SkvjpsZpqLeaJfcDR1lXfGoPl8+5/TVuB4qXcrcoO3
vm5w78LwDNkn7Vrf1TBnrQanXq2mFKrPLTt2uhyD4Su7ehQcjbae6lLhFwqb7T5jYLPYtdqTZdIn
h1UrQa4XJ+6NARPl6kNYy5+Bnho77/eNK9njRrEKxg7pnMy0FIyOlJcaG1c3a4UQWv6crMxslzzb
KeCSobxuF2mzc0NM0upXali119trpaMJI018z/jTTjps7Fhv4CqbI3JtFVSkEuAON+xgQTqS5Hal
bR2UTiJaDOVM2nnKwCKVDsVZrodgBf3cVFgT4ZLc/wBneN3y9amdnC9XEalSGtKhbVzxuMLKs+1F
xlHUZsCHcSAIF7+GdDpOkyYfCBf/Czuwkos4MK2ynb0ko3TwgLtCraRywhH13f2DyprtzVQttgdR
FsTWBY+sgGFoJpw5pszdZ7E/uQmgNLAvllGrRrGM/PTZFx2bCpnnaNfGIrVm2ZU7GwC/HPGteLHC
YxgWY2MJKj4Dh2mj3zzpab68z39X41grl2sL42jRzrBF8RLiz9CZuo4uW66/qb61Fsh4N8I+iWhS
A0Mr+g89vyUx3n+LUzCkulSHQHW2LhHGXOwR1qhX7wI+C5GbxUQk6G/nXzC7l8+WcnzWeA7FrNtZ
dtcE5+eAEVourge+gHCCKO6UJocS9LBWCQ0U2OysazuvFs5MHyBcMBvCM6k+gjhlmp+25UYy1/27
XpKR5JjFUOM2HLkK31rv/X9xgQnI4p670044kCNFMMZ6TfFCCTvD04pYZdZf/20ghbPxgzbPCz8b
TWDbVszzWyvkHTZsZbuC7NadaGQdtzpk+XKGSWiggEONyDkriG81q7VjUBi8FisKk6VPqZ+TpwA1
BsUkROS8yagmKIO9+Eh5EmjNcvB/+T7WYAoVlinZcbr1JyoDCREitzZTlcW4sEcRL4dUlXl5baHP
c8jIg7q5A3ggp5Vf5CPjJZbQ7X6tAN3RA1qGGTUjLLqnsLFwQqKiusrKEbGl50IKqKZVhhzK7EPK
/rnR2nG8aJwtTSAEBjGnDLDU2Ws2Vp5O3O+z6vsb0awQDvOv5++ERonFeayTAo2c7XFc5K+dYcoG
PA9PfQbUme0Al17wj6vt8nI8kQZo5XNdADh0QM0Kt4UsQFtpfSw9ASlfKs35KVbRGVsR1sZZIb3N
sDdVrZ0OC2oiD6lnNlEfhN9Vz0M5t50+rLKsIQCp/PCSpAHv2K5X+0IIwOhL2ApNhweGgY8iYdmh
RqTkegkO4z/4UJfzBpyI1hpzbMf9OolFwUIyWTiExB97N2gLFBsWsqzcDT659/sqvhTr8GApYnRd
EnMi2xZb5cOPdW6cfxiaZRhFgviZagZe/Kfjr3jRMTUxFRXSiARHIOxiWGA712QCkyTNX6WshYEQ
eGPS76tSrH9zjbOnaDiS+FH++hIHyAcvHPoiX8p/fNqUxosipCw++gHyKLOfgOvFV+gAgcX43Ek3
SXYxZvYCBSXqdK9u7U/OV728QuFvu25hU+HujSZSZeJF8VoESzt6UqXk32ABXG6JRgxqTqInBKlN
+JLnWZNMxApQeIxeiYi7CcMfmphzs1IMrfIROktAzSSXQeHmv+nZ9jL8eh1nkDmKfkksjfSwtLdG
/lAQ6I9cUA/4CHU326/Qx6NvBmzevV/LQnerGsP9R9pU/19FFjCK+9hHZHbPcjMv7DIUZnBK2a8t
x4mDYjMSOBDCnQYgZbs/XkxTT/CRDNuVaM/nMx8jq2WPhvjkJL3zdrBVu/ct5rkkGotId/bdQzf8
zADusqJnYDJD7IPRJSU2EivIc28nTmagZ3HBYAE4jO4S3GyZ9NKbEtvllYb88rBTktWh3YfuOCef
9NNHYxBYhpfMsgwEjn/B6ZHPme0MTpr+ZaNjcdWdYWW7fJTS0M3vMouMvm8lwjewytvHjuH3lWwd
aQFWLaFUo/X59agHaMlu1wSeoLeXzARd9ovl2bjg/LMUteqS0jTeSeqwQfaUGb4gt2Iw5kEoZPN3
TdsBY7JrV4K5SBZAn9ONosCFS74fz8B63ar2dhdWM6rP/0PeHVLJkOItHbR8L+dT9NK3Xwp71/kL
FzHmjBDiJ67JnI9lzIXBvtDTvEVvjwUeFLoehTjBlOiHn+sCzC7F8EeXuVE1bVWmUD5bDid2QYmj
KkJQrNIOIYcC3RdmPWkxFQkdCWuMxxWLGSBf2/4dOLyiaFHzZ6kzX3p3ns2l08TO06xOuKQPy1ca
JEtyJ0lfuv+Sq0HRjTqbrDBE61E8mrwEKjc2iFv97P4NM8iMKwq4HzzQwre3g0EJyqu2wPASztZf
KixrH9hYL9lIFRXlQDd4P53n6EgHAajS/MqoEkC08W3KjfO4e9+iSdss1LtMyFT01jdPdhhXTpmI
t5rmaHHlDvv3um3oqWW71EaNREfbAshkGxXnJSeIVRYUjZMPoWcseggD3jCumWILxadlBWTRfgrS
Aeh+VSt6fef+xyAnCR9BNxwhj2NVVA3tF3dJAa3rua1Zox7Yy/43gQeBuYWMiaGw83p+tsiJfCKH
CMtGYYeAsYkiY2ZmvSxgrg4HAENBuwqtonj41iHrwoe9120iO8LQu4+t0iNtW5hXvsUhpV32YNyn
DZQfWRUXfrjmeGapP8uz7X7AlVcw2qYNjxXvanBwb/dpZE7W1+FGJUVv6Zgz9w30FEwLH8rl9JDM
vyyAzIxYq98yDmjistEgbmaLHMvIndm14EWqbnGnm1CYtmQjgqJNcnj+MLuexOlsrhhv79haArhL
wqHKZ5CkGbcaGlg5a1eElNYj151ugx+nU+2E1zoemhR+5Y20t/VsSh8gRFTg0DG/o6RzE8dUoe5F
sz4gjLumWpC9uNwchtI3qup4S9Wk0BMNEI0ybleLW2lekPc3q2CYiU23jgszB0b/eDE4fX5Pt7jD
KizGSGg/Ah73/IDOIHIEIobow4XBy2O4plIERJHO3vNdTjEI7Xkxb27J5BHPdZ/qwYo7yx5sGNqN
jwBNEnCkh3G0Y7wNmVbokn2s9TbZeM8XcAVmsT0jSO+FPwTFMCFkPmjTZPPgup05zvU5lr9TE2M2
h8QKm8lOUl6vgYw/MxnH4CwwPdTLIHhvXTtCdpXTMgswZ2upPyzX3kHIoQT8XrLB0a6bI6khg2GK
0xF4dXGwHfjlt/1v1JmiNvIV+sybblXo2uEXI54tpfyaRnSXf6jpS8sD8iniWG35TWlWKWq5booG
WYKKxxO6yrcfhfSSZtnd3WIKWE12SUU9llrqaYVMaySmncK3qc3ei714rbRa5dAtKBTZ6jGvSD1J
ERwM8HjOle36DJ4pNkBb8iVQU6OMYfhX5ZQDjyfjDeCdGus3lg3x8etIgEJaj1w7aCD4s1HjQkc4
sjR+UM95uloLLKv+O+s0jM+5rWuvJaWEinj41Oz3ORqJiNQd/ffh3poJZ9FLisuTVzAJFEbAPYwW
+kAMXlhKwq9vdCN1tuU2SPKCHUuB94XIN/uQ+EpkzLTTp9e6BjcU29KDxyuI56I3539sG62Zoaa2
beHUgGOQfdAPD2TLKAjE40jfLEdEvcYDu73akfXcPjt32QZm5WeyBhMIrrGsXyA/gbCE2mueH8CU
oKBGOsLdf3BV48OilEVdxIFFFeakJJPI9w2Sw+Qe94quPwNAUWFkCH0ceuUkUekdyfRLi6Ofdzmt
Oz2WIfBfYiBbQoNlJ3GxjwUWDB/lzErrF0EGRKXCISKc30PVUH5vIA+DDb+afzEk6w1116IOnFVK
ba/fIidxE1ePX2F5Q8cwkh4uxH+2Sjxv8eH1SdHynXrOzrEFYp6Kq2gT33xr0nNp/KVbXy3XUj04
Qh+Iz1oDh/iU6SeZhcKZGDzatL7NuSCa3n0J0ejfkBkAFz/1JcKI3waoDasiwF0jtiJEZr3ipHBV
zjxoxBFLzGRcak9BfSQuygoLS7mcV0orEVp+VS5RJGyA8ysI6j7XWkYtEUiRVdyqJ1S5mxREczwB
6aXWqx3204qJTBDWazenpyhHtpxvCKgvFne+xZBYfvqahfa+aTNnNTSwgDc4o0xZ5sp11TFtrhms
FYryj3HGzVT1CvvmdZyY+ypRerOrOHG4vo/mCO7pc+Ix2FJvpEeEmueh2CVUpQJRktQPAWEp5HvT
B5aZjIGzcupm2Pabkv8K37jhZUdTySaW2Fdxensd3444LTv6Pw8PXluNgqE0doLKqSsFy5m/Odax
ZgTzFQJLy0td5GXP51O+WTTgQOApNhY1PpOQNUGfo/lxF9FzYSbeYnW78kaGbDjFi7XSQC7oxt+L
4kDG40jbhX4t7P6JV4b1loX2jyfCd2cltXfVM1upnhqJ9XtApOPoFqVwn8+ZIT6r0fzLUkZXoA/w
hHFHF8Y2jSLhXVkWu/1lO+n7G0hDqGVXII4bDy5b/Tzf1GZnRikVYJJwxkeG7wh+4FLc2EXG5inh
MAFW8v9IulBSrPzu8+FhlN+LAGpmVw6HlXnAcUfD6PPyGkQ+jFHWlRAmV5cTzUr1leSMBLg0KAEZ
w+i9JRrG7oVb+9woUE2ygo+Y2/UBPLyhFXZvn8Ppr3+o0NbS1ScVI+wlXPy9rvDBYNGRsPTZTbW+
mFou1JvG+u6GN5ebnok+JCr3q5vuJGbN52wKsnDGKipt5RWacf8jk8Yi9ytkp+f06HtCVXbDvb+X
+D3TM11UDULoxiq1dxJ9gn0c0M8eCbJFwwusc2QCHhGBCTceCjeTLgEnWOmmVBZ+gH+hJ1cq7n4Z
hemcQqU7UaYPLHiTMehkpgLe3Guj5B0ctkRJNTCS/63lj/Ob1TU7aEKCt28751/PC0yS3wk6JkZ+
PmMVAMiNB9ykJOXo02CZIL5wn8gqS47tLH0sio1vzW/9ccS31f44er43jPtKLo/r7xA3FPY/Yrmk
dyc22URcI3vGdfTJtrctnc4Qj1tKZlhQuB9d4G7XKMZPjKm+b1c5awKNny2e9ie3f+sTM00Din21
KlS4VU+veU8o5Wphn2bMwda7pfkRvYn5C4P/0y4pAO8c+L+7RdGw0Javd6WuitZ/HGDnkJ0tpi7U
sWeNVr2DQz8de/kJ+hZBALWRfEhAs7asqCmOp5ZxFMgFgMUYOdkRTY7Zi9q38QwUkhzXsppuV542
B0Y8UwPnsDUVyu9V3n6K25pPGdV1fV7aVGv/JT8+uZUm+Q8s7RtuJ/fCo1M1OYueEfRHF+2QMKSo
5zQqqvWbVH6CfDG/aEXepxjvBgnWgHl0BS4MgQIiNYF7pXn4V4HpQy3HhqVXkKPFuIo11qi43Css
AICwMrCq3DD9g4SV7QCh9iGAkVsI3m0n8CgYI87yMZoQfciBq6p4mzc2/gYzjvK+uNoqZvAXwrCW
3ztB9SIcAVhJMwPfjNHZxujBIPSCZFw2Lt5wbs6uy5eysw9y98qqPycxNkgJRY4DbtNbuTPmXEQR
7P0C6Ox48WsYHEGQjAhZr9bmFOti8XrQLm4HG/SmT0iInhPtgB9EAAlaezvEyoD4+GwdJmQ3NCtF
rHeaMjM1JL+JABjhlVFLUyW5BmJhp20/AsobGFp+QNHxeAZ0pom4ZdjiuqFONL5BEQNVJ/9J79IJ
WztYMi2c8RYp9o8I5M/W7mQfqlpsDPiNPrAGO+xbc44AWtzhUbXnVML9JC8OgdZidLDzhiG4TnqD
NlUWZukCL3X2DjSS19CyMyHIHGtl60pO8ilKIS4dmQNwbyX8L0UaoScgMrueMxyE5qNh8vShamPZ
y2ufGoZG5yMgEp6aE15NnjkG543LCRCi4qaSICSONnw6S3hHYCZ1lhwT3k/ziq+O5GEogJV+PsR3
5xtFFBureKy0p7tvmhOBW2GCI6gEQEOLAuNtPHiMCgfdTNEQjJa4iabU6vQveST5SpXG0u8kJt2u
k0II0TfMEDCcoX6TWyz9moUDKDVHiZbDAWkCKc1wUWiWSG5bHtNrNDHzZlVh5gDKk+XcKUsvLljV
dXHDS1Llk0XQYpX0Yrp9l9VBwyoEL3y2wEPA4o7ukJdiOmMJg9QoqhkJ3g1bUTExVmU6USYIlZ6r
AxDk+GOIqso50QDK7b04xHhn6qR3xxpQwWCjuKD7qAp1gz+0RYKLMVmE5tkuIWe57ruuSw6VfYNN
Mzyks76/LsiB4KKp51uTqg+0hEIvHBB/zmQB5gC5zKzQKWqkUoy/2bLb23XcgJS7DRO+BVhgdi/Y
cQ58YxnxD7o/trhwYbB0lKxc1mVRAhbjM6+cybjP4Mr+Ara5NBrEbFP4qGbanN3euqDqts9+Dx4O
hMMUz5Kas8Gdj7XE+MpgZrVUbOH0iIS7Or0cERSIU2sorYWE6glq2ssB7cIGLNPEDhkLJBSK7MRV
es0AagGknPAzNvFePWqWBIMUKAn6CGA7LJDHsR9ZSRpVjtYz1elYCZ7KpTD/3tP9tyRD/CvkA54G
QUsai07WHqoZCqqp/gPxmcJwO9+BVUbHwAHtElZi2iSiIbPCs6AB9AxhV75LYTM6zm2/FYSw7p06
pbqXOMZZqxkutu5zIakKgvT/qidorbtAb+RLDFANWLIx5+sbdHXF9q7u91YNAaHEufAg3tpaPTWh
GYE3TWio1kzh74VfejkhG/8KSZmYNNBmiVzIio5FLMBzf+odsnvituHuTsOL1yxsY57Z567KakoU
vzo71IlJVyotSY44wyhjhAv+TNOVjjV3ukKFCZXMneqc2dlcv9/9waVawi9O6lDj9qud6va6OKe0
jKLJXnE+LnFc/XzYFp+9DFGPow2ZCoT7yHkgQWnCpmKMaNyJnv0lKDiOuFXW5hPnVX/odSWkr3kQ
ttC0KhI1jUEB3Y/KUGipe3RzWlr777jFVK9yGzcRBOqyzsSGTFWV53t4Zdeg3HdLwgcQG+KUzuCy
gzlbbvCNRs5SSFcD+gP8roaYDrlJKTVIHt2mkL+MT25IvajGkMUKCEqFZQKVD1DjhFLpW6nZlNzQ
5xq9k3bjSW1ATyUeYdv8oXIVN+x51RxQJ6jPD4VWGMhrI9hfJf+q7b8U/DT8HspJ1/LwBuVc3j+f
CD2rkCdxHwk/wsGJlaHo42NszbycxbJoqeOJvq8u7NcXvSDt0nVH0u9PsLlK39yNPkykHxmjRqKE
97vl9qMYgMC3fCJn9TJyN3FE6AgEbrya9u8oogXvSyjC2Bmay2RyWkqjYQ/afwwnidOtpP+7Xf69
oCeT4JDzRjVwMd2cwf/M2se5O6LmXugrIPWaMIE1JYnAx9c3mjw+PFHj83dUTnxdvGoaoFGrS8OV
n2FFWDUY2bZE93s4Benm/xf6Ux+s0blBrBGW3Z/KK2FHiWVBxeDdjhR46WX8QCQjQKXZsyYyTF37
cz2MXB8iUd16skIjhc3Zi23yblYKa4xL0Au0XUv1bFt3gbs1eY3Wq6UJXA4yjs0V2VT/IC7DOn99
diohfK4rAOPlvlAnXYPsByp7cFLlph4e+3OpPDVLbX63/JZy+X4oRZO+qiEjF+kWD9IeFHrwFoAr
ibaovtq1kuVZho6FHy5wXLRjtzR+2FopBFwnoZrhBXNNHpLA1lWBStCc8nktzLT9/Ih+xGdT5oaJ
Hjxn3u+2hczXzKJ5cLj7pNdklCINybjEg7GwS268Naz5LHPnRGvWx98pR3lE0KbYB2sspijmb/yG
AMXuuTiZc/WxFqEeCYZovVwpBO7aMyyvpr9yOsdkucnz4ZzACkPjx1drEJtZRLpaLBLnZFuF1uQj
SKTn+jKp7+2VxgXQ/HNyJl4NjqiTX02f+v7BW5DxgAqkx2g8/A/nI2Og07EVO/teNT0n20u+s+tv
fRoy+fm7JTQPAzg4ra8toVytkQLXMQIXuHqOd/19gjyqke8uGxdgmDCiNg6Kfpo6L8Ji7wRSWVyJ
nAwZeMXgynEHn0umiBw1P2+DEllh/+zTRLCd2Zcap9PDTvyLiossUvg1BDViA4qLrTOUrNbPJdT4
mK5hsMFbnPEhj3MAPaS8XvHmSXcgpvp2uYFbD3Ec+x7DXGqLkzDkbH33I43Xd6UlCvTMMACUDiIw
KAc1EuGCOrX3Tf2W8nbRUK+qAVMHos3mjZ0OqV1/aju/ycENJSxLFPu11pE2Ho4fiUMQ4CwbEgZA
0rlgHyDM2ScVSkapiL0hxQL+UXpji4KeXF0iFnKc6Bf0QoINsL++GYXVI5VHBHG9wCwgycKB7PNq
wbziyPpoaZBjYJK6WgGidWEAD9mAu09rxCaiXvwafl801ZVDJRjRpW/H8nTFug1XtPFya30z+niO
+ThZSqikjPdrnJScnLEG0m5DTmKCXrfe7xQ89y4gwqKbwIIAFluVxdg0eGJa7BAGcrXetORPupQH
gg6w6KaD0PL84SCBd7dBRtddn63t0tp0RNvBdQcXlUQSGGDL0s1tyy9Ot1dcn7lbGy+jLxypi1Um
8IuO4MdSmtVcL+/fmU3WZS7/MBxKaoawRtkCDZESIsYwVvOJIUZn91UEDTXCvCd9IpVVVq2y2ftT
L35rRtHBHW1UOG3p3gzPpjxy0FMtRPxOuUCuuWxwpIRDv3rXGKBAfKpzKu+VnjZMrPWOgfamlrV7
FmztgXC+nms3GoQj1MUJFOYo7wHdyB2wNwaUEutnDNkxINzeAklwjQH9+lJ8dVWw2ZxraYZXxttD
ScDI+upxj+4CjRyemHUz/ca6ajBC67eRT/QA1UPqiK62sLcqXHXZwMbD0dubdtfWiIPiHtIV+zXu
c+YiAjcnd4aegVAq77e9Txw+VKEHThSydia1xEGgSQVPlO83tvfRv2MVKQsdPmLKCWtrzU5fBakU
zuGN28RR205yOvhyKD/G9QMmY2gcyLfCJOwRuLWxGXB99nGlaXpxLkLn8HtnVranGrl/YIF+867P
Xf2AkCPTvjqowabjQxRm7Fi5YagUaJUK3+a534/MbWwsykk4r8qvgP5Lx51zw+FgJdbZOsKXGyqi
31jQLbDB4jjlCu6cVCsvhjsp6xFahsMLwEubpLUXQlsTXYYMjYZFfEOh1EuNf909FRWXVSKtQMvo
iZgfSQWzxMZwrjBfLstxg9nLIaPMqoXYokmd7AHUhhks7WIX3B0MLCsgQO/htxirTIHd+d4cwTmL
JHa6dv+sQAH9dcemryU1rv0wiKFtUf9o1GZAl9f33dwlFnGVN8o8vCXEcXB0cFyX4GM8dACbQjjo
k2yrDn6pLCSlBkdw/qjBDtQZP+Ac3yhEp4fidE7/IPPIgopQG3Aan4smXVOua1NmRfqTHBkERyKk
sD5ra1zmMhDpNGhsqpMKhfOwVUIa3j26mjLDPXvusL2BNAo24McPOfLNW8ctBLkdldAXVUEYULNO
51ez2tO1a+/s9HFeFHq8RrcokYoY2y2RVWeSCrtVKu5UlyFZgoKmaF7CpUIU+pDrbk0oDDRKMiko
6k35ooLWQLwhG9LhvJC10kEeCODpkcjzytB5biO4DVBJ9qoVJuum7GcNn6i9YITH+m1+LkTBpWbp
s/POaQ8DLJYdPhLwbRoY4Wf5FULAJzTk2LnfggkErZXEI9o3c4ZTksuDGUOxJrkpKO4kSBNR/lbC
rCwHrMSTs2uI4B2wzgESaZDauWzsAyTf0rSzbEJBJRHqdcoDLkoJaNp75DWW6fn4G9mq8TWjsUmp
ZVwWZCBl5r/6JLOlbudhNppPjasEp0Jyj0Q9uLhN/e9GUYYGOBZbmgM1CAbL4XVoIeWNUexR/U2Z
mTOQMut4pAiopepG0RC77xE8VWam4fLHR1HpwFDXHB+L3QkS3gc/pwu6n94vXGNuKjSDCDFVMTzG
GdVUxRXmBYH50WAutUBZaHLGQWSKlljlPIXpEamVl7flQjEybBwYncP/C/H9Ji8MjZG+QpQCYLfs
1UjNumXYnOYledLn9QctHx8ygxb58nJ8Rl09M98Ch5kx7qIxvSt9AQh9lXSa/pQUVVqIIFil+c9e
Lj1WPbB0d3U9z+ISswQ1Vl2ds00fwjkOLyixKNl9r/Tb6MvxWtCO8dOLUOhyHt7vGVupxOHWOuI6
n+ch321cUGwZY16LvFbXQ+xmj2aqO/BIuNhml4VGGEgIu9Y47KlPeJ4GrF6AQXc6POvvUn85zqhf
eubdz34KlOFcq6wmd2jWNm70rwweCItd6CWXvalf2pJv60Ob1cSM/IfDOCZ6+21wHrddwH1AzCEv
M1cKUpWc1YvKjeYbZE09bO2+6+EPvtv10UkyH+JlgoJh8g6HHlkCPVRRrByDQnNd/nQ0ANUAoPKF
5rzLgjIdVmEvWXY+FIQWlpfFrfizBJZ+fLglpbjZ6pv6RbBEmINETX200P2wTHKIUUunO/lN7St1
EQdw9NCHX4XEUs9PykrQsfi4tdgm51X5oiWoC+yhizjQPkF1DsQ2YnR056mzUlAti7tuQWszRXLX
4UdecqJTK2UjXu78hudUJkh3dB2rvqsNycKaEiaricDNcrHRO3ieK1gniosh7RVyOHd6f/mCDmP5
B2mOrP97oWk4Mdjm3aV5qwmzYOk1DZd0LmwqLzU8tPVYXJTg5en0lTVycf4t5cz8Y/G2L83IOJT+
BuHhjBXqDWCx40rYNrIlYtktWDHBVeIVgF5NcsdB4OMHeHmViymdK+q4Y8zTWS2+TqGtWCCj/WVP
49/pMa5+Xj86sg2b1metIlDeOtRRzot/n7wSiG398JhndW4A0ZjDu91A1rGaT7m9vR/kLxTfZivh
3EkvfPZvlBMgi2KK7YP6HgO7O0JfmX2QK16ij9HzbqK2NzI7jiHZBi9isP0xTY9MOBg0HG6DupFF
30ntLx/K0KhTH1PxIy+690JDpNgetYIEWPk4gYQfMAHHhcwsv0MGL20E39uIwCHT9PQMejpcF5Qu
Of+FHF97YBh9y4gE1PDO6yw35NjwYC3Y5s9+Xw+X/sadIy8wdhCmrm69Kc/N8VHtbDT73C6P+zqt
kIhFZe1MGFNUW/8vkUUspBngKrHN0R3E/xOA4PmySJVk6Y3JUERSRjHj1ANldRYz3d2Ic3eynEtr
DJX6glBD1UYNT9eWaDWIZOUodv3so7Mpx3fXxwQlYIwME0X8hUvtJtBosyTiO8pWenNruOGKAQWI
JZCVYnHL62vdCI/V0qnPm5x+bZZ2zzav9xCUNnO/xg7ckB8u+eBd2O8Vi6kLnsnIp02CTgc5ZAzH
KHyxBEc8NlQC+p0DjgkhIbtNl6gP1ILDUxVFB3DWPe+500aICCWOe641a6adZcg+CS3dxwNe94ok
MwRJyGB4Dvg72LqE9RDN4hjVHggk29wiYZmogWa1CY118TOQLHfMeqNe99HPN/RFTP7V4uSkJtPZ
U3OpXolHkGopd0hMgRrRfrm2TbpMnUP6B0oXgAMLAfODwwipo4Uj7K4qeqq1KEKlztv4dJAJgvLY
5EoJ7QYvg4CnNDcsRGP8EgNyzq/TVNCRnfQ6P53a0n5DQSVtq/Cvs3jUULh+TabZTPqhjNzZYZYU
64Pd6bA1vtZQrLTQvjj4p6VgkW12VrJ6JOl+yurp8aDGxwQ0VFfsX/8K4e1JPHXvgokvMMrZlhES
a3aPRmszmyfvmrRNAdh3QXIVuh2QeRKAsUEIaW9thKdA6S/sOSkGdAR2h5GFjtmqoW29Hypn57dC
pC0xSerRUVPTMkp11svE8A32Sqox7mVoUUm5i2MKxjpTKzGTJXZaqbJTSlNemoMMXSsOPHa+3O7y
ST79pSwa9HkCMd75/lW2ezSXxd3qjQEVmwdYUdxIDaSW1Y8/rgBnFV+y7sYlANHFFuWRzFZ0ckIL
L9uVh7kQ+qDfJ+0v/7tBc2Pohy04FLr7xJjGJW8A8BZZSMeCDUMuD2IZtH7O+LaGLC96vLc0DHTp
dal7Wfd2U8tPmRDnYwIdnD7dmvWrJfibNgx7xSNH42SppO0kWJtHgeGwLPBzu+tRL3nfg8wsJjfx
lvvuAHqSIsgruvSXgBvULt+4Q5T09/esnYGc23x5tb3h2/RctUUbBfftFOacPrjE8hxIjmc0yUzz
/fOS5LgNCPL80PeZeASXRAO4kYWJreV5k++zUy3LqDdL+tLNCVJzm1W38OLOe7zLV+K7/kkr+3UG
aqGkjYKBzwa1zACE41t4hW0g6VizUJiU2RNK/ZXVraIVuqHpzp4jxzkv7fKw2ogml+QtTv4GGtWN
0MxGsjDoV2CifHpCUg3JEOxitEwWsDy86e3LaDUpr7oRf0UgI8pQThq1DpwBgCKuZkJyyxV5qwOT
MTmgEdztloUkS4nrr4gaQAC0yuin8wDOTaL3/AuhL4b/vzzSlqx46fUAL9zkQPJbaVYwLDtQ/L6T
BYGHi7mWkvvXCzAcYCNdu4njf/xSCzF1jUGEH6Ksw18VwKivAwsJ+X2Q6idwWjs5j8VeeQhSj8vh
3QBgenfUZbrmZVueBl5km6ewzN6xZx0qGVKyhuQ/6hDmw9nBGy7vw36bj4dOPr4sEccBy8CrejUw
l/K1bMRmKAHUJS7qYlmvG5u88iPAtywbUzwQn9xctZ8bEWmwA2F9hRy5erDKjvuu9zMQBJ0PvVJs
vhiJkgnFQYxlxKqamnGxGB/H5ap01LwJqtmTHlsQQCZHUYk/TczrXZDin+8+gwI08QZuTBiEIsAs
3oaNwK/6fnSd7wMmcRkr1cCACH7Ojb2njJHAAftJ/jK+Z4hGm1FraXq4zjNhgxN7WwtVIOW/PrCK
YRmuiBw41Fy1Vkm9BSZHzaHxo7F5jitCfzI1zh3WcGNx+KiL6VHjolcWeRvd1y4cBNfMjvbh0O6D
0Y9doixqxR8kTQwVXNyzl16DfO9Ktp49iqoHuPkAflBn/rI+EvHzcGeVTwU28XNdy9YQqklIA+5v
DOZm3SAwoc1/MpokmHWW/kaJQ9WbCrKWwB1vT6rcHQ6t1WF/gYCphl9RhFg0yGRRu/vkLfp45Irj
sB34P49jQd2SlTsU5/KorIsz9IHFVhWHQEhDFyydnDbWvcrPbJZr5z7vN2w8BHYKd+oFI01QODh2
aJsZ4TvAwHRnBM7NaikYdijjl7KcWFqYJhtJKksX+txEl0o0QkwfKqAkqg9VevDb69Nlr4z41cyj
6pNHL4oqdIv2ilgyp8LF6AgRRdsz4y5QsOx2U+V+92U5V6dJJd1WNlS0grVpv+85Ed+gSWwGcFIl
XEKnRZHLHzdCSkNTtI0qe32vZQRklnx2dKKa1qHHRtfAs5aUPilnlma7IQUD+Y41hQYFekjkU4da
tC6D4btwH8WLl4P3/7Z5uIaVoHi9GUDAsn3iCxAH6CsBNUiAC87JVzSkq+E/RrQVgxBP6nuM87HJ
JXDgKCEo5RDFkcoa6tTqM9KrFh6TOEqRdDN6rLXP1ZAwNep0NpeJYcuWYkKFxfBq26qmZlFWAhX8
h2OQv/aKc/7zs+JBlx5FSuIjO/lTrbHsAyJ4jvkEJBDfjWxR6js02C/nMdCItUeNpAJCVknXJDCj
tMeEM7ZyGfLMjSdRfYeYFvw7tXUu9icaM+Y1PktP/OwaRhpJK+jkmUfLXp497x9CjIbzs3xiAznS
YQEaUt3FrJaAXZteiyY08jSsUDPaykDCLpS968m9KzKb2besMx+nOajACuXi3yq/bGFbKfuPTxb4
7F7w13sqLmkfSdlI7gKFRttUZqtKvTMOJJjb4RxasEvqbynp7UtgCOll8sW55FWosrXYv/uymJmJ
5M2F1CWn79YRPvEodwYlewvL0RGRjGev+Fz1qSvwidmNPojO/Po05WcUjikx0iqV703rBjKUlxj+
jwEeEtGQp2mYqr8M4w00JdMcyxQc5+1RsqvagMCV3/AaDcpQdCRpqid8jcDgIzhRJn2+JRaW54z1
JWv8dlqnl213ASu8sMyqMG2iQ2XJYUiz7hvTw0kIPMUHGsATmmT2lH4fTz8Ssxeozjv4fqWRYuOZ
qZr618WqYQSVlvB9nANtaPZVE+QvjwyQsIl0cSKO59UbAcHGT4Yz8ip1gQ7cfpAgYwX6IcuOUjn4
+MIKTEkUETfnn7ecT2cu8RMuEyMcoI5FZ7Q9xUg31XaULO+zkspmkXcyo/koD/7TX9xgRiGOLGj7
NM2in7Yh+bUjrgMMGbK/R5lVdvWmTA+zb+DJ/z9c3PF9iuMJQLfNh/hBdTm8obWGCfBrWIiX0kND
zEtgSm+kIdnfLifxhDJXjjWLozrNam01R6A/xVLBLIB4rUmht6183CbzEo+NrY7IjQd0fiijUcgd
Ka++ZNojLPoLMFnDrAU0hEkLaBlRMiNKSNzVz2h+9DNe0KA0UQsUjQg7OhCc9ULxfwIf69I6xgqR
SK4PzxrL9Pxb+z6Q6OCko+s5GCE8YMRaQ+Jw2XCIoptIsW6HYOoGEibr9CfIr6djyhuZUNtY9Ze7
DZuPExY5q9JxCIjsVQ+gtkXZi5TCSDGh025cX71mtyql5RgTM7GidnIWMprB9E3tK2J1W/KB5S5j
bTA6N29KONIU4IMYzAoN6ZHTZnkxBLSgtQ6S38oZk/1RVmW9FmkNuMpGuH9WVDSeN2AcUBoEo1lX
x4r9Au1FKfedNpPPDi9ZIeeKf7L3Bs3Wrnz7NkOYDcEnjq4TFsNQWVg7YW8STrU4XF9y9/72W5/C
jGAIo1DSJaxqMWTvu3PYW0RxrEys1Ag8nTlW1pLBQgbqrm+B3D/Et51aoHKZCfh1B2aaPDc/fqhC
GsP281JyHq2F1MzWExbY/fieKTpT4A/OtLW88hJyFa80aZKNooDiILZaV6KNydSz8Y4QtgLR9oDp
wh1H4TUDIFydVkqo+3Saw4PwVMte21U2agF0ZG95laJ50ajIDSJS6sdI7OmghEKJcL0pC+Pb88VB
u7mMwREQH8/gUlVyIIBDzg38gQEEeyyzNtfRIAgPGOMkM3aIDXHHHWx4eYjfCVZV6RbHiWWjb7RN
OEbSaZRhzb4eTAxwir9wcEc9OG3ZLDwJ/y57HvmPbdDM6Gf7SjqKqvF3/2LH+uULyWhhhLN501fY
thdGp6MqruiyRgj8H2cCC8nT5uBp9BG4phfBupIlFH6qPzCdJog6ipze2eQ9OGJbB04cvipIELRy
8dQlP19uvnaJUwJXFFEzHBb4yUDZ9eyPUaO+edkRpSbfXLOxG2vnIZVM8b5BL8AI+iiRQCyVuBuw
cxlBlob7Ib4Yy6skFVdUR5J2i2AFBPlM9HHEEJjQz0m/hq5LgqKn6I5o4VyA+XE2QpSx0Ws/1urj
FjZhhl3gqxiLe64gdooBS/9LUqzHH1moHlS5mux9wtKFCM699jjfJxt7PRg6PkrgFrithWB+t5d3
GCIFxfFA1NqvzJ/VE6BHRMWrFJDrt7RPL/ADXHxzBjsfFmzG3cCYnFqrPhGnFajTBN8sTwOJciDZ
nohgBIirrY5v+Sc0Tx/hd/jQtUrZXM7ctnzxwI55Y6YjdoGsZVklFLzoRRe7ZafrJbpKcZ8HDIBP
v8bfniGOOQuONHzLGEphQZkht8xXwXzFTMEVK2ADmLxWTEK2y8ew2zNilDpFlGoeg7o0HIhD54lB
tl1dtaMapbOykXwweNEpAWF1kzSnHx9V2eVAJpwnUPSJYFqjSVneXEG9L9xwfIObCdBDgvraDAPI
cMmuivzp3BHkgw1jfPpKKY6dweiXrQXI0mttMSy2QYxEVZTXLWihTCf97ijVVRXwht/7qUq9jupU
514509l+y8VdeSlBcHKmWTqUcV046OWjoPh8CQf2k3/vUmdv1oYuJ3o597RfdtQYl3MAm6/NK9Sf
zhEPf9SCOGKeuyZo6ie4tuQHZ9ljF906a/LflVyZAPPD5HUlVefBJ0SiieGUqshIvHYwai/S8qZ0
g7w3FR2BUO1mD04Cv2q6zHNrqNgnRqxvEdtBsDxZ3kCeW99kFHN/tlh95gWQphdgO65yowHIkxM6
A0N3unoAvX/pDl10Fx8esQSyIEkeXo6kd8fw3L4jAQ4xzfgxrHiJim+zSI4TOReQ1SHNJm46F7Ce
3pu4QHFA9xNNfzwjjqsKooW5b/SEw5FXiMbjRBSPPN9VCng/Rw8vi/FXZoH8Qoc7KORgRJkXX6ZT
SBTvHeOdEPeL2Lm/LY+6OB47UAkUBqsnFyJ+kimfNcZnbdASQr89k33vFdIZI9/YHN23P+0lYT3A
Iqc0axwi0bFo4PNz4OLGcy9ONyC33+DSgMtkL+vgfbvbva/uI2r/IQZUtb4l76t3BRTwZzN0ckZc
CbOIqV5IFoonBrGn3vFAW6jknc9L2bQwcx7QRQw9Yh1+K4eWd95DZUvNsW+QYJnkJynLa2PQE0Hq
JBUQ627a8AyWahjIGGfJBrkc+ZQLsDoL/EQhB2+Zum0bjsFmZJYhJe4zwVNkeNi/OcECF9T0bdw6
B68LiRlC2CZKCXHLPS8rySkfjvVEDmGHOuiYNW0Gb3rlrv9uu29Ca0Ywh1KLuppvW2WpNvk7p5Ny
kQJJXEKF2bpBah229+9DlR2+5XSDl7nCF2bOPUppPbIAE5R2nVf/bpSouy5sCCmteYhhZ+Gl6qFe
Kq/zolTdtQxywkwRbln6fUZvXEfrfypC+lAbDFppc8/EU/HtnbB4YDR23JXCCYaB0jBuIp9fNTOS
BVlqPoNcqMyZgfR1f6cWy9E4paVQNe75EemleiEYOE8TS1lLY6RrHEZx3BXfLnA4hYML41TvT1jP
OzQrJxjW7d+kQ4REDZPvT6rxZYLELcWIkAoiXvO0zcp8go0Gfl5recFVVzgJXTmByqRLks4CuEBR
oK8mi0J6KCZLpmrtaCXix6xaMlqUXT9Ug+8QD4w+xKmI6PhXUyfaiwbdm54tOwFR+tWe8Gldwxbf
Z0rwIV2uyqsi8CCLWw9tcfeHVMBklB2/1QNVj66iKOpX6e6LYgEESIun+whl3HOuaoGuknX2rj0s
e/JpEdcon8ZIhFP+TNdKG/JWi2mD98h3HtndFiwrHLJmbGJFpDDCtP2sVMdTM2zE3rgSVpbyelol
ZSPTti9bzQVkAsHamz4pl0UiyfrdDf9wuCg7QWgdykP8f6u+FnYOsnZ3s6ZKobSYjOOEbY64Gqck
TboN3sR6pbC79xqa9akD8C7wrjGhTK19cBRgzLzM+OPBYsFP4DKqsbaXzbanD4ZDHn4bu7f4Twhj
30qSt1o9FEGLCVz+8RznwFE1+JTjngIRh7UGFMvzBwnubX9mIL1ZGPXrxKpIw1VF83kc+xjr3UGO
5pPf4VMAbpGPQOYSyMuiA94lGQTbOJNXdYfgcVoPeHXOq+JBMsCBfXuZpSqTLQXGj0xJp1YKBaH5
h4jm0/nOsxCYDYrHwZCvkH/HMJyXeNuonnaqqxyqAk5O+BcXNGoaRSivQ7uaBbCkBroKlJaPh+PX
Qd72MRaI9SG/EaccEudS7JFDNswKnbJgSXxWvjO+IPr52w164P0or/RhsW9zJ1PrwuTNVXiJcjYg
mOj26tQYewLg6FGcy51GYR0nQADEF5/Sr10uV/jjos+rE969SjIR9hcER+jrPKg7Yf3/tb3x6vfs
+FuHP5j5B6lDlP5c4UJVSgdPIYEX6HLYccsTZJjBGF5FX/eFU3wvWt1APwGNmkPi3z1E4woBfYRB
bM0WHKqz2vMTJ3d/o1eT0/QQ/GdjTnOB00IgcprjkgYWLDhwKwYqfnFmUvl+FVwds8/IdoxjrTl9
78lmwr+LwXeQwsWJJvkNwY6lvE457sAQ3DrnOuahLAD3xfQIxiG5mA2cp/xbbMEiXPjLQdQu0XFK
Zpv4POmlpRgxLhq9LuV4QjxsDh9UfEBYNg2sViF7nJGZ85ArtcBa0eMDY4CXbAH3f4zaVxa32QrI
gbSKyd8ShwFQ01iDrj9Bhv4RmGs8Y6xu5iwNrVAZIqYWwHwonwXWIZpLfkvMNaghHklp31cGCnwo
GgYassoounCqT51DgUXMXLnPlp/zmk346E1fHu2iN4Rp1vhhuDzK4cL4hHcmIYdQHiWmhyrCmYWT
vug27qRCvlZ8ontKBFGqf2bSSA1Rlg3/F9D7SU8shWV45SU0WVb5ELDKT4pFmkVmMa3ePNMU3bge
aWOTbLSUMpRXlSCtATcWaACI6IMwydShQc7Bv/RFMJ/PWDUOh0ysxuxnXygPvmhvIr3dsS+TGbLN
PhfGWnatBKESsqi0J+TBe6DkDvdp9fMJfq9WB1YKEb3tdni8UPwt3G326JW4OqkOEnlgbnm/aanv
4F59kfrYNwOtsbLimipboHxlMvxixxrszxVne0mqJqswsdAWI+9osg3RDzUJis0sDDrnuE1vFHge
iUXRguK43xe/lH9EM4VXIlhfS9+7XIb/Mg9NlUcUOtUuBsL5LiI6zWCyCuk6vbg70K5t3Nq6hMbY
rq9LEuAaVBmKqe4+jo4zszOUolIMomDZeDjCFgw1//O+t3EAfbmqplofAaJodafWAnEq8g0t42aN
gihvv4K1nDoabaE+BkL/lmUN5NPPx6vlgBImizma8MoQ+DPwPrZrIgU+kuHA5zqID4qLAKH6e6Cu
j5p9bwY2oGGg39hV7TZodU4LpVjRpxFhryPuyK7R3FzWHdOJGYfVMIDPJO+o0FNJIUKWCqxNPF5E
93uNJc2UfQaXp8rZg40toX23B/EMJ07mSNIWNDz+F05k3CI5x1+/um6wblbOurJcrXRbULiJqlK2
X1ml+XIWhkvHHQZNx9T/aKrA86BeCKGRcd12CnMnqJzrJKbtF4ABQZepBG/RvoLv5oXOr+9apDY6
xR8sjwrzW4EvT63fSzWL67s156HnCveTfAsD/idmMufS/NamSLY9iKiaYxazAVlI/CypJnGuhrwz
hWwCKdqA7y40KGFCQddp1YBkZMrYtmoGWzKRYfgvrvKfJ6zuhKXsEUzwb7d/JV84fkgRqZwz3T3o
m6aJ1plPq1K9iP+hBBnx8uLiS248cO0aeZYjVQ+XZkS7xblHyNeyjIXWiAYvg4TrRBAt2bs+pt8L
4FWlLK2BB5sOQxnU7wEvBTcNzjpG6QgGgJulcUD6Sq8qCH9mhq7vRHKCk/fvPjN1ivNo/3BCy0ui
arH9YY+avCqy50Glue+lsAiWwuTsX4KPUTQXkoyy92HiSrmoPImJIeE2EB9AdgQl0KB7JJpxVQ30
bTgHIQTVtJC+E2eQ8TyTVN0BJrfiGhJEJaQrELo7HUNsuquQWHTYsSj9LzDdXrhVk+85BUo3A+Rq
7SuVOEW2mCMSjgLRmuMlE0yIr+qT3YFZgGFFpqMd/4aFjY6eG/oZt+Ri8rnSOz+3io92ek8BzYTI
ZwbWf1H6anFfuXS9Z9lF6qb4MgWja0/NhiA0YQpw8O+Mq4BrGHRsnXJt9kCfLb/xH6rG2cB/RU0B
B/HV4FuIKVwXan8og5Ghk1VChv8Osyfb+rR1wtX3n6og+7wiRXWE/74zrAFA66gh2kxTiK46FDUm
RnTQJ9tQcmVLitIuBM3RrowEWCj0xlTVEnuM+AaaYbc+7FKku5tJnJPvTN9n30ucZcN1RcIpEe1T
DEY7QXP4z8vUgmYCsueWcYZBE7W2/SZNSeoJPW1AVTFxeu65J/y6DUw1sGacuW4gaxnd+gm8sf/i
OTu+PwsdDCUGyo6RUInM79ScC85pftB/Ylw+Qc/Oelqthgk+7Xj/nbLIyCdPboFg9uuR8xxPGF7g
JwTNm8CUj53JmF0bnHoyO6NH/2GlUMklQ5itsz+/Ivp/aSxjyi4qtuTKuFo3ReKAmHVATeC6Jt0M
/Owbyb8HzuXBK+KiwclXmmcIEJ4cE+M7+aREe/16B/xKd+iuCajBRbM0l4KX7FJ61rHltW4oSHE0
VmeoyJra8M5qYSSNxE5m2azOLwzn9GGAHlthr0wTIvSDDA5u+2Q0e72gPeNUTv5rkagcFnovzDft
cyAq+1X+D9WAmlPkC4dU8g+9J0d4Jq8YHGoKmFmN1cPcTXLLkxmFldThw161bt5T055pt8TN/9Od
Bhg/S//WH32iRuGLQe4P55nMgQP3uA4nuPqsyvRjCBsI1LQnL2JEKHlLVcHEeNRSL3ufskjo7Zai
eoKmX3/jcC0WB1EamcWWzi+3F4LRkPe54W5p3NgkjTOBq6ULstiDFqsFDBG+cBXetL6CpArIgTq+
GLhnoi3liJyE3VPtLJyzz1Frj0jdmKATdyySRLEUd7NjnfLCKJClGo2piRa0HyQClHC/+1ihoTkW
GGNzFky/0cvMTelsTRy1L1EV463BMERcS/Tl9R2Y7F+1jgc3BP1yq4olEKkghli/SNZKClogNq7e
ZfTz2Dg5vUl/UcOplyC3gKMq9NOECDvuYe6/Awhn+FU7GD/FLtqDccztGAKEpnsQgSPHz8Tg+DW/
xV9unE8/QaQNMFPzKi0/fh0hztF3BdkZGGZmR/DMWrii+kcb8iYbDJ6TO8sKAtvw5ey7/5wYNPmk
3SYHhRlDkdPGF0gQk6yYE5GW88RiiDRM4kx1/AdAv9tdGQCGBtkZLtREsI3PeJpRN8YQOdo3Tyu3
sBZjkMfTrfpQkFc9kK5O893/KGP+pvVYMzNr3ARgiyxwDOY70K7HVmXdQIoRumAYKoiMK9EQfdk6
UVA8oMwZ1ykAj9v07iUx4nq6WocQVoBJeUC5UGGQTXbI+g5OFsnj60tQVaxs/JUsQVjQrYus0Yn9
uzme7RLOXO0LFZhZtsHPWc8ERpp3BuIIkTBa6PTiuyY8E3BKZIf8mH/CJ2ztbl3frU6U0BzhJbOw
PFJbV9AaLvhUquh2gRecDBwCIbJsCrSJ1ERXMj0NkBEWyW+DQu4Pkm7nq3EsGEZcQX1QWmRcEp7c
/RAAUTmVkgmPUXAht0s7APyjx7zigpsFG8dygglk0MyKvuCvwXewyHE7MYHNSR+spt6vZFwqPjFf
ypTlIui0nLcFE9gBePWToRkw03yeX/0Kw6VinGhYeox8UIU1+OZtjX6u4BUVRHaJuek3vmvznalp
OJpsY9ZetSMSmlNWcxRRIUtz96JQQYsYCSA9Owe/1pYje5lDahFyiDRF8RHnMoKfzeo9EdPXaoXp
7RiNL+wtBvZS94eqdopWkJsSUp0UiMQC/i6YQE7qhX6o0CePBpyhP1A82oJ/0J5IWi4jFqpEku3V
NHmtnrJ1F5NkI9HK9U8h2MKoF8skyJhYAL2vee2wlcAcy6Sr1PrNlLL08HqffnWn8wCKdGTWhidS
kpJ+f09srAwXDPKmf2xwB+lyFA66rnThc1rMKZWMsOPz3ybKzA69v1JhkWbXo/WF0t/hmIjxKMf/
o4BI0kOzMTo0hDod4QrIhG1kVJdG+0tXJOybHLIYB/dzJUS1xpH+TTClzmMxiICatGhwCjk4ad0b
QTpag0AX2E667TCG6YkDp7CBqt3FVRMjRtQrFqBtXZZJ9mjIJqHlhq6AH2VYIrtCjxb7/U1AANw7
yqzNIsykWp0/s+gr53xGpNVMCKtdNoNzSnv27kXvaj2SVO7jIC4Z0URahwFWcupCatYEGrvoNKad
rF7lwbChKzuSi4Ccg9/1WokmDzAxqTUuGIgl6sed08voOBHgh4wP7Spmr7e4VXWYZ0lo67YAo9a0
B66gnd7vNzPIhi5eDJK66J2gRXOJ0M4IjcIMYek83uH1NH77xPgyzXy+C9J40mSy/5fPUdNxVpbF
8IwfEiXUdVrI5wJ1nBS2p/BUq3EIltPJoK803o6X4x0H5ntiKXYZx3NtLQih1ismXAEKoEMWlIBL
h1oQ10dIDwRjKxpBrdzst+9ULN7ATSMMcwf9DhbOiW35g68rfn/VqHAnnoHD/gpa0VXkGjTf9orK
QPZNlMxm+dx8Lozt3m2+FdO0jRjciCIPrO5UF+YHuEKiRWeDo9RFdGHzkIME7eXNZi57lS6mSmbr
kF7DTCMdVULf5FtEFEutsSfGWmmjk2ho2PWYwf9o+IXyXicFjqjvCkCTqF7rt9MfEdYF+w0Ny9t9
PKMArtfbk1Wk5Mgq9CXO3cMGjdp5sz24x/GgeaTDV4zgeTWuvzutxeiuzg5r1uATeJ7r5+K5DIDi
UaT7DzMiAtHL0QxbqAgSg/q/GHgQvWtF6D/9Ou/WjjBBp/tEJio6qXE0RGvlF/PrZ1MVpd97BhTS
Ny8DiSKLNIIRKybpuYYDkoasqDbV9f+VRgtTY2ouSo37h2Em7ctvAH3L/aKS3gbW9D578Q36GXrS
Tlzq5e/3DT3/tDcNpHKTHBXfbSg3wJKx4Wje51gw3uJwV8xm+z6M9npfvg5NB3roGWUS3IOhVhmG
t0xotMTrLN7dcJ3iCgvKacHJc47izNgStawVWFckBMqxtTzvAuO3bILV+U/sjiTnYX8MnGUYEKkC
EOk+eZuHfaE4DiEMep30g50Dlhygsm1PWMptt5zAdzOi2BCiEShGf5YhmGPZR/2o4urPSIH4Gh0Q
cll1hrOCNKdxxSLEOKNv1ic0vmESTTWNG7x2wQDZqfPZDK/QubK3yf9u/2VePqmK+PBOVelPgZaO
URd5WXgSc89iq2gJ0CTLroX+NziNr/s1+PzbMW/aIyjmH0epaQHyIPloIWnFG7Qy2IzuzbTgj0KV
5uAi+YUIlFDv3Lc2MtmwLkOBqFnwj9mQMrtb69kRL8YquQjlPpliIOn2qR5D5L0BfOht2or63/fk
gs9uClOWPAtS9spQ9r90zAi8t2XGtbXe3xOrE8Xfx0Q/4BkH9cM1Qz8eRYSSPKFG0SWXBWN1X89m
eavnFNzELMv9oDccfhXxuE3/SvGfMgHyLItAy9eMGGGmIGr4Hx2wi6R9IPic275DJldiPLGAbxZ6
e7oph8mJvuMTgEdHIhrT0hrB7vySIgVZo5NoWaoF3UyKhXpJoY9kiBbKyH0VZ25gRy8eSnti1cmK
K8NUN2vPM/HUV1s1GTUAc/EgU4Ibs53BR76xg8wWcl/3W1p1lJtQn9xwRZq8xxc0nUCEQqyikUyb
oEwtu7wZMDvZ3L8Q6rSgrsCenB7T0JjhhL/kvwqf7R/vACaAb1sNFo6+ZDryfnhoSRxhGcUAXjWY
4WfBynJffoDCYtjqntENwEvlAShnoYpc+KQMz8QlFLZ/OrTkN4ZVvfv2kqlkUY/fwNK31JIpd/gQ
IH3QgochCCNADbg/fNQwzzMJcWdadSXyi6sEIutMDD4rXXLMQt16RtwwYCPoKOs/ALKFxNClQGmP
rQXItOUc1SCALYxTRe7Ky3W4GHHnJbS9hAjtH4UaIVCgYObfFC9fBJMprq5z8Du7Qs0uOC99dfBJ
gfC1cM4VLGVcj45yN9IEUu6MlofMwil0PV2xWEvKqaLQ/rkbj5Dj/1rvtblQIIbWKGNLkPkPNK52
jUnaj+FUo8w5AxUzHggETW8VFlryGERELyo35JmHUKxItGnBHKm7bs+Ut+feeYs4oqLDBCzsf1vn
IBfLxx+qw4BmE+jZC5pS+hEAtXxgx1UNLh/ptxYwZLh7jxY0+xT3XBekr1pM8gPyb6sLQLvburrU
eJd1VWNakGsDI4njYAmteNiQteA1xR0oXTpBKl3Ty+qZCbNSoBKRTIKvY8jOHp1WRkszssTFV05F
cxwiHQgqEZc/puS3iC+kCSf/d0cEZ6FCp3cQJVf2ISlt7R/k8OyibkE4+h38CDoLVKeaRwhiJsGu
FXIA/UWgO0l/Q2H/CVSecIvCVORzVD7R/CvoszQY5K+OeuEjUy+q6CqIQBbduqy2Ltjh7ZrmHi4h
rH73V3R1oUkNMXJvMaLAFfLboBF7+WLgltxdj9xGe/ESGwGOYJry+4d/4/rCrB1FLYXBaNWuR4RO
Kyj8cXAjID3DahFFdpk1NsNgrHPj7KISpmiPiaLMwRdIf46yGRJUxhTy8N7EkDt2NwhjmaCE/fqo
vjV4WRqkifjViW2F6UYwekZJooXhK/tcUhHEAib4g+RpDTf+xvGjWIPQ4MDzu9SjWz15uIZNdYbW
iqmNjy8dW/FemSGeB4cGkbAH9wlqRSAgrGANyKLeAZaVJ+Zw18zzBrcr87EDiGzdaANg023ODRLa
yEN7MtfwdXZcrG8HcJbw5M15zvxxBulXMSrhb/Ev3FEbnpDCOPN4FZitsCkTg1N3ptKS/SIMUslN
F9RXTrnv+wJahGlNWWzOnOmM/MyqqoPnFprR2Of1cAYamSCsrUY8ZN4WN7NT5UMXRHT4QxP4Ak3N
EW6j0uANYThujvxUsTcfxg8e3LV4z1Ho/nFKa8C4DVLJ+leO0Tjm9VEYeoY3GfTgbdSOjfhKoyC/
ZtFFEIoMhdmSzfmamBkxgKpY1qDUfxA2dx9t9CRNL+XiiAkTON4GVhj6rxyYTsygWEYBWGa+gWmV
gLwvxiv5Ok6peXvunD1tweWXtr+y7IwPU1F754yA7EERt6AgGr+e/5jA3wQDQIQhestErestFCYU
BbYmeWc7zCzeKFZpWWMoHPaukw8mZ1YdaOgvNDg7vPn5lh/3ubwH/XNu8vDPnpAqT2s544SAS9TV
4Q9thJNQ9NNUcR86Kx6n57cTUddoiTy23WNLPYnsTE21P/uYyYmkadvFPhyXQ1wKNLFDBwJ9TPsY
AzDH2g0WyrFrdsIFjaNOHPPmwR6WZSGY4n1n4k13rnj3SWsmOvUKDdxq18npnD5W1HCKYL173DD5
l1OYwRIAlw7/MAppcfdo/wy6zS6QZIMheaTIyrPodV7VEPoRzuYyhVNUpxvN7Vl+nfHNtq8LBsVn
CmZ2Vg5lODxu6Fkpm5o8iGU6zbWb1b2jjJU4ifF4x3+IgQ2FRWXHpXOf+SUFMteb15gMBHsIfIKk
PcLPOwzSxd+fXFoaLghML8KU3wO1wG1PrQ8HTjP7acNFzhjRQMXYGMZvJhJEvK0n0ScSOSJwikea
5fJoCeer/eoKiQQiqRaGLmD0tOtF3bO8obCKs3vptEHoZwvrq0pQGVzuVucHfdKVZBAdvPTeiEtb
2V0cxSwGz95t57O7L3r3xkxWj1vHnpyM9Q2+8iItuq0G+liBgNUhPkZ+wlS/miagjAUwpZ7qWhyJ
G1RMs3d5QvhnDgXPKEjOVGrinH6hvmj57D3Ry1WjITs+KIQJhShTf0kpuuORLtGQ71YUHZntfGay
Al6fHtFIBwlInRbesoyP+WTGGZndSRrJGC6FV9jFbSs8oPrMNFTD5KmmCZHxjCX26Q2mKq5puIPv
N9sWy5IouYu4Hqut6mMrVW5Q0R5R5UV9t1/nExbkPB6CnAAeiSsODLSNzBzBgU9msdRbdnQ3O+zM
sEQyN0ruTAQPrO38pnIbxvTpo3e7shCqhhh+GyTMzNXT/dEdusmkNrVrcS31mU7oXtMVtUwnvDI5
9/6nwUYa+Clb8hFVdD0RWqDIiYJRuwdbn6SBBUMGKmLEMSJkczcSJjNNNBDCv1+4836t26M8SOop
Mh6Q4boF6MHW3f1qgZg/otNEPlEpiMueP4Jhtb/ZEs1Eu6Fa6rklQnImkEHMI/Cc674A2Acp0oE3
VzVfIUJq0cVZfJCj6UncRIeO84CMrhD22wC11KDtZlcLTrHhDriB4mlxK9cnIYgPddSzDhHcmTrc
J9lWK2eQG7ksydl3wKs+j6bX+VQmajxqT4QXDSWrF9iVfpTODuhNuidyXDjD4YVRvWPfs6Hq5QL2
PXA523HvB3cNlG80yH41TxlsUkCvBqjXxUHFj6LFNBqfycXmwgSLlWh2SM/WMBxC6mfP40bCuznL
P4AM4/KdfjfVjUdsrWyHBhYvAzAbmLXgccXtbt5hG++7pi7RYawUmt6o5Tfjy6KuMr0zXMASBbRL
VcmogTJJdR5blmm9QHcJ7p7ZcEIiYagHwrlhZpAsCsE0QCPvnVNq/9yIb1L29UmU9CyYG3CG3Lgk
XhVhEzHUyuVexCT28bCX340pAkQtljHqXiLLhgV/Hc/X1JvvxIRbkfVd+V4TLCeMg1IBziU1E13r
P6y19JIdWuSTNaEZk/8hHEnSiVV5++ayM0poaTkLkk4CsqKJA4rZGUgjzuLsHsBB7EzdaVV6nIIC
B+jmweEbh+bl62ndgiBTSU5V4ELzkLeJnCsY59ImRnAhvlHPX44f5j8cgnQIU6bcVyh3QVgBNchA
ff0rBt1JM0g1hAkM2QU2R3gYYUY/3KxLoclTv5X0eQTlir9jRHPVKEqw5pdIb+dzXWY4eNVXoX93
LoprgQjFYQBZdHpWn7YJy/B9MlVYlQ2Zb2wCQ4Iq1+Gfb9hiauhMXrU57VEGEPF0t07xpcpxY6x1
bBs/eUhRXCH0mKhGdpV5zBK+xOaFDME3+uZv8mbhDHpuTUG4vCsrL47K0VAWVw5f/e01Zh6ecVCP
5+E+kZ4XctPa9GgRmtsrxPNz/Jc1cTjG9CLZ3Vi9RJTvZeVRSbClLKVmeKFD8eJ3jMt2IzgRnodv
+U3A6igpxvGoX1weg6ETtNLfDVjooZ8+I3RGZRnNNHIVQR9j71YG3+i2qj8pa75+PxkejfG0nl8y
TDqb3F8AZxOA3+CR6dcNqEFIVbDyDUHRYnv5ZCGyo1AmBj+Jw+GFlDdn5X44TYnlPn8CtS28OgPq
9l7uyb0+P0lEKUhokKd7pwIcfpMIke9qvrWUXU4gJP2i6i+44HT6ES23Rq677OKor4UdJg3xGtKL
fjqVDZlPbZKJhJLRvO6EuSDPSVNEoX+Y/+Ch/po0ZDHa8QdeU5+f9UkUQGq4irSbN1byqDKR15Gm
7pIxS3oRMb4UvupBrXKp9NuEMcsTKxJO1Ze5851fZJBjNoVICH9rtx7jNv+oITn8s4l654d3otRB
UNUlYf5+UTK6GmH7chMOx16pJ1EI1tJY047q4u0o4Y3FXsrwaOOlfuM0zUEYpeeLby1w7MqNt4ik
YMxoKRXfrblL22uCBusVzqPaI4hffa5fLHdvmnGhE/56p0l3VVjG1YlGzDy1Tdhube50o+HYVzQk
sT4qmO6X0EHPrcxy4aIZw9cihDYUHn6N5GbEZP3wVPdKTL4XC6mkOOAiwqcAKbGVcg5x0id1KV3u
FPn4zV0VqPkoUp/CCUmAfUpCnyjZgp7zGOILzJtpYEaCjhPFrwhCwUXkPFW3bewAb6ZjPKZCSYH1
e2L1PsEVL7PQXsbTeVhfOzEepa8WD/Geoa2KOBKSXmSk1oNtJYCsvN4MWqEVMXZdg+Vng53JK8es
ZX8LlRz0iKx65WT8ehRUut7bPvAkddemX+5NRfcHGTZRZwPsOHdHT8DRe5UbeYMYPWnN1cvq3UxL
o3AN8xX8Iz4HNqWVoybUqM4/zeNE2taJKXro+AMa7jXqmimHMVdMyH1nBbPGMO2Cm7TSfoTSxGcJ
07ItlJVMdZGWVUlx3Eqm9sxJRvj8/XEFZ/81NthvyFlpZKquaB2iTZNrQhYO0J1YgGXW9gAN8Rt2
A5o4/0D6tL8ghF7NcmFgHhx3dhrGnPen/uQom/V+6gwLhngiyAdt0jRBwjXbdBBogxrIKVSV+j+P
vmtuSd/uB9Gt3vhZCueNs23Vgj21gd6EA1rmXjvyTuy1hpnAiGnlkPYlIldboMpH/Of9DtZKtFG9
nqHC8R7F7Pv44Z7KuIs6toKTmmhxQncM0J+hm9IKmHzlejIpD1eZ+BoGBY4l4SMgSYhmv0oVLsVL
s4qn6FV0BLl4V56JZ213NeppoJwFxlOrMPw2zqJxKpkFjgAS8c0tlitZB0B+yaFLCKjU015mxgCX
0bIllMG25E93mfuOWiZ1Sf2jRejyV6QgTIw3FZIf2g6Sjh2ewCOhHGKV7I4vDdiAw8qsKlETrhnQ
vOWVukFxvG/rXMzEtfj8emucBAik6DGacvOuS8KuyNryjNiqnaWBRT31rF8HhcGqFp5q8t+x9YQK
IlQ6ytwoWMqO28JUnqxyQ17CZhLNpcMHrTT2aT5gtK/YsBwrQpb4RNhvjr0CzT/DT75NjiU/cXZj
qkbCIchbP8aCLU1pEoGWjagqLHnlwzVwXvhvcyJK1KYPSemQ56I0+1/rO/Gt3HsN7lslIkwyhP25
eEB0PylW8kcLJauZkPxApjR/V10RaqNOO0gJpeZiIsdg4GIT70NZOk9NCcK/0zxvoBHcm2N+jjjT
qPMU4txY9VhG7vS6NzxugY1hY1LUQ+YHc1dvTXKyPB334/4BH0dhnvjyVwuLaYDLC38/ygh56plX
MODd8vdvM3UAQcfkgivnU+sgpvig2miUlXYJTCdmXcnw1XDMhK2J6bXlYTIah7J9ZmcZUPuq6qH8
xz3c/uDPIM2cgi+mpKVaCswN+sBLeF7ZVwSQLWvZlxz5b2TzM3+BuU+YqX5Fck3iUXI/KMMUFkXg
/oUs2pgMnwiROFBLWYbmB1AAYLC7zoVrsYOffIMBTQSY4/796bETemts1++1HiAKho8uR+4Ey5Wp
H/4TgSJLenvXuZvYkJ7abTwiECevZt0GUL7fM0zdGpTgKgIdW0muFf4ACb50TUqCV/ft1eb3htD/
sClH8AdU+CBOf+HFGx3GTBrHyvkgKXsb90gPkugwNFrankI9CsBQ+vkNLZroKPrLMB07r0txWqjf
lSTNQqMz48Kt9B853ddet9LNNZpbJ3tRduwLCFDr3PgKnv5tqsx1M5LcuH+URZAxP+XRRtRaJF/+
4njjUTr8D4cgZuXGS+E03aXzEhVEztQu7Uc7WpKMKUjcLEG0FHrOguL9q9IlO8f2acMjLp2u6qGg
myuiCid6FSltyy8ee6Gp/52ew4VSXqWBrB3epRXnSyfUIKGuX6Bl4wFrze6LIUiDgKPGp5DU8klo
mtji2TihbPtiLDzO5ZYGzGscLC6oeRgyrkm/o0xZjpT6pdb/wjJk5fC4NacJoonIfyo5gF78Zzyj
gz8G56bN2z4W1nV3DoyItVpQuUO8wN8c/x259IlRhOIa6UvdvY7U4JFP4PAH9lcELtlzRLbvBMkd
g5jExNtDfGg6P6WQ3ZtUtURy1OB9uvbMS2IW20TFZJ30DpAvBYsIZxrWtC93nXKexV5iT+VBjyws
o88ko5ofQRWDxND4zB8GZMgR6lVJvH0Sh3YAKKE4nxe9K1QXMrBKxk9l3OtZgvkURgSg6gOZ1RwA
1NM6L3BJ9vYKRtLqifQh8v27/azMbUhs8IR5C+60Fk7UAtjMu8zhNPJ6WgxyHLTHZLhVH8vG73XC
jh28GMZKiNkSzPo2ue6/9rmymUvWboOHVAohu5jPKAnaPCCzkCr0vcxuWNs7LM4qBG/w1uhvRYRU
ssHinmygl/grFnBrZuLGWGbjVAotYlvk8ZKu/zM5zr6GONbHrrdaH3xqBkp/ejPpD4cr6KBNECZu
leffuIAQuT5NfIIPsvYAJ+iQPD0Bc6OIFxyM22f8nKTieOqF0ByQrxz97GqmofV7KC3jiEzXpKlS
zVGKxgSt8sBK66SBlPq5CvsklgRSgf7h+v9VKiJnA6ukaOG51gtG7pt5nRU6jcK9f9gmg54hvmqn
/sAdQ8n+RcZqDUJjFpkEGYsaT42e6BVRYGcShv4GqVt26koYvK68TSfYPOD7ovAv2RHlnMnm43+h
l60qVSwVHT785CXeSEwTDW4FwnsP49O159d7h3AcodM23l2vYIywG9cjTqbPJFfsSnEXFXSlpgTl
0vfmP0WTo16EI9SoX8CtQqN/U8kyoBLAPchl/Vn8mt8f1EaSepBa1gyMlkZBbgRWVKRL7Cq1uAIE
ttd5FzmoLLbuONSfE+tnpEpiX2DWnrGD4QiVm87VHpDDsWwLEUeMDv0uuzhdKddSStacbsO+d0/t
0ovvIvc0QqAuHyOcL5etZ2Zds3BmWwcN9kpQP0YD4TFYv/vrM9eum2Nr9v0VcS+eKxFIauNKT+bF
D1YL6KNktbFPhDhPwxA/nMbDhA5Eog8WfKUpyx6wbwmex3D4muc5btlExVrAhceQyrDFkBlBJcWP
QY5aUfzFUjVTtPnBq/8X0N3TodaLUu60hX/ZwxGVWoH5OjbC8OhhNyZiBD+uzCuIxwG06xIGXwRD
Jd61+jOJqhbVweSvp+ifJieIYMZWjqI2V+yrpxTO7YIsIRQ1LSc4gdWOb8xu1xN6l+nZLNNBHyJn
GCxZ3tFinrnPxej2qhgDFBl3uGN3TixSgIthjezct1CnSpwsyqwT6xXi4CGUokTQwWEi5Ix52fwJ
Im36AUbj4oid1hzT5XITVVQ4urRNyOz2EpVYTKft1yxcXmiqoNFWCm5UYgS8oAA9WxDOnk9e0FVD
c6FkDEAKrIEV+q8gDVd8a8qOXL5ugLsNnQIU/Bz6JL5QxldbJskxDqhx/6HhpZTXVAWjuRRTP9Kd
ymOrlNdY4rm0BEiaELxQI/wdCUTzSpawxfevFKUmml3ZOcdPzQz1Td8psFCBecVZQ6tLedbpyqw2
hhqXnh4yMQu2wG4XGuf1WeLqlSmbP7Q/2/dI3T/AuH2s9GNyyL4YEiDAUGZoyzttZTf8fgpIKV9b
69eLJf+lZTDSW1glkQEYpdDCfj41sXpGKmhZZqzGv7WbS8iMBjbHDIM31ApN5wAu65EzOXKEEDIa
/svI6pSKCryxVzGP8vZ7FbEuIjXe6yFnSXCf1CeCJlBsYXsNjn+rcXHEc5XKaoo9qnn/CscUdz6l
O5j2+voT748v8A+lpWYeqvAMXlSbuFIcgORfyNSTPTNRu8F5+bdhEcWD9uoJG7ZZJ8Zbse7n1jyo
prLZEUG4olwFXpVjFOkenBbCJTrhCrYrYeTWfKWWxqnAjUowqN5Z5wZeHU0BpGASo6ItpUAGwral
+asvIMVLpXpxGX2r3O9uVHwcx5JIuCWy4ectOIcCzY7vUe80ZiEw1OtL9DmS9g0FXcafhuCb7bLE
Eeos7BrRAmyCT1QXf/rYjyX1burW6N90guuZ0ZbsXZ6wdbLJaPbtJ0i+Dgn8plDnfpo2MpUBJa0l
zTXbelt9knjcEVl2nU++jzKfz/NYEa1cHEk9Nc7u35SqFOdKsWN+MdZ2w14pooCHDJ2uI/Z51szc
ikAJKDYXvAc6rmA/CUOr7RBBEjIRUSqKry0EoGS7++1XkkOxdsbvc12Tx+7vTuQ4mZbp7RVl8yGT
1b9W0rT3GbD/7tSL0uDYiNTrZApkf4nAe6iqYNm92Q82x9arRrB/vabGuIG302C88xedIrK5guKa
JNAV4Hu8WM/hOj6K8Ne1INHG3F69cYHEREn12BlBZCMktdGNDXk1EAjmujrH/UjrhQ8EBe8pBUxn
CBGapM7XK+vUxEzjHEm8SNDPm7KwTAzY4AV1zuWGlA3ba2ZTiMzh8vIXBcjcUj8dkooitai29Krr
/8xPUQKaD4d/7lfETcoI0TaghSz+fm5Efx38IW+V+q7UOIUc7CyEs8YAcT30clNKVqTcJfVYh4XX
rDDZOAbJb60nita5Da422BVLucIM+1BrRl8K/p8IK60Z3lU/Y/Nqyo3JgowmMFamelORtUNQlrNv
mCqJhUHPR8YJZnSYuzKhHrJ9zHAjZwMg9G3B8Bq97uTmaAfN6623AW5eu5J1/aUhWY57VUSgY62N
OQEW9CAhI6MXRcurYo6c1ZIOARZO6J39Wt/zUw6gYlhES+JDK0VFc8iTBVPoRRdLGzb7nRSiBXWU
ar7w6/Kix3ap5PWQRuSPw7SS+fIsg0w355eaa5zkoJ1MkZiu/1PdLJWQ6UOSupqVsRWTaolW2kOh
7TI5a0o/tZYUxAT/hvKqxJkEGlKnRy3xHmwxFoE3INsqXoM5pGeqy6uwYTKvUZ+/TVT8B4pbMaC7
c6Sl8K+owQGQeMbZyUuyi9+D5NNEQiKcQy68J7anDcQOrSFFR+7uIzmKUOM+/xELQB1isQzCfbx4
HJoapnp1BQAvRruB0JDulL7dWFUY0KEzkn0Iz3QGrR/kFc+lfberMk8/8+5F+Kt/zU2Q4AFVAlU3
KPGgNHFkpzA1txH3FmfalpiVk2P8DwC6X3hUCi1MY2O6djiTmCJ4fQbsh7mSJnX2SIcpnkr+gcOU
UqExdTx5f64Kfz7HARZkZdksk/ozmO/Mrm8Nc0L1ZdSQecQGm+WJQBgrgBZ9dnmaOcljJqW/6HFZ
IRhIgwvrfji9f0fSLryTU0ESOlAa0GRwokqWEiUWh40Csx+VifxSVRBj8d4U+uKBgLdnrH8y0l0F
zacLRGn/yzdOHQEvypwdY9u6awEi4E93BWbtXzCViSsi+5lfpxK+sJei68NcMrb6MJdaFIPq+gnf
sI6N4m1KJrL3fs3fl0zbc+m+dJzScVuezx/XLDhIShWZV00+bBvGaHBczOvdUyzA8gg4M6IQO1AS
TpoOBA7Jxf6TB2uPni7WNepiXKIEyVHpvQRF9joYnckvI+VvfPFKjUUS7C179qj6HVxlS9KFNAR4
zQmYrNWot6oA5mgMww42boMntmbiYEZ8k9JJFqpNKszbqqLUnTZj61/d/PDQjIhsTRVq9SMVaFGz
1jY6OOmU5C1+eWrXigVTTqvEzRf6Z/euzSSpHeMWGOitVgNnj6q5xRMsJrAfVU0mMyyPPK+FYDqi
MgAm2kKSzsw+sqC6ovR8HRQoacvD8ok6OP+oVnUTBwKEMDO5cLjKLAtPU40YBCfttAd9271B4Trs
h9YZLIn7lRcPuHGC/9qK7VyqR1KqOTbDx4MPaqbf+XdapChj4qz1K3Hbic1gxdNaetZWa6G/FAVK
xp36btoKbDKmrmyufy/3NIs0Iz4SrNtt8t1HT4O1SHa9wvKbouu2IvMK1BYEQzu2+LYx/EuVoII0
sB4HBVTz0c45gJ6NJzFZbcqNmJAn2A+8lFOtkMWE4GXQtqUgLC7I4SYEJU+KHLF+8zqA2P/xIUAi
d6wb8QAehQ5zLwAOeXxrfTpPdiYIWBQZ3RELwOe+oQ24yFtrr9CVEjPkPRuzYux2C4keywnf8wYp
Uw3S+tol6pIPqJg/YrTyDUIF+g3+2A1b0wozBboLFfAOa9PlkzDl+EJ4PGrqnK+6qS2wy23Go6t5
ajmWySMHWsVzYFWAC8xzhAzVXCVoxWBiID4+xM6hx2vMbavduBArI6mhDI+Xne/EJfcsG0DmcvMg
eMV59hWGHgWhuPAQjA0Ug8Z+fP1Vvf1xigTnX+5T2z0BnxX8v9LDprQZVF/yiMzAt+1/tDbKUsdf
99ff30YnqZPgEqEojk74Q72HH3siyy9TNa8RRBQFTc6N2ac2ivfGjFZRFti+CJ6BHBfQLMc+dIry
IokkzzAhhIzJVIcGavdcte6b+IlaJulBdr7r+gzwnSCc/FfEuB7btRbQ/NmaB/6Y3ZsGOfMQ3M7J
77qCF+1rV4PSDHq/PheI50ggR4d4dR1/qcF3NiLR+DAjaLE84k9StRgnORMcEIt1wipI85YmFiyl
JD4C09JwZtfeewJUCrDZM9xkDQ2zbHrJeotqmD9/1h3LxgYFm5Csf3cFDF5UmQZff7jI4tK+ta4y
xjuXpRAKFYobcCjDxUz9tHOcQ4MI5Dt51tu1qlJy6BWbDgFBlmw+ZJQGKBK1JJydZDeifBVknGac
1woTVXELiwzjLUB7G3Hcl0vbC4QLn+inTMnriB5J6l/CZctPrxxLG8oGvkhf23JQzLr/bW3ww7Lb
+lWXnHXINz0M5SzgCJsV+QPu+3qRU3aI+Ndxu6rojcI0Aaji12RALV94UzwfKdIFHv1eI33QgAMW
OqVC3MLbDVPsEQpDP2+Gg6vlQXGc2BJZzgLz4BuDATL7Wa+sK3iWes58FBXD948jlOuyL61lCutj
6NQql7dE0rAWLUVe/Wjlmk5DvsmTGsgztGBHe/8EDGm5jZj5WeyIq4sU7T5UmXw+1W7MIpAXXTOc
BgPwqjDxGFqkVIXyigmLUcI+5E6mtStsmTdPg895B4eXzC0pDrq3bKo0DJTHymMUzQYen6fdWILJ
ZqHZFasjHRXVEP4p7wfYaMzT66rZbKO6bpUj0x6iCxZlG46XurmEmuqV2oWzK45PMVZrrTye+BNu
demJBQjDV6hAkrMozXgncW0qTLpO6L+BG44/o9C+CEgm0WaNyNS4LP2PizLyxpCbtbCGLJtvhftn
gr4q6gJfzKCvmuqW/MedUfKzS/GTg64AypJ4/aOm8zxW1YDJFbrDv+JN/vjJyA8koMoMRxHXIj5y
n06THhRoZzl/r+AYkjZvdcw191omeC5P7C69bhiwF6evvw2/saOv8QYHkcuoaBe7ujsvWFYgJkE9
dLWe1EBrChTrGVUeCACDEvmCajcpg32oVqpgwetxF971f0Q3StYL8xggr2UR/5s1yxMjKuxoFCQS
q6F2Ljxrv6/sr47E7ZTLXjQMxJQjI0fnltqZStUjDAL5Jg4YtvSfShgcDZlO0LSpkQRjNc9Yn+rG
qtco0aaUlo5VxqpV5yGq+Bh/M+f77hEoZJ5+n69H1++4CNfX8UVwo/bbTJ49fIoTqHT53qQWTFHX
SJXebLN0YVavJZ6wCYWK91v7yYLsRRWynVI+FNO5QZCilr181G4c9KepGMY3z2Fz3CGGcwbUtYf7
dGj7e3Ie14NIvvYYRBnpisf/NrHpDUEAZvSKxKxpdSRThKsAjz7t8h/g0SNK5l+0yjWCFleIL2uk
7CBrd9ROGvBi+Wgc7TxvF2xG2rgJB0k38BdsOaH+6tkEjNPSgKWLk1+Pmi6bW6UZnprwy3mVhW7M
UDJ2S3wx9ardRtKi00IE84P6pHu1e6O0AcXCgT7UAS/0TZLR9vrJnMJg7PdEOSr3z6lNBgfLVfzo
DwUJgg53NYErh5q2WAqzVDkKed8PIC8m7QEYyJHMR3nrYAqMm7Yq7cdfWpDClcNU9NLSIUTJmnIJ
opRmegxev2HszqzYBEq3Wh7oIODdX9QK6WCLowS5i/bf0Dvcc/ltemZld9EImCCJ9A466682GmHg
TFo7gqwP7/gzv7ZWSpbfoSm54YP6RWtYe+0f1kXoSdHU1Ky7SQNi31jNLafk6NVjywYsNYh1Gi0k
l5ri0pQs/o6udjTbxRDe71QUouV9nmrsvxweYvarvN+Ya26HciULPpQdH5kQ8p5lT8pt1RbxHJZS
mksZaK5qjsyicEi7L3RrQpcuXZfDD4B2qXoq3V6QRwmBflmyyU1Hi30gTvO5hajhWMTUkcntMT7e
K2KPaiM196mzBGPN72iLRogQA0F8BjzA653M7/hxS01sRwJismwaqY/E9iFCVYFDbX9jZ5Vf2GLj
I7rB8k7rz02y4qcWEo92d0274cG043yToZFG2Q8US6TeZXcf7zh4u8tvDVNGZ++RL42MznGsutc7
0JzkDa1IEmUm98S2YmpMowNnpcKteMeR95CSYAHDnP7N2CA/cAgb6gta7rz9yJsIXmmnVOJETlmw
UpCdA/6yVDh4hRokLCA86aYTmuJ3t3xvnwXhpneEOOvA2qjMSmxB1M6uGtQb07ilKvt/x4vpBJ55
XQ0E15jY2WvdeUx+Fp2XTn6YYh3jgNpbWGEiTwa0eys04n27igUXsR1tchrXDrfbGD9lt+GqJmK9
FXwebcZqx22DcPQUgRO43V6sLJren1u6H6ZzvYbnnUHK/8m4UWNr6G18tiNPFBQ5b5geGBCTTBzc
oNGDia24GCj/L+hGoC55GBUxJeGLTF48vtdG1uPIwg0ueke1VkJsgjZYsY99LzJNlb1hYHEORg0A
bgjRed9UiLbUGQbuQxwK84ehgmvfikU/u3CEKdz1G+Zf+J1XafKTgXV8kT7M0mL1mYYBA2ZU1Fq5
7VC91fsPRuOabkdgZQsMASDmX21YXQiALlNCdyRU0ECayCXLFjlRJQ55bYApJNwmc9yoRb6St6G5
rQTD/930Al5h64jrDy3izHMNcXGRcRfCNal/b84cN3gq6K2esXluMetMBmUgA+BnOZglf2NyfvBH
RrGvpCXA35laGxTJoCGaAAshqDxqut+edaChO1oJIJmEcQEyZtijY8VC0KJRPi+GjmsJpnWOAPkb
YkdtXyNKdjMun4ndK6A7cRktuRiJtHE8tpataCWQts0OLOQO9PCf8JvJRtapnNv5HqTnyuOrtMU2
Rk8aQcgBB4mKztlm4r2lURfPDlrbm552p9vHNcSf7As535id0JR40MWadL6f1M9YCE2iVdXFQvgR
98eg3rMSstEc3Twxe0CsWvFuhWwa2nNSGgWgm/ZMTYEus8ADFUevyKANJLJCrgiaoWEhJ4VkbsvL
DiRTiREYMfB2DBlbgvn3+N4dcPQ38ylQ4YCDiL4Zaqp4EZiCpFfh8VI9TP7Qky2fk+nymwBKP2of
o8Uo29LMNe81fXbo66glfJD89R1NUvd2ssrctwPXdBJXb950bPlRWh3GUbMAFgSjiXxPuxXOOlR0
wrHw3W8XdVH7ZqEjhy5JmKN8KhkEF5RLV9ISKheLKUhFJ5aSv2YyCTRaXOZ43wQ/V3aeTSKwzg+6
vqwrcoEiY0vOs9fXhVkG0zZspcR46Go1YOh4ugaVujQemchA5Bn/gKim5d8JRqmnYlWXFaiin9DN
PkGcUOE2Vkz8RmsjznMdPB2WzMED+GQa1xGzn6ZGSyiFgFrKDOwxME7h25N/IydSiWHBs9uNjn/5
X5eeR9EdNRlS7EWdb6v+Ct6uYLPdfSsVClg33iwsaA+tObrAFThMGzC974mdHBgKR7cRb6oroWfs
rY0bEQYL+Z+j3327H4Mv3zZWDZo586Zo0CipgBnCt6TvdyP+AZN0aug+p9EmbaGQ5V+8Z+zY71gk
8YEaVluumUjbYOugUcGbnWa6pq/GFN2sDxi5jlmZmTm3Of4G1JZUkGQSqJXZR29WHYRBH4O7Ecjv
o7+3GgHYaHz+lHv2OV8nKY6feFjr1YBUq5AbqcB+6uKlpe+kbth2MPLorqM9oagKf54osRT7ALTW
0m8aX94NKL7fwCphKZzsDdRiGjn1WZsxPDk+wN7XrpdbxMxz8CNQT5IMcz0LEbZMQSc7Ey14NO2j
3cTkwDb8vqwL2uBg8+1i7cfIz2sK4475TZoNirN9PP/A6ZUW+CQyQRpl2IMNZGv8dVUcGdmEA4fT
Ul+G6TRlDPYp8jeGfDhGstuYNULAGGuDopg4tH5TgGLlPYwKkS1UBA2z9YShZJQlfhXIkz1z1hvl
DO+5np/jJ9BvX4Qu2LpYP26CcS/g85KhFV6Z2mJfBjL+w27oAz/nPXLE/Q0uyHIX0PMWEhBrzzLL
V9TLFsF29iRGhhanYhOG5RsAhCZhRV9g/bPzzbjG2sYhonpFB1jFy4EnGUne7XkI6QtvfAL97/zw
EVrCJ9frQv/iY5Huz8CC50R4K/CiTGRxG4HVsWEEH0RYqjWNBb+kpXhkBDVbCNJGlQPygUpB9Tj4
1/Yr+GZaBOymf3il2yxs8c6CVigfwq8TjvC1tCLEaL59IfR1tJ7OLkAvics12XXhC3tr+UfvD/UQ
TZzVrpzZ+eK0JkUjCXJAiSXrS7kpxZ3XZ5t47IET7YCgeOH1rVisZEST0VbBPiAv5E2NgvzRMKP5
4qMYx9P61kbckfNV4StWdw/kRSFlODp/VlqDDdbdZOVdSvhDXY4vY+7qz7TLrUZIctUc4oXZdvuN
Ct/gF440IXAESSawJz0ujVmXAqctyjtNT6IvvnaCfS70dUNjnvJd+GKiPQjWFLO4pqtJoxiPYRGD
LlGGxyB4tL5il0PowF3/WNYN9rlga03OdQpRQu4WnX5QQbxZvmJ05+I2HmK6HETTTOhe+fdrEYKc
HjxzHbc/aheNcRBBm59zGAt5aiQLp6B/pk3lx/zniHAfDsklvlwYsVGNgKwXj/JQJfcxwdvq6+z3
GZrIEnA2dwP65oFdklXph1kliv+Ne4QWi/zWRnLfpyY1w97LcizBjhmInMdHCfrVVx0MMIdtSYst
dN49SW7yHUgrW1LdRAZ6ewXnmBgAbdqa2ftY1kOhDVstPOPD/li4Uji4kjroTChCvrdD1Y/I4djU
4qVH9Qpo74dd86t62o/uPIkFxuOqsEnStS5eehXEw6p/wtmraxC0mEK07x5UpKylJsTzy2xLJRtU
dyBcQBfGtj8tsi/OlgAWowk5gwsqh+Iim15VlcdW9WvKvp2VPpRDGXFmz1v6KHu3CBNiczg7BJWW
JnLadsRwBSqo3bzDNsjov5eDI/9pyCMzAqDRiUi72Fbbg1rljfBujEX6JCvkiFgZPAwFiiBSGOPO
hhLxSTmbzCT65XdsKCC669LLCaeTxQj/8GaFWtEQk1+ActhNQpETbWtYblKqW5/6rrT7jr71ulXR
BRKbaaYp/s0HHnEmK3TLc++ljQBVUMbgBoylqELk+XlUYFThZVt0XriTB8ZKwsQeQyIi9NFsYAA/
/H215qLEvSOLEHwePJF4T3W3FqlW4FvBAH/OcZH28ekz+WjU+gFas+6NwKYM48IA7F+k9W30JZIf
tVw83wwrmJmcalyWMLRUzphJBsk1D4QfqJMllOd3Ah01mQK8pLc9HCyKwBIx56B18Qe797qeutDt
ZBVO0NfvFbbQnW1KSsRVcEvp7ewMhfTwbIWBMzzEYQNLbJhWEMIhqybK0PfgxPN6mpjyVmMfvYcR
AaGNK6U1Lsy4Kyd7bRlreho4HZZGUi3UtXJJ9GYH0C9qyAEYbcEnpFjVqylgjT5Sffhc2HxRs8vp
tW2iyvP5RejUkBap05dEj2C9397n3ohxlcDt6brjdcXCfNez6K5dHBKbnZaw61OgSHd1kG1NPTP3
FVboO5y9D/Q0l7NFDufi1NEL1RH/hwvr0Jzox0EjmeKUm70boqWNBfx+C5R0x928eig/PKYWhV6z
2nfdwMWmw41rrus1tbfe8QmmiB0ilrpVuyIX6G7AIdYXfnK/vKcU32jsWMnZPTMyBQYjSBUmaHik
jh0ixmUJdGU9CAG13SQIv5TJU2Mp1skTeEidIbFQacT5pZ2FYD5eBvoZgcNli6LuShSsu+Qles5Q
aa4TQ7GgrlrhqtceNhfW+1ub9uJbfOH1p6pB9SqNZyUmBsFLZLAn2x/WxuyB9YHQSca3XHg8q3/h
gAOO5qWEKidT1QCksU611BnoGiu2b8WovtfZ72fPaYfMmeEb7b8NJGvcT0wJDeOoB8Hzx0hX0/q3
XBqOJiKt/dNLd7DMmqvUHqQSRRjCZEUPWwWh2sDr28TFB8Zw+9lkRPKaJn+jA1LdDsHqnqsjsRSR
+6lz+4z/i3teh4sCUC6f5VDoqrPyTB/hw4mE0+GgoLB/PTAVx0pFlzc4/MjO+n0zbQJkYD8Se9J/
MTD7kk1BVg40UP1KtO4vryYSAj+XdpK6CcWMeCUhDEqLggiWlm+IffI6ctuYesLnu63qTK0b3FrG
i5ZgmmJalgORhd/ZbKjA+WqglieCQhgWxxoraJ/pgVM1VjXcpLzVweb6k0gmondXkOhrF6Xc8zKs
PhZXtoRwIG7o2G6Fi/Grsgxk7/ZdaIzn+9hX9WHafhZq1xFlGFw4GvUXwoycoeog2TQqVpr++QTd
2mhApNuMFEUM2UvFGTBEuAq0AecL+aVZlAysBYHjAzgIJltJ///YQzqc8gMa2jMDw11GGdLPQc3w
13TkALIgWlRs6cPcZtE+hs9kz7MlyyOhWsdRKt2n+x1Wee40s1TpMF6/+d3ZcE+n0Zpqnid3+Bae
Hf6xF58mBvH318gacqApVCF1VJp8CO39Yz7Hm7imccbmax/2J5EBlAUjE2HAKheHcmbVpbF4UjRb
btHbvFdHKyJ1XvhTqQmeeAbKWPbihX/hH7G+64MkBET3i2FIWyLaoitGVR7p16klxbh9UuKI5KfF
9Aaj0GTowPAxnzWtINRrTVH8WYLBzy6USe41q7QadRuAGUsOyzg1ZLXm3yhMgi8d9N9dtlp1JbIl
yVp+kNGiKIMvLImtmca2FSzBu1XK/bsoOvn/AVyohojDW79O8vDemGgRfwf+7Kh60Du/o0S7mM6R
yzXTmbUf7msAvCgDKg0PA3dNeb1YInyHhYTbZ5oRnd9kVASEO02dzhyV3lAnWF88LgK3q5Oswhj1
3YaDnFUlUrp6yC2J5ZjrQP/KtGcOpSrc/B3vVFYXDk0KlxnsXK6+nT8ZuVNfJV6X/2qleMpi47Zf
+imbEMXQseyJDoqT34hB1vQDBhkRBFLi7h3OHWYn3sCWbLTWRf5L9Gcfg3tmKeCfPd8v1eopDes+
ey8gIpqPVfzM4A5/8oqTTfFZtPrSxLTjBHR+jV7QxATXnwL9Xposom0lq3ClOBvtBOXuRlSFn/fj
BvbcELwcBSt/dgLImfNT8mw9NnggpNutzlft9snC0yONoBeFFLw09hdlzWnhFWmR8th2l7mQP18t
gT+n/ItT7I0NVgAtXNoYWAIFnhLjDfvIcBou8azGxF2DxqVKuoQke9vetFk77SzReeofH2GjYSTn
Tg53NvyBJTwu5fRlqKoGAWAmB/SHdGRWIUlVGZ/z5z7IYVyI8hI5a/xItO6ah4BcHAgpbNa2c5vj
c3grg7b+8Tjs61ZhBv+Bw0rgQITXUUwprW3y0BOhGgbuhc/JOww01Ova5rYZPCpo0jPkbZGj3Ja/
vF7XN3jqiJEVQ/tLsBXaNYysS3hy2Xz+zgbQ6Nr3gpLLdkJm+Tbw/OJMmtEFwxuIflHf2WLOveOS
9PxARGed8HltXp+vbFpNpNgRTeKQtA0pgakXt0Vfp0eMT39rTVlRsegdCqM2drHhTIQfczuI6PpQ
sf9kvyMP8zAxvDFPPwocYKvxoKr3NGkG0U7tn4yvx1sSMeYZcuc0zrHcff6WaLpkDEW0EV7oVSyD
7A7ETzA6nRQCUva1augyIdQftP/Z1hxE7PW8u1Ii5zBp9GUal5hQf1olqsp97LIA7x6WQxCSFOz6
oNj7vpQ6oWyOkOZIq4//ev8L7EjC2j/6laN5BYgVUQ0staJioAWick1dkLvZ2lBhDbaJb112VNs4
CH12tJS5JoVO2LdLB3AhHigXzmaJkdHcMb3t1ShIm3zB2QHRPAvoBc4BXaktYWo8Ayj6V7Qei6RK
NigkLULYzrQ/f63Ic5MU1hX3aBgEuP5aq0In7SYLstYfjyzPYq1YgNFPJxJRUOaT4Rt8iWaUUF0y
M/TzsTduva8CiTkV8g8mJeDZnk7UCCbhXudHiCNv8oUo0oBDSapRpoF2zwYgTmCNhT+Aycapcpmm
EhbSVwUmfpxD3Qzi3ytoE88vtbovVAOcbRKcpl1JdP2HyFez4S1qZFcELLpv9aprk+C/fHFtf4Jo
atImgu6/6fa13SJodnrRi31eKTmkHLAgsSk3bfbK/xlEAEXpjuU5Wjim89sXUTBiMb/eKc1gwJP2
yqTRMwsHX6o8vluf+O51gwQF+RCxUhql8hO0t8uocGfwz2cuaUb/vBpVTjQXfYHP23/noI5J0QDN
unCwF/mBP4O+UcOVhp4Zp74BJ4YpdjMOJxaU57URNQJk+zyRGJnT5cGsUt+GMiRs3nzIPXO52vcP
ihEKTLpLZB+UJtOltLfmSNTi4wOnjGmSQN7ps+zE4ZpC4JxVmwIVjW2TWk3II1kiBmXaWEirLGDB
BdhCUxEkLJGmMiQf3H2HwnuPiQgdVm/dDWP8FOUIz6QvDstXbBR1DIVJKeIcbx7ko37bMnnPN/Pa
5ZbdO1wzWH64m5HZDyH1F4+FF45UOVSmpweq8atFDrJledJsreT2l0Rbx4DLKMllA884JsOiATJB
2ADGAHK8P6WB5WO72rX6c8hIRmOpZyKmFcrReH24zg/Z2RgYqg5sMd8Sas0Z4wl9kuGc3fUUf/Fq
B6YnJHA+en7wTOXX73VF8OSJwpHe7xQqkujPl2zL8FX4KaqwT6ASkiaUDoNEe9C+UQeedK1J9lwM
xOy0nAs/F+Vj8PFjgVHWoIrUelt0K7BcCLrFB9C5lvwo2CDrCKiZbonC05rWGdxYybNrLyCNU2Kv
1h4tWfRtbtcSrU0wbiOoJ8tmJeysXA+O8aWsFNQvcyLYQnguWrSxVYZKk3PMhSI4geeDNOHKNJvr
GNPu+rZlW9rAUA1qoXuN8UVD7OiJOy8h8oIrNqB1uzbabRESypnOxEOD/NbO4cQJqpzD1dZv+MQG
aDWpJ+3wAJmXoGfi7LQpLkhNEkVLmwQujsD5ya5HIzMx53DOKtFXKkev3drbmuWwOxBlJs2l2wOp
tHwdOLJHI341lu2/bkJv1f0QTCYTxuRqNbQdHq6E4B09E6WJvBgkz656AtXvI9B0IVEG99EbE71V
a73ULatdhJ6w/km4c1rjLf8np5XrUUuCcPaGvu/Z7isIPGNyhg7fgraKlNNwqF4yujFOXIFfSW8f
gutHCtHoPtPXRE/D2/H+Qes73Xf5HynZfWlzDEfFvZ2+xuzRRe66b5GNJ9NtamPJY2DMeH1aQ+iN
Oea1q8z+snF6gP09fY7UubnXGu22ic6YvwNbbzI2d4K3BKKeU8qwT5Yg8Ky63D03nDBLYUvQEe35
Pyk+DANpMvhBgb7fuqRsFXpKfIa7TFhiL/3dlEqVpQ/Ssn9+E8fM41JUudzCuAS9kivJC0IDNgl+
FlbqN1Xu/Yd+lxj7FFJWS2i3+KnOIeer0UtlTfLmwKUoELfKg/i7+5uqubynoxhgW78LRKKLIXai
Bt+aNJmZJxXrffyjXxy4tfPehdeh061OZszjUA5vkf16Qyvi9S5XAI9xPYv32XJcpRB3Pbem4QlH
aArfKAetk8d6OpkrFmo5zArmKpt8nr+Sjt8pdx5BwIAuwlGvHmksVKQpTtGpEHoBDLn3w+jUvcOm
yQFDurMMh2tChp8yFw3n5fzasmRNKTP8wtN1PpHbbmbenUIhC89AFIFlLCTBaXXHWeZNNYd5lQfu
7rFb6OR4b2hd/0adwwJpjAE1qZShVsJJX3CnqYSGb5l/7SBGglVhYuO46TnahqgzqdQZ9A8JpANo
ESiARh5kGjGfpYtSJmlTfvE3/ViD07/XLy22ANBiLLayYALVwLadWZOFy1NpyujNMPbr1fKnqsum
2tf96KD0dUNVaZZKkuEc0LVy5Lfuh5yNcA9lVkO0kOXPIsjWfQQxg5p5NFQpBJhcIXlG21x3cMGr
qs3uDco5fOUb3U4QTije0oIi2I9g+G08R8ftsGR9J9RXM+DsquOKk4NSivrzckXL1grzu+y3gdOm
OWnrGtrGp9hINJlUn9MokQitP6djn4wg9OHIsur+LpvPSmNOKAMemwa6m3SL8av1bAOL7TeptARb
1ljNnBcFKBpRw1uGHJzLdWv2w2EukBFO3/zJYu9eACGAgDxBl/TCoUSW57rN1jFe0WST7876mWmJ
odzFiC/B9JChmOUvd4oOcLmWn5F0MUjZ0tPEkIlYLr6Y9kPwXy5sCPEkc8VNb9Yu2Ce2f8qlBAiC
wZFqOQ6Q8zrKxi2eaBLAHl7o64jchNy4FkEV/ogK/PKZTuRdiJ6QMDNH/YstuhSaGLGh17QH+o9P
Jf8/Du0xMa8yWElxs5UNwTBkvW8hzHh3cqI70qUSqgx6CUfPgPlks+8Lh0OQ3kUmwMzOMv/3xA8/
qPZNCLzRDrH/j2KeIiMhpy/osaKTynqhb/o7Eu0R4kKmVVD2fOdGHkDqLreLaBs0S+W/nf47WoJS
9LUQxshtqwaYRZK4UCt1WE8T5jcaLhutjUepf3yN/zojSGLqszE/eSrju9hdyHcFwwZW5mV2ltLd
cECWIJNumoSs9BAbiujY6r/yCnu4y8boGuj9nnRL3RyCRa/p+r6dzN9fnYEm30K+SEtPmuikTMBb
eAP6EY63Z7cl3cSeYh3ajQumnzVu5ZsWgvsrVkh6bJoHBR3G4jytcXgYopWnkn4ufCMOgs39+ker
k0Rb1iovetsfjl6INq5Qh98nvytebARcOWm+RRt3L5x5hMCLYqoyH/ERvFlrO5+I4Re80cjmePiH
KyR+ASxlK8ejsFy4Trrkhg04VnNgs6x7bT2ZIQRAXcBDql078gi3JapFvdyrpdiJuIupoQuGbGNY
o+OIVzjQrvlzAAYRJXd8pAUfq+Qr3jJIaZdJJcmtM6wdP56U+rsNDuCB1ewYWLP2ndLA6Aanj+zA
viJpfAfe+nIyUakY/CLTv2AFzxjcGxqZ17BKCmg2LrjposFLnpihdtK7RUk5bVVixbRp86xyCsOd
xcFnbgkC0Un9eW1kpyxzBV+OdholJWpPPjHFuL95TJv9qqqj1yd1HVlDDWaqap2eF2qOCC+9Pu12
RBZr8fBzjK5ok1OltapRD4r0xyCke9lUnk4aGK0/BPs70C3PCPsIxLgKPzv300JT0iDi/Mgzta6x
usLQMJhRFrf1oif/gKVEjguZ0L4QSLsjlrOn7LrLwnHJ3oGX2gaJsouLwSAlCFWAugr1ZRBfm3Oo
Jk+kQwFcu2IwoJ7FX/iIXS9LK4dwYDP7IaOULvIipkN41EaxlYHUq7t0JH6s2EXJJ2G1ke/KpeNJ
aoX8vmmLrZE9gnmYC0WE5U8L4MaRtvVqxhBKe6avnCHiWo6gOREjF35wwXS5V3GacvE/bNuXGHfj
RxMzv+PUNWxPdo1JzlvnXOpLiAbYnFSnbqV2l0pgV7aItpRt2bzczoo3PJF3Plh2Cgd3UexBNvvO
i2bVBc86B73VPzzegUFdMLrpdmydYdh0+JW/SyfTFAJA83uQP1t9+/0M1sroooHGyDluDqQINum8
brA6QjREoGcknDeeZ0D+y3RSDwblXVGLy28VC3aeKgrRYTy5CkQyrnJMGWi5FDEN+zgnyaCF2m/o
ZW7xfsheepdmwWKvdbuX9tu5fdjxt4xGd9ktsSF1dZAq5Bh+IKxfh0sDNByVs7e8aaRquMJiccN9
fPYh0xKkEBBYE3f6gZZvrZrcfLTZqB//j1VhtgSxE8yUWIljYD7l8cchxxleZCIRWtO7jXU9bSbK
H11CmqD0kM6syaokCLnVTUY7SBNxMpRHIUCYq62d4+bqB2tB1N+MLDL1Vrk38Ghzc4EnOq1qsPmM
w87gwvyAXkGa+72EFsyrNyqVHwT9YOj7TC1XUJuoGMF3EHIF7IesllrMTSTMQgvxbKsdGusuj7Ie
1+QL/npefFMmdzL1VMo/1Jk8uAMH2atz5m5uQRonji64vTlSPxHlPiyvdlEkikmlwcC223yeU7Zc
Tuqn2J8L/sATwJofC5XodC7rLRSJPUOAgPmbVkk8IQH7qOEZYq3Z425y4VpA7EENZKyY21gLOT6U
3jM3wRun7gKrp4Nyimu8bqHws8v6pE9AZMoLzLKlQolPZThfM7b6Ioxygll+8j5eYd4+XnbHU1K8
JZ/75xTZ4m5wEeEqduGOFLuBj8s2IJMg8kHkGyic9Rq8cnBVIJjzrf4H8AwRJQs1s4WsgnwC0aiv
ZT8D28kd9zDdN4JuX3idQpmaCDeDdtI2Gt6hJPQh56lw0p3S0zQSu95TsJQrfomdh9gC6h8PCS6L
cuUY0APZXyJcQUH95rhvSLHbv/eBhjXg9LVJVbH+c9zwBNhNWmAGEiZdkBZfuc7mix8ZI0pLgU3e
nDM8Zyy1bXDNfYuVE+CVQal+rBG/TXofwqnlLkjHkXcSEBwQeKVmKqtA1Fu/SyOPX0MuoCrgGOgY
0cNg8dGCIIWwXvwrsU05oiNyuGroAWGYF3VzxqSpSce2AU5k8VC3mZmwa69HLTsfXVP3wz8vxHwX
zYrQBwRzsq8v9LhAAj6Q2smVgL34vpqUwh0MLx/sRjeF1llpxGttCXZ0jLzz40TobtI2nGgodzoR
YkdTIDEx6tscYUXIy+SS8YrrdhgBWaJVHBNInDS7efvwwNa8gRggjW3b5q/TXbLJKcK0WRxHXnsF
K9LbYJ75LqdehwmvCP3NFv2bGRPLw7Jl9mwdtATbDEvjRcMwjdJoDmQFnT96MoLcQvz4CV6porhE
E1bkwx+94RSmTP9wxjqZAkQPUIXNE4kuoAK6mbLrBn7EkI1EtLVFRGkr+YnT0DSTfODRefloG9PY
szOWcNTxyfN20W5jvaVFB6TMDqgOm4zXpl0wrzrSjeCYh0t8WNBiVBTwf1kmNEKT9dcZVRhESQ86
K9zbczw3DsU1trnC2UUPhf2JsobrbL+1ugRcIws2/9r0/4fHEdW/qohAkFOsEGEgQWAUScNvKpVk
8jf7jYQz2KDDFnvcuVAgu+RFoieKftMlUMmw3ZqG7N40wfO6WoRTjxQDAGLn+C2kp5dLoonxFQGR
KffsbWSDbJ8W++3UlwtlsqQhNKw8J5J4Jek4tbU+HYQvyHZRnI/EuHfANrywvHbeUtG/7o5rxW1/
V4Z1SguBuqkn8YWBHRrlScoRCsy4pQHz2Q2QsvxHgst8dNpx2FgQUo58XK3/VrZ0T8ww7wckwGRA
KCDpzssbEmvvuFkERz8jqB6m1RGGkFE5s1Sw4JBrzDgC4DewgvWCFjzb/rt3sga4IjU3a/N5a3WD
oosU2bwsmbHBIKaQ+fLOS+EVFlI2/tDtLFMm6MsO+ZAEb4rxCQRy0Ni5X1cnPED2s+ucYG5d8Q4v
qwsn+fOybHwdboTRctiEwJljAj6HGPt/I50qp8G+XYduF0xhcUAit8YKcHl/3dUEslgVjLXKxlHW
I4wHEL8T+SHu5f7c8JpxpP31ppyJyCBoQchTmxqVk9gWb1rXGJbXe09UBk9UuHUTOACnwOXsoFcY
FJljmYLKV+Y0Ah8oUuQ9+mgstfdVd6+OVzyg9WLIcMf5rSPYoy7Gi9GRpHkmbm93UNqgUhG53A4t
sUwDTAt071i2bfq841bk29TkwKQGQR8AR0l3KEEp27PIrPNY5GWz29fEVwfYtyYgJAXPJXpo9jh7
1pR4c3eKCDBbWSxEQtyT/8s/8QfZXSgQoDM8PaikLPB2MMh9J7KNzRWoMUXu0S9RWpCsKGq2I1V7
gf/SKRsVsR+pAiU+KKrGUJS51VbwIO2yLAm/TXU+FYzkV6Uh1bR1irkX3Coxe449jbL5FdLE0G+z
A2zJ+lTPCsqRaFzAF/6vfBpm64uPKfXZXRZAewURrMCecZxcfZCvAOzIJUKLGFpEVvE+agsoccwO
R1FlytCF0xv114M/x6wbYR4tD/Gq0PGae6b7w9+BOKP69+BTILovBTA7NK0mSLosWbmL2rypgj6n
uV3xGtNMYaZmXtpCsOCgxL0CGBbiF4WkFP8FJVAy8nbOBTO2hBsLNj55vv/vyBGaQzXXH1H09gSt
gGTP5MazaIwkmhJJ0W/HSUp7xZxs53VuTyqN+oJuY/3bwWlljpfJPXxQTnn9ohTDrf/aHaF8hRmR
SRHOf7LEob+nblzrmXTSFo3JxfiF3vikvAJJU8W7eEicYmyB3hqOLRQ0oU10AroXwKKO6Ndg0WSq
RHsHBCMVgeC1U+xAC8lpNezqiAMn2Hi0kxy9sgPvrWofwdpQxlJk41RdJ4E7kxQZMmZjBTNLMn4T
KlatyrGBRsKWWOHyWs7gE8peXZfmeHD1JtNRxbkK2UyndKVDoFuLaR3qxiLdZIORPTvHDXSGNep3
cB7+3jBZgu2+QKYd1MqrfgF9NJj4/R81jremxsMNtEgIwfjV9n18R2myf1CbwsqcovaHdPDVkdT5
EhjkUCjavi6RabzLUAXLv8IpH8BeTZ4x/sqKIpLNZ9kJNw4TX7fMSTcbE482P63DQCf1J7A5vFhK
fxDXHNWBQKMLzSakUwzZbnq/9+pGtQdm3zC3eHwquqbFONHlJ6iPDrjqMYrBxEDlGW7szAsMaEbp
9lakm+oWdu8lfi2aazkJBd6TIYR7H7P+Hp78Pgp1UhokddayuZ102gTjr3+EazW+w+IAcLjhiImL
RI6NvWrtcVO8CA3HE8PsTHcFDxgg8m1vSJxMt7+LAltNLtvJsi3vAgtVdfPzMjdn8SeypI1PW+J9
tpMPU2ST/F/b3TKLDTYDhM6Ql7j4AOIbXX4HzVt2ZSkGxdjZ8u8p/tmgys9FFM/MSTpsX7YXqIlN
XKIDIyz/BuXmE4yS4G/ke+6D5WGaT228SXpasMzU5vrB/dKxO+JAbaSS5g+9DhO9P8fRHEriKpYw
4qEHtN4QPbit8+B6H6Gv76dBGTMAydx5Sq5gS8QKpcthO6s5tR83uWjzFqqsk/umoFRdgH8wryEK
2KRAWbODa9pNjq7prxbtPzA+774zb5+VWEZZs5mMBILAtq5TLSTx1LCUU1t0Ay4ce2SmJYdJXWhi
KB5yX/eXsDBYF5+f83aZgrjzBPO9//mpd7+SGtFyo687VirUM64iEOfmJjGLYWwJgrAu72N5Tq/+
HclF4SAG2Cfxej1vvByQ+L3wJ3zeXVLV1DfcjjyBWx8/WNARhqtZ6CXPu+JoCmc656AEAhrYc48y
7qamMRNn3pdMY+L9fxO7Y8SArMyRBlGtIHJDqi+pQmpLw5cmG43PrbW4biI4qzi9S6qs9sbd6Pgq
GPz4O6yK2GdH8vV/bWJJV+X6A6gvTZy2ndwx9zdNZc/fYF25U86Zf8bER723bskddyYZypN83Gvb
CChISbqFrmj0jTKqD1IWq1bhWu3+Y3+Gg7jhhjfqjKKrcYe8qIpWWCh13DVTFNpiW0Zkg07yhLwL
sbyMzxYlQJh8RVEWVgQxkeqX/b2WdrXhXtuKAAxZQe7lUQJXPPzWqmhl+kB+EzX6MZGEtDS2NBnG
YTeqfDpAYhBkSBvbG5jKEW1eVhHa23IVkHCX+AHWyNRjeYZnTAI7FY4+ckG7lTE+GGibS5S0h108
3lmtT1O3f80FVH+1aR5+ZpEIvmtU6YujoiNv9sIhX7BocGdqh5FFRawGW39T4BkcxlR6Ekshmqtg
XvWpopCT/s08M97sdTmth41W+fP2UN76QpBrMPZhM/61/jqvFpz+XTwOwOSYSpcVdmGAUDAhljlM
Er3VnXO3NhEgV9rRJ+u7XAJua/cwyq+zJZazkbuYm4ZolD0A+NXV6hCnC6bKAYHFLKIUEU6d5K6w
+7Vdm6ml7SLji3UuPmzd1JX33sx857NFBFEfIjy4+5x/rJVWbqqKiqA/nowdzQNj0eR3r7s+a87L
4Q5Nqx40Thdsia1pKPG0WO9s2N2f1MyQ9zNysf1+wxPHQkCn1r4/2xA46n3kVgRFWXsYurLzurUj
IfqMhCk754yetBdwfIu+Zbrk94DaDSKHE5Eudmf5VJ+U5ml2Ni82JN/WSquoiu34DmtIDn3anoQW
6LrOs08cyUcccb4wiAYfzIBYwrCLzYYHVoIoI9B/UH8zcJ/VM1Qwjj9ICp0P1eFSoxhG8mYwFgdu
Qh3YG+aJPG6Y5kq60MWFuhhStb7GwLx6CO6dITlUHg1lMWql0dJMaySBnOoTSo6K5rMFamlF1oGp
8JnbwSWihvkgfgVOY9nbzvyUaGO4JI8bWJiZR0w1cg2PRjRfKYkL0z73uA9Dg6pZbY35XyjDiXqN
WxfAc1xI7hZhIfSFb+IkFgEQDMu1vxu6kodsZwRtsajwktxVEaT/rUyuMlRpER0NGHXR++rr4WhR
6qWcCY80pVG08ETFCIk0sqFLuPoUje1nHlk/mvgzOKy2IXnyx8YuhuAAsK10MWxjCvbZ7nLLQzIa
eC85xwjCAiXecgwYpKjmCjnQAaLR3CUfAEtltWNX5y0EfG47zxV2kzSmkRYjatJNQkhhOhwROjRi
2cJsQW83wXlqI3D3SlaQvKsJTXSoisOEHGo3iNRN1UQnCBckB7gyBKNvAyZyI8HIKwJWxeUi88dx
BPYea+ML+A4TcsiGer7Ve9iPe2wmKUubGKLxDQsEgBbfTEa7pi4fYCEjTdDQw2FfJFNjP9FViGwG
Z1GmflJnX8RUIfsb8Pl911E1latRve30+iV4I4WgozbYEpR0k/zzrsKMyQN6lnZTCX2if+PvMvVe
KjH+Cta7hsSajGTXysWzamYyaSOg7OH0ZGkqCDKdOFUvJAfi8o6cAvpl3iYfq7pHnxMBvVSpxrD6
wNkW+F5E4tFEhjHEi/EKBC89heZwafAxoKGAHithi3vsJuRQMJOwkSbFcVxzZd4cddHSS5Xru020
ymY5xjkTWxvMeSJdZDctDsJ+3Hy+unEUPLOzPNHufkqKDYxoLDuu74hRBeDaeOtsgHeGhqfYF1Ki
5luSWQvA20Co8jHVB7ZRmNQ6F+BhqMW9gcRySqrQB0TOx6jLV1LDVkWwJcLjBoKM6czb3fnOsuUV
qIJmMCdkcCpUqdxgwxA5tfFUpAHESSVZloX8sDEuBqNjOg1CK0+aLLaTORQpXS/tkMSR1yDFb8kJ
vrTmYGHxYi2u6GZGPDOvlAGnW1cWCbiHoW6kKOozRN4bK44rCy0UAHi1krxKYPQYVanlpakdrTG9
s+VBC2pizZwETnexuq57lW6L6y6d4nLMou98dpPZP5As/R9iT0uqBn0x3zSyPNN1RmugpTf1aM3b
6zcpaQGfTv+o6P182XDDD8QXAdY2fSzZJGrx5PcGwhDVozg72au0uotLFCTD6eDT9J+2vNv2WySZ
bS/N/tzIMmdiMjPtOzYyHejkKOv1mgWj8hwUfiITKfMLrsqlFQM5QEi2K0Ql8vmUbTOdD+XNwcJn
S8iFgRVTaMokQQZmJaG3z48N69LMVXgVNSxKNndQIAoZdxfTamIZQGH5oj1ha6LyfeAKNaw8qw5m
liWuX+nHzyWNjfdk2dpmlpswkao1LH8Zz4OIuMAWn65dV20dWvgLUEjH8uqbo1F7ntktJXF/D6zf
A+SF3wZF9UrJ0TlKYEMMsgnZVhJxmeBZlaQPGF3U+5WQM1AV9FwlrBaeLxbAQC74jwQNpgdIlI7H
IuYsv/4ff+uKYIGputHm3LiTDdaj6noZ5HOKwy/TGqUbU37t1USaVbz0CV/8W4p5hMG5YqzVrMMw
f/Rte/EV9BInsvdCfvIctyuWPuUxnFWii0lH/8v4HZiVhzYWBoqTiRtLsPOgx8mRBmPyqbEOZcCr
P27sp1j5bcrhoQwLeYqMD8xn/gbNzxIM17B2LnGUMYNvDflzPLugBULxL2zz2amUQ9yDfyNnWSXu
euU7uczpf4FX1NKjFAtVATP4Sv/mLWIlLfIAeGGhdxmDLi6uUOr/IgucajtpLt1NkUU+LcXXk1Vr
lAxzfcmL4zp6lZv7l6XIsRxL3xj8gRypMLQ+RLGOzdxNRMBcHJ15bj6uzT8saXEy4sQUb3ah6QfR
TIbEco7c6caryAUDsINryHV8n7ymx6a7ATYpjlZ+rJwWCuR9NkX5KGnthBpHrluaW5KqCywgiPDH
Reo7yaL3TPIX1jehldjk0T73OuHvXg27iOuww2cAVdFUNxpDibm/Hn4rdG+wYUbODFiWvdjk6odW
km/75MqK9Nf963+uGTahWJJIrbbylITg9I6OAJkVZUaZPCjauxJQ+OBsibJslyX3LTiZXhbIi2sX
TjEIZrC2kTj6VSCAftzNLJlwjSnWjU+9g3+t8EM8FJ8Eo/UqeVIY1/D5O2MQ17QcHNBEPMuX4MeR
gSoCCFduOLaLSqTDU1d9JYulwhdYiWB2APIy5lVaOQoLoo17i++d9LGcUjV244nxqDAAe+TmO38U
chKStA87I+v4GMH+WoOvm5Uk1uCbk/GgOS9pTuKvakBC9H8vfyg6b5YHcL6xY+pY9chOUilTSjo6
yYcLRAJS6JphgqdAzzbCls3coIwCCD738E1iuJZTrJ87y5AkfC37EPNP6jmF1MEnXaIgAS4UGG3w
WL9CLpx/c9YUJkBuJO8aGqY6ZOFuelPxql0lwJ+WeEFyquJOYHwiK5HanaGs/7Va+otAow/sP0yI
YiOQHln6FvasyZQhxXHFnhvnUpyxzf4zvWVoKKgGCcEH/wjvGYTG89W3TLK2MbUMlTXFCNsKehtY
DYcY/LTIj+HerJKYqjqBL+0kpPgNMYTB4ep1HQAkRhH1KSldA/AeZdZgb8GuxTSBM5jfRMK6RMyX
HrzbNznyiOw5nEyAQYUHjiSDbp5pyagW/qI3uglBOcXtXy7TCJYFNfPNJaaLcVNR6Qz2EADfaYYT
8DXGJslAW092OY5K89GvgIjR18ADtD0KlijqGgz+EhNFJya5R28nr1i9yM+UuLFxNO56JvXnBat8
eydaAzXoWXD4gFGOucWqD++twQ1F6LJvYXhq+uPh9J02PPq1t6KmSI9Lwx/vXt960Rhk/LCGZqxd
tg3bfcuVUu8tcj7KG3C7gqswPpRnKdFLBJoTTFvKNkLEw+GQEjCViPLxYYlERdHPvMvHR2MibnPF
+3x70fEb0RmhL7Wvxkgn8m+7NCQSMHFUtvrPQ8xJnhDCfG+yLz10WZoWIcN+k9AoxSl+MYvJDXfm
u+UT574IXgV3cha0ypU4xC84lLkF7WwbsNg+kPn7Vy9is2+kQTcjAw73e/keubTPSvjEGvObmuXo
3UahtDEd5YN0mTPVY7MMNHC9bsB1rkXEmG5hgGKgl3onRXRmz7W8XxR1dGTdv9AzweIyhh9sPP4k
MRtWyt0tPHT/ApNChtj0ZiUMyTFRYqFlsJSnm4ZGzdY4AYdai0eD+fW9zvF7KY93nL4UBjhUxuiq
t+/8z8t3lX1ZjKHM9bnBgaRYYoqqsnt/iSRkAtLufa7rIHAuaPEorr/K24YRBLQn0mYFh9NP3fP2
tC8pDCyiKWVBO1X/Pd22y/6Kr8G8WJmmCUpVhe/4WwlFbJkQlCfDg2gdMYWsaDe9LQ389l+guTYd
cOeVEP8wjImR7nIMeOuxEk886/0ahVTCC+bh0AHrDdsv+Gwe+S4e4tbILsX+TxmsjOTEV2g8M6PG
szXUKcutmDrUriDA9zowbY8QF0zD4D+6qstDAD8+CGtZdTBPxhDxHqY1R4HCASNyk7pSJd4whjZe
p4Yts8v5hy29QBrdFBxg1JWnRhoQexzPeYEhuTS+9rlU/IeDjOUgsmQq9e1srR0p3o5XkOvTlu8J
bygXvco2rhBp3KXd5/EJXGPKz91TNy82qOO0q+RDbucvAlcDZg9VzWurpyuYHvrTSVH3vmkYG+KT
aN9yXOhaodeOHj53iTRbkA1xOd95XAINmu1FuKYdvw4CAjhf7WFval/4ca4sqqkKtyZJVW0chQTk
FNxjjGhD3U/vCgHNsj+PPouRksRH2qSuIk2Pk89aCGTkBsVJgZ0XL8dR/NYNbQvQKjIVH4LB2Fz5
SoIy8ce24fi+fDppC1S3ow8Jo926C6lpo3u3cMNFBqgsw8V1KkXopRlMEIRsP1nrQArm8MNT0zjD
rDlFwsmFgMcp/QvMFp3IAGFi0G3cGYY7C6k0uic7I/Tr+8/vBMxW4UZjkXekGALBtFyBCVOXenly
o86oEi5bcqYpfTfbMT0AnwEplzAVYOoFMzTw5jYouRL7qy0i1Xo1aR/HPJEKWD5hWKxQlMdjX2jg
v83NP1DS/cKy5emwIcJa0bhAaJbSbQo4veASBN03ClVRMiZ1qhTTgICUZtQoVGAVNL038054CmFY
uNLYibWAu5QlbhxhIuCWJn5l0QPBeaC84BD41dfRad99fpLToYr1xYbMN6d/Y+heaHfpsIzKA5tZ
Ac8EyeTAGSRiK9okR9+qCJ6Rc9IpZZidxP8T4JyfbhVCqkA0BCr8ehYymcSlxbnahcc4CvEHZC7S
/ecXUfieKWaIRwk48l3XYV2MK8E/VD2JzOFSUBSeKVwYI/z1d2qDwhtLpX6qnX1whZFIF/L+as2j
xlDPEMWvb38JMWgP7D6Z+yH1OeUvDz9Jc26Erpv/v6XXB514ZA+fC8s7uGh5bzb61Q4iftPw909k
ebw72RucMOnHpCdomp6sWoZDambEKbo1Syb5QLMUnfrTd/eFJR2d+Ae3rtxpnZG+50FP/y8RQivL
RLSC/XnKi8AzNkwYlRoMew83FXwI6M/1xS+DrbiKzX5+oUkzEuiD0BShujY5IPRPcGbdQrrt1l2H
aAeU9xBMYH7DqnhtdKx0LGYbLwehizuS8dDC1pRqnfyNEq6vlqSnVbwDjfa4J7xk8uvYXfhEUafL
o/1puIA3xvkYkdbwd4diguDHH9hGrNpAKZCxKvAXMT1YQ/AEPSL6ElfhxzTlP6KVAfo9j9l46Bw4
eExUi+beZRlZ1JsolDudgKYzsv9BmW4FOJq1XiwFp8pmpzdlKXcyHsZX3RtYM+WPgTfouoJfLrnu
3P9lErYkem1uqppzTGI0yMi1wL1v6D23jSadGYrIs/dO44FLgeLZ91F3DTYx5DAQvDQUmWFBpTk8
iWjyNQs+POHhMKDFWvK/HVuRR18E3Nfv37enanCzWRmQvUBFZXVF2WQZZgr2ObzPtFhabogitF96
i2wGh9Ek1NmGhGaBm0jp2z8NINa7vDzT8V2PfHZMMoObweuqobF4CIRKAukUy1b+XnUInGXwLsMQ
gIL5DNvMfO4NsSMv7eGYVu/oaMZINY4PYRv7xioUTx9dTgF5K7LBifMjmtNEj2iVQ/Vkk3WR+u46
TZrhzlI06RPadaqpEK0qoKbSJhzRmPDsqykdNDdqAKmpRnZM/huv3nuajWSsk2TteEHp7F9UxUDt
Ac5JUPqqmejJyDXmTqsLQ6I8R93PSStuPswlaItvATWIX6a+RhjTOrXTl/a1pnqRN7NxfEVT5db5
gj9M72Yn8FxmKz5s5EvSK9DQqcU6PvCBC8sWcbbkcAvsR3c49ljUPUwIHB+0IjgTjfAZMlbYCuWl
AdVXwY/pnMRASUPVkKLoB84QOveflP5t5Dwn8old2X9c9Y8DEQ07oNRe8+vBJ19JKZN9/rokl3hZ
1EGtTw0Dp4kxabx61DaugpVTGHobykef3o+tad56RA7WwziyaX8jZSGaOz9FKHzj3ZajwUFBrk1d
Jz15m729gvpA0Mv5PndoFb51jxFmfO+SdBa47ZKdItFHd2t2gvATk1SUP4qG9XXcWlfXzJz4ICfF
QaJUx8uaxQMKizqBzJzdHnXWk7lrB5/Agc3Oo/ZgTfe0GUiBNvhpVBRdz7UrdfpAnh1evekRvmlJ
MAfsLtc2bNq8/F0uJkAQMByChb50lsXImR6qmYhF7djJio5qJvLkWYqSiWiugcrHB5WmkCtgHcvs
PMr0J+MgKU0lu8dtWIHx2A0So61tqvIhCIQUjP/6AIk3F5IQMFGK6bhvX6GXqbCotEw2cwY5B8mm
H8OU3IaH9wX6kNf9NZUik/1Crlo0lwdV0hhkxL29Yjcm1FfmL7ueStsDZGJ/afDATOgpE2cTNuUJ
Vu200vpBWb6v0Ho8t9VSA1IVGwO3rxEY3YPpWwqbLNRCYAnfWOjU7NK49xfmN8m446xzZRUkZ/gU
QHgI6qK35hlPrl2KJ42JnNBhPrl2Yo9Xv1FjADzVc2GEPecFQ8RtIijXCRx19THPBygP/7lyYCfL
PyW8Wnr3XGAMlYgXywhoEDa0OyNQZ1LYKIU1g09+Y1enHAMvhkMZsrsar1RLxwRBYfmlTB6w1ruZ
fGMZ0i2EGCMyRpyxyAxZMqA/H79I8ktIpQX6n914MofjgGR6ovjrOfFfJcODpvGoCdz7aI/SgL7G
zkh3JUWKq6Rrpwic2Pp75cdl8yH88t1mGU4j1hH0d/eyZY/q2+psep3Fi/vP+bPkGHX6M2QRXyNJ
1ZWe2mAvImTZX3gxA6OuzgWxqlrpYqcE1YJ1SC2DLcG6NWbrHAaXKGhswcmS06dWfKWr8WG5CeCz
Wu7jfuEJxHQhlMXuHqVrMq0KppWwGkcpi/GzB7r9d2zS5tP6zX558tAH5xD6c2bPrNJVER9Ku3HY
HdyYs4Zs9Cfju3Zq8tM3OEhNIJk6uY6z6BaJuC2V2d+bkZYtnsfTMay+yr3BHtWcWRGR0kCM87ko
tnN68DidnauYcmGj6jOxXpSJXWKYGR4v6W1glhgDWvdkMX7jksamGVWD0neywDkfAkaZpN9GO2bO
ihC4WZxCyxkH4zEhaqLKHRRW6b3XR09RougAcRIgykztyOzTiuYS62fA9fTjz1FpnkLsgQtGO9V/
F1I0cGfvmZlcODwUveeCVLkbxHbOZ4wseu3pc8KjKkI6SVtEv7gzi/AobaNTVD9fmcY3ZFBrXKJA
e7QLYCA1+laZgz87C3R6z+wp/ClYS4nsshd08ZG2jJxYc/mFpZQid2fpsy8fqMcR664diKDrRpcy
dXikXm829CLjjS/wKGLveVo7wWBL0Zg+R4rSxuXg8KuJEDLq5PZERgKpnGf2Hf/jl7vpyErFCeFJ
ohZcylrcWExlfDEKcVuePoLutsl0Ad1CsfI825qxtRabyWRZMWIXPvtGLb3bLFffP5TMsMBaKdfX
wd9AvVrDIzZOF3fmRdgZ8fMw5J4zO6c+RZiyCsmaemh6edYtWxqXcG37TcToKGnb82e/yhEJgW2g
e64WEiVYcFPmaCELvRhEJrXwfPbw98m9065dbR/tbO73TqA0VSkeyfy+sWm1QNWBrYDHMaqeJFl9
w6dx+CD9ZC66UI79iwlxez2hIm2LfS5uQybmFJQEp7SAIPTvkUyBKtO/TqXmLhkP3gjThL90CtsU
8hbzmAhHxQUC2Yt9YoayBpXI06r72oftB/O/veMvyvlTt9suOC4ik2liDgS8sypRSSGgJyZtuHrW
lwUh2LqQti5vkBo4YXOGm/qITQGLiAiJTyNgSg+RPKmWdvdSFs1Iaq/zjhjYb1Po4PFHnBx9/Ogr
g1TpfPsCUuniVRoA/rs5rd2/8hv9Z03FAwijlMK8jaPtRfJkuev2E1B4a/SPXbTQOLIP4i0Cs5aH
xzd7RidgXyIdEcsV2ewpvSkbacLocquUtAXy8WCVKu392J/2CiC0ozCsCu8UJQ8gTJMJGBPMR5kz
x4Cq0q2HC+MxiJBPlGHOnbYJ0QRjesws67PBt3G1umKv6sH7ms0pjNE+cYOJ0UolxKUf0Fgetzo8
Aw84L1kpq53yi1MOt9mY0/w1mwWVeq1Iki9nZuhO/4PasWk9pj50uOFpO2ex5iaSaJGBQcsAQCax
IP1xYWZ0i14MhAEQo7f07EBNwcYWP/aItI2AZigNIq7tEkyXOHjX3cX0kkF6RH2LRDn6N6BkrCvw
iJ2Nz9jbTLLyJdMH0nLCRMjCfM8wwdlhDQsr94FhiT6N4nFWSvNyH4VhwpWG+EFaerIPNK+z0Y4g
dAdRly8BcsR3qQ9Pk2a12QQcSnQRu9/OvJnTuj8F0rOKzaMJrjB2c6pwcQ29luacIleWXxR0Ydy9
LAEsYraVxfML+ubexcFoYKj/LDD98vk4NTek4PXUiYmBOiEtPvO837kmi3wlxX3z+dgXATPPoz4O
2FcMa3+J6M95btZ2R0lRu16M8gGYFqn1HMJiuiPGqaZuwzrw4Q57srMb6tm6dfqqSJ4KSwzE8e+7
2lHgCbqaqnT/TiQVlwctoxQu0NyNyahPe9U41tm7uNRTUxOsyHmuICBUBClPQGPpGYTsTxg67N+6
UXFTk0icIc2s5uloeP3nnJXdVuXQabsQxQnXsU9fo6aKuBgbZHBWRWcyg9hHDLV5nVNqBcXd58j4
qjPtwYzBEikeDEjZWf3hsg9S5K5m+gG5m3ULnCyn7Nf+FLN45yWq4ip/ttsUq8RFbYShXr6xYaGI
Kmw+Gz3l7nLCRKNieZ+uryAZC5IfXob+/Kl5SJZ0bCRJ0MGtRAlbTGdXAljTv+PuXXqgNlturAO1
kEULtPdbTVhHrhMQBuQKgn5Ip0GmuhyvMVOUYd87KChcHHKlrI0QEO7m+M48NGmUOqUN0Yw02pSp
aqfiJYSYGEBMRtvos5sct5+OG9lOegIt4hzF4gTepwODkSQlqSbE42Tk1i4o64i9aWO0WH2XEBAN
9oPUg9Q0mdyVpj85f9bzjqPmyQbYmPOA6pYQyGqyhi8I9cgobnC+ZZDxhZ4oiZ8n4nKpqF7UyGht
esbh5m1xXRPjLkmn2CHh33gpzgdDPANgr+M8YTqWcWS15L2pPN+7AsB88N4VlMnoSXHmbCf/jO6d
/fq9taDLHWVcHfPbWfZ7ea8ZcmZYj6nUzsGiL6gOrXcIZTcJ2wOFjgyC0AaC+5AuyTzy0Fh1afiQ
jGaEBZZIm+SB2FCzHLoAvz7WS9AkHvmgWQOGsv1b5k0bXIBwKpHV/VmpwSyJSxLHRWZWnFFoTS11
Qu+EAuFALeaLbNkvirwEjIwmONyewgKiTn4PCGWoCLkBf/FAN9IknrXp+zZAznP2BXXeLOvujtID
6oZU/cC2xFXuDD7MDJ6whJWFcAddT9Cj0fvI248lyh0pcKurnsjkjVv8gpqnxlj9vgTCFPwc7rRz
Y7vgR41XqsTMuEWD4BgNfcerc6hmi0XrQ0rSqY4+aXBVv6drOMhVknybLeXS2f6sDzXjzWOK6lLh
YcN5GRx8CpJ6ULNHujRQSoyEmTWnF95omcvbEwFYGzqK59z+dAqaCMkF8vHWTqutaj/J2z0QWIeH
J6F6fiDQ37aNxQCCB5PWqjf03aH8UhMZPp4A/u1Y2TfG7p9HsCyFlnHOwaD14nBR5MqCAfwzkSri
gUw7hVArzzIL9Vt0cxdV5n6Z0kjsYpjC951Ueo0jYJQmxju9rqYwTxJaNZP/Nos7oB4kcuZ/GLIL
RfbGBCNBFUBcwzbgMaTUtqKr34W2qtkiVeXBoLp0I7957gpXTRLWNdGYHb+GFCF9OUMMzvM71VV8
i2HPmH15wM/wt2O25W27xoJWaXgqD2hxhKk/XVbntF+G9fWC+SVMne0/u4v8V5P/6L0HmZ74HEGv
S1X0XRnZSqNKVxljCiJb7p5Yp/XgYZ3OccO/nAmEd8ow69c/SPMf1Wzu+j/mRr+esxOvj8jjbFBu
iqP2MTzhhVvMMIL4ctKT9J45fHQN7nSI1WuzFG81FBI87VX26OWrbVHKvW8IX/a3OywWKRMG5Gs9
x9cfMHAe5/MJOazCSnLKILY+Px7U5tPEHBwACXM1gypUpmxc4j160KuBVKgaqi+YkKDSlE43ZM1f
rKk4mD8s6f5V/R8aVTCG/tf8Kr+TrFNe6IHSigJrdoQul+icC0xrkdiUbNHB31s7cnxNOnl6CzAp
l7OZDm/OH6lCROAOkOQRv2FZOiTOoqUVcXqU3bheuKq2pAuS6T0rwBofNccb078TIA0MDvz3+8C1
yfhIX/4p3C4ong8r2wNNiDrooXiaAXnQk3A84eZGcvXMc/oKmt0WVJz1ZFQ7dgPTOYIqztRusK4M
IzJFJIvvQ0E59zBwfKgVVHk+Aw3i2xSDzgfeyCR9dhhV3NOKR92GpJzuI6ylVjplinptYFhGe+Mh
hk4NQAzsiFN/5gW7OcBqwQ12/37+D53PT+mXbANrlEqsmgI/4Ocnqnv/lPnrykjdYgcBBNdvPtC4
bOHmsfJ3STU5V6+oQsSImhuKR/xGFdjLrQFNbkfofbMIE6lDp50j9hmjyRpoZ1eS+DDpmYLgiaBO
0XvAQnHxGK0kMCf1STBmPt2SsdARtjp+f7OXFiQ22YzE6k3hAFDOViPZhjYDypXaNuaPnypT/6R3
aXQrfacAIZph4FCfzNOGmblKpTeKuXhvQgjaU+gFvzF7eFpKLovcK4o3t/Sv/YefeVwWFNcfQSz+
3zhlLe+fYmhXdqwIvf8Eghf0EU0mrvXKsl1wMDEPN2xTI9/0zWe/tC+UJcvs/hSnRI8wCkeb9Olb
9cQ/A6Cv9Gwj7sAtTRgT3xuDahVRF7OAvycRmKzY+kLlVXuhAoDJebvAbTpl3EnlsQlKKWUoOtbS
J3G41c5sQvDVVPF2iJIYMZ00IBuAbAL8M+5fLPunUnqo7Vb5zR1DnFV6Ytoi9gZaWBI/lpLnuUiq
dj7aA3uD5JZThnXRQ1tQEBpHMBsmMpj0HM7Pb6RCFRFHK72LuJQoGvTWkLQSAEpIYfvPlanT7NfG
v4RIVkWuUMzq8NHVt/yatjgE5GILZr+2E+MbrlHwUl00LQvwgeFJrBfwC3f6yXUmu4ltZ/Xcz5EQ
+szKOiWiKajrJnYVt5TS4TGsQq25+wztrVKjcm1NPkM9xvv6LiodLfBfpLrYwELJXvaakcJBrwGa
C98YXv5+6vinXF/2lUCWniB2wE1uly7+lps9mId+MlHA3gPxaLEKxl19TmbfuD1Lsw6Ozyjix18Z
wKmEgpAx7uZTlOif+BcrxuGJ2gp8vdn57gKq/moSEifIV0EeBSZgXAnsV2ArqJaWYpzPV2a8cYqR
Yu5fn0SRwBQkBo4wXu3ruq5bU2mJUC+jrxdNBRgh+2s1gyGsMpb93azAQUQs9kgZfeUR5Qmr1gQm
QX5NaFRc9U0wBwwHxFhx4aHKtoxOQ5WPKjIzwOpzLyz+n/V/qD4jNjq+Z+EOb2vB2Vlwv5jeJqSx
m96AnIOE/DRBbWEcCxNd5jgRrilIAUae+Z7bF3GOnFS94JkQ5fjUpBqCyB4BxWYjFQ7ftoB/Bl4K
viAfAhv6t9ArPnefRY+1F3STHX3P/YEPY/sBHEX0ijPxm3v/mhA2ktz6v4pVDkFP/u36h8D9+g7N
bvGIXMr1U44kmlCHWMT7nGhCXKnBP8AJeWQEe2cprDGKSoK9zYoUG3hLps3CA4+Eprz6uaKC7AXl
jgAZZdbROJ56ZJ53Odqak7sMoNUPVQoTh+La6XRXZn4K1KIJ2U2sIO1ZCT+TtVImSzNboQDIpHX0
AbYfMSYpW0VYUjxpJTrOrWo9OdujEioUZqVS3k9v4fDz5h/2b7DHv3gnANSFBTQZwvB9FfPol9vu
Tg1v3YmX18uTiTSrGNNInUAYYJa12u+c6jXmcCcMg4967T3FsTW7Y/XEsGrLe5TGsaxIQ4yzo18r
sR+ZlQgvo2UFF7xetnePB+W/kJFRWg03+JGU+9oVOcnm+fT/f/jVVCkQIj4VKMKKxC3V+00qxqR4
ElJaXEA3ooEQ2Q1cEH+ON2eFhh78nE8J6etIXgVPtFHnOScj6n1pY7bKAGwIABVso05fl7g721j6
LxwNUs4MXwCNOPnvYzd+2T4QTWDVSm17zoMFsY59PAZLBlLu/IB99LuYz613NChZrnxKqYnWZiQd
6/dnrb6vV+nEdGcvkJrElqwJN8een3kgtGRRiG4YVyvZdhvtbkTRsFokzhYqqeHdtJ7g3g96Sv1S
kGXAc0cg5JWI62wHvlpQN9ksqUZpn0mEweE+qxFV49Nfw9IW77J8wfAAxqCgiAT59+MowBwCWkF6
hnt5EAGAYW4Cx94f5QChFqTIHfrV4bn8I5JJTNYb0hCYFTRncDSTl5PZjdJYi/44aNEwWu05Gv5o
0sb2va/Hd79UJjO82yq76BPqpagyGjYBkHVz6kRNz6sR1/g5tci4RRjrbLHbjdJuJ2bfTYYKEI2D
Ku4R/zYATBMyeCSQCYk9EQaErGu/6p+xnbXzNcrMIYuomlpXA4wn4HFDsbI7Po4IGyYAGNDGLWc6
sTfOd0PVwb/4OYInbasUsrWAn2z9VXAZwJvhvS/96rdCfrmaq7XBZSQGB9NO2D2aPYgWXOHx/4/F
gJSCGdzopPaKVH83uNlQ+RtGqiPPXGJVYTMbwVUb8fMbA9ovjMQgUVa9B5Xe5QX0C9/hUqbNs2ui
Le7KgYBgaQJJCLst0icX7EIY5geS8eGdZ6evjYCUQodnd4fpl5g0U5+hSkLXX+nAbgiKujdSgA62
s0r//LCVAMj2UdmFmQ/tyS4plzxYMQ+IgGt24/c5EhYS0MNeG2rkTih3hEwivk06NDzCI7uvNxA3
0cCO43eQGc/QRfRdvqew02+jDmyrtsIVSfDfLXRB2sAgZPes7/5FMwt4ByurtWyvGdDQ4FKbu7ly
ihhN2DRqMxrs3Ys/YkW/VidkfM5JyA/Xf/1wpdwr6V3z0kkTe1mrmBdjDiQ+eGrAdX7HfJBLgfXe
qnqRqGkTeAV9NttQVDMLDp+GxNjz/cZqxDo1/iEeMUMlHD7LiHdr6fP+sisBoaDZk4EhDcneWzCv
Pi2XOg0gX3dvHWSrfE8o3zB2nJRO7y/RPfUjygbwDFy+GiFagN3DcxKXKHyYo0vxiEfa2/L4bHH5
5J5i4QEc8oU6GnwBBQmqSMClkSgrXcue2vpEdltkjw6d4vZbXaIPBZdDK/cYGPcrwV+QpO/vDDA7
pBdvnAvHXXm8nzpnG4Z7cvo98RCAcikJGZfwQjMrhveOvAJzmpnND1j2VdkJhTSxkGMJZ5NHDmAJ
HGzX5Z0WXQQjqY7vyHIL1yrcM7h29gcg2lyzGcLzRHEtxCPpWdU2IRzU5ykMO80fZZd069YxfnbD
sx9zoskxGxOtjIbciM3Q1iyV7oQqR2hh7ksSOQcHSRnv0cunq/Lj5romKYQKXc1KcA/8npt/KY6r
dQ6fPKbka2MpFotQWhrjVIZmAawIiDScRmd3HtJyy4A0AEH31bAAQigZDrqDZR27MTroXigDs/IE
T+n7o+BTuFeGZcgeqpzG0ndNil2xNSWQhX+RB+8VUXtkNqg/GAgXlCA4E6dIo/9ZAJvdpfGuRGhW
odSiku5jgWMRGdEZ9MDYAsbuEsmCD6LlEKDJceC/Yp/lhixscW/og+up37JCMzkFCRgHqjz/hQK0
rAKicu/EV8z0O888gKSd5FqU++dIqM/iUWA8SYEABGBtD211j3FRaLa+eqxalkiKoUI5QSiymhZx
uOCZmdBwi/MB+qJt3CPwRO/IpZjSl/nWWRjFr19OIiK9TYO+kRJoeAHAVTfbTLKNWVPUYU1paeSS
h4spjRB0DMhOhrZeJtZHpMDA06vJV+Wu42aBTLf04aedUloZbcze6oTuyn6kf4gre2RjGOE6g9Rf
iacN/Zk/0tXMk/JlejS5TSagJV5Dw6dbX53Ku6pYidiQUAnn+g9z1x+3+9DrVfL/NWz2TIG5OQce
mcCR7XV6ViS/w1ElVlZwIinGDuUWPkM70iWKpmObNc7z02IhodbiS1g48FHxjPDn6o5kJzJgOKxK
NNoyclqbbckaJRKEaIBB5whv/xnElfjxMI5x5SynY2FB6pknws4MxFCm/kYfJKIRctSAmQv7tGWf
2WZX9pwdMGYcRcgHVxpdVN4+xz1e1E9vB06rEJTskO7g66/j82qHETDEHqmUPg9iJ4r/RRAzXRze
xlhut8k47tLq1CwclwIA8Y9RZVXTFt99mIzTRBQx8Pl3uDdTfENBJU4Z6BuTs5WpzHJabYbV+twh
Y/np7lF/X3BBlW7XNvv7J5L18AprAwpzGrZD9ijaHJLAZPGM8JG+QES5q53NMqJ0R+KG84j0y/C9
y41zz/6V3z2gAOI4buU3gl4f+0Xs8DXfPhb1AgUi/R7gY1jZTdxRSrwQdz5gT1yVQ4paNMDUzatZ
+QsHWkFbaujp4+bJbN6O4UNd/BOflg1xJJ4cnIoiH5q51dcOSVYUlmvXEfnjdfcRmVz8b7GqamLw
Kb41umbzdy/0xquUifuDtgo4PPFNVSlEIJxv/OahtqZnLTRrexhatAX2jEJO8rW58hAtHAb6v0XF
HtRTKD6Kkgej9ynb9wuFP92dTsaHVsS7timYhzWQuBg1g/bZUPV8Na9zr4njBL8doV7lLB4sEXQO
DKxiCQB5KO4kgNBNz8uEeku8lBA43gkH4syiEqhLah+iWHpTJjpETPV6GD+Z5uKvV7LiXtX3pRvv
2Ww/Hp2+JfIZGwyVAAt/1KN3REukoifBRYFnUkbqy04FdbSZCRv7+Fi69S53SnQUUUgxv0cMhwCq
NLnr5mMr5NKg7F3A0DFP60BknxCqWMVIXaae0FFKvHJ+P1I8uPnt5VB/tV5Owj9zijU2zfVRIXu0
hvP3k9193oBSIBq0KovzKvfBOLs7kFztLxxwjk+FW4CgbRbkCJxWMeK2CnrAx4SngL3dca+WHmkv
xXr0xeluLHhDTMuMorvFw3P+UpYS326FBRdZdTWWte2EJeYG08E7CSzSaPWjkiwS9W4DnqOaEiCG
GKafhpXS3+E0vXpi2PMY0RnjX811sv5RUeRU9CGOWgqy8Ab++0syJ2GcMQKdDP6pq9wHQ9a0aBAq
HiwUjmjjDZ3XcA9n8x4+bMiUiroj2PsUf/GSNaWPrXfO5RqXemnOqbJ9vqH3tqghmAJQuZVnqMo+
4XLy4GZofdSQm44Z7eaLb1nn459ppDxlfKNLBS9zELbKRIdGJQMP4g/UmcRlxiae9hV/p+wzK/RU
oDf6IktZPcsPznyw3lMqK1vbsIBsmGmL2180fWZOs4i2iZnpOTSyWkyILwpuFu8ZUS62bUlWDiGh
V24vzU/E2+ytwgt9V7ew9CDmFIQsZIKZ9fcIv8gDia6r3a5DQDIUcx0sJTLrpqJzWN1JUNO4ljIf
CnV17soYuM9z3p81NJkM5sD86sGj/jlX2JvZdVvRzQGKBOUH3UA8k/NKJI34ap337eqBBTJmqFZM
e+9NBymNcMe/hi43LLGZTeoUbOpNLtHtBY88FNJcuLZoP9N7eNhWvgDw0pRugR0efv+nw2J6EFHb
evDA54WPmp5k+zQVYZHepHxgwLgpeV4/sRcc/NBcGBc5fZV9B9TKef4yzfsUw2BfwT5c4yGPDOMm
cLhGRrdBYtd6ZIOEeZPDaF8xOl5WCmE7ZrTcUX1hRRpOxCC7khrgWDXKYxHYHZihpzyKcJr4G3T0
ROlSXqlf15aVXczsXly+C01MOqPswiGNTRUO++W+06s+zXkWV6jRRmXK5X0Gdbe6+YMNgI2wuD3T
xK820LLgXxe//u65ODTu73K0+L1oXRb1A5oJtfrklfv0S4tet5RzgfjyGCzeHNS618eelnJNZcj4
X1dVo4HIgXYKNzYAABACKHO5fEYKU5fpUWgbgnIUHod1n6ElGh4vTmKA0qRIuB7efjC4v3DGSI60
1MWrS4qcdipsXDoUqB/pmHKzEAcZA+E1yPgS1rT2RiYQNigoBFpZdimxDUNnTGgJU93fRlFnbj7u
pNnauhPB6JdqzuW3mgt5nCodPrOUJXgfabxm180SfobipqpVBpC6w+IHP+rJiuChJ41yKOYIDviN
jYM9RliKbN2tGcjT6LtggfI3uQ4se+t5xGwT3OBxuEgwuVmIOUHz5BB4C4A//noExtBcjZb+xDWX
E3jqHD1tzS7GLnfKL/7KoFXhBqHVqKwD5DCPBQdczbe6YH60Fua84J6f40WRmux13Xq9voKobqU4
9zXm9E+hIpfsj4UbBx79VpYN8a5Y+8C4sdQWorBdu18yPdKIxCNzpR0V5irXGXm4HDiGtgKg0ged
yQ8gul15yzNb9497G250KRsmZQaBUHVttJOQ1zhxdF8UmVqSO6mce7ceaTGecJyihako3f0RZFWM
EjiEuR/F+2Uf0sEQH1R4nhm67GK5Yv4XqEN6aESMn3QQAKGlO6s7froZertLc4OThVs7kJDeTcM5
IjrHVYW9gCrUia7/adi9A7f741b/c5DMmDqYpEYV6ywiDPG17I9ahYj63S7tk8iHxRs+CxdAzWEh
10MxHmtzXaViKdR+o1IQglQag54fhq4tqzjFKPW+4WuzfZPR+QkysooWyo98d3Tho5mmNjT0NjM+
wxhPg2C0/KdqW7IhDuOQ3GxtKkelDqdrg7YOZjRe0H6SZzFzGjXiPn+gtwdXQ0W4MJfsky1/BOAf
/1AgHDrwKeTuXXjbRDy4jwv1ZLY2T11KSjcGgmJJFrpkrFt/WqXY2vv0sr+L003JW+JPrt4Kiyec
/W3Rw75SuKnFpl31W5tdeNfrjBYVnylIj5l6c8K0Yqtay1ry3x6eyGKYtSRYGoyMQJNDrveVvAg3
+ygQBmcqK1JAmtS63cGYsxOr4KJvmZ0uWMsuWejVIIcqo3GuyKW4wkse0ifTd4m7MVwNikLGV2WM
YFMgOtkr66lfF4uct2bVCgB9ik4vwO6RFnRSM51A+H5mW1i6kUxK8xBX1a+KtGbftdFCobJTIHCA
SJ8sF5g+ldL0eQ16xixDC42euM0uD5gXM59tn4/QF11/UNx/CUVCs2hpJmGE4rXV/ZZiNJEb6adK
iVa5zi8gBN/VqZVMjCurWx7TOyE3eKvXKO8WbDEXDP+iWoK4mGomIkyJt/IMuobY7VIky2WZ5v/U
J+CSlpmZULcS3Oad79HfNetamgDghR6w9I+IfrjB301mNnInr/egm45+y/wdlFOy+EUUXBGRKF1q
0j4kfxkg8w+kp7AmOIwdQ54UBL5nB87EnJo6pOZUFOzX7sTqDeRf1E5nUwc4tacN2R+Svd/5LIN7
kSCa86n+qjEnWd0zGQQN5k/Uti7Yo7LAnLKEjQpuRcRMA5SNleuKd9kEfERnUdVGQo0MA5LVGaNc
NvgfrMc+3pdEjZ4NWaG2TxCZl+pFYBlH5VuBAUvDH+zAg4+veDzXyZHBaRa5HsjsS8SD1p/0GMrz
Td05DIzAQYoIMP6M0NthzwzZO8wOmusHoncFAWMZbsHkKNzpY5BLAc/nJd2vU/lqn7qtTfyVDEHX
brCHly7dZVc6AlqZnivOxFjkabVwOnGdIsiab3xpQWcMxxpTlhWax7aq84lnIrYkR4veg+8anP+D
5dkV5XEwc03TyFhGmh0ELkyl3hsFxZ7bDKNbZrCmVZeJ4Au/czhAf1DQ2iyI2kEuoLpggc5kZuVo
+UVhoxpT6jpnEEBzLzjQ7z+BQ8EZANThBgtecmNNDtX6YRmPz65DUtmkExq/Xf1FzcrN8PjL7D5x
9mIcMyu+KqvnJHPvJKnpOFXeh4rZudCTvPswRcAAiJdvdFMoIOmnb0wfzp9+lpGb9s13Ifpb/MlZ
OIIk+HO40sB4EoowArZqqZx0UB9wmwFv5AKg2gsCAjLcUW0o+Z6I9JNhaKh6oIpRB9D0cRui2hzG
aPE56cdLaSqh7nqpbg9eSme7SrT9zwVTbPskKT0WXDt+lZVBSNC7IDaLMxj1yngqkHe5ehy8hrKd
a/nuE89za7T1QfMlgm1f7nRzq8jvMJ0oX5gYjRosKiUXgqZLFjVRKAudqRq8O3ZrZzGeNIL4qXJE
xFBmph9XJjLHS7CaUsFKAr425jJ1lSNAI9PnEiRyhmmDubxNIUe0pKH6HuBGEhddBTsLQfHlR+7j
JJK3wGqL4AmMXIWu1PVetRV4B9+IWdoxyAZcZfWxQElJQdeAcnfWbLsE0TBVyiiTe49CUVjNtr2B
wtxFPINMsIzvuqlilngixHGXSBMfDeqO3WRKs7NpieZIvVlH5CUUvJGUU/vzJhuIkEGTNcqrmK/U
zWWSe/zS6PpZnm3Syn88tv2dxSjPn8iE/ULs7gfFXxLomDjhr1YnbW27PfXfwh+Jwa+Ri7W5Qio7
sXe2a+NC3rs24m6+igge2t4XOYhzLPTfKf4CZIeIHZgRE+Yo02lTjYravJz3nsdCnwc9a7XUMAn+
z2RkZIVyAppPEBaM4itSfhjIEkcCFimQvFfrjHGOUv7i8rw7EMHGBQoYadnaWV7VJlOsWvgzInBc
wsaC2bKXeutZxZgCXVVkv7tlTmQ6pJFUru4iLD7yGzVIUEpm8myOUsoHghRcRCTkQd+tT03y539v
7ciPkXhfMlOxWCaTQK+cU19iP0dS1QL+bc9etiOMfa7KOXPI0ZQ5XUb4CIb+Kx51UFxnauxI7u92
eGhUrXRpqDJOyRPG/jMqpX/3kczWjOLMgVxkGWtx8A810Ns3jpSupqn3dlN6839FjzOWn9CldrR2
Q3zugX3NdbZV29R/tx4ai29SnQDR6/CBYwY/gfBZBJRcdU2x7oYWAopMseqOtOj9P+N/ZRcT/1q0
Gcs9dgAGtdq+gZt1VPKLgCF1F7svdtz0j/NykKVF5ImC6sJTc60PymOIF7k1CuPhEfuamvb04OCK
tZrhUMg8ybu+GuKXuz8ez5W8oFTZamScJsMCUypePm3Jr2uc9RQYESJUTpXcQ6uX1f2JukPBT5Ed
JG89N7jiJJI6ZbQ+C/XSRHCxeTEeUqkY4yO+VA1DA4yJkHIK/VIymC4mICZHil6PU+mj4IWvXxaA
Y4DJkt76j4ezH041zy/FzUrOjOBnfa2hZ44IAkCfigJ8xhvjJT5H90buKDmVNmD2L6WbNNjBl0MA
Hi6uF3sbNAtmrcMfhy7hVBIlpdstt4D5GJEqD4dLt1SSUvjgeKTNBZF60/wvdUrUcGPho1OelR5m
tyQTEynuuNVR2J6IbWN5tWFo50XeEUXghijesgXsDOdOfSQzcZ/tsA5aHoC/nEdImWg+3xhuGgHZ
Q96/YNDJ6ccd+PO8sgfUrDBmJtCpZAUrLeuuczHWKppSMK4Husgj8FaT1WoOHzoleCVgE/7JXPSO
fjZ1Z7dkN/CNnbVtZ85AAac+mAq8NrsCpj1dw0JjqgpRU9XtJGbWa74XXSEwVQ47GY7bn4XgFvPl
4xkhss2L5+upEllytC/lMPmqRGTH5Qxuc/xthpxEqZp12FlKmIAskgiHRVPy/zZUOZz0qLMjEcr7
sEQByUtZXTMceJeAgighHhDksCZFINxTGkCtK3wCuThxm0raMvOq03/bDEY1HovQuLhLM8F6LiPx
Ph5nItmHJw28eUCI9eEq4bL4V+4AWYqp7S8OBQFkqnIaLxDOqkThFBCU9cSwILJHlATYI/dJaU6p
eCbk4J4RqD5+Bet/7qQ3loeXwGtPT5x8RFskv7f2119oXjsCTyyDwVxRvmnqrP5ijSnbnhCdupEV
7MvtFmYDepii5qCB7rb5Q08E9stRpJRHRUmWXnOCV/zW69hKxMrORV3BScXLj3ibyWZ3pCCfoqQA
EfD7rllaV3HzHFki/SQbOE59OYBcz+/mA7ypDA11BhxLd4l+nJ3RFblXkXEVtgiMUFdXJ9vc51zr
1j4h6f+Mc0TuChsbgE6rRF1NGBTTtOeXQMOOaKeC73qFCxnPQBFgdbaSaS018VeJLO2OVhu2bxzV
UJWmtdNnBhotMx9WbhAw8i1vFdHwp1YHSTE+6uxStZSrcQoj6Q2L15RfCLCikDj4HvWomQvLeYLs
1mNjdthif1u4UgzIgtAQs39L5g4trTjFaRWs6TYypFai2BqMRGMjAKwKLZxWMOb72ZOp1biHo/bY
dXTobg+oG5ww/+qI1wkae8ENykE9DHMuzOnYoLqI8PIbpX1AW4tYWaUjg7DRot7+UDKg/JdoUDx4
VR+oBOzS6+Zma7CurMEgOsCdnq7fMIrMXybMF1x8stLKijiNZkvtMLWxVSffBsSW/lGACaVuqyjf
HRFfX7G5tGV6Q7wmHcUT0p1PkwdpZPuS8gYRzQ+oAEbMw3AqFmKaefX6IrbR/kZbzV7Igb1aV8ui
t60swNQdD2t/AFXATeH6xNuRDxHS+VbtgQTv6+0I5bK6EBDZwFUGL9UPlLVV/0f1zEImyCrA2g/S
DcCBKsqDSQK8vHxvNXA3StPR+pTxv4GrVGeUAuFP7fzuklAHK5FwVI+bQrIa6t1mbep8grpCJinX
aqaNnirOJtWrVItokTRA24RRRHQc+GNiqX9oy6cU8apuLwpvD3ihhQkRHe6gsiJUXpYQpkWCbr8X
jLhtOYUZJIljdevPSvoHVzj/Ib/LNsajQcBsSLNKGe9jMyGZJ0xldtClZgQZOWXdFsgEsrPomFBq
w1Jy6hSoL8dJ3DoYuRX4MhBL1LkNwxS/FwbXkA0meqftqrLK+cdcbL5Ce57pAw2xOESElLog9xn2
VHO41fXHpIbfgP0/EoMov99gak9E1EtPpwd8KCxbNm3jWooV74SddgI4vGy0LcX+9VsSxHww3jcb
k7AoiDiZms1q9+64c2EzaJVEUTyFiu3hhsxyVGnwGV2P1U93K8Q8ZKvMRG+poR/RtT9VKHRHznMU
+3TzyG372KUnmvwL5aTq+a3UqhnIfKNINr/KjA7osRDS2jDO9yg1DdMbNCuwF7dJQpNQyV2wYvPF
dWVbYshNXXM/bW1FP1/bt1EZOh+QkK5AWUgBFPMTiQxGm5uD/L2KbCHcWHlM0M9AhvmYBi6AJcAo
BeU+1ZbZAgFP93bCYmZEVSLA+zvlK1QTSV/Ya/qSeZKkPAU/9ZSSftSeHdVeyETBqhjFTtrwkIRb
2vkZLrDnDHMOwfZO6H/7R9igUO3OCw0wNU1RkVoUeMV4Ka5qIM6VoXFh23PkJqlLSQXr4YljDhAE
hw55Lyc/rLqdn3idS++TzFki4bjcwyOiOhMR/q71YOkqsL7/W7RhZ9E2sQERoOdmrNdWNJsvPNZS
jeqhm2Wa1ec1DfQ8AFwi80j7P9lCw88vhgcHQxXb7iTiJ6XOwQy1CdbsuP3Ina0J0aITU5LbK4BT
hcDicfFIpUZpXg9cwiBGGMez3+2Lbz3o6c6TtVCGn2Y1pWLeybsAnkDJcMH6ZTp7XSwtk/XvHGOd
qKf/9Lkw/Tsx9XvfhsF7WpPAlpPxsjEYqjXdf3CXpmWlHlQfaLcdcLkhE5f17zQ4ZQYnpkzzYAv4
J5YpyYeEgzAJGebzHXp68rzhnVGi0P13IeZwGJsltliqjbfr2PktDh2WFUYo7ugkFTdEub6pIV49
3EhkeDOGx5hURV204oc+jf5QWS3W5HDTzokCZnlrKoBz+eXsRi7bqDhbIkS5cAD7MJ+hPVEkvB6i
ITqauFToGuJQ9Og3OH/Q0Oc8I1ZYJ+rh1QdW/grx8hBRhUZq6rcgUYwRsPoTFs4gxPJZtOoTW2FS
0BlltRyLYZbuWgzePwzyJdWKMLoBz9tP8AhVfCC2TOl0PQPD19Cl6MEqm/bSh+RRSLjCcJJmeZH0
HuHakGfi/9cczQz3V78kOd68L5GCMIRfl39aj9AstCZk0LRD4JfKxTXktavppDlqzxKghRCEawcS
cpMXnDPWJG7PstB3saEZsqBoUaAi02zWBhB2duo12lxuYJonBhTzc2JeKZtpcaHgLTCZfBg7W/Z7
xgHp3X9YIwpgGfDjIrJnsLipCVdD5Ev+DyaRPK+4gWTCdz3+qMdTOyePc6b8MrAI5ChQnfbenjgp
OnrhY72aIrUCfHsPJTWO8Uy9KHnJlIcjPAAzcG42xLcH5oKKi35EsmsY7yJhToa9sA8aQfx48q/+
/rwP9XhpJ/g8M9LXssOwe+c/9ttfWgPUvBrqMp3Qiy/cDRoCYUWpdUX3j8hczdrmzL4r/g5W+jPm
dxr9ZRem3kr2PJ3mxcUN+dWHMVGez7e3TNKDbbrcmi5U6bO73Zrlpw0vFf+KSY6cP8jxwRn+hv2K
jAMcpx+Nc4yGaHgyaExvqwlrCRF2B/Dfn+pRIX1ZbYUYtQ7EtbdGrUQ7OW/enHqYoD3QbYQRqBsS
QqYwRQMeqNrn78Q9RPw/b6qqwMBViHWacJ9FEoOFx/bgT0GJ0DWUTUkvI//FtIqFK3HC0eT5ws/q
RjB/ZnYmSUz3LNO/p0QXppucP87rtmlzCqHJPWGxdZRrpMXiU/N/j2iPljESqbOPn6sanOcH7Zqq
O2uIXPLYmfms1NzDgyH2jqhKTgwSAH/jVZuXjViXj8NMih7VWMtTrg5cQdxXo6+45yejqsPnOkyG
qNtB2qOwhLIkGTgx3tI8RIKgSv1GJ/H+J9mph3b0edys9hQ7t1c7RofSnrKnJp/ops8gEP9vAxD+
FPddw0/DQ1Z290PY+1OLNaH22tZNC93Iu916wHPDlePBWIjyTofhAyMYrFAligOncFpzenM6dho3
532ZJgwWZzKBnPxhSAdd5YRvH4KkooOKOrGhGqQ91l1Vg3bZts0/CXkwe5HWjlVA7YtRX35jgGww
e7ZLdKsnkK+w07yfz2uDbPlcZCMjHhSfHJvmorUoydvUtddjz3Obv/jYVLJxPVZ4Js2jKFjFXSwZ
CfKXKZIKLW1qW3bgx/xxQVbSTDVZSyzvViNCcl8LeVcM4yBpVCxH4pXZ9fNkhCFY62CuccI+4u+L
oqiqXQCN+jjqqNIhszQ9cUf12wFqV9x2EjsTbAUOKvu5PzDv//26uNnZsf3hgbNt2JUkImiqpxy6
JzEqm1c+lFLD0yKW+gCz9P2kiyIsBBtyyMF+tsvosIij0sy/Sux5Etk+oK2YC7EVqq+cSa4hJnYS
Ke+D9F7gE45o/H7qVNVGAFg6rJohBzhebY0/pfHRWtsa0yeKRpPYqCuDuZ5yc/qTvAW2VBqP0yux
p8BvSHrX7kVfFF6IoABSO0ZPoWCxHOQjA7NgJDAmaVANiutBGvlu/K0vNIO8LW8BWnHVyCGquISb
THrvM8VSFkfx3pr0zZXBkMGiWSj7yOhfdYOVdCnqpIZ0ICTEDZdcIRK3Ko/xVjiSGYmQ2TStyRFj
XDEYI14fyZQqcxQJ8W4xbqo6IedRZJ4QjK4QscuadUT1zcdku8+2DgWen7ReHo5wHrGwU8iXW6TU
O5p9HvqtTgXA5pbrdCPqHgKRVYxGAFWLBKeWK0KHEoUc09aS5LdS7L4fOExGrRKtzuZKzZ8nUDKw
KocXG7L54T1NN2V4QE6K5lixBCoTAP2HK4J9C/cECyfCDWMzBPei455pvMLp6V8FJnHhQSBdpr0z
9GI2ue0T8qYnYsCasHZ0iMR2XDKCw8hTvBHbM51hH+S+GHpE0JBd/AZVyoGpU2L4wohs29N2FYnk
VRMS/hJmyGHn+ZGHuA0EAPxauLS2+bYjUleARFrlSdH+AdZDPb6MXkqM+J6r26ukrsOiACpPp8ca
pHTeu6Tn54YlLbkcF3Oua033WPS6214RYH/aAexwPf8fRwWHLZkSMMdv5+4FjFfvvUAlUvVCghsR
4VOmWXVNPdLDtEO+QcDkkYDzdQVchoFip2ZRES1jP2lpGIDDnZT3d81JGS63iQYtKP5S6okWzBhp
Sys0YfaF81mZxidI+yFywlJcPAT26M6ToAqIT+F5hO7o9eJzWN8wtoter8o+cDcmk/KpknHM1KtP
FDRUcRiADNchOjf2pCpb93Ezxvao6iJWmC/9U4qLkhO1OxdvzfMpqPqNgw1QbLghJYtTZXM1rjKI
J4tFXuPLosz9oCIzbeCYAJaYOWWDgQ+/g2t8kMebabjiaY9xRamPMfbDuQr4Daqx0krXiIFKpWCX
PPCqV4jPu0aXt8QTU8XYnrRgP95YftyTy3SuSkcXAKLH6JbgELxCSuGCZqmtH0lQMqX2b8Bp31AG
vm8mIv4bQlp8+MQKBlhdRoCrcS9MDPj2HNMGXeIMDtoCUSZzKgAEgx1y/LW8K4UPyM/DG6zcNxSA
0wvCQzawbVtamTGcNutr/emHd3TxTYGLpbBW2oTZtbQAa92meKDkWN1XYQBJ4yUhCAaGcszNYsiA
KmPbmJdEPs6aXl0s1OzAIZJ0vt6WR6LGN/oIoUn8QtBUipnW9u6sKk5j0gadjYqtQcuj5JUijWRJ
jYWnfeoBu6LIiGge56Ldj4b6dx+CI5iqXNRy2B/dXeNCvXmT8DQKBUnd3OzxeW8RbdMhMdfCzsSG
u/vbm7cja2tvJqgmVBVzYrZFXO2UvgxbDvQgRGvOPjIL/8TBsdkLC50Jk5n3pAmk/oGR5kG2lDgy
/YVe/5KAi553RY84s2dspZGM7yCj+ZuxyxG9t1s20oWhQKZEJr9LcBlq4LJ4o6GhPd9h5GZFpNhq
M0pGt4UVAK8ggWPl9+Do9d8szZt2nLdDh10TT3rIB3052xtuniB60I38ylRYnRDHsLqjvORf11Ha
2Yqvp5NzqECOup/nGzwOaRZOVG0O4ws8iLgRowaFGW5//3cGjg35Eg0qYhtyLJC6Qp90/kUECzdS
3BDdpVLRsdrndvB0uxequF/hPsNSE6yA11T8EGtZyzAbazTb7krUT1NTOeFYx7ufzoIWKWvCYVv6
xrbyKOvtGYNyIR1Nu12LfZYYU0TJyuDnuHcth6zlulCC9ltORCgTC5r/n2qe4mDpE1XB3buR1sh2
aj0YMJyrlAOzeaaETA4QUce35IxuW1QJXlLE+FLxzdn2vqdzl7pq4Ew0sweFWD4OwQi0f8O94CNW
KgpZz3luViChWXpC4PgmQyLzsnrtTa9KU7FGHabHor7LE6p9iPLyMbbJxE6zqaLlFFvpSNW8B6Ra
rP6gL/l+K3R6L1dvUhlL3HbnSfG0W7lB5Iv7KXI7uZeF/p7uHmc+5RaZNlA7EwwOERHEWeMIPLcJ
btu++Bgdni/4SumuE6zUDRq+F1uyDpYfbr23NeM3GJV8nNgO0iitTLS/PN4QE4jJY3+S3pmX2/6u
xmcB147BQJCo6RdJoKtdA2zFUxf8UNPGxnMyA+C0ksk85fxXq6I7Km5SXXLvHwmPLzNb47w11fY9
IlLA8EdKZZpolfOZ6jFi3Bvx5NW5TZEYnBkwoqXw9J81zICMHvD6DoUJJXEzRl6+gsyTHJzVCZQB
qmrHw9Derp9VnTJB2+cBoaTU4KvjyIm2qPmFjvykQuRLI00Hgj8GIWiIIR1mqWVJ3iMhurrhWiPE
4ULo6F/D7AQeLmSlvAmOBGF9buSYzGpGT/lk0FXvaQ4qDcuXv3PPl8luJX8xpm0KhxiXPblQuS5V
hmT2XcXjS0mw8xDxrDxMeCCr3dh79trSdcFdoJ5++Lp/r9LIqt/Y9xpT1uad64q44nr5KrIAq+Pc
v5NY06rgMTbqKZ2L1B1WSO6VRFTHTtoaQTq+GTNoSrUVC6fqbBf7sQ4F2Zd/QYyhI7+r3TnYxNy9
CfXlht1sGWXjbygWBjLUwJSYD7CqSSeC1tLZw6ZJFvpunYYouxtCiR/XPNpe3jgYPZOyLWsYADjc
e+AeUv4aZha6oEIhNJfTPCF0zLRez3dKOk+T3wql8PCmBsVmSdTfiZ3sNvnm8b42NTc+7pPawvbM
MyJJ/2xLhFvLoog7ieDotHzHryQCkEgYfJ9BIW9n5a8r2+v0C/PG+2XzGVjbIcJPornE33uc1oYS
ojxXyWm1iEOZP0EZOcLux9SeZGLW+mUkyDzmmF/rMYIFILSZKChsAe+HBAgJAAKSV2PCCRCF0BYU
VKf+T9XlHtN3YpiqX7ZKdyx0p7E78QkQ2OTFkjqynxz37AxrJWivHCePj17wnF40tfT443gB/Tdk
SjQKZ4ITiDTT+J5ldcLL1fU3eeofqE5kZF4cawGIz/uIX86+pwMuvzd6ROB/6zm1sVncT1PvM/ZM
U/zNATsDJdFNRLxyh4bZPE/xiNKZB+kwV+rYTagSlOFTuI3U8md9CjvSVty6oMvqbAbhJ42jvLMY
tGfZrKteDBZjwBSQt1dktoRickxVNNlSq8ycm7l7k0XpNexLMpK5HyQFzxD6zHr1I/KhW6PWzdWv
Al5+Tx5YNdwnluvMMLzsKMY3QO612xwNPFNaw3G2CwNhOAnS7g5lb7iIb2cOQQ2yUxlHpu9Kc3wv
wYaONYFMg04m60J6S3U+agVhUpMnofAuSBDQTZEjf94Q1VIMuiO5Fusr/5ItIyrWccajEuXpJoCJ
tF15OUAhg0bhqkjJ7yWi3JY8chy9zB0Jtg7dlhahm+6i+ny4AHjbBzRvIpJ0ZJfXHj2N+0wM1cH5
7eBQMXTZHKfvPxRcBt617VktfqVZLl2lJvYNy1U48Xemft+W7Umf1vOT95J2tGavqSwH7xCxR2eE
db6XYx4oEXIUPaN/FHPAYceIoNgrPrawnrPsVZcSjoj+VsU72HtWZGLgHdCzjZWj9FiBQuHRXti6
DZD4QYHYXpOZ6xjgRSSUxdRpj620XKyrxzlXJPJBujOlZlo9bI307PK1HSNv0JJlfWfmH96+s20D
prMNF9h0wys/xWQGYd/RtpoB5ZITU0fTud3OdbhE0G3/8Y7IgcWMcgVpSrFEnKjdMyxQrlKS/3gY
RGGujq38QbX4y6oljathLAPgItSmxPqc7hJmMB18eiGT+VXh0s1WxH4yTjHUDPrYzaV6k+5ifrgC
ZJs4RpDkM4NQoSamtc1c0vfZL11pgBXTmd+nfr7j63qExvGXufgWjYmLQHd6dTSrr1ZoNsfcghvc
eB3itHjOeSnYifUjKfOJ/aTQviF57UuDrX5bJNlFPFgVmYNV2bBwDR7X3I7R4dzYKt7hm0JoJXMf
eXXmE13ztUaVskcRH+9H5kEfkOCkdbl8944TWK448MCmtcIegQ9Pc+0+Z2L5i7EqnjYQnZFInPg1
W4C6QpX2P0lPefjgrBBjVJJPnfzWR0UntpZZcGO9mUqhTo2TEZWKkEmiAi9FfktUv6S0F0tE8YIE
Nzh8r7IGuQDInpkpW4i4Cz5VVFZH9ISKiwoSWBQqaFXePrlGfUMRMSo8hMtWzox5xbStECY3OWvH
vHW4HU6gI2RF9DUTsyO0rH7RbLCAFx7HkX7PJC1SzBmNz3ULZNifSXbrj/zJsjD02u5es3aAWvmM
iTaMf/WHjWtsxfgi4MWrqMyxRx9qZcZDnXhX92UHP3GJIR59kutbDdNm26WE87Q62xorkZgW5J//
93dJCogojZMPYZFDDX2ZRfsEYLXIWHr+CQPstNdRl58kQGYKekwPXpdb22V1jCgmDZpWKq2X311z
jthtUNXb3RWbosE6MVb343m8TgY5bB+onZwJf+Z7DX8GVWeHG+3zmm8x1/yu9Dpyty5AnoaETj3a
f5mhLH3ky/19YxcBk1xhq0APm33lrN8NMSYyujamjTVVFJcMfquvKhJ23LJzhuwy8df8cJiK0GMQ
z71Dv5uVfPCzCDgZS9kP95nAa8efmrapW9qBvwUTcIvkAsPJNTGgZlfr3gJ2yM8XCsFIAnzSPcLz
pNZ3/aeKTn9Ws7ZG56vDM/07Q5LaZlB90TdpQtfo14P9pRYkDADdHRC41pvyeC/+xt0pBUKZn4w7
HkvoKvwW8Nv//EOM4Gy7o0x7los4MST/iza8n3Irt3l9VbYn5iVmRM3tZ8cwuB2cT0eSNYatyi4R
eLwuVIyq/MELzzUIcmd4Bldq4qIjoQf2YPqIF9CIhF7EDsIutxP8DCvRIgpMFfgIaYaleNmVq1QU
vSLvCGHZkADH9OzGfuqLWpFsWB1/bgoDLB8PEsqcCcJSrIR3O52+Xypn8O9iWvKfSL163NEnTM32
GgY0pbG/uVTPZgcjJKRKtde6vJKEYZKw3fFIRTDdayX/UFeom1zYIB6Fhf00KAa6cJJvj6f09j3Z
yo3CbiQfKrPnXMtNfFjtwK1xWtL7qTYBCH7uewvuTYKNX1iOG4khkne6byNqP3I0wRUiT8W3wln4
vrO4nzjUOfkJLj5kaI9i9n3XuK3sKVouZJaZ2OBzWRFhUeLdYM/CiqB/4xO+mjmAALGhGCKtDcji
GKLONtyNkJjVjnVFXgCtAeEWBgF8v3tPg5pa8b0r7bZ6zgTsogpZhJ8NUJHkoA14k+JzTszeQn0j
xm6KnltTbnyjKmxngTuloCkrF7isg9f2z1YYyCo2mKJs/fGZqeHE8EOlWuCGjcruodWAp2+MLuMD
OcD9W+nzfCW72TlqXpqn+q5iIi3CuZnxfg6eotBqbPirF4/h7JSEEPr3m5utidJqNnVclCOA7qHQ
HomeTW1VOFpNs/wShdy4KVTqwVnSH2DOyq4GU2SuCMEbumTWqvn0EccfiKEpX+tzgXFfTUahHuen
YNussB7zt0Ahe5lJiqr0hu2Frd1cR96/sgoH4vkSo3pB+4NmT4tlTZ9sqsu+lPa6jCeYRM6onDw7
xrgppRCmfg2ZxuKclLIUqQl8fL4nWBkarYxi4SdSSH6qrnTmWNOgCt1QJCiHqE+1BMIbG6SMVjKz
u5j1JlukuOc2wWCS5I4ThtmtWIkKWj8LPOa3HR1JyHqRBAHJllQAm2PkFst/3J9/3/U1gMAgalYs
/oXCDkbm41iUiugSEQf+Ern0/pgtZr/sGvd2LnenJytpUnHIyfzmv1yngKChhLmHUZG5frXUIx7H
VBBqgfQwq8ZdvPGZZXbbcPwoPO9vU3VMPPsb/pGSG35HxIQzAaIPp+tVilJa5cx4WPYdpSSfTKi9
eIsd9Et7neIxu4haPl5YFcHuy61P+KNUSnrfkMEO2H11z2FgqjWQ8ZetuOUgnl4O9cleRcPUCK9p
e2mrneR1njAZPanRUZlPvxRc1LU04sy4EAgM0B+08xQMxGOeIN9nhVRCTdFTdMcD6Q2r7baC+PUu
PAt1SiSQlf90ROd6xMXIbsgH4U3pCAUuvAr/5Z1rdSDzbZJn1Ya0srPz+1XzHJML8W7vksRrIiFf
MUkCCijn/qD4Cx357fT/HBs4Zx2yKi+chb7t3uALzM5LNhfuZO9ZJwdhpH2jeookVfzb6fEZeBpy
LGMDm550IAizjXpzLyi309GQtLpSBy+7Bw3zjA0PuDyJAVOPiR5UFNH3EDdCdy7Td1ODtcMBPsA+
fJ1LzcbtfeMIB34MT6PkG5xwdwe35oavVlW3LKhw85i1Qw1H0HsP9JxCNJtQvxHYsxt9M3L5O9Ad
XGuDHhKhLIqzFJC5ZYeg+VpMdmzQ0PFM7TIVQxdoLUYuyzrW3FdI2LeJ/dgs2gCyY0gnxkaVpbN8
q5PMqFkUkdd99qiHk9LO5TY7+L2+Rhm/w8X0ZUncrThWVUXUMlPf1xJIyqytlL+VgZiYsLk1YfrA
99VrzuSBv8rbQxV1y1b9ylEqjGqlbt7rHJnzjh4byesnFW7en/DTExRH9sSZzouqjBpWPXdBZlD7
mAOFPK+J2LQ/Zcxb6ihQXJDnABXLG9BjDr8x2+ovdsOCSHYfShweqOEIXOHSedZ+AKBxTgcLPa5g
Z07WQW5hPsK5Y6TTnjQ6Jh0dwNuiwr6YuDk7Jd+sX/AyLuvM6+Cj566D9YigbJ6pvZXd2fvMU4Vt
SNN7gOrpDFVFPTWqgq3g7xIP+v+gWBaeeIb4Hx6tLhl57/23lSHpwiCoocJG3BWZ5WRifwWe299w
938dOpzn8gnoz8xUeXW9V6uew2H/yITMIHWvPtoZ39EePNNpbqsRgO+jxzjJSYhP4V10je0NUCox
nuE0O2gH0koEGYymjQ7EZskDS1+y9CsMUTYxBqcx8zLs2GnYA0WkJ/k9MxqV5iXbMguxGUrTT96S
SIxseidwoXKPzUiiTqnc+US2ecMfioyLBnt5V2GscG6lEiLO0K7HWA/kqK7SRU6d+DF67o/OrFDY
ktgzubfrR+TVozwuDVe6BB71orYtrLAba2Vbwe+SiMX7IIt8IVIIZ5j/jpb45Q5eJY0W6XJ1XOt1
ss23vo7c/YxY9DgYS7sWZdcNU8ag+lqxSTRKghIIKvj3APoi+fWmK6fM74RGc19M5Q4wiavxu904
6zUPpRWh41rXgeqah1kkigJdlDyC5VTLEylQ6ak/DxzgckvMcJJ7KWDmLxJ1EadWhWF1BdaNknkV
lKrlzZ081pCARajD51S5/zzOlp3qb+1UFDmwW4uChr2ssNe/09lGVxMFh2H8jjwcGXCoNyz1Cjpw
oiUdelebQalryQTtI+koXRZO5HLSANAYYWAiwAm3Xbr0jI18OT3fNEhE2OkFu2FxVVUsrXyIesvi
iyLlG+sQHHcttsg2N/dOyPieS1VZw3RFdECaZ/nIiNEOW445j7jhNvF9SiIGjLyZYdN28Z2nypMW
XoxDtNnu+BLAVBqbyJFlZShaMEXmT0/+RGBCD46lvx3C2FnhlG3AwMv56xrBb6Yh4kimq8gpLoi7
pMaI3neEpWPGeIw89gNnMeMHYK8TO55d6cn6xHS/q1zvyxpQELVV93TOULeWZu+jDpoEzT2FDQY8
eWgxniQ/xeHXkeB2n5NZeEREG3h+5QOHr84JDFE4y1PUaYVE/rnXqUcMrBzzNhUmGfx5ViyRKReb
o5MySTyRu/H7DY4zQFzOpFw/fTZ8RzA9h5+9rnmN5Ap1C5Dswev/A+ZCtkAg/9npXCjbWCPHxVbg
gIvTYGVt3LzKEgLJaW1xWxdReWgXShgDo9Qc2aENv6Dtkh9IO4V3gZaeUG1/WKoTG5lW88Nf7nqb
qqBLqe3d6Js4/p4sEIpBPH7HjEjy26umRlYGZdKFqKrjo/ejynMGnf2t5+Aoc6mqoyanG5RW1rEF
83yrxecfPhEcbPn+bFvriSP+gHfHb+8x5cgHx96EsVHqJdaoIe4ScgaVkSUFkxghNg/c+pnwtVaN
q2MjGwTYyd7oE3HQS2FIOW/rdQUOPvhxgYvN1xj5jef9polHHP9c9cDHxvKr0BwHsVmnu/ykeNon
WGQJBkc6DMkkL56wf9osEFxcf8kAIGJZFOFvbEiOdlFUYhxDmQ93w/yQVXpzgRI7Lx6IKHQpdqC5
ua4M7hiUQ5iKcH06C/Hwsj1owdJsNdqeio7WFx6Pj9TTuEq3SSNMQzaGhQProMJx/0LbQ6NY87Lq
5Fw8nfACHP9MEFg62TfW1HnY62OLXAXWqJ73yCMfpl0TRwZkqg872tF8F8aY0P/HWor3/jgSc7fw
5jCbJhFpOxBLUCcKFAcUgxKadKdTZkyrB9rNewuOVmQJeUAn1dm24bEcvp+mbqN5LspgHBaSA5KH
vfy1V8OtuPk+3TW54KAACMwdn0LL6MHiWYhYeGA9eyzQpZcwxsYGudrVVCMB13wElX3u+VzHuRlw
qSjVE2LFbmHiviufEITmYgRRKdgYYxYCOrJSQFYRP3e6arYyq9E/0DQrnrmpm0SgoG7ZEQaleZxl
iANB+idUbo1AAvcGwL+os+5ui//WQ/ylfMh6aqepisH5On6gPdqLibSFpPU7rq2yQjwH8/NQdm66
RRuahIffaXWF8xU43LbOvgzls4+/ETl0NFwJ+zpS5HoXe8m8ILYJcLdBTXRip+NcfPtTYvrE8WAD
47noFsqZFJOdC2ncrOCL8dLo73aj1/ApH51wWclNvIJ2Bu8/DyZ912EAiPZniP9QjmfoWzhijv5J
UiFPegUz/lxQr55YhwAvKMU+DghpICAdNOdoOMnJwTfJ5o+btGiaPLMdWLnoAx6DeTQuEVnUKgd+
6HABGfE+p4bel0Y8c9nIczKBqN/3Jk3Oa+ZpvXgNDGmBW2J6+aostPF0A3b6iUuBR7zIC+sM3mh1
uexYYpfIcT8IeZnZ/48//zGvOs3ONY7WddcjJymSWrejn8u0drFeQPdoR0t/4cIkjl+bq1Sp9rM2
LF1NnouZr5NmCLI/MsN/6uH6UpT5QkvsCqGnCoRiRmbL60VLb1nEQSKqa36F5e3Zb2Evkj6fMHSU
RrCJxkPeFsIdD1GSEPANcfvS3OmmWblp7nX8Ta6jF7d/ZsmQzc/guc3bzbmMa+xUNb0w48cLJJzA
K0c0NgFAjoRltLq/jb0glwUVEU6m3F7CZ7dQGoUpV9OIy6wNBJVU3l3buMQkJxV1Bj1KQLb21c+/
8eM4uULWAXmagvKdq9b7JS3leD4Fo1BfB7oa4GKQj2EXmePaWVJf/8I3VI65ZcStphx4cRY1RQpF
shsRc3fLQNLJWWObzEFcEFTTSwerTUA9zPAdVZIZBthRQyIYXi0QQEwNpLgESfGp7wWRE59rEgGu
OYkOCIulFExUMlZt+8TnWIrHnQYvyxA+iqZ2SeqWzE+frZM1+Yel1ykeJpMEeB1wrpKhK9AH/P2u
YB9b6GlXDqU6KiuD0dQDJZHNIuqauv0nLafhT8gFn6/SXDYK9QNJts4HOFwba0D+qhUZEjj++hOb
fMJ8Qetwo6V0torcsyPYJcaG36tQbV972HRgyiKIy9kg07smIbE/M/COgu8xcnYc4nCl3EyKFOx1
t/H8tH09E6JybLBYvKS7BLlpy/pOtSovDApGTA9IyReuuVG7c+pGv/HH9Dk2j5YyC93Ow1R7CVyy
DX8KIar4pq6lAXSpQJ09zPMv4hzenQDTl7H/HnVDKPUyBuooM7D1x+kI5da9toum12HQHR79nLsr
OmyskM4vofaAQ0wRhn3EWUurT7PbgBDQjXvYamQbKBk8FfqZ+3Gxak8NLIDeYLPOhny8YkUJw/aE
G9mOu1D6NsPGFb4x6u+NrGdJETdMaGWaHm2jBZd8dkOIyZQ8OPGl0Utsu+M+g/26l5iBFH2EcCpy
I3yDwMXEEkQfZZic3tMKRG1MujdZylisyT3w9icCknMLBq6hjJt7Zn46VTjagjLngHfW74VagSIx
Fb8ezfZgAurA/ZfnAv70U0l2zExJdEhn5xgawsOWnmnglstZJSbOwIKusd+FE1m/FK1Lwt9Lv142
/5aro7P3cbCUQUURqmm0Ru3yWS3MZVlrp7cKTDLR6jDJfHveFYHnPnuJDxDjqjxF0q2EH4o2aZs0
Gapinbs1o6XCxRyC/vbLPzyogeC86sJAMukC3Xy7zeA6EgEw7Vxv4SEct/7/dPtS3GGPhWA91jq2
sSrKOdIHQUxwvwufuPZ5pS/g6xdaM+yIPIAH2M9pdtwHCT+0FvZN1iR+z/yTrvlSUF76E7p44uEg
JtIgwHq3CJ3APIN++rkKStSznEk9Kx17exjBimHL/0Yal27Hx9ejAV22bb3rpohyDlfF8XoLB+Pb
7uVKoXiHQwqYaSKv0z9ZaRSL5jJBiodxQuEXtoi4D/QMynaj3HH1fKJjcAjM2xPnUtiwMC6kYju8
cVsARddTpzbDvHOU3S9I7DKXHeR+OUtttIRz53dWCYUZ7Gc35avoPzBkIfGVgVqh3wMmDPa95qf8
t697itnUus1fDpau7dgxstFyUwYQNXBrRoK4fM0BKIOo8uXk/Fi50SwAuYhU0/H+dMJq7MgJmwBA
c+4veCdpYvkMu0SAjXkjCl7hNDdz8GLzjT+sRw8M4k8omxoHUlEAkpxq5BMJV5HGNDRg/xYs2Owd
0W662bazq3OU6P1TqSG8SQfoBeA+Yozc8viIZXgaeuhWBSVXiGhYVidJotrFORcuBKkvEHNBVyMx
4GaV4l2dIkgCZmoa5Vq4r8T2o9aLM4wLl7YUCrDFxZyniy5B1u4BbjeKKc5kHnnhzX7Rf5jNiBlQ
VnmkudUDQ9/mknkKpIHe7kJe/Q5wYLX2REXiJTutVV704XSRN8g2c7+OdDKU0MMdclF1VcBsU/FL
wN6ZNrbYwqxA9kzKlo2HCSyOO06i++/q0FA9Y9WXNDhvhg1cjjMjSf84dLLjvGQlyyJagfBC61pe
Xdrj3KvUgKPv7R9wOle09Se7KYR3zDFZrHRncodt2N3rdOVqAxbdNcXcd/6BAhW1fg1h4xYzgjpA
3croWGL7r8M3FvQtndxlNriRI4weJagPOmi0AJsS6XaEB2zO/M08MS/vgd8K6ZjhhOVVxeIjF4x+
TlVey+szweSqwbdxixoJSXUaj+BYLLwVefPlkZ7eIC2Bdk2NH/Vml3T5VeaCGFwnZLl0NLHPjFQF
1T4q04cUnRwE4rRg0iEo60NPbv9sjCYbOrCkeU92EFC2b8YZ/CDxrV/zIOe++EWok2cpk769uD6D
zO0OhZ57dzAAM3ycwFvxNlIeRNIFff9/lYiD07BvQ4dShtHYLKundV9eiAi0lz/6ftyEQsupyQ0u
Puwgu6A+lBbmPoTKbtdctQg6pzXAkaDg7EKPk1fIGD30mP+4D56VdBmgUKfGolUZN1pBhPodfq1M
s/HF+N0ASDX+ESVuLdKWINC3Puvngi4fkiNBAE9MSXC7FIUm55qA9rnuGSuquLHHBnuKiXOZeBeu
PXuxF8zOxjdob8cjdtN/k5vd/te0k93fM/nnk02ClZ8C2ebl5FgZtzvXVhyM+88d2WiT5VljcZvV
Nhy1PIKX8kE6HjY282zO9GAjm3KPbF9wKiN5JOL2Yv1bxX5nuXBCcbGF5h3bd/4E65WVt7pphEm4
V7WyzFjZUvnUGGxDyDGkQusuPYp2gEz82wXCOfSI699zm9NrX/ryFzZyviktJe+DV85ivn2rfqMJ
3TumNzlcnVlu7pj5BqR14yDca+pWxpefYfhJRGgnCLJACDLfUrFvXlqiPYPSF3jFQhahd+FZ4LM/
fPIjJaHkI/l8HWsPGO0r/r9/QO1gsQ1V45VqJvWD9mnRw7a8Nl5E1XuR+7aMR9LZFfx38xPX1Bog
sINisb/DRYEC4myf9jdZlRdhEMeeL1QmLUKZUyQyWqT7vmGbMHNSl6KNex2NIzB52kHydnLh9rBr
dyEXVxjhD7xVl0Y0Mz//fzvsM4nHGA3+0Hzs2t+NN0xY6lGSWcXpy6wLGCCir7eFeYGhTm57qsz4
qwAh72pFFJzcqwHpd9pfGq6/AaUvgDsIcIjL+jdNGzmmHjHdZtfs1Gspsk8sS1QGne9stWE6wEmg
9VlAc0PRIs/kDzDwUnwFqT5qqxbIbTIi185LT6n2EVTAaFZ3Kzd6rioYrmdVX/KY3xmpvwy+rESg
bQwMECUCgWWMT5nYKvRN+11QQFQF2Gf4vlz86un6AxYRTrAVfrLQVY2JHTkFYeKFVGhWz00yIb9t
8ByY8iQMeslrW3hHQKvuRonLqL6j5QsuymH1Dxq3lvrg2zFi9S77bcRfFL39+fbLrWvbIq9KQaDa
98osnDybtsOcUzzFpvs8iSB9m/D4vPc0hP2vaQnqHrrKOlgzL2+F9W5PdKMPxrm2r2YImExG/FvU
1M1ru8viwvnPPvju42pwfKpwfumF1rfHBGW8zjnLwrzVzvIes8vaH0yKOWmYiSLwCNVhifRd0HJM
FZ/lXo7LWwdGAzGZgqsOJpPGUIGtqkRN7b41Pdk058GQYnK658J421MmWXXfIfHg9KWaGMJrm8uL
OX3APNos5ei9wwbviiYS2bBf06tQepYzJ9qXgKL2DnLQqMMjlAd9LOtL4BnwIXsVTdaRfvj3Ga2q
sFE9Lyd09ffQvSUT/PkIN1P4wzkFWXcg35r/fTVd28YzMPZ3wntgvWviZ7vTR/R5Ov6ln6emfRVq
HCm4CMbQ0wcNomujl+c9e/g6LlGFVa6FyQzPtrzShohkJlj4uPYOpjEov6gXiWID0Ol6NN+QCbVl
UNpoAQkIQZu/Qsl55t5DiVu/dW9kU5c5he1vKlid/uoxHmq3IrnEyHWCz3q4X/8z9sMJpVvDUB2/
ZOH7oF5Zv+eNjMAQBMu3dThe5TZxPE+kyTAsrHm+o73PbzD3LHJqbNTy78gd9e2Y/xnFXYXP9Uy4
qAVnTSWA5mz+oEV7KWOghiziBzGjoM43lA222ufdC18aPOX3IXBADLSd+FJVsntD9rf1THyDWbXI
tElmGKzZWS2PwWDi0MmGcZTQdPjDjZMH4b7w1cuK8Q/G4YstKJ55eC53JtuePqR8blD1ihpXGiMg
3KPQljXnbAXOWPR3oHBJrKls5Z+vDcd5Jd1ubbt1WttXpRX2EVVwCetNDGALHPAEMJ5jx2Wums5i
nP37luOPJjgrGTz5D3kK9ltT3HTTxU913do85knDjCT7rYAvQcX6UEsiS/e+/pU1e+vpONPWbGIT
WpwRj8nTh10++8ScXpGimHRRrPXb3ghRq6+Pnt7mttpqYXGcszYNBgdRKPtVCgdmQamJFrpp9jdl
D97dSCpea5HyseEZbtO0yCMPD7uQNU1v8lKDad9FWC3ezssPZQNGvsM1RRYIWm8aad6W9hsQe5BW
67JYpjM1dkmE21Wq2fgUQ8cUfuQTowFyXjqvIZ3IuS0nPoxHmaIy4INe3o2b6AXk2YNYy4Rz4I6z
L3uDyQ9Jk2TLpdqEkBfX+0NC8X1uXhWcTgGImMRPDLem5iCW7iBofjteHFNnISLq0ug10gNZpdI4
mj37m66bCssvxguKlsfI0+PXCDpO5G46ZYRkRLuwt5fkCwPWsZEX8OUus01/tiNbnGbLu64bCjrd
XKzRV+F5pzl4GQVHpdlI0o+zSpKtR4yH1u07y7wLuEBgiNNca0WxX/AMKSlNwi2OVbzUWB8HmSA1
9PHucmvyiPZOo7UMUVg6VP0pUkFKkQKXdrjwwUjsioe6ekCKSvNUCeLl2zBTJLxyY9na1UFPiH2/
YhD9w7lgg1/AV7QG0u5IR6b3/JRWbjERMVTwDdMKlsAapMKLVy6GCoIjyOE+YS0lsDgySOqIyRvL
Kx4dYEZSwI75x+ogtBSf3zb7yaUV6NmFDOK56x9EDPQeP4j/ufi/F30u/z6+yWpq7B3PT+FMiGmC
gv9k0WjV5pcDwP1nRHPGK8hDGx7vzN0X8zGUhwbJH2j9LJzljJx+NqiCvjviyxQn2V7GAiqdubHC
AzQEaDFXHg/nQejCRrMG0wHLQEfcl0XmzNqnyCMGKhW1XAgD7EL6IcoJAQqgK+ci4DUABKNGbueB
wkPpyC5qqOvxDNSOdI99VUcF7X80GKHIm3+Zsa65LRdFKVBIb16e0HXgDZH5x90RazxIie31L7Eh
z+QgVmVesib9F0Xx3neU7nBl0ZF8sGZrfiHiKcDOdWtcFbn56TmEx3MIwWPZf/bG/MoCfvVTPFZm
6TpBSP8FJtNEUC/qZlvbul9ElD0veE+kx7DYxiUUReTQ5TgE9soSgfTESVNROzecc9UT1hbwTX62
1f+Y5iSYg3QBe3As49WJ0T8kWLZmnet/Ew3Xlp4PxOwprmE8P4Rjd7rbZsbGRF/f0hCOg147vJtA
bIdMgpwtvcn5ENY7ftn8Wq5qlWOYKa2CkDTt586ySxJXOpUWaJMI3opH6Xij29WiUZ8MARb25Lmk
D9vTRhKdIHKpZX6pa9CKesnkmFyE8C9BAooSYa35SGWe3xRE1PR1P5CvVOABikJifuuM5rkFpbBw
a2Zvq4WeRghvb9hYYNqiAbmwfdrKBnSVctLl6AwCZH7R91X92qCKDOW4b4q6uRuWB+NylpfFKcYc
MVQn55OCD13mudy53PpEhVJAqLPKXOIygoPt1oJDZg0Duk6BzqsKBlNxwS/uzRUHlvq1+MOBcd9d
YMiI+zPd7l0EojGgICdFi042dwAXhdLU1xyTZ0AE8HwNPj4V5NU1qCJ1r52Kq9VFylAzc5dAuXWd
cEbFS06CvmHa+JrtjL0uIWa26b+GKBJeAGTXQubGCgT+hk0CP1lH1le8wl3wxwySpj0nGgOwwHS7
fgtdKTFSKXwclf8pCGN2hEzvaxgLAkpg1PG/6tTRVf4uf5RRSGQlRE54MlL1apZKyD5bcAdRQ+1c
/3mhhJYMoNViiDQYMU4o2rnquwmsNdbnzp8/bEppBk+X1o8FuNh4pPR0Jlwyrrdpc/9Y6vqjTRgS
04Q8KF4DVUmv7WOvqMtcOdikbb9dKN2utm/ybEIunXq8NxQudaLS8faOc2g/HBIuccM4C+5sOSDl
II5aCzghlHdS4jEh2eUUSIl2/hS5+t4ZBumO5xFmXD48jM3BLhAHkssE8EJzPdAeN0Vajq6UsswC
DaGYdITfsbrkTZO8/AuhGaU6R5u5U3VtVIA7AJHghPFq7mzn/w2k97nruoHdVNP4JS+z4riigOlw
Wb5hZKVpdYpwVDqny0LYPgJLw9W03T8hon/y45JK4rTXfThHCq9G86jZZJXjMk/MTjhR/1OxTbQb
j5u4+So39rjmaN4/SoWOfohJ4WUHAKrzhaBsHgVMbgYut+Cr6zOF6xJtEfbfX4QgsPAr3g8RbKAY
nMxws7Zbm2ap4+6U7+HlbXPKUnUoD9IXAuNLOSzSw8diXs8MbYAgRFefPNzuKuB7Ye2xWyKXczf0
TY02rayK8b7BH9QjYKFZjWP8jL8S93azFvjFVY7N+n4HTpDPlFXocyFptSxjKXNew1WFbz6v8A02
OScPFFIzD3WaqmDe20hqB3qein46Td576kBi6GmRUq28k4VoCUOMy7WW4E2TsJHKV47ZE8iJgZpn
8MsUWqFUABBepGv8bBYoqFqwGbouGX3NeUKqyW1CIndC92Uk6x7v/TW8EdZHck/qx/GKKWCmuXe7
+8q/yqkRpzXjBnoO5Ya6FHF46DDOLvczKT/DMBnfimsFBIwYsc/sONHetv9fJh0pMw7sZwwKMEE5
mI5yxLHoj1+cVysyxtvzvyXFsJ/xTX5LdXj0iOoACXWJPnyLfFL5+dTGjqSKpOU5NtbbP4cWDV38
gLdnMpOCYfkc6hll4s24D7JGAJ8ofG3q0MQbwe/GmJptsyFpLpgznjpujVsVzX8/17SHsKYJlMA+
ZcJIhLhkgrwpsEtJF/9NTf9Wu4TNsoVKqjGBFA8iy/GBQojZYNKdeNlfNsGIiDYh5MCwer2aBZcD
Khh2YTEWc5tvpuMlQUjXK3nElm5bpjrQMSOvn24p8lZnlq3+p6PYNEJnxTLPias8/Kt/AgVaRVtZ
Q6PU0aSnNK7IIfXqTas8z/Q/oasqGB8S0x0Mm2ly9FIg4TlPTRWn37pvb4BWI15qxmans9rmBeWI
/0BWrs/WjbtNNvmRqmxz/GkSLSeMrfalAzpHrdb1LhGK3eXv9P+9uC1sX+qTzXPoBRY3Fh7zY5Hn
hn8HLy0rr4HzH7UY/Ip5sVZmCiiCLSCPF9e4ZeNfb7AM3CPYiBItBzxGiMRvGgwC0O4LtR6sOE58
0yJWUiQLKKkBld1bDQ/HU6qLR0inZvBvq5C4xNISo/plRODrHXTObVCAa2vPJcosbbw4/8RZVDYB
j7XIJz1PxxL+S+A9KIW8cOlwL+CMV7NBTk9m/o5Q9CJZi7G3BZLrslAWj4hzfNfx4W0THreQ9XZC
dMckiQL1qTCJwp16z+7ehkPPvpxvvxZSC6rHnOVd4L2uug1zPf6MZRvwamht+wi2o4l1KufxpB3q
FfFyz50i41lXb612W+GS4yg6Al4PRMKt+BnB/sdv+vHKN5IDJQsfzgpqXvnSu3b5GQAxZn8e9Zhx
vhorf68zarz2BqZM9aruCz0PtU/j3eXLvxKl/z3BU3AfIeGxrdPPcN/9NMbpdBSnM2ZR5F2yyPmc
KWunKRF5HK3oiUnh44mws7+MyV1Pb82TgLRnQ15I+Zo87bAeuXRXJ6Z7OuRefgGI1x1m8nrADnRA
JRE4iT8o7DosziG/5HHKY4PF+M2W0AnG0O3xq+a/WGWxlRu/nGqYzvtYqUig3SBvdf9pWTnytyfH
vNYxwTYvwsyL7Evd8ToJKpWk+26Z+F1lAbKxeVNbMZywxx138FkO/Qz+BSWFzFabTbeOWwyEod8a
s1eBCCBstYD1tn3kDlDQPoTpDJdZKz43sFy0TTDj5a1D4rXRrfdnTxbUKqfgsKI94MIY8E1eyTY3
GkNurvZM7HyeBevaybZ4YWf0FQyzRob38CsrtGzeRaElntnIX+E1v4+N3EDX5/xeyY4GUBWaqfZ6
VR5fAtAli/t+VzLlE2qZM3GtBEmJ9EJ2SOXcPUloKRf9Tq3/Kc+Lz4BD9DtMjaU6xXcaZ7B1vhw9
amfEoh/4dyyTTgylrqac5Z+BYYFRkD2lOJNI4l2Mp8HnUQhYJO6X0xrzKJI+0iK9dMy90tMfTeHK
SfYfVWQtm0DAsD9ldqLDha+7qB/KCzr6s2EpT3tgCJwuItE8lSU4V/uY5kVmkZvFKIlGMM9wiDMA
hjPJPRV3Y9xRLYRalTF6N8yKQairq90NQHFTRt6Wlqf32js5iC4Pl4fs8n67Zqw9zjtuKFozy+Wa
fydaGpVjutfAas8/p42nDNpLy1Cl63XLOtLQAm2if5YojYP3tD4Aglth2Nf6OJKV9pipoLsHiEHm
XnZ6DiCt/Y77zhLSVt0SsDUNfr5nGYNCiukqd6rT7CPT/9j/sCcPD+x+PQ64W3SgFSkh0uLSDk4b
w5lDvAtvBrPAtAu+1g9OWVrFnRIlWUINvAYOIu89bvQCoaVPz8I1HFin5dduL9sN7jRw6cY1S+c4
gz0D2PhmTBgfPl2EtK7nLcaGzaS4hnw0RpuP1kYkZet1kLribm3+NfBpmfV3x6F/9FQRhwnbfHIp
wKt61kdq8+zWpcOvFyNvsVKjlXWzU/4ga4iV9pCWO3MIx+OQAjDM8acO8KZKIOAFB+iqCmagDSeK
zE6A1owY6wxgg4baSSJZAHaUWwK7QwzmRBUkPRaQO339M2DWYoF+OSjZHVy0oeGakGRvQu7Fk2CR
Qeo/+m2rCHdeXeybnCzJVw0I3eLDXW1utdPvvsqvtTf488cM4aZh4HxSBVGEre43WPUBURr39Xf+
mrlL4yJxhRvuQQH2mAdNGLJwzBFKp9mGcJMhy54tsx0BUAlfE1fvkR4td+izLmG3byP/mPs0yA/z
1Xu9GA0QA4soyogBHJ3mAk010hjSZLGzsd1zUAxMpJ0GF/XryxZMUv4Ap0spqqsZa8sI9aJFIxpt
yCkAu8avMQX+moKKymYhanqUSOly/7ZXJ6nVDIuW1SuIAazn0mvw4gQb3ChKMf40S+raDSOIQIjO
9cwiMOkdD9wAIuE6HUQbk0OHaLWiNttDbrlFkaTPhjGM/9v8WhHJck8CPVgkmhqldexJQ6Fxwxib
/CuBk1OvFI+3NnE7nT9beeZ02ubVZlYhg0dNSEqHK4CG7XIe5mt+MRPhVKTASntslCaTcVYn7v+i
3+K0LHfWo3OskkowBbgXcgu0MaABO/NEsIesU83xWjAl+MRM8xVCjv/dBh/wQ0bVmbqBquPuYElg
wHHySrq/RWurJ1D4u4wtNIbWq6MVIV+hOEo2A6eCpI0j4YAwEw8TY1Gm880Y5/x/diS7IVZnf25r
MprIjCq4ZuPlvSIAOGoFO3V+M2AkhSaBLLYcJEIrF1PnYJWLo1DUE9Dy3frMAdXd/NfPPl6f2a2z
yjuYbbkYOl5+NO5UK16K2eVibHG2+XR6QGEGZJ+qnydLHWTGA3rn3OswHtkSBYRRv6DL+eLh2MXY
2mWFZ8cqPp4G2Nz/BzZWqUm5ro/XoAGQLTHVFX1UXO3Ng5Eihgl5oNibKbxrPDMOJrluvENpb7sj
seVwpEGeormhcT4/V8gzhWVw5IMw+uKlkxKfiYfP9dY7SjOLTCUrcQmH+CvGx/Xk1xXTtohMoils
mNt0OV9LcjHNmbkONwPjPtLEZ7uHaK6SvgGbufc6uNn2APZjKWp/q/dycuD0vW1KsszE1+GdwSys
ZmYpy/xbNlhPn/Wv6FNKtTm3O0WkrpSiVx2i2K7YD1+h67UKicCU2gB+tXaL4R8eim9v8br/V+6j
TUcH2NE7ZRUXY0ZXQvQ01qsM20K6bsg+Jcguxnl8PBiIJfKR+nQEFhi6XLPP2v/Cj3icPXBiUI97
EXxd4TovgVOmUQntiffdV5p81Es1p6NpkWpK0xycKdF3g7CqHQswmyvjosf2E2OmftFepEPnVOnn
oQH8/DBE8SPJBQNKe4F+FgRePwQuEz6o9j3yyFGOGMEsuVtQW2dZBMxWXCk2KmW5YcM0H67+srvp
euR5SnnxUKN710JQZ2erfIa9ZteUcy5OGyexGjbwFOhSk8hhOJYQ5f0YPcBqYUlrqpMalqt4wj+B
+TlTstWaxAGXcMdoIIpqpnLTpsLkGhz5gmVxVpUujoPIuaOUWWr4LMWmoyUXGLFjtYoro3Q706tM
9/Va/8FBwRDP7TnpnpmubqVHYikU0ufTBQSdmPXeksPlcWoobVmFQPoN5fmAQ7KCSJrXj+iWaQJt
NhNxlaB9eoiRnMxm8U5NogGqYhDOhnoGmWbZlK5mvE8+0jVpZiCb9UUQdzeRppgENi7Vm/Ne/9ki
tHwWhov0cE7b3MYrPzxQXpbeG+pV5mpeMdN18DZ6fs6W7uBCIxq5yy6B2hEft8ExlUx13srOO4RQ
HQpi0me0DTFDRdFjxnNFBf18AqqFRapgbuiMLB/6lKG8+gMfaYpQv9Vyx5kcrC3HRHTFjCIb+M7T
uGSpw/EP1JqFoGmmN7ksv9LWPEqI5FM6mB7OytM6o9XqN4Wn8MFDw/vWD5Mi+Gi1rICv+ZyhFOfI
BEVwS46leL951C1fWobadl6N4XwlXiKfa/NGFDiab5cBOVmnjtSSwNnVKcpXjNiCTqaZkuapC3Of
r4IfETrm3ipWA5V5phJ/dXYU0Q5MO4qSUUYhyl+FD9jD6Rdg/4CITmiMLGwzHXfu27CMpbupF7EK
Iomn8JWiTbGsNPPa1KnFq04DVwQxy0yY3+vuyGJZuZibHqFL/9DWGsbyt4TZZyKNPk6qgdONPLZh
Hh56qvt1iPb30JNKfqUoL0ruJayhZHG3bDMUw8RRS5A/4HU2SfzMq0at7RSNvjHRldRNHMSrcKpy
hPVT3wYuwf4S+RdHa+cGSHgORELVLqj+0OWz/qlZXUU61vkLIP1vmmTnHveySLDu6E9oYhngoTEB
JUoKxE3w84Ot12BVRnmXVfLcpzK84dyjzaRJxXxeBNLzLyk17YryddR6/ADxi1ZhMM+tBpx/0ZW1
EsSHmQZhodtl9rjs6tQXwk8CVTH6KiXLYtX2hKoSAaPvYEBOg2Bp7NMhzdIPdxoGlFUMViXWLzVS
rOOlgL5kA6uBjlr7y40oR16dM5Xg871l4AtM2VPoffyBxqayGjkSeBxixL+T7V46gJDk4PB/D4B7
wAx0QV+3tlyW7s1BvwEk1FjKW8e9Skt9OxKjHXuCRAVQT2VbfOjBdEOY9XwFfeUfiIcz8yt76Eke
AqA7PelW0y3UaM4ygU4Yb6XGh/Yi/+0CkI/DahjuGKGWKW/GDNhd1B2tHMrioGfnRVBhoU2AOVZq
6SuD2dKDotLZBgw3N2q/w3af+b0x4c8I4FaFX/jPD9rnJiFF2nfy8TCWaChGeyL/RhfhQE1UQFzC
1Gihu+C+zqLAntQ6CiwWkMY5HgbvhZBHTZAQpl9w/XaKA9oo1+UR6+ddyah/9/IJDLmYBwUOX9au
6HQGLzUhbkFpTHMgf29ZYBay9G+GKEL4U0BtF5H/vPELNrDdEA5aZLn/UGWtPHLCFBx8Gij06/0H
GbiQ82v5bKh1BzBs+DAVoayAo62LOIbE4qcSPbFuq/eTYmYMG/Dw+Z3rYqJLZf6YSnqsShrtx4ZJ
JCSMPNwKPTMdi9alfS3taaK99ADx5EwWXjvNp3JBmd57Bg6RUvzon/dKT3jB/xKHJGZ5oUGFq+NH
Q7TI6Mn+tO9sqmSPp3k9QDCiXFZ/GfVFDiuJ6gf6mJ25ppi1/Bj4KY/6s87pmi9tjAS0zK2UNqot
n7IDcZLnVCcwIdZsvDoQPIwJlZdXIjYnSgh1nkRDX9fwrwaME7OZJ2FgQKVr+8/CaVcSWbpPLW+d
pasHtZS78q7ra2uK7TmMH/geC6RmsotHRkml5xnXkvK1sX7ZLoPwxfrdNWQrTfL/RH+axrtLEoW4
nCe2iWG3y3RS4DvRIfckdO5pRPtEc+3HzEUA9QKHlkDQb0qV7D8Zm2VNAkEpNcNgaMF9xhpJc3hY
d/W4euqjE3IeRXmN5tr29L1FpDksGSPU4OO/J65TthWDr9DFregQzrtqnih9kSxr3r6GKvkNEwQf
QJrMtjLYG+ZVJmwsyfvwzL4M9Ts343b/1OPy4kJa19YbN7PDEHtAtz3lAtUn8VVHdzkPke/y0mfA
2nZFGfNT8jun6mkVf4KR/rt5IytphRM4IJrthjLW0i2ixQ3itz80BsINveHYXQJa8piaejbLIm+y
UeUQxZeHT70Y24RcmG+6xRmPNFC7JgwCw2tOi1YBIkzvRV9Ei15CHWX/gkfE+0Ygq4ss3HAYkxkO
mWbruv4SE8b0rS1nO3IyvQyQgh8fJlgHn7FL5EmnbgR4Gm+TUWyyJieo7/H511OEAi9TyyovdRF1
jFvmX+7NSAmSLkfnp3myR80oHHYI9CWcbcvwDCGZJeW56+TzFmk4dscH1kUqtXZ0sOXsd2Tr4pWZ
ZxbwC1Lwr4UQoBxla1NIUL6T8/DmWQtrSRnYBDwUZUUBSQb7X6iJ4fAA4WTG5VBiJytZra176oAa
sHS4Q1/vvxKxbsI4geHoLcjMV6HuGMlGVrZVG5P1dxi4mhWqgOTXOcsidQPEHzd+JNfZDcDMo2Ar
ICkwuPHIU9EBer3TWx0BFsrVN7kMyC5fr54EXy9HHQ5TZpjl818iG2VMqIgeNZe+AW9aAid65H+z
G6itNWpfBVO05iBGprwZAF9ykbPNGZHsOK2xdXJlkUlqJcjpaeXyH/G64OHSy0o1YteNMfONKVUp
OwgkkNsf1dHgcGlyMyY5/bnNpo5AZi0+6rnnq6ACKLKdm600Jl7kcNsWWUybxWweNpkzB+l73ezE
kzGy+/0Hzrb5x2nH8MJJhV3PmV0sGQY3UGN0AV2QhLYsPl4/RAJWqQih/Wdu84WdAGpDHYZMfufO
iTmF++JgOvzdpMGqyjFRwuaB0+gN4Z44Pvuiu98xC+0ipAblfXHa0jNeeIwa8sXasG0OjfMrcxIz
H2VJVJJAp56dE1WJiFJWyZEVq6a0Ie4garsKBCiFTSSzlnBh754+r71DnL8QaQqY9AW9WVmdUZiV
rl5tAipp4uToB0lHK5T/5BddOesBCIwv6716JvHqvLDeY8zm49du3AnNuuZ1DLS3FwTE3rhfJ1OT
8WLKztxGzcJQ3Q+N7rSfZ06QFOoGrxlqO7FlGQFhdI+gQSYpSIff9YIH0xhCvIIKnYkv3tmERih7
FSNcLweXa+F00Uy89WDCFuyknE+VXy+aaUhv0M0c6H9GTriEePJu0eHlxHbzDQzAfENo2nk79W1X
J+vkiHZFN5n1UwOEIthzdzpqWOfa1q/K2DWWYQv1VBjiTCIHkQzGkqBgZsLaGq4lYoyrEExuQ5vc
T9Nbr2vPxUqWqsz967ffTj6vSw72Wze/TimQuaTJqT7og9vkp0ZFffA8xL8C5gCe5+UcSNZ0tLKZ
tJ0CoLRL62rYR7qBZ3r8p7Hu4UQ9rDQHyp/GYIzxPAEHUzpVpU9QkYPdxpITN7eKPj5ZFrp7KrKn
OXw4cvdTJil93c7W9ppijF/9vwT3/dkTGm4muaGADRs5TQyCrTX6sRl+pnUNPch2zm+NiK/Ql7Fi
3tRP6zZu3vhJcKdeuwrtwo0QJQkUB9bHnQ4wnOYe/mkckrD/XOVT4mCrgJ1CZcK08rXqS+yX4jhq
Jrm1Wzzq5BgQ83YG8aqNaWLyvMOx1jgdiNM0++UPlPT7HH3wZL7F+E5yKNt2BqfDPQ9DsRqZey6c
BWukpvuNk2AU+cEd33SNCGcDYEGwDpH4hK5+z6jGtAg44gzbjb3aaOjeHZX3aLIUxBTWAM3vmrM5
vZOvOqHtHm9sKYnNRmkOe3qtUSEn/VNrNbLnkYq1saBZPsYAwK2XGPioy91q/6WONgRfekT0Z3+G
fkQ2NaRTD+i+CXN6gfviN7flRQdS339TB/J3JQaeH5vbumvZsnlW+pPcg/NXVTg4FLXaWh6IFI9/
a0/nDOqUI5DxxxO4n4h6I49Z3QRx5rsBAljgvGc6BNvsriw+c98C+TWuH6FX6YiUq0dz3qPg4QIm
gtPbHBP249OLOhIlgFAjWCXyUUwDdRwR1TaJ/lyjuilPI6MCuHmCLA83ao+JJ3d7qBtwcRWP684u
1mjnw9HG+6pHkDBuzrwZAOBktkhdRAzU5fFFi6l55ZGld8m6w9mUlWjOfLC77p60x3MMNi1Kp0FZ
mv0alDfVojwBBfzZcEjLR3OHwjDeiOAzBL0HKWgGOpCjxCz3VtsT60v2orZofV6+IOTCmSBuxf+k
e53xYO/vmYCGhszsqI5gM5cE3poqJgLqmAe1iqmKfVhDhGOmVoEmCP1hy79xEp53lLFpaTjHUbvV
nSESvXQdXvY7bOj8oQ7hJXdPP2kM5IxD/HWo/J6YKErcV3cCeBsf8KveMFqbPT/NHmqb5FNGVo38
xjEmy5WW11ZEKm7XwyQyWxVrU7mwyE/ROArH0XbTRIQL5l1TS+2JoXQZgnCfp5eQKVyc78EpRc57
8irbKgMjHN93/tdaG0a+snh7lsWf3oR7+ovlieLuV8nuTn08DM0ksRah93VxQo+Q/SddkGqnCbwS
/9UdX3WdK0tHlODKkfHBwXXVIFErDX7GVyc9r9O+5LLMkYl/KtHb2rxnScKrsi196YZsbi3p5o2l
Qnm4VZJBRrlnAuhpqzIv/oQ5IxD7NZEMpwTASig4UTikveXSIgyptTGb9zpSMGJTUoq/ZbOzgxyD
N8oLsYVm01wB4ktoNF8ES/Q2dPfjVxs2ZTNTHduYftiLG0ebVDkmwEG1K0/76CDyEjxD5pkgD4az
kG4kRLyMvRFDJH4rDshjVPUAD6yMEAmobqLLWtWY8NlHXmdx5ZB7a4FGHrMhw+HcYrpguSqDCTCK
U9jJi98IJbmJG4XKImz8lt26XCWwcw+V+4X2seLAjgVigmoJ71XQZD6j9j+lXdWVZK7bEDHRzspO
FcE3rC0K8VZhg/Dkfx3qredxyMtdG6H1QtcptJ/0eqjNO3somb9E8a516H2GDbT8Hrzwd7Iq0pYz
yNuK9bgsEutr0SJRIOdApFYtl0bzQktgT6dmK1gSJfVL+ZoSlWFrrRmaS+6zEhWOJC76Gl2WVYP2
eZy7LC0hFYvrGI4zj/wRK2mznbFBObewXw9WLzxAruGX+SCycWFEiYLleKC+68hyxhf/wHJRLuME
30UiHh8BdRPIordRxbbdg34tCss8Vs3YuS2HcCAlXXiIz36NNRnOP/doF6lUlq14bMNKaNeOxm1u
SvbUIOBWo1hJBgZVlXcafsBUaJpLupccXCICqX+uaXgWV0jV8okI/Gu8frgrFAYNyqNArTNyoe3z
B/lrHolMdSlkTId9UgbRohYd63ABtDR0t7nUKLUvYhfm+WIORNhhoIygZ8WBsaWBO2JKoTvt9nsV
4XeFWfood0qqfk2hSFbGPuTMcE/xaZ9c+9nKyWjUVGPiqE7E2Xg/IhZtEZq8jDrGQRLor8UtS8NU
4qD7y3Z+5by8zfIE3isyBgVFmnOkdTTEm+Uhl0PnrKWWiV/NxzbZ6Rzwi8PYpFokHiSZOZ19e/jz
rBpRWzmX4FhT0VvGYCocDkbQoZ8m8SZJHJyJuTMTIbaA7IYN3887E86SgY6H8tWri2bJ45XkRNlK
r0K5mZFYhoZSiulNqO7XNNQ0sHmrVBCYUMS+o/xprnCJIFrbeLUMW34oUBQapejb/z63ALx4MOkd
UYuhBi0mnHfbVLPXSz/ZwNlPVPI628yqHWvep+WoTt6CJlkduHFKf5sDBBu6j5M1stZWclV+dC27
0mImw1AMB5v8yYtv4oC+StAWq4pzNy/6937PkwbvZHjzm4mFFcWi0qz9zX2bVpOoVIT5nzGNYUgM
pKDcZf1kSmwRxY/PDFf6OJv80LVaLsYuUs6ch6hhrE9K8CQBVel37MBINauz3UaYE2BcCG0rxDEg
cuIT0Kl9gWoIAi9PP1qKz9s4ZDdjIpxM7Tq8HMbTaRRzZzlyabF3TI5ldClOvjhyw6ljivOINxJM
oOioUD1Ui7OdtkaXs3/878uY8aBvrbiHJ8gZz+o8xpYPMc7kNO5GCg1FrlY2Qhb2Kiw4GrDDIN8r
plOC7uK/QCONMWYvKc9KOMZHtgLxgdEuKhin2oYrzuxX6N+hOFCdRmPZd510877s5/5zQlmIKGFL
+/4/FeA84Fw1R11Sisv0GNb8fQq0W4EraPNU4xA7R+SpO9/evgmCy5exYetKkJQywb9YbWsDRKdd
RVI6XA7yvZYPzOtWJgSjDLSHzryANfANdBqqN71UzwElN97Bu1dB89dBqmm03zev/b+mSEKcv2bE
CdWG0hrINaiHhNIHo1Kq72yS6qiyqFjVZ0X0F7snDBNd3aQ4+JTro+QYGBQZRZuLUE0NtVlF8aFM
WiziRnWynDnfC+R27O62sVG+qIlkLvyvGiJCc2AiI37xWDc/CJYWS0niDRszhDHz1RhIDfhzoxz2
wG3XLIRL1lZ3PylIzUFCJZZqbng6ASkoMHMF7U9QHg/hPdc0wir3Xb8xJg4+ZcuGNFBDkmzmLW0O
3EGdf6/09ei7ZKBDvTNex41tqNNtmmi1isBZYIz7TsW61GO+G8SX+2yqzeVxsh1VlSIAqg6WOpqU
iXi1SRixilF9vkzpgbJ6TGvz3+07bQHSvvNgmclnMfoJ+Y0/7KNz/tz36pSkXvYKNXPoFmra7Ztd
ChGkwAE2P+BpF+eOnYP6qLVTI1H+cYsVuhxUSr9J9n8tpn+wNroqps/jOFGZ6tN3UuOGWq67RgWD
Zvr30f8xK47eSc/Hu36maUaTj1ob77nfnAAiAJGMIVNTCIVj5pQMw6fPJQ5E0Aqsl+Qrh6IGFI3c
HYKA15ccxPQLEQzLwoQ+1gLzvdOQqCGX/Equ8MnwwCyGKjkXDtI/BsBwk5Lm0Gftrrp0XqvJuvZZ
n0hRKEHD/k+0+5PUyeWWTqcRb7Xcgc2dLtlilIg21nIdUNP3zIeUKq/whs0D9vYgszl6HWfnEJeG
vlxJ+0ZhjxyR889FN8ai+QhjFIE7sVqufFAa1H9+WvjmOzTllixTL1BGdnS2SMXIefCyDiWkOgnx
P6QozEUYvy/I0otFoJUTBhsI2ggr2ZR1vRgYBBuWEw9MHTDJA4lduLbEL8SmlMErQeQadzgC+OdC
LNBa/iImLQG/m1oXguwT7dacSNq8k6TvHztRNcpI4mNUx7Gda2bKRptEk30rvOvzFX/7TYYWYLwU
bAXLp4Y7SCl+8J6hz7RvXFyngxp/6r3STJyjxjvI8ySnRH0BPI7+vvCPydaiIdINF8Vs/Mra0yvY
0zM10XZ1XaCXFwUDhtenlYRfTVP+0gJeH8zU6CrfYSbnrZn9iCD7jeRX+Glt6Zjtsv3rJ1ZvB9/C
g9DEEdIoNbX2cSHa8oRSiUmJy1P4VrVa+5K0Z7BwhKYwl9LbOFc4ff/O8bU/4TWpoFsyMjVtt1M0
fk4OmJGC0bhQ/RcfZNwrGvVo8QKsdfEsT+MNwv1exIL5cXMX/w7qKLzZope2eLt4yDKylWP8N9s5
dy/Yk6IBLTL8us2HOJCkKaGRKhROIdo0RNwUQKpHdTOubl8iJjmFPpvgbW9wE34TVMz98ipLIOBS
ZYxAd5suydHcfSUGRz1JUMLqtJQxl6xK6cRpfbqijjinh101aQ1gKiQ6bS5ZavwSBYbNCM+xrszh
pmTRDxzDXHLSSj1TSlLJGsvMdwAPDh/Tee2Gp3ITaeF7PlUhX1ORdjksSjJCZ3RdapSF8DY5tpLn
Ri+5+0+LXhQ7kKCCp0gSjTWXhKU8Eay8rPVD8/zMK4BD8W3CAxdJbjY0Z70pgbUC1Kpb/8NXEv+V
+MP+7b3GcuJw2UGuv9MEL0c0kvh1zBpgx1fFo98imjgOa6LtnJubAiWNYofy3NRWma2dD4nNL1hm
0KJpDCLFkFmbB21b7vjdAp5adpTjRx4+EmxRhYusmVkIRdEChIiKDV89Omgxfn9913ItCaS8nJ9j
oIYCm0jM0B+x38PooY8cvR9Ou68/yh7s8XgTpIdlsAH9/bTT+8MhvLJLPMKiAeQ8xqvJI8xsr69i
DnVfZjwvdudGtayAVcUrbGF4FgYF0ff42KpKJbU5fe5WqPXWlPO+oR/YXncosgVMCL0lrOM7KPzb
aQF5xIq5Pl0USVIm32tLrNK7xVLBycOnGbrt/HhdYtIa+P1UZOfLAzM3WIYEQKad5xWjM8Ptmdpd
tD9JNSF90oBK/UjowMKHgQuqikB8Y4utnzrYniMu6vWK0GnHO5HnU07mnZu4wZANSiW2jtB5ocfz
S9noiFwPWNjfpk+ULNp78I3cKsDRm3kPF2uGOwsNfjNbVWpxWfI022bQQsjk3U5szPPpWHTDZCH+
arRXKOTv5aQb4iJ01dOckpCQgRvKw+tHCizv3Xtt8lCstIRsOw0sT5hg2fF6aRZO8uKAyMWXImbt
ukgvQp/pgsyBsHvNrIGzwkL4Kvzcfj24QeoFbilbx3JuN4HSaeGUjUgVNJJoFGm8q+sR4QqFnIGI
v7oqnCERJx6AZtH0we1Y5ir2H8EmtI4U2M/7KuBtGL2s81Ae176AMgRtj0Lb9lTQQxs3Eg1fhbRG
gtxRYhLj99QXY7Cc7my8jfBXvVq4y7NbiktrrB+wiXP/qcrpqL9aX5B3FxVGBcLNItoMeJYOs/VN
Z+XblWW9yK85i2VUwRJxokM176oMYodEZGjoQp8QHmvlqlQ0Z1poiZCu+vJbytTcBIXb39ecslAE
Q0qA9M7xDseITA80NPlzl+axlfKqda7RME6MzWeHLZ/eaYgwfGw/Yq8InNiLV39oOaHE1DWbnUEo
ikvDfJFtfF93xGfKVKyPgIFiqULyElXca3Tm4+XWsKGTfXNdnERO/j5WV/OuMoPzRxqbvCPsvoBE
JqFD6u3eXVO2oqa79TFNsJhNI4fp357GJWwYBmZ8XaODK7fZoxAzkfHej2kp2rm83LsBTBofTgOe
SLM76HSrsp7Z7NldQXISDNpHnWlt49wKoioPUo5wrYD49eaNoxg4G0ZwfwpmqXvbPKsnjeWJV2jt
b24sByGHFbdFY+OjTyHfDTTT2nGSgKrY7cfbhRMXRY9o5kX+ETcgMJ4bJ3DRTM+/5+1flgM3zgmc
6/f25Z9/BJ+b08SBrEejbKYhVdisg3pHoqrBHZ9DDNO49VwqzkPIw8D45xi4q2ofCOa6SuYA3r4q
CvNLE6twnuIo/xTAq3QZiFKhoEUQz5XOKv3I4ng5fR4u4S/AxErTHNpnO6wVd9Swn7iMhBdM9X5H
XUVABugucEhAlNCsDRuGaCd7K5q/wpxzJgiqdKcqxJoVAveaXG25puzvvejxjhBg8XsvIaHeGA5N
91+9fZzoFSJrDJO2B61ssLXcQJZ7qrquhs5ek4ilVz5Suymc6ys47JqFEEWodP8Wyz40E7XVLsqR
s+jTVOpg3nUHLhjp9BTyaDZM8RzHTgDFKwxFcxwarzV4BH1Lesa8IpbrMy3MsZfRrTkvW2HVAwlW
k3g3vd5p53tCBZ85JDbcOoq4bh3MVn6am+xgat39lKrvs3xMtFtWEzjwSx634qsiv58zVB37BeE8
OeZBxHoRahvuOZe6Xxy5Lp355cde9ntPxJ8O6J38IEac6zvHgRgfJA2AFf9bBar+vXCwblI5F3n6
CAdgeZRtanyZJMkS2nvVlLjVYvzLQowqa7ogVBWf9iJdtkboEuJAFXjMuIP330MPw1BqrP0nFBCK
hHw+3k1SNwGCGYeX/F1Utlk7gH6SiM+iuQdgV3fhZghuy5I6XVeLl8TvgBGxmv145zvUOG2JLAxT
CB3Ws8ND5NpmlrgGKpTBS/G77GQLAM3UNvkLnsPtbW2403nWDm+7uEsQ/sKXMJmVDWRk+5VZ6Od4
ldRqA3Lmc5ljnpnqw1TFVprZJUaEFJ+8+tpogAWIFFlbkioz/NyLVCee6vHCUtaq7qgGjYAgbVVI
dLSH/PZ09Pkru15hCkaEeFYVn0dMBzvsUohQTUayEm+t9d/xM+BuxU/+t0FMMafqkAOsrfKdxgnC
YVweHayRxTWeyODbTyoP+zqNvaYWSgY0tnRaonNZDlqXebk4NHWPXkJAwRoor2/r5gB/e+nQDcfu
5DuNuI7y5No6vtcLxYYy9LQ01SyKe29BU5AA0Q7FhV8N+PdrH2zfE4sxt1fsJHEkTmyCAIAon5ZM
4Fli8qteIQncRo0+G8M8OspZLarGMeM1Tz0/NP0Q7lS8cxa3AUI/1VQnFaGvaNNBZ5FEulJCKlg5
eXfRGAF29LGoGqwKwK00GLd4IdcZRFHP36Way2MUfCacINC/ddX4Pmn1L96S1rNNqgEwCy6yeW5B
I1OyRqW2YGBg13vjGu/5GDCTlSeblNnm14l6qCdyCLuEHJ9aXaSzA8+U2u5d0M9ocUBHAWIQqx2z
WvRVcKaFJYdHP4xbDqlK4sv4UHwGtCiTg+aRitFMN8Lzi9EI5GeY32f9VWyzuGbbwlI51xH76T16
9xUZYEZrZRGaMAm+r8hfVs40/G6qHwIpi801UApk1NO/dAWxZlHEo46obRGedVHDEnmclcEUqn0U
IVSxS1LaClZQ64ApMUQvV5q6HIysJdRVMM2W5F0QTQH43rEVp3uwMMxzCJAmLJWelifDzpxPzclp
l/X4U0GWg3657yr/LnnmYzPvmQZ4Ra2GIo7TUKLWDAPbfcA2b3gkOT53/1/SPJ0KoDHTaFuOae7i
yQrjFbWj1+EEFUQwH+lnRLFOW61w2sZAe9R4YHACWrtJQPhn3Q1J0Q08j102JSjAo753RvCOxGfg
Z6DeGn6GMhqv4sio4Xd1TvNOISK2o3UmSiasdjtz3acvKuS0H3DGEfp4r3l9ErAyhSgp+zEeNg3r
A2EoNo9RsFyF2I96Rnw3Rs6x62dYnFhYLw9EVsXmZ587wqmkTG2ws7iPVHVIf5wfuTxD48ypYab0
1Rksg12bPIR5ZMeyUyhF688g/fN4aKg7fHLE3oj+Kxtbcz60SpMeel9SzArNOEERiJm/UENVOw+/
QBRcX0gO2X7XLk/g5RduLV/A+Lii9cI6h2J8n677GTEQesfchOQL2eWxbK838O8F636p9WHnx4EW
Gh1QlL+hpVNAmv0dwnGGjdmT4YzPR2Z3SlZZceoAoQbQcUqE7OL/OQyTSPGmROD5nR25bhT8NUb7
TQpmJfrvL6L7ATwQlMqv4Z71bgqnJl/dT8H9vU/UDk8TLHYc1vEcW1hTsK5UcSFyByDinfPrxSV5
aREY8Gaix/l4umHojNz9CJPobShhypx72E2Mf/0vaLB8nbF9moqXUrrmdW2h1j8E6TFtwuBWC7Uj
XgPTt5D4TyiDrn+5xwlNOXQ1luXafSwwxkzdg+zNKPmdqDVkceXvuqYXmOF7n4kK91ckD/rajQ0T
sLEwXXnPqXO9t095id5unoP5EHxuiE05E6KfK5HyJUuxhdhjwJYM9nCHtDjRRk9JY47XGPbHZJn4
q9m8vUsDG9REX08Pw4OHU8HPuK/JtBoZeD6EAau5Zf8AUdHm5YNFCJa6JxNqn7/MJ4FfnzyYQ6my
DAzSW4/nC0kXMODkty1eBXnmizEkjRk1sAFfNYTgVET6dVq8G5bnCl+fzB6wIWlkOs08TRnMenDr
XJ4ZVXwA/55tg/YCgL8p7DdiwwCs+EHh0R5Cr0u/nX6912CnzUNpytz29NUesmFU96l8r/C6OKvX
+lx7yF3zqrrjfME2A5ewfz6R0VQk7IqDZeNKlOvDhRlHHxy1VOSpROxZLm6HRfbfdeHhLGlZ3CwM
dC4tNZ/A1CTjiYXJC8TXWFmHDv7SU70G5LPgwmVXc7erfS1MXoE12lv3hRViJb2n+raIhCkI2hmS
rSklEtinpyztJKwwlCDzGHRuMKFVAQ28+0vhASO7CJHqGaVb1iQ1Nwn6yi1o+4VWzZC/V9VV23CE
aOpp0HFiRF7B2INvhsViWsCZOJFwz6z/Ue46Wsw1WFcDk9pDYS05o+9DBZlQLTY0AgpF/wbEI+L7
zf/m1gfmhlXg0WtnvtylAnCEHktM6MRNoJshSg/CNR9Uc28lScukgl9AfQtywNDOND7CVYAXEcFL
pQ1jCUQIqqvEkG3z/zemRSwx1HaxTz93ADxR/O3LTW8ca/W3h1mjos1io2Y830TG/yKo+Kj3hRog
s5ENKkBRVTPEvpyPfB4zAmbQ03vUZ4qWMeQobvAffIwRx28lmyV331FNeuzxVST33F/W4S3Zi10u
TsCiKom5vDMKoD+HmBMKAOOMxavuZA5q2o/FGzK5qvqLiGSQw9m6asGaQCz+TYspEkYPA1novlF3
mchKH3qkw/9j0bjs8D6rylGdChYzVl0n1oA8qevHgyIKCwSf2FpTb55GoEFCdnRKu1VaVgpqlZAu
8BtUvHfZ54LUEnNwwuAd580vTgFXPckIUFLzKmPdEe+KaMFeh7O9ycN25WZh1cHo5b98KNU49BGx
4kyY/xPX3ujmDw78NKoyA1y41sP57Q070zjJIXhgRr+YZQBp8/kDa5Eoubc9nYmAjRK7UwgfdxYE
xJ87tFVO15XWm99RDXxkLu7n0mWrZFNz88VwwQCQdxCpoYPa2yo8uUyKNQaVHZjTlgD2k/Kaf41A
epElQfxvV7rzS5m1nRW8rPZjpMnj9H0LRySwPEzqipVpx4fQ6UuH8phcztq6uIN7GIQpFsy1rOtV
rlxQXDqjrNH4WHp4oMQ1X/3MESjXrXPkWQfLoYw5CzNPuwU3gAcWrkFPv8VJbygwWMClUqZw+n6a
vmrD7MyFluCj4meYynGN3FRYD2xO2o7qPqVV0jTBPhR5BZFyx1DBmMCfBXsqfpoSql4zauR/pcgC
kGL93KGeDApfUgla5ORgias/6SHMbHyKq/2p99IBgS3cRJS+bGT78sjO/IzWFPQWxbGrCU30wdg9
/+qqa/eOYz0HOK6SRG5cCUCYSa+iBZMyKVprktWRDeuhyGElkfMI0Vkya7AJF6TsHlOwxnSost+Z
7EF/GJRxEM2EOWqR+ttR3fTNyXDMTbP2TvJBpRodd/0ghmDocTy1lzFogDKdA9RgfFXpsvSJN4mV
jbTfE2JHlFQhCIEAEBbg6lRmhMuTvGET2xCbWaiGjnnJKtkd1aWzr0+CiarBgfKy40ctKVNxjKEd
5XM1FqOT9+r0YoQb05QrmrPt63dRBNBzJ4fJZUeQhDMsEHs7lkAuqbaEXPhniLCxIr12SphWbtzQ
lZhb1FOsGRM7Di52EFRb2QWqHQhygjfxJjeNJrXaepxPcrYYAr1935JOxMkoEDuSeMFaLswVifRJ
nNBsuQ3NhlEVZ+iCLOt0vRH37nUySafdKBPYklQU1lxEoIdv0GA3CXtxhAN7Z/BUKb+8alH1/gLH
iidHVer9LDwR4RWFPg3an2g8RcSyoH3KJK53kdfXqKa9RSjuSIkA1VszG04Ev0t2QLcfXIlwU3D7
waSR+bBTcNOA3zzQCxvFDgqkM5eypTdWCAsQbzsTujjkOwc3VORIdTPQ68QdkqzojRonoFXSiiwI
G58x6gXN95IWEUMr1gX0cvUGCiyFpH3b00VesdqtMkRskUnjZ/OsEhgX4VZex1LuAqIm4alGUuuL
Rlf7ol1BhKqCSYWtGoJ421qTBLSb8dg7pwpna7LlfRF8tjbD/WZWPEwKBKJH1L/j2tCWBRG1C5ef
sDBn/lnyo14BY+7lnvCyDhUS6p3XDHnmmysfHy0patatXTj6X7rh27qXwP1cwzyRuO5cX3yaLWJg
cC9I1yetwSbTuqRcdxBKv6tE5IM0tAJ6gFBooXc5alJni/RM7ZM6klSCSN0+s7m7uXqwFyaByP6S
4lP7wP7m0Zbd/opnBBkJ11yGjpVXL9mf5ZZCqJWjeYwQTuhod7znsxVWTXldpqNYsUKMF4+bmOfu
Q7k9YGH1J8N4wHEimqRmxpN8Kfi6QRS0qQpk8nIf58rXx6l4gPuS9Nav5ZAW4CR03l4P1iRu+GwN
+Vb2tiYYofF62aONghVFIV0flmr78Fs+Z5JFm2AdiB3vejOFtHkbXPgN4KXlkjzkDLI000CIL/hD
h8JmOUGJ7BHqwXXT7iDjaZKUDq7N46DS8W5GOLTyRxMnS+sS1WPd0JRYYFpFrGT9VldtoRhL+/i3
f8NA+zd5m2w8SgBlNWuAUSPcDjd7Gelk+FDmzvscBGr3/V9toHNCixLLfWXGpvxfI5nLEzqprVOZ
pt6oUAL19gf4a28LGjmwnpW7wl/28i360SfHLYvQaLtzpVfbp35h6HkbWgKx84v1H63VnOC5Pl81
/KtOd98qlETVDgDE5MuJIxjkL+7MV061JXaRbnm+z/on5S6GdNsJyL3/Gb4zYkyPOvXOFmLE4f10
kEa/Tz8YWo8wIq/PkkiRl92h87V1mZ4S7MhuW7Aq06UfQdzw5c3lz+GZ5+mx83/TP8nWhlFIFwXN
jx9YR6IDTHJ0rKcqPlcz5W87N1imWggwhFuvXbNy1FhRQb6+LO14YxsDoxCkYEOFqeE3JL55kKae
AYE82v1vifm8XybkP7HEE9gx9Ue/fvb/VNMaS4LfzM1ftghPt0816t9FKSrg7DUdpUHwiAkfl4WN
KqOtWcHTL3Ax7hObYFJPkt4vN0DF0KsncYdkLYMXke/zzEaM7RftOzTSM5x9HWQk9XCZ7zb7KF7e
6yJZQmWS5vSAgje3qgjuHUfIPdc15/pbXhpMMAGFos2c8+prrJge/afa7zYaMhJiV9tNTc9DOhSO
VR8hBp7EtrJ3y25SujcTqmtRkfeTJ+moU8v7VezxxWlHou9pDR3yqm5tvmcU+4pT9zuT1Hfn3YRK
pIre03tJrSAnoLROjZXIoaqHv5KiU7WVQg3R4qDlN+xYNkEzfAow8+fdWablTwXPXx/QphF63j/E
v0kuuYv2tS6UeqOeFoXLECmDqOkT+0lTPGhYj4LkClyW49ImKtO71XuSBbPqUqus+ohSyUmqbFkw
rpiJda0Lk9/7onR/86IRTaZYQ6q8pt2WtZkcw5IK8abzOMvUqPlX4DPuP0H9+2RY7Ll9UF7tputn
g7xm0vTAkpu54T7KrV9a4ijkWHbjudB05J3/418RN9o2701QS8KpCSdQN3ZhIvoZA20rk2NTGtDV
xvCUJQq7XMLhufmZtgHveIzuQSVDbcm4Szng4XaFUj/ZoaOq8kgcUJuTFa8GnY6fudY8jnn/OoCo
xDlOQCjeEsZrI5CHMjd86uCedY/dnRHoZgxm+JIBMYFFdWoT6vn2M93QhJLQICZeWpcF8NuBcSaE
lcZb0tTDA97UfFpbf5ovkV/9CQIYAo4o1Ex+hmDUC3RnV09bLfRdZpUb/efPH0o87L4PcuKYe6Xn
48PrPTSqdJ2+yhN+6grr4cQWRFCm2G9waB56BT/CnWWikDZzKhHP+f7rcRcgmGWN6BsPHjqCg02e
0/uKg1CDUJeFqvaxKkL+Y++YGCMQQp1p+F/c42KCqQiaRjlnHZgRJmbQLKMOQMY7Gs1FNUyMWKCz
Q0tWKwVjnwaDvcdj/FQKQKEFaUBwdAXpx5+sd8kMyYo++o4ZYpxiEWjRDCwq6Owlpm6jJRuFNaf9
UnVoXAqRiGndAweVPjS4Q1ONlq76GgbMNqEKZkoxh6/Qv+0DMrnNL10AVylZP6Ams7YtZ4PMW4Ws
j8btipgiuOGNzuG3Nwmy2lOFbj5/84I/Ghei/o4vBmKXkfidv2G8wgDAX6a8hato0F1J4S2J/D5k
p/PoOjcT57sT/5pKzggJ5pY2jzs7htoPoRev9YVHPCPGaokEszNbFZpHIvuNvIbrFDNyzOjq1H3M
vNQrag/QX2ZVRYh2ki/xHo5ifgIu+Scm9t5bZ+5IX2My8UFtvbs26u4TKsR/D9izpcNk3XNSA/fv
O1ztAJXVzlZAGQDAxA4A5GK7jW3BSArTWHW9QHJRxYiDiCZsJZOsN3cSqlkr0oTRSRxQmOjcsWfv
r6PONldxJyAHpHfgAQWW9Ul+YVuTe6q6fzx64+0kP4YxUu68r63iOGiTFWv8x7D8Wtflv5RjIx3q
GPJpvDfZYbO7mAFN8Wz0SDjOlegLFmoxj+uZ0eE+t5TderXPeYCRc6E8jffvt7rZlYAxCpDolPdM
KzCXAT5ncHVFM5QioOgES5CTthDLzoc6yQrmfhbmfzuWrbC9Cz38la4S89ZCvGaoHiEYljH86+Ac
M8RfuzPUyEFidLQt4tO8tXDgRh5kSKX0Cg6cnnXtLiZVK6IJfMQOuXEkOjdPDjyAwraPF/uHGrhl
yFEu+Ed4jxYI2kqTBk9mLbuVwR3G9cDEC2aJLBzrDxcYblgOlivvMfQKPXWVzedMzbeju6egcxsk
DcpIVJWy7hDh2AGGsfoZYD0v6g+CYit9dLTDyEMxCZFJ8hhSwhf6R6yrHt+4oFLRoaISPBlu/fOI
q6XRE45OtiqzL2G8wAUcBhEzz65aQAPpk29IZM1EAi3ZTldjeeudu7AVHAkpkPaKI6NWvAYlLMRB
bvNSKdCtNAWTWKRwK0RohlYAj9XKlew5KtdBesHpiAPDC9pNzlLJneLT6xjwlhHkpLquIFDWt6pR
p/NxxEDt95JLN4dxU+6T9NxkMPKCqREUbNl9MemQx5NEHhJk7yEPjsFX+b0gNN2bvf21m+Tr+07q
nVFB5B/uKMxUsskZSUQI8UZpGTRknDySZAb/WV8DKRLWrbSo/SERfPbSOYH56J0nJIwVE1M0+H/Q
kEDHNS+sQdBqKNfouwktjcEG8GLIURb2s5h/qPbenIf1sTtLEHAoUGbDZJTgD547WCoj4wbDhfuO
ok5++i7Dvn6nJON0jl2/+wTHVcjlhVa1SFhbZiWAsf2F49D0OyEUGHBZeom0Cwt+Cl67THy8+gSy
JaLlYUjvV1LDqx/Q6Uo/NicFKcHEho2IaBwhmd5tRwDMPUn6bSkroPQSOFXPgUgFpZQHUXURvGce
Y1gQ4vzvS3CZ8ErKWhYNTENizDY2DMJSQz9DB9NMAqAS7xLkpuyquyk0++FWXkQnYpW6VYt+sadd
bULxYM4Ou1Bq1QydAsShigJC0ijgClsP/7+tv0a6wgnfIwSwUh9yA4PTmpe9rjrLS9uJoJ2LDI9t
5avUfHwKTHUT5c6/2nIOcWiogrqq2IAQIviH5VHZrOBo4g1QWC2mVgzUiRNSA/8W5SjIu92KMEDI
2G4QxRwOtxpy1DtMHchqsvEr5EIFcsSLZuCmK6jOYK6yPEhjC1cPkOlZlhq3stm5gd/3uit7+F7i
7a/OLXls1d0lb+ItuVSv01gG3gggV76M8xjBsNjiwJZfNv/x1AGVQuw0/r3/dP6nmM/0icsKtTel
MO3pYzamVOC0HPoM+wtU2KPagWxa5IOJr0koRYS5syjqOaYVZRWmYK0wjIJDgTpe4wp7MkUvlD5Q
Ms8ad5hyXhxHeDSUe72WhfuHkdisApDijh+0r7Hm7lG7MWHsfBO+dq2I64eVlCnlRj9e6lPOUP2L
gkAw1kEciZbqaPixSV1Hsc1QtDAjq+KzaG5IS8vjIZngyBDX9aBGuncnhU2Jf1x5rO+8wAFdN6W7
cFgXvAEeyO5W7Ft0238dZa1KNb98WVf7F9eurfdSwxRLpM+wlCHnzXliT5KMO89WBdMvcr9VQ5Z5
7xzrvtgVoqyJ5GH+W4CqvuY6ICe1kxnAK5VnyRJbFQizVvdmO9/zl3j62jywZVMjerOsUtpejf0L
ICHlH2lAwpYugfApSiPfdR7SDdYWejELFi6ZlGbMKffEZuyETFraph08s7ZdF59YbhftmERqZB7v
yRWoMNKmUzccTNyO2WjwtF9vYpNVN+ie5nJknMEcDa4jNzTbIiNvsb6SCp6tK4UNTUgxpn2Wkz6m
aMAIm1Nut6kRm4Mq3PE3tlPz0HxXWxa6tc+N3pqerO3d83B93Cyiu761HCdb77LsfgLNRuYa5KYG
hTt/+pTYftB751+JAJ923qK2faJCQD7o5MpbeeHXuwdL8mgjR9pVQNvm/LTAm7su8w8HbdsTeeza
SPkXke+7TZP3G5+Tm4aWWn3QK4rarb2ePikbXqxx/5lM4z+6IAYsuhFu7ZB+dIWEeoG2RUEbR75V
dAzENqUfMP6h54EI0Om1UySZo3jhd7YtZlDoVWZanOw/Yl+d9OF2RXh7vqGnbmiB0qUDleP4k1y0
1UBYe9fjOCAtZc3w385J5RHOzGFD43QiWHGM7G+EwRMJflU8ud/ojgCkHTlnR+PYCOWTr3x9Z33M
s1zDEzzQVBgPNdcCYHoaWYckczTNi7JelVR5BpGNLLECAsueV+t5NC1Q2vv3KbbssUdF6icmtJGr
q4wPdZsf0mMYwcJsq7CWU/+wB0pKFXob8B9BCJoxdZtOYo+2OdzTNGMVu4QVZCqrGCF4Yy01FWzc
tHZTnQ++x8GaSRdSfJHUvYx6Mf6zLUw17EPxfWzisW08j0UO0hPL0zuXEDeJrF7FabC2DUFD7ZAz
BCaWbx0rTMs6V5dqKOOVuj8BZEgAif5+AxwHnSmpcAPV5o5uqx7ZBmtJ/+8Mu+Iu6Xq/HBjd9/Qo
NG0GzppWmZfoeUmGB48Opi4+Xe+6tSxblzhYo8m1x16NbDa8mKM5HrYC3zFq+GHd96EhVlOXRgOU
jLYfw3tnktCXE/az2xt2Q+x3+dTJRVELyLxQphzaRa8CORaiVDYrYLRViXcE/wl7XOYyW0Z8geDe
lE7CDLq5ipxPNIrJF4P9aCmD9sYz01hyK1nc7l06+oYDvVcx58b9KGc98TZXg4IOjftj6p02j6wl
xDJiUOW9+YymuKwPBy4BRxHNJ5zXpa1zXlFjSnMHgtfskWyaUyc5xAD9RO1tph+5FOR6Usdq3ho+
i0Ms5hCXekKPjUBpLdTwHxtPCxdleIQUROf12I9xHnJ7WwR2cjpuvCib4lsn/OKEzJ3fxnsIskkt
2YF5HgJZGfDbzr07B36nAyKnlaYRtVETqBLcQPesBr5pkkWirec1hvMANwAScJoXwJMQ/1PjlV7o
8BgqobtwPmldNwpWyWZejPz6Gp+89yOGnW4VTi/Jl/o3nv/SZOC9h44zwOK4291ri9AASqUWkuY9
Bd08kPsLRjAsZEBM9PZtliyMQrIzjrZHvzjH70v6xyEyqgUwAGvklfUiSK5+i4YxDEEmhUk5fjVT
u0zBLfb5fu9DYZ5q0jawq6VejOcwA9/SlfXfYNinRMbNKvKSF/r5jNAb1AFkKlCmk4ci1+yJPRkq
PIogi/V7+TiryAop79aTPOb5N+kI9+JnpjLquBMQbEbPth7Dj9PaQ+X73MVbhDdjkpj5FvuuSDNc
5s8T5FO/Mvt6zCnB5rnnlxAELmynI48FjjO5ye+mkmJ2rg6hFiKB5thx+D8QA08FfzfSUJDNR5fr
dud3tPQFHa7hLc74fWvYnFn4pYqTL2q9uexosOfjYp9tPQDfPsNA0ZVR5f5vXug2LKpJVau2fvyV
dvJQ2LhxreEzJ9w4UyETnV7CzcW2o0Ad4j2GnskIocqkIO+faS9UuRX5+vq6U+h1fhJJherwHzKw
luZaO2Njq0YxiK5rLhsH5NOxRq5BPIhK/JjDtq35lFGNuRu3Wza4LEuA8qAttUfkHXU/yWvVaTLZ
LzFx8aHPWc7iSFmzx27A3+F/W1nhPLc/DJJ3emAMRzzo9hFi8sU4Bdx9FhZ96CDRJjbfER+YFROA
RoYh2HK+b/PY59tND3V967xvlwFCR4PP9oIU9nGCtKUwMJRi4zN4yKG8MtZSUgshjrFSWDELgGgf
2j6tHR7Q5+JdRG6GIQ+YfO7J/Q+doKefjXQFqA+wtj7PeYUGvp9X0Epz+9hOc3ETk9Nzqh+/wiCr
VIrpdFUwMieJQsIQGv4QNaKgutuIy8C8GsuZZ0wzqGDyFZfm7dXpYGpUyMCELdjD+/beDCmNepZc
e5AwKyIltHdei6x7EvslR+G3AC2wOArP0RwEoIC/HwF8fkYWLooUUfx/1Fa7Yo2FWLexzPyHGhpx
iZLuMWd6YJ/TJPRLR5+PY9uhptx64NtMIT3SfQ9KE94HtdcKItjT7q174LfGH/maRzUYToiFlhS5
Pi82tSArNcU3eKUTXANDyfipy6COBt/gwc2HzlwJicoJTe3XRn4n6rEfvEZk9bC9v0/laP1Lauhj
cJkJlOW9EN/LIYjH9SBJpmZDSa05ZZoo2v0EmIC1uELnwXDHNEfCDdnRgFiLuP2y7Eq1PNWtNlbt
W4bp7OAA7HDz5TG1hxPKDvP7pW8hRaFBzo5IeJQ/NuUjLlCSy2VEUmDr/lLGKED25rbxXsLgtivV
mjv2gd6lpCI7wnrGVsMdTCORIKDwPoCOJ2OsU/kcee6IAkXJOvBOIYdqyCzqe1QR6GmY6Arz1tZJ
KG+bjjr9rafNwQJNVJ+uytXKKZmyfavv/VMjPxFN2QiaCP9x87ZazHuUhMnAQqI5OPxlR+ts/pX1
RVc8jwDLD83znbzOOieb//d/90wtYIWEcNAPfK9kRgUQySYzsLIKJYtiIFdg9WLPWsJVqe9BEHmy
Vc100rikt83NobmDE/mqj3NMwvaj86oixWfp7bSYhxoOHBnX76jL27mUC3ZKliG+L6gaVg3+LexG
ShMJKTq+Q0JXBBTwanxzmQaSf5Prl+wtS2g38L6dKrIF9ysv/UUmn3CtBLkDktqTT7YUJiVu7/HT
xEr8Py9li5yyIndxnC7HLBo6f2s3soH/tMD1rL+vOPrscVYridhSCHMjp9szA740FaNPWJ/Wby5i
J6x78d54RzFYEL2n1N3BjtbJnswKeCll+bQx8PUXoORlZVuaQPhdyn03pLQhZZlxKXCTG/mm1D4e
gujp+Pzdwi/AiBVQ0x4LkCxKYeQqqedy3+gcBhF3+6GN5pYvGUvToed9Xdb4KXqepL2Ha4OVemFA
Zud7OcOVeffumpteppoeuGFbyElU6prH5gcyUY3z24KEegqIoxGFgzHrjtRu2S5Tv+0U3Tknzk04
C4ioQ008yXfrFcy78483dWNk6T7yqfOM1X8xxnv35urFVMnkwSzp8a2cO6WXWcZHzsxt2lNBML6F
4O9r4Llvp/e8k4UnpSWGP/cpG1mBrGDlbC+4KXRyKkLbbLo3Adaa5ZHnDiZDI2d3ah8YJDhikspk
p3OzqAA8auqwtD+FNvxj06QYFHUM8mCfrS4g6iBjgJ9G6Godrraf/yQI7+E2KxgjAG3Q5faULS5X
ghiONKQxWj+xW9FgU2KHXoRMqXDVWc9lQe2qr96jSbkI1LdVNErGiGy5kx+KhULfnNEN/PTz5xZz
JMBHdiUW+r1FeFUGiTM5x+FDd0iFvpWxxvXUe63mns8YcRZsh8LF1wXn+3gyLBSuliiAyUxaY3ej
WGQhCSDvnFsx8rlRJJARZVFaRBXZkC+uj1CQFEDpDac9kmpF4IzNJlU9OpvqIxcj3hccB/7G+uds
vj7/qRdy8RA54PnWDcgGBNBwtXpU8a5D4MbnN5zr3gMzKSPkLHcOeCVBR18IsTLirzYh/kBx9js/
grMkT4cntDReBLseY7jXfaQgPosNrcKtLpsWXkE1wjuDSIym25m+gl421slHX0aBUwVB3Er0Tow9
qLOcWUdOBGI63s8UOL201yF0IYUkuB82dEuZffLmLCwj4Zt/aoKvP53xaogHPRu66YLIh8b7bHD2
62IVwxTst7keTaUELrLHHKYn3usGbzZ/k8TSRE4kl6gn8BbgjdPOJU1V6Qa8UYIOW+yM/QKy0HXi
ZipmLra6cJO8KqcxU0tBG5vFRByJ8PMr2hqNEIiEkpPxCf/4abLRwzmljN43kYDxXqa/p95SsCRa
raM+hPYOIZ3O4UNojZ8tlPdaHf4imvR8mff7X+DP6T6tKiFPkFywSBJLtrDr5rya7+eUezKqu64i
jYUO3hrlK/mDHOhuo+3DTFiUEwOPgStPTZt2/DYPvqcQxIAiFlfJEJOxGo41BtAxLa7qN60SvWqI
nvjlSlgxSvROx9qBadMF3Wcd1HbyhxuxMq5XgA6jxcudqwQouA9JUlhukbuo3n+QPGSlPk5LihgS
xJyhe2qo/KnqH1FV1+FVBHtAzLJKL7672SclbdgBVw0lk5QeNlY5zDN5ezLEfgxGbblSqkaDMOHW
Db60SDGYh8qRQQo+wDC7hPEg+jHaMGoJcJmwTmJpoNJhAw1F4pXYxpDg3ofY95zdUdR9yYeK+MHb
3UjP9U3lcA7b/yEatA+blAUdljfd4C14f4hRO0bPXo4zRQ/NJcff1/CzvfqxHUnrPZ0qHtsDj1ig
DOGdJvz1YQH8z2vFZ8sP7ARYWkqfn6o6ac8oCcpLV/LJFQC186zh0j2FlyJFVxck3xKh1eFUS158
oVqUsPbByqe35m/9mBMZVfjgDZG9A5CJodiVb2ldO/jvNg4RRRLFkuLEUQATksxa/fJdcyuNKEPv
OE5av8VaXg6/OoEftKJoN9vdTCpQdRcWrFTbBTXJqbLRuOaxGljHqnlQADvGRf6VLfifpFJ8F841
rAHlZbaFNbXNCfBsSviXWinI/NgXrPS2UkDUktw0qdIU7HJO4Slnv7yiu2kK8xxEdIp3WXlCJG+M
0da4QuvE82Otu+AnzYaDK1reV8P8CEJ2RKpyrvh57FrFeUG8U2EQS8fvBE001defvGFc0x4Jp6ps
fGdjaqEXM5eeSewCkLV81IBh12tGirpZvjwqbHibeLipObgNkM9/SN1moUSXS9ITXtgEGNfERdGF
0SZ1P/obkOMJ3cRZ49IiF7nqf9F9Nx0/rkyrTgdsKlwd34W+h9AnVbVHLU2zHDaFiCxKaEwVXt2m
A87QUUsigPLnPk5clRHekvy1/mtnmWVn0JKiIncAqjQVuMgvSL3kNrgoBoSEleDIeInjnYRpKTtu
1UJTer2NNAsHVNoEROdLdIP4HAjul0Izp6SURFyU6/MkNmK8pctJzecvWSL2zJnIW4BKB+g+YGjw
npub6X64LaO0s+TwhI0GLfeg8VYlgqM/WR28T+0QQPR7fZyLc+nM03As5FVSPqIjfUiqC9WOGj12
CMzLIqTPtbPQ65bTQGQh6Wvqp3aMsLeePeTrGUEcZgXrhP1EnyICV6YRhmwS/FN2M/EB+8nyUXsp
Hn2Ig45yThH6c3/P75bRxUlw3QU6y4zoZT7mgoeNM0TA5yeps0kB8PDcYAdUXa1WixmBUHJAYRME
nx/LytHsOV2Dt5tbzqTyQuPL5pMju42vXB7gBk/40/zF21dUEdACWB6SBNXV7i/JcurUsnwMAhOD
EGMRbUQmEKwLk+WsecPKulyjmBLiN4GaNHsdaudUARRd4wrcBLxbBWkI6rsnIrVQ5gf9HZkdRdbG
Wxc6Krt6RSZiqU6QDoo80J681BcmnOz1YLXzb9Y4HoH5MPM40rPL12FMKJXM1J1tcdwiu7DyPDFn
eqLbW4pH2cULZSC9TmqJFKhMA0t5gKFa5GhAVsRD7Y37m7A4+XCruYmxkWggdrNtf7B0IaK9XrPG
YakK7qRSsB7KAflzko4gve7HwrcyQvApQVpCAkXJG4h32uapRvmPKlJ2fnAUUj193IiIj7Gq3TTX
lHkVHLDe4JovszmGnrRYoDoYRkyNR51YsmmFv/M2eWin6lAYmhyVN5yNF25vwY760rWhPiBHGXkG
dRK0XTJjo730PWvyWpmvUOqRTj3Xb6bGNTyooFpDnwWStYcUKyYK/xYlSUSjiblCsZKdeWlVmRbp
4ZyblmIl0qN9qmTQRarVvyKSCN3rmnd0UMFuDg/PpBfqqY8mlg8ujZKpO6KS+4dyMqcsAfjY6k6U
sW59FbTsGZBfNDlLex/OLEOcxet/nTmUxDkMwXE9/ne+DAMhZ8WkE4/Ea5vraDjSWCjw9a2AGqZt
h1a6ERHTJ2EZSIuNias6TN4f1535x29dYKMzkai1HYLCJbx8rTB+sbev2LZTPaUUrurm9phcJESO
YFSLZ0tCcs9ISn4MvfED5oDv5h5PoRea7S0rlrvXray5tL12ROg7VMKk/KOgDovTqBjmv0U0/a9Z
eLu1HqR4+Yrv4DXJ/HH7f5rQsXhlAaU9CxKQxvcq9xeTRfXk6fIiq6MwJ3IhoiCIJGuMIbl5IQAl
yD9l/xqABapdYPEiN2J+csPhAV4U8v2CvYKD9gZJW9ZbDT8yXlEZZubnDxlpbczK3/1er/PR/KUt
GBdgcu7LVK1g9IfHuhiVWV1gqXczkptQuDH1+h+B8vr9ZCU9dnOZl2KHnl3t6KhRXmQ/qv+bwgEL
j9m15TbyYQDyD06Q8Y4+nX1SPPDkzr9D0URRXitlFec6sigk0WfHm4ozWWsySjux8YRzfXkD7IJG
yzVBFZSnWFoOfSrrd/qxWE9zXHHADPUlm+md4JKvvW3qFQG6qZbS80ocugeCGjkblvHf285GmOQ8
9t1DGJVkGRCAWYB+MTTdPLkxGciENPv5XinwqUCz7eSQlmyZY2ebB5fFIfcAUxDLcXulLNNn8RRd
5nLXTcy+oe326Jc0rG6o1T4lvCwCyJZc2XOCQr8tqqSL+jqPICXAKdAwYswkKwYCRHn7trYUGqbo
Q0Rf1KubHO4Ngact9MuQzkffVjxocBb2FxGSYPt9n4UGdN/HF6gz/93XA7QCt/Y88G8JlpMN/r/n
0IjErotLJJTJ+ARgrB+hDrnat5ASzh0koexWfkfANyB3MOrdO1JaYolfAL9nmuoDPiu1UsDn3Aq3
zJAJYq1q4BJXwK/vQjDmC4Rp6HTXuHQI+JTmP+NKBUkYncPj7k/3YmwDlZM6He5lFlgmlRUDVnj7
zEiE3zksX3OrdRj+zAhngfQn6MY49UcQlOQsovQF+LOPYWPLINuFxqAHuqYla4S/QStPnUxqJ3ln
MU+FOAdr4J4Uy8lIP/EziNXx13uST/igkyJz0s2zOqkAFi6M/3sakQramCKaQRHvxdCLg1FBsVTi
qHciza0PK0pkqe1OOgm7bViqQ61U3j4tawxD6J/E+0fTpoAdrDTdG9bPEbl9hXJGhNGRVu/zWRY9
QAKYsRMKfUp1LDf5MRJk3syvVyOXwGcsbfRginl9RnZ/hL4rVQojkWLrq2TrsbhXKJqOHyhtvUoG
woQcvXnDZ3THjLugs1PZnv3fNrBNLRKKFPyvoP7cekWAScRUtHWQGa6J9C0f3AA2BTXCFH5ISG7n
gP5VlonlWCAvwN0BaM2CMCZ2qbqvCgf5n4b3r0AqHqbI+UrT1dpXPlINBSMDTQ5G7neuRKMMAEs+
IddVHkDZ1GQzMNAm5GuqPmgbALNHiKiyRfPe+PvuiTRPe66w6pqj8StHE2kvD3j2exe9fGaBnyw6
9PIos17pNImC8dxwYbWZag7PTcHc7clvBul0C1lsPYP0kv0yLtNoUIP2DjK1kaRtEKBJhmBAin3t
G8QFvtx5CK6BcTcBDD6sLHkze5pvIYMkndvmgPUO8/szGlDTGbMzOI8CHNPtMXnLyYp6d3Hsx5aL
W8GBoOL78a2JXXzDN0/6T89Z7IuZTRHioTkSiNVwus7hDiBVDkYoXq2A4TZ7KIi8W4H1HehkAZ1s
eytctcoDXbpqjvrD0rEsAqFjMCNbez+ZL4sGiRkL3PGDqo4t4S24XIwcYtb1W0JAgDNAY0HieqMl
he1wAT+kFcflpkNhbK3J28tdwmpNZSkcvFEj3f5qcY2b/IMSicmNR+IIwbOaaD0ILiaNOjIlRhjm
Ia4YCUQqDgz8klUzycqTzwIJZMz+krkR2iNJ0B7YhTWGNHNJuf6RmdGvgfQziZBO5MU6hCttkP8F
t5nkJdL7m7VrkRYSpEZQNaqKELzULfRyQX1bmbwC9rWCC7I132U3uyGsF9M9CHeEZNgqJLznk065
vMvnWkJUWsQYrWaCWRX2jRBw3N3dQNu3xhDbCNiteuiO+bRnwnuX9vyHt7gwnzdNk2VylsLrMVC0
xSS+28fo8KxN2kAXszWoh/nNyfrw9pPAvZK0leetuiPoGlMCZH/rq+rd+cleU6tu+OR3oVN8kVQj
1fombYxC5hsVd3I1qTNVvFsjrh0KS1NT0ZyrGKuR2k6St1s4n/WJ/OmLf0xbFZPXSPlyZtfkNh0N
ZPmTYV1FOhKbe/NSs212dmWuargpoIp0pCt1khZfcLYVsbIRxgaW3M9rnoLl4/eqcyJCQv1wI2P9
w3yt+GTHXKpIxxc4r/nzqkZ+P/5qnX+S+1OxqHlfn1eh+Be4jjKgePw/opnuWdfJLmvX3yNx7dpg
3V5z+K2sSkUNPRIEDc8WbDR1Pav2g6R/3SEEDnoM162v+/nsgE8vjvFuCi3snnE9uOcd90jzTAMu
H+Uq+4YGhr5qCbzNDJwvWTiARO5lX/Iyh6K16aeyLdy3TDd8mmOOJALN0igaJ1ZADQ7wyj08bOiO
aBslHGRnjNmBSHfmGqYZK8relWIOj8XTl1n39g9CVyB3EIazZ5MZfqTWMkKt/2bCemZHgpEJxKTL
XNTyAT3VVDeNjylqAG/q06f2Y21xt+39Wawl2kvDKBSUSVndSvH4W3AFsufpoyENrUtKaGSkTRbv
3wdFvZsKKDAxWR8z2/FwyHquBefSbRWVNmZzxXghVruKtyiZWt5N719uLIDvMMuOGmC59iVsqMDf
n3HUZwEWlmvEi48gvPYwFg80F7VCd7Eg8jowEq4WFsMKmdxfUevtyxq7x6Th2SivTB1gkdH2HQsq
3MUDwuwRUaYXFUMuQWujkN6llRl5M1UJJvZHfopsof2Z9p9tm9tIMj7E3YHIhi/Neykld8XuYyHl
C54KNVOVnElQPlKujH5R/d4UMW0S2gYTXBZTmZHE4GNdAABTRMHtr73rXK6PgFcGTMZwVDuI7JJb
FI2KsmRUkbmuClBgUT8bTHy/2t+cW1/0XKRbAzIm2x17UkhkhrDda7b/OmpFOL1cfybrJCwKyqF8
mpJAnXqofhWaz7w9cM6bJXkNy+lgL3uLTsp/CYrvfOvbn/I5UgOPh3iW7Z4m2zvR1kGHqN/ULqVr
77HAwgBZfmnZm+JV2mPXq/m6c7Ueijs6h6yKXvxO0KFaSStDvxQ/6L0yyBWf1Hxdrp3Zjre1FZEI
Qt7n/OcITQJlXb6T/c0XX5TNscoWaijTxtLVmczY0Df9rFs9iLigQY6aMQ9yCWUTcIEUiTdvq06D
ErXQalNrHNUxsnGkWUgbqrgeSJbyXJDzuji0F424EmJg5aAWJgs2pHCjSFCl93exasX+hRVMoaSR
Hu2QsPeE9ko+s2uWoBBqZ3HghmeF5RJZw9sRrCwkHcQvA0pgtzzDkWhQJgHMMq6Jpyl5F2dHzozY
wUuKyyc4RPVP2rA/ZsxDksG2s0IDNJ4fVzWYDy94Vf3P59mKBUXwCKrsI9Op6s1piVRYAp0SXHqH
12IgD0m+Y1UnBAzxpRbZ9m1xypKtz1psX1jYVG0EhSk8QakXQEH/nvr6zabMnY9gZqK94Q3qNR5s
QqNZ6OeZgxf2gfc1IDfcEcQCNp4Ilpi3oGhrOvbhuKn3XZ2fPS8PiSrLRuXXh0DLjdiZW1aUgGVl
pw9+KZsKjV6GZb5W7XZNVsMGKAI9FtSYqSDNyt684aASijVRKX+gSUiRZIe/zACV97QkTN2NdWr+
ge9+fQZj61RPKFcg1rCWTEYeI6PuoxpYIXAuOb6L762GMIXPh9fzenMYyCUsONssXUQBf3T73oMP
dDkijb5Y/DYjJ9pVEGjTfrnK3TPBG0tdopPa1iPjNDZZabol88iKgYIW3tAKmUK+1tgFv/HTrMKk
2R7Igr4dhzCexdL+Ym2TpW38bGiRNYAmlQ+3nD+p+Hu9llYL0cy4lO9DWlmQSykSHWzIZfD+F90j
klbwRmIUA294sN0WX4qC0uhZT7wG6Lxr/XqDcubqkJqsT04kMB12+DcYdyGuTm3+rsv27hFypGCx
YLFA2I4K7CCiyOdovfCS4exgRolWT0VHT+8Peb891447Rf313c27Z6fuvm1tA1NDr7i29RSVqMtf
5dC2N+NkQkjGABas5EpCY8S+OLrDzhTF1Lp0RE46NH98WK5MbIfKmBjnkIio6qTuuvbLNsIQXvrc
GBVDInPFxoquwXEWWFLCm7L75aiCCOhYrrgupznmp9d2J84IgPFTnA8vhRkn62HKiGiQsHfUp3+7
pjPeIoh+sliriITUs2Hy1C525rsGEz8rSuURzufhnaOa+p4S1rs+1npaLbGreVdGEUpduWjxg4bY
r/TK6ZL4KwZMZ/ARZYrHz/FgmO6I3YVB6ZbyzLMf4Y++vhu6tLbee+Ke2o6rhM8Li5hGE9nRn1zx
9n0kgQptDF1KCl7vBqyqvIdFrCDRB7HJyO9cFl9HFjUD5nckoi9LCVRGTNZOt3J5H+kvE25R3+LT
ATzVPEVbRwXOOtKryLMBkKYzRbgsWzqD3bePXJHffJ8y24kHI1tF2rYOSxaRCzya3xmtAS3CYB+/
3wofPEo5WYUNiWDsbSyK1IzisR3Uoh0pfP2Ja41b4g/zr5yuGX0HcTjx3yBagvjPH2H0oAjE04eZ
LXl0f9cbzZsFgD79elPt8g/nOzDp0KTdpcEGGjs4Ft/uF/19MFYcXuyFPePG39075Gp20EbR/f3m
B7e/3bo43x+VZvVcRK5b6iXt9YiJ7lRKvloWDTtegIvNg8tdfgzmKefRvyoEPvInJ6OwIqe04zYn
JoiYqXpwlzhIIds5nRe9y05UfSlfeWL3FWZIAGGQXabE3HhIWzohE1IwjPkKBZ3neO22T1LSEC86
YSfWsUvF7nbqSAwwFPEEwJ8A0nAQSom8v9f30lWLgGpKOBnfcBs0uoP2m9i3fCNu3QhqlnzsKCuL
lq//U6QxSp7fgcFQmIAEzA/7sOubUbQIYxB/g39r/tyHU3dcQ7HND1xq9tAUqi0vRscmlKyDWHbv
8tlQGugQkjDT2NlYBAKwS/ZU+YzochSj5fGG21N8hiBBbw0rIPjaXUpzmw3OpWbs+PTsrueVXMxu
u4foQRunq4A8+Hf0IJxCb4siuXInRcs+eHnamC6fu4dwde23aw/FihLHrHBRNs+BGe75Jq5C5GJr
YLbqAFYGt2WqSKJIj2pYMYZU4TgEz/YYMUOb8AoQPcGb3kxZK0d6HcfDXqJvb0eUk7bSye69/b2u
CJjIIKjD57dwOt+pETbdIHq69msY/HDyTRx2XoYJ+xjOmUCmqlkYRVLaTW59u94i1WbWp6W2DOO5
UXQtlYDK1dIgFfRUaYBj0/RMwb6a8Zq0sP9xOe+L7ZYzcwogALPq87wV90SkkOvrnkALLQBZqEF3
DHer9Ct/koHEfuKl6LtAmk8utH2EJYrAf0bq6p56aDWFuccUty+KoI5wMeiDW0UGJAyxgL4TeTH9
rmBMpVQKtE6UayUcKyQUlZYF1AAf4yTbqxGsuhm7SZcQAuIqjzxootuB1z7uUK6LFpLjXf7xYFm8
fr/riqpd+M/bj9JTdUisP307biVcDmiq38h/JPggDYxne19ACx8o5CCqSKFfJrBaNCRRJeEKYNSf
WTiYLMVdUFjn/ZnUR+kBwqvkYQnAtXhs3Zy34I882Wd0bRqiDwW+oUaOXxbSe9j3ujlUhTCzzMdj
UsT6OnelNDzjs6WFrw0d/e3Ur+yY7mlaZtqNr+Fnx+D8fDE5WnvCih2AX4F6/Cu8x2lgXvSuBZMU
Frik7F3Vql0sPXxFJ96cuFAiqZk+RDIOQC/YLf5zyoUjaDsHVntGdxJo5kGM1DNs42OgKvi0TF2A
NYM2MyOtYK4FmWwIxCX5V+16eJcZBwkM5YMpWASqEtlScl2E6s1AjT1krSV+I7dGD79mg9Yr4YII
O4rGg3pIydxKJETgUY2G3MQNmblfA1VVo/A8olBTi73PIk+7P8KgaVJEeX01w+RhCaKxgDHHZeL1
EE50TjnSXBbgaWbsT3LORrCuK5vdUb3A94PL+aGUSYZ6RnYrcLtaPCeVMYKlApFnQRfhNZom4Bsp
5NW0N2pO7pzXhTMcubgZKuMz8kySrz03m5Eej454uhs42norAZSrmeiJjnUkauLB9vAZnmFDhUwM
T+6Z1SZjvg8cb1GccyxuWg2wgsEeviuMnTlpkIjv6vgPY6vI0uxeaAvdIdWxXlRFaRGOVUSAOZUY
0GL5wDCqRURJFvAWcTUpDozK0ulycnFOyqyZzu0hRJ6wPnmp+evxGOIaAuM1Y3AJReFuaUm7HJ/e
oSdIjb2f0hKRviEn+426Bjfvxw4HK0/1PiAO8naVTFDYSQQ146lsYGb0PV6CeOUn4H8Btei6BFIi
UWBpytlvx+pHhtc6PTjuwsyxRhK8LAgJFJDS4Sl03eTC3gTMEMovfK4AS9Rc5VtXJWGu0t8WRfEF
4nAcYgllF9zmY7DDiSCmmVQRNuR0F2tcgSIk6+TBngXLDNaGXNoUMoqOhPhXXHubuve22N02Hedm
xzqxFm2UrPvv27/p6JEK7IWn11gn9wjvQQBDl54HitHE+7aYJUgrXSkLxKqiTe+Jug1BLVx1pbvN
AjAps9fWHkeDtttu5Pa5By4KO8OSOKpdGupf9XpFFq9lDUmr6u0lwJHsnws9e4qwJOcyyKjXhjzb
PoogWvCHBx05C4r2tMHkL3hVVDoZveEi4gkh2FXuECU5iJtAN60vEZZOR+sq8xA7EkTQ0bbLmxbF
nBa7Pku36c5mboQVFzoYNSmJ9mTocozAcLpmP8HVQbWslfYNfnqy9alJ95MoV2rTFdHPf4BiXl8X
MvnHSt4m+EXGPMqVXPGtJpk/5nvkNDNx4OfBdQ7dDq/gYofSIatUs0YYVC7LMThwwgvaBE8AsprG
jDtq0C972XqZuWdKtasIAYwOvG2o65eK7S43JF9QEs6U/37X43iPB2CBApl8QifzPgat4jfgBweL
BAd0xEEafZ2FX1nYGtQlT5Ob6h1k1aQFh5EeT66kSzs3sftOIydj2/Fd2nhe/n1/DiTUXkTEizkk
2oJxQSM2cVhSyTfxV2jt/iPvFXk1oGM3DWhL2qIgSYT0/neqlGPB9esRWedv5kXvq/aHe041QWcP
qK0rtLnOu1cdsZHz+5c8xLWA5Dd4n62hsbsFaaTR4I6O3zBv14bKXq88iJUG9nGNCNqdbRO3C4BN
SGxb1FPQfDNcsC7gvSPWl3QfMj5cqpjGkFVhK+/tQ+uz6MJgGeUYmZgXPWV2V4DhDaTLFcz0w6LZ
xnS7gng8NBxEiPLHAKJj7jHZhrJNvp/2ACp/CTbxBJn9fAvsX/S4WJHY8/zv7pM4X9P1wYPfFVTZ
pzH9XBWzNP0ZDltn2bOetVq+3qiHsLHtsPOHEpc0IePEwcH3feqBr+Zzz+3pdBVLHiKULC4pH59U
4FPfLSoatxBtcARAJzhi0Nm1u+ZsupSV/QDH33KWKK+w6bGkl7gzrHQtYqDwv7sR7YUeeOsR+TMN
VunB2myXMsPGuSBGWuyBRz6NGXfCpYn9eo5xSA+otIjvPC3mhXARRejA8XsVp6L0F/OHjY+27St3
pf9F/xqmNcL8Amjqc7Dof2Hg24Pxx6+7jExDf30uyjBGwAj15jPVRIJGBShVEa1xWBgPQcl/kXiz
uyz+JPkQjx6cQyNqrU2GDwrHnitmwtr8D1bc889gJYoWnaO5+17/F56PJ2fxE41p8G7lDOmicAje
qvOlnMynBDENSFjnT5dYLeuQV+hAcD7y08RflTBsiE57TBkiHUuA9Np9dt7x+JkZc/KyP4lHYnNI
klHwgk8MQ8gEAygGPsYb1pGSvzH0rVgp1RaY6nZkNfYNvpAvDavB8hWmBhtStupDADHVVN6aIqH3
n3UQVXE2gCpvthqU9Ou82ySJ23Jgldcw4p1gb1Fe3FxbTIOn52WvD2KbFhh09fL47j0QhLz9gxdp
4S0wa5J8+qhCimAnwgx7hBrGudL/1ip8hI8Aia92e+06Ex5MByCKqoBhQpr9w13X//DLdgn5PV1U
CYrpkwsXQLHCL/Dp96H3XLcU4xIRjsxuzreYcGYwBeOKQQLUZQnjLOUdR/pRoiLc+9bBp2h/HLt6
oT5e4DZHP1eZLn/NS4hAya9hQUJG6EpQQgVl5XjGTo6xKhPwnHYXdIbpJnNU5Gu6MrcSMAYtgKvQ
rz9kJ+yULY9jv59q+akCx18uDZw00wUWGL6G5k3GVv+khmEsdAnkP2kr8Ve375PxpxWHEUNUEWw7
1YU9TsWkFWfEgv62ghZeos3+UmcM3F8TqL7fysVlavTwZLFhH6TV6bKDPUyn+Lud3KPZcW1RvaIC
71vOhvv4UKQMhEWusFPA9N2VSb853JngiT8u95PjotdJkrH6QVOPaBk5AS6d2lh3yRk15FSWWx1T
Cm6ELxBePmfnCMOWZBUF1c+gXFnNSFQsZSGpBlSXtka23XwZdxE+gAfRZ+24AbEKyF5V2ykQCFGO
vVNum+DTfb2YvUUL5daBWDyOSRARNss1YZ33dG7ThvimC2bYYztqE8uJKI80RBTgBb7quA+T8P/C
cItAQqmxbyePNvcmVpdflIdbfET5jPHsBzzWP7JY1PmTSJwOCZgj//yP1hKUZK/avXk93pFstOZs
SvEGsVro2pVV3S/IyVslGd9gQpc4taNCaTN+hPVWjybTIPOQ27L0aeK7U9WL2Z5HDXjUhZzrcAYD
uOwsAPWWDXKoMV+OathFN/yZTAexB61fIAAsrIFaN64HMHKft6NSyqgoWLgAS1G8PjVhzWJNWuZB
7Kfo6Wee/55xlxWbZPa1AT3pQrNvYCFlWW2m828lpTdQHBnl5KocuzEv8Xx2Z2BRKxz9Ll3kiAKl
Lh+z8cv1ypEKke20iUP6ju1g6nKT9ZltJ6FIGx/DD2oTEj2MZwMF3eYjiWMMzhxddb1XPaMpHVVh
FEiLcIUPy4McbIl5pMuPcIP5O732PX3kw1YCCNtxIfgD6amNz44GdL6q5lUHRum9zGFXbndpL9u/
ONNL+pmrToz2RQs4bcSUXNOQ+kzOvcd+lNnrACZCHM226qsxhnC/59wwY5Qt9Gt9uAAVbLb2OXkp
/RghMaXI6sm8/Ubtm3qGUZL2fdQbgwpW++Z73mhSaTuQ/7ibyyZRLWcSaCPNxG18VOkeNzDdDHvz
tZD24vuWw7rIyg+COqCb12X+TK6fYgBBq6ytwuykiYIMso3tFcVktqmndvlepJG69w3eUD5F/N40
UDtB7WkHgE8pGwWz2yccks7oI89FClu29a5FTOAX2Ct7cLDOnrvLr6tia78YEDo7NUY5viT9heyR
/Xxi52dLXzb0oFYwdsyaHdBW8Y5x9s77yrjWJIDV7HHsNRP/tYLPDvGt3HM2BUkNwju4lSRhlQIS
yJubRU0L43kQG9EnecYoE0qqDTNsNl4zHHjdPW8PTOy8e06EQZ/KXznSLjFasvNGSqxkx04UZiHJ
fofguTGEbW1bNGths+5R2LVl8Ecyw1VfpKIyC/Eb+R2+J9/kWIJRPUilp/ZMPhV19nuwi/rE4AMt
NK3N+PmbIQC7ZiycixqYzYhaPWhXHia0D3HQV2Ow+LOjc4brvBrKqlVuy3RPTl1kuY/FemP0oyoC
MLiSX87IWtmUIEeLKz0jNUnwckKvyNyHensBSgUPN934GomEFMGzS6p+O0KG8nOGqn72WI4F3Nur
2+M6wK4HecUYH4+IZB5Ur+0Pc/xpv8oRbVT3OsWXavyqTmStjcZx+XT3n0fZe7WYTjZc6uobHn4h
ROdFaNq0odZdFmaaPfEOrIzm/ZwLbDCblfHI5ZmUdw/+YTbOXx9wXDQeAJop6YoG+m09Uja3Ceen
ar5OMW13bCsf2KmZrBYuCSNz/j8z2hZeYZkXmIQAYEshAOkgIZ30LQNKTQrhDdCVIKDjW86VLGek
BQcTDtMqxF97KD7sRDuj34Jd/huuC2/Iph5GzAXCNCgDx7caCLwg7UhGfPdrzu0lI4T9rdqGgzaM
G+XYqN5C3Z+0P/vHYMdZAsxC2AhFi2I4cNjCJFK6SlCPJrZLljWs4LQVdlzzBw77mMgXDOtSBt0j
nAd/VuKPUfmfkiqM6l4XLgpYqGxQgFeBc2eT+wzOR3coF2B+ftBJ6jJgEEknBQYqhVd+KgSnGWF2
zW9GttSg1TbVJdiYRc+X5WrFI8PnfWint6oVvSF2S8dvpLiAzh41wU4Qz9udFAag2+LSXe66Ypra
Dire2K9W8p3PaZzFWvcFPJTfOo7HekfIQLm/NFyS2TsJscBFv7xKq7yBWg2sKm82KdZPcAf1Wxpz
OKyBAytDhERLqKVMNkMyNjW3Bzzm1q1CnMqnjDiVjdovISlPcP5+4aRKp0qG+fLzPnt267ss6f7O
d2O2MWE7sXAmzDnQJtJVkBXpYFiGool9yx9ajoZzcgbPmt26lr/KXrcUYDSaOOU+lbxVE3Nvirq/
H3hvNKNFu+1GnWkrw9171YO9zQTJWUJQMIiwxcEO+4tYKOO77oMksD9HI5QGEWqvOWcIzEIyPiyU
GOE33/Xibz9eM67fdVA7v0uQo72mudWs1Pj1lGoqVYxdr1OvcTpXQZOEuHeozYRAgIZ7FlJkWoXm
Ui61Qr8buEY+NM9GLVxWoPA+n22TQcK2u1rRCpCwX8irbIQEBJyBSNM4MgKU8dXXD0fPyqO9HCe2
uQTTQFbWoVu/7AKzfECgCf38mxRgGZn056I9eXi+F/tHHRH/VWCTEMmOahojCVLPmj8foM08dqoA
hznGfKnf7sBwR4jjjXwbNViCM9SybXXf3OnS1aVIlsCeR4GwZlFN5VAgVpJE+Nj8d2QOSG14KMYy
+WSibgig/AG+JGdpCU4k11iNXb1Uv3PwCoCpBd+kJ8SdAJP9ODEyOAyGzkhQ5pTbS4tOHUCJGjLT
X32pmwysXRwRLrudoABOlJSqHI/soNGiGkWptTW6zZSIpZQh6SX6uCVCHBrs9pqambAsubZJQh+/
km2q5AG8vLMffzWLuY4G8n/ndsXtHImlON8faOezj68yl4SCjEXQjzmMBLlf3c+VNp4LW8MUliwZ
hOTP+ZIJYitln3J8M8dA0jcSdYGCAMfh3nZ5nCyP5w9VtaVp1QLo2BQ2I+gMg4ExmzNB3gSwcvf0
AdQkCfKD55bJquGZLLe0veFsxZMQYNlEmc3B7CIfSBp/Rl5NDVTF32+sBSzuAFkbTyaSqwE9EU24
GUQsLF7yvMnXZNsf6mmT7cqoCzX/wclZesnvqRQlQZoFvmzX/YFrrnnrf3roHWQnTHCjpuBk2nZA
6NEWLgsmRiCsyHhjT38q+SeXsUrzVCqSPpCqaG666Y9TAxzqtV8p3lNRyutFEXDewte/mS7jKV4h
NMoVYhRAclzYCQ8i03myWTHNJiMNDOdm/i4nHqYRY84EWK4AGn2CrkE96n5VRIVJFkfRzpcVl8xn
acPPqFGa0iHSDIrtChlpQLG1IKh4JiZT9u7/OXbqfhoxN02PqGT+CsA70wW0FfwA91c0tZ7Kx86x
BLJ+xqzFzH5VufjpukMbDdsW7y4ldvU8ZuufIYn4e9T7HvNkgrUIMHWjo6b+teldDOAcRqOfcWCs
7s6FgLlLNkGpQLvgL629APavOF7ZZEBRIgt6p7SUXFG2j8Nd6u9grI4um3Z1/b8v1UIjmv5UUI3B
iT80ConayKq5ZyYPOtvY2zKkokqRvst/C/k8JWdtvvT6KJvffWuzErP1J5hLkezWBdyxfVugyyAS
iIV9nMOUCwdNQMJc7+VQVQkD6bQcS8UQzzOCKtGgCku3hlpweYVJNNwbVqL6KZQUVrMUjioQDe29
Zs7IkWmrU/XCR7CsBOBbteNvfvWddaKQ4qE5S9X2CQRIEN/Loy+baLzoNks2nLArQ+fgmFl5+me3
5wxlhokKKKsAD7b3YEeOfKj7X9x0sXpkv+88yagkcrC3Zk0UhICKZp+DykZPD/Enq7wh+Abev45b
BLd199fISBoVog0QzLeXhzd/EzBzjn32XEf5gXkUIJ27xs28JVA3Cem4TR4F8MA/Cgdw2zg12dyK
Odx/7WetzOgAIjlY07ulE8xV3CJpU3fTVeMyyeiRBnB3EEVjW6km73uG3vCw22Y8D+UAEGAfjZDH
1Act5uVJ7us3tZS1Ga0cc/JuAmuJdSdUD/yXDXU5bVw9S1EFAchDyudj8vzikdMPoKUu5sAMC5YZ
uRlAVU0mm1cplhr9PNJN7dPrkVeZlf1NBeTubx23ZJbupLvCFyB/zfT87j95jPAE/Pvcn5W2UyIy
FTSGuKmBkXb6s/8IGueAn72fM7T7yDF1avwynSIXy4nPx1xjsRPqOmOG7AVL0ejrO63sea3WR/Ya
TxvPIxZMIgVJ1T6ZQxXciw2ZmV3zTsk4IQfx+m8TuDGVoeNKadqPC7L0VZPBXiN9lgDIwDJnx8cs
F0gSsmYIjqqUOLWnni1gbapoELbsuCXMhhv8FT5BhAmkT39xBcst7O0aGVy2As+hJvTpeD9kTK9z
b5qHhnra1yc4AmZRSuvSLaN3+BMpDmqiOgplUxmnE24Jg45Kb1eOrKXzPYJUZxHjfRYmv5PZ16gb
knhTqpLWAtmj0nvfdCLbpYyFZfuvo0fJJKDlLvf9QGFcgRr32pua1MGNkpKGYrYXnO6l74xATS3g
Pj4GLaHUcRaqhncA4OtEEYxkwrw+Srgj11Iq5BdOePtGrMm6JRKms2UauTw5XiN2JmQgDgUVdsAM
SV8+aTMsU/rwDqUyKqct6PF+S+Mr3mUryvoOK72NuqMh/z44TXv6wta8lj15XRmfdlNxOtE6n2Ih
FTPmpBvU4sX6/58341XsfAxjUAZNc1GmaFCANGUf6erjia4GHJ2AimtlIt726oSQej34sZszkji6
DXHuuxkSui49jqKuFUl095g0XtyhYETa0Cp7LYCyhTs5rjhMfHLGN+monPfaTSY2y2+g19yCbGLZ
fioeCTGxpEr/fMoZ06yxH6sYpjFvKSm0atLBq/4HpBtfOhSTKOBUvIuPrFKbZQM5fQ5OrMvVjrE5
SNuP+ezjzyWs0X5PhAwFhPsJU7uKiVtg6sdxWDkcxLAA6lanNWftmHv6zIVbvbOfkrBUZcG2yvH8
1vS6KUsHYat744q+Tq1KYtl/weci1iy0QKsZCDkzTlesruQg+YcmtP6sERdUDnuI0FZzZKtn+M1L
jAMXdr0Uv0gznvy9EaWJic+I4+b1FIMby/TQCreXxIAMQsn22LyOf6B9+HOBA3htYitcNN1tWU0q
eRfp6FKDuCbGC+I6cKs3CNcbuGRG0+51UpxvyxHAqqqbtVSXPe7jYp5CsTv4JuMy9+Sqhu4w3KG0
k8uLn/OXorTqWggUUQj0vEqyRwN+f1yfM1/trKR2RB8affhlyAQTQU4ugm8tsPkMzRtWH/6JvJ6O
9TN+Rho06B5ytGkoTjijABRXoZy8qi1fPxOossuXDvHk0IYX//C1tNzOo2ap1plNtoXSvgzovW7+
1/XxV+71SpdC2c1Wpf4YEkBIuzAIKBxrbuHOHVOAKoSfZ5bC84+4+IFuCoINLvtxGNZOr8hyNg3+
gR8GXvJvZ+3Rm565tZ6XoLtCgDkXcRq/dsOos5Iq7owi6ti0DauH75TgF+pxLNvEfU2gB9FFO1A0
fn9xFWnu0o+0KPwfvZlHO9pvAfD1yhBRhQSrXSQBim0WwhA5bbu7H5OPhuAhqyd3m2YSuIo3P6PA
46h7EeOvjFcvMlMNabFrlksGxL5SY8JQteEBiWYkIclZO/uGhISBu0Jnq48R/PTatz/xfZ4QZCS/
fqe3pjLRdpmJGOShBr1/obQyL8b5RQPtzg/0sMKlf2LVHOtbxvPgpJkYLbxNpgKVtQD2wiu91YjO
tgCLC5Kobm6izIJ0ueJDE8KplYmNXOAVTypp/gNNV9SlnojCLR/6BeCEWZdsdLW2JRET8eLFmCXM
BBvBqlXySufuhL6rB+rT4xIoljfQK2rt9S+j5RNyrb+gv+tjAX1yk8vI1qL3WbUeLcaZbXPUc2I3
1zOJobyDv3HzF40UdzjD1FZY2O4yKtZn5Wal/MR64rjQ8ndtxlCn39DnhM5x8rA0pbVhZfkD7FME
Hl6KXfI//0NzIapPj7FY+jcU1NfaD/ZqcLhdiKYanXj4CFpzK/I6M3582R9kV39vjsGVbKePvuST
mlg+7AybihEUBOd/qLt0iFEKh7NGSai/UIgYxoldCOADWIxfSn7sRaYmDXUYp7U5no5jjD/yn/gT
SW1RNJxKg1g6azKxQ8KUR1DYzb6FslERKO9BdO6ubmp3NKqMhMoZWhEfOdoERUUtMLUzThVrX/hU
cEQTlDcJtctUVh3wJpeMWZXOB89KiuGMqEg9Fdm+L2wybykk/6UagTRCGgK3oLH62rOj38WCO31y
PcdfEAtVz3XgYNnLduveYCT0kz9TKwgmmtQcgm9s10VyAPyonuoT1E+XBgr15jv5TPVRzHCD6U8Y
NyJ+39Bx7HlGWxfS40AYUAnpCwI28y555BcK0iAmH8klTi+vT3sANhxuEvV4CZDyFv/D5Kw1+xAk
6lNP/IwKAV6xds6JMGgMacJhxXX7a9M+VDC1GqQ0uznlGD7BA5lMQcdk4GJMfN+IvETZ1Y2ojM0Q
HwG9YSBzWtik35cGw+Xr4LkYnqIkgQZ68Qzv9EvEAwm4ZBrqFq61QhHTDiEQDzdeneikdt6HBPUy
T7GmKujJeK28M/Z/5JnZRCQk93pJyVDA1Zr6aZwpY2HRhxOqCvDkDssKB2qNTkWKQ4BuMtsqM92r
lvt7UpUFW+EC9M1gs6Ro1wpEaY5tfY91on+qJ4mmBzXUgXrBNTJZ3VUf9W3SmofWerTgkeBwAgtj
1IGMQvyNOB7EzPG95Why0i+LX0er1Pcv6Geau7UoDyOi6iso0wlPOKZvzGkUDPJcCB2yjh+Z6O71
XeITRPx5TcGhRsFDmy89ox4XelfdJuFHAj4IrVbUPlNCv8kwxMlwr6gIXHWOnC8veUmcgcYhCMi2
vWvuOrIRWVMRmCRjYi7OBGurnQiwbFgSFgP6Jo5umFLLPvsLTrgqMWngMIEXzGAF3nKvk0r9UeKP
qVaBPvISuldZRz2CBBeILRmcGH1en41zYYyRixN2LMR0dZnDetCwGUyG/ZK+9wVixuN5cAa9GoWI
wmQilBKQX/S53DQ1Q2birywU1odqHGLB09ZYVd6ZQQh3WkOpv6+KH3qtKPo0wU/ih8ruoRrpDD9Q
zjhSTl9AUQ+p1tAwRtVOLJu3PD73z4ylzysOntpxoSPPvfmervl9VPH9IXGlK7qpmOEhhV6G15sb
T7X3tUdobEbjB+vR7JXIM3YPfPxWNdI1M4bXv00+xFZLBkM6AFo+eDx/NBwD5jKPbxkk6gs/fD1a
Gk82pG0owB0kBxuWf8DuGluC+AHqYHV3nFetF8ZwmTYpk81KCdOG7jMgD6lehwxzTnjzVWyX/qlY
uEjbOttugSGM+0DkaBQQrjTMxDZxaR/8v4ejIajbPhDPMLSXy6xGRfGjCt9x8wQIOnGCIunC3jbV
F+D+KonTKWk4qZQ3Kjvr051yP44XhuRcIAoLfSVqIM8fp3SVc+MGCbSjgpeZuFRWgp85JaFwnCMz
nvjkesam51KtmGR7FlcAqNiYVjojz5Ydq9be8apCjPF2WagUc5iaN6PODi+1ghdvuVRUkevSihHX
exme16Y4D9/bLlkTY2ojJHV4YfDU0fXBwJzjghL0ETi0hCYs3k+XedKr7E30JPkbcGFdsUUKVTrq
5VMTHen6BhwPkNtAEt3df1Yj1pvUswSgMh2TsdtPg7mSwnA7cw0AtaxIIT7EKgzM1jrkKRPr7GBE
j0cD+BU6wLJV6vxYp3J1tBbpUYX2B49o1vYCfJI6C2Z1Jje/gsbKBQEt6Jc3IzC+UEJDzEIERXOz
VRd6kjCqA+BXnwV1ZFkPtsj5GSFr3waG7IKHgQnon9HoOQWZYAkeA3Hn0ij9NWhDDFZHDoMPX6ko
8OlHpgf1lsWCgjsncq+DJxSxkl3Oezuy2w3NOn9yIueXac+mTPMZ71fEVUwkg33EMa0/giRI6pzH
RaUJBC3xzUGGIMWP3q0leKYRT2qox2k4k8WkcJm3muErYql+F4I+ZXABbTLgRNYfvCnqxlWjg0r1
TA4/sVU7xaGdxaBwt2fLtTW3z/iFs8VajYG0Ks8k7BMIjuRL1SLgF9+oKR85R1XyFLSarx7BMiF1
GVvTfZZANKw83ABp5Gpo5aPQ+fzjuUX2dHj7mh5vv4G/8nO99ddGz/bscgYMyKYBJX+0jKn24xVU
Lq7Vqz9qD06Ja0mnGvruRpcs3FecY/N18hVFVh3Hw4e8jzcFg1vO93FY88Bg9Np8HhLer3RuVxSr
fZZvhpJIBwmEOzzvo9o+a1qwysfFSX2tuSAleWrf6rNGXR8ymo4paj8yEh8UD7Q2Pu3mKv7lRr5N
mkRJ+WUy1a9FZvwVx/1P8E00ZGusZeKn2BpDVKdD4unlOqgut0cvHz+z97GYix+ifDkCfWpErtqa
J1N+Oji5UPQUE+xLDhhWlSTZAz9xwl9twxWomuI0c2yugpJg/7kyg/yb1TgwZeWdGxCxE3axXaLP
xyK6W80qq3ajTkNrUEEJ5Tl6viUoqiCE50YIUPnDiVMmFnEYRabe77TzNefNJCINbzy/PseRZLnx
0T56AkEqDk21J7OamjEhyLO/fFaLvOykpQ/u+d2p6I7nJ5T2dagCPyWY45y1Vg0lmOMHyW607zgz
XdHAhrpKmU2MwOC23Ovedur7ihFHfLt54h4QR2x0pgIfcDymVa7bVHpIIjMKUv6sJjgDdVxrZwf4
SSdAVqmivB7sYbsdWw9Kpug0SdpuNCasWYLZuBTPhsFVvglGg3o3SPoNQqM/ZdA8V8MBPfgL8ov4
mDvQeYiHTh0FVV8xy+M+1ax/UPnhLqfJf8GEtjxdhVa4oB17aYnxINPMU8e1bxjeinWThyDkmIlN
tHvgK1j6RKrYa0Zj/TPOYYsK+dt+Gy43W14AacVHJo9JaJ2zuRCh2IOaOhCHIEV1BythqKPjegr5
BwhvZSBTIpvZfN+67O/feNxzw/fRFaHi77T/o0SAFWZQsfgnJigi6evq0FPkyc+X+IsYUgzhjmYa
KCNthbCHDAnlyaHvkjC+6Sb8pkzvNxxcl98sm+tkBKSk7Nj32/EAR1VRns5AiCjT0XFvj5shzD4U
wXWAsQZ0ieJjWCZRvTXt8TY2M6O0iwGsJ2FE7ubyfvb/9KRe+e+AZlX5Y8J/VkmuCGQe2j+acJTX
duF8H5XAaA46tXmM1Iani///YFNaU1aXXN3S80JX1kk/4BuUOpGAMO07vFbh2mvTnDRyU7rHiHeQ
kqSLuDrCqhas+fRIVCg5nVkU4GcCYxIsqVOU/WO7TPZznjJOYKA2pXD1jMhFq91WIEVX0iQ3rdVC
SOMpFpTtU47EKKvMGfHK+nsaFtbsHIgk2pRXn+JN6jaymgfzs2WOHRxXU9DQd4+1ewGhFFGhrplc
Z82q09c1aA1nE3qCrE/SYhL/PtXhuL8b329tmkrLwyo3kf//rYwETJMfUuKzFdujoVNmoxuSzpZE
0OYPhgYuuLhR/RxzLa5Hx586MBaFHdZYWh7kC4INMuxz8XIcpzHU8/FgtUY65I13Z31y+xXDfYYt
1eTEyVpRaIkvq8bCkzjuZ9iU0sx4KwaLyj1CAcjMvug/MBxFHtElDJg5p1vrPElaa1Za9A1MpsTI
rijXUB0lDsZAnMu0ZUsDt4S0XDSzPLi1JDMDNO8TYpBxvd87+wLn+G+CA+ULfoJstbzaMdel4gLC
2VHnGKRKvFTW5grx0YBZcb3QnDOfc+f0Jo51dZ7RKfFfHvd5PAXDRduoZDH3mBncBhMxENyUC7qZ
PIZPpufhfoQS57Z6QOE00FMp9+5mPYMyj6rJQGVhg2hRFgtAogCjV/WyoUW3iXUV8zC4rhRpa4Yr
UEJxQiFdlcvIMJLL+B7OV5e9Hx2jaZwiSUwfb72QdzZG72DhXjfgcfqNLWsEXOtRyvi11mZb7U9d
2cd4CJv07MFasRsmus4/7jJL+f8wtfZ/3K9b3aKmHtufuRGmbGriLcNize76WEKOAsBKWIL/bVYf
MGuLM88cNA+4Q5BE/79xgLPOnOWdRPAgHsn94oI+pJqNHA+p9DiKyt0/Sp+gSiDxjE3bSCoJamia
C9TeWMcUX63c7/BF80Qw4vPgDi0MtNItNWQwmmKCS0TIvdNv+28nIi+V/LAxHHc9a+LCwm4ZA1at
AeI63HHlUZvnYkmi/1UOEfw32JRFbpFCifOXP8yO0emmP7UCE099Ii44agUvPDSvf95a9Pgl459H
KOBA3IjV/DF0KibZphkryD2nFt55zqd19EISsxeElcHRn9NinkSVcf5iY5fD122dWkALZkSL6B/8
+r5Uh/DQp0jSx3OOJw66Zrp9ADkd6umEBe50CrlcTrn88J1krYz1mANJ9xRxmGHNJFY4ErF8QjYR
BabMb5r96V9NOnjjNAuRShrTq+yYkwRcba+N+irseg2V5hoCax6K0ai3NNzromEMZ6YKWDs7lGOK
qWK/Z3g0K49SvF1YvLZS8K2GdSVJ6Bb5E/eZMG3vlZB2FZvWbWOaCziIaAGmrMu4njgkTyToqD7h
cv8fvZccaJZlyoPc7HXv605mr+hIUJlIHTqEP0NWBOd49EA21mdLzPIcg/X3j1iFuzL7nnC7lueJ
ue+dauFKmW5EPZw4oRuqQt+OQkXXZxRw+tU91x15Q2MuWf2FDVQD/YrElSc1y3w6dv2znrWJ9E51
iyE7KoaPCGNvod27MnYWFcEVgDBPIxdyAdef1jbRebPyw7odKfRHBIOGaoAvxkx+5YAHcrmsjmBK
Kl77oBScsZLQHdU++T/BnvST17hmCnLA3gAl/i/c43wVo+8jBwUdQUEoTaMs6rfHDTuTRcp1P/bX
89nAAAJtHKS4rPe4IAZAzsETLcJkNP2QNkqg+OtjFur70lg9Gn6fSCAD1/C4YuUL7zOEBFHSWe/c
nU0Tj8D+9kYnxAcOk8f//3lYuSoPepaW9cp1Kv9Cn/VkTdeYCGn4q+5pD//2sHxBVuk9M5mtIiif
jdeZaw35d4B5pqTfuO1lmHZNP3ZvxVVbmF0lhRs4S3qkTIP6kn/Vn9ppJt3FchGEm4rfr05y1fKA
bkVUNaCqsk3273Hy2cix3sXH0T2O6qua0Y8HIbvz2sJHiC6nieYWrZihA4vyE9awLNanZiVMb+ET
FoEvDWTwO9pB+Nb2S6lWWueec+mRgjJUVPtKcO6b7/3Ki5oZGKvIeEbddX2M1RovLLD1QJBZ8yAp
3ygf2ZRBLyknkXpgwX47WZsALJ8XhWUcIhcSlrXzCdEj135tuAZ0PmGg9b4Q4Dn6ipoZGD5bqrUa
4nkVX52Xev/GbnsLpuBNAsTtkqtI/Zu+aaXpJ0C9f2DzHmLThCH2Vd72oP+UsLFXVWosor4GZwAm
sNsjp952pFtbJYLvq3PaFHE4TvexXwJ4sX4l3CUMGjlWBXNlJQwMSvNtGBAbW3CmLlnfNdC7EpTJ
OS0V2qMl3KYNTEdCazondSePyTNQXOsNYGHwXKGjB3Glko6uWjfC1qsAKOlsGNT6o6XQTM1dFBMr
jQVWm570cbht3XRQeVtBz3I5vaWvV4VAeFnZPTz7rbQ/4DyC2yrz6l5E/0VeKNWE9uPPyPMQNFQq
mpn2xToOFswBGT3K2T0yh6NlJ0rKC22NEHy912R+OB6hwE+80NYiFnimnYhy+eu9GLM+hZrdH8Cf
abrHt8KmFIKfJSjSAheK4atUdG5v+XnljmxiHzY67u7UGO9/f2qjUZL8QpOCWcow5yAovZqPQ+Iq
qyBGQQSnmOSd4EhuGURTzVen/7CrHWWlAO54uso9DYQqUwyO8tJ/qWBMXJoBtw8a9+9uhhCfJb2T
OMFH5i7SmBpLCphSJehN/eO9Po+q9nCd+9rWaE3WWwH7ptDA7XgwYQnUCu865s3FXaKciF7Y2O9Y
fsNwvaSlNOskW4+KlA9O2omQC/K+UWMU4+dBvYYw286dbJchcJEAYiREBYtb/abwYAGCvdqu15Jy
TUwQXRCSXWJ0ZB8Z5r3hmrH1p1pIBBIX7yskwy/dy8HCScotoKUDnYeTwk4T8BKxSwCrP9Agjz9f
hY4dJjMKj8cf4ZQgemjfXa21Xi7XDrXOGVHX81gIDY2+Yhrbys5/Agnwo/IwWhEaCGkXNvSNiZ0j
J0Xr3AwinMYJ5bL3JPVPMJ+/RHM6gaQmJ9uKFPxHunzBVbSesWsqfWHdFLinzeRZx4FbF9/4S2DE
MACdzSwvduDY1UvMc4YyvDoFnDbvVjfoCuVfB96fbg0AmTAVmGEfQLyMKP+jZAjArrKi20hzY1wW
104HyQVX+iUutHCvqdqCmhIBnL9qS6L2TxQO6UEL98J/bSC8rQh11oGFeNBD4y9Fjw9izX5QXyvU
VgMOPV+7NeUQyoKy5bhhVbLEypYmxYo86DKkMWflBYvpkBmCaFXLWVDFu0gbJWANft/LTKFcmFrw
MaQ3jGrna25Gl+gWt9MWDfq94A+Y4fm8VnKnVtwyURwzAft9e/PpQUsckMqlALH9D6XITr+4DODi
nAoc2d5uEtDTzlackOBsEeWbbvMNP6iIHznuMgaXZbC60QQ5YdOzQGCsAQP4pEmxOb6diunS9zRh
rI/J4Tq4fKbVvmCCAkQG/0r4MAwKJJTcC0iPbC1WMh3GajQM/uWE1qGjyvM3y/sl8sLOjffFpSeE
0855nV31NUOMQk57vZGvOVzNZPOpKUxXNROVUQKGkMWIXq8UoM9wbKS64PtcTVOWhUEbCoBrsKRV
sVjWxbAWyU4em5ykF2Bi4wMM9lOMVEYBeZEOgWa8oRVLAdMlMEuZpq5mDaiaTX8WdptTBddfn3/m
EbH1fmPsFlRP5rzrlWFCZJaEtjfTVs8I6/JKjUMGaFsBxjTkL3JLaWojrekeWXrsIHxUi/H3ldj4
NqjWqqv7wtFOfikEk97xNTB2SO4j/XUJZwZ2+Gj5E7RdeS84jWUwxJvUUcfzKPHzrQhvJfT94G6Q
D+K8qGC9dhrT2KmRRAq8pbfqCyAwJ8KyaZiReF2w2rIQunXoiawKE6WdTpOOk5BcAFqeHRjyNLRA
LRq8TcuijqszonS5jmGkJQdYQy3/8wL65v/bbfUoj73GerZy/I2ReOVdGM6EE3HEJbuBNjU9tEKn
09m5Rpt+LN2F+beaFWThG6FDh5bZYvFf+u7Fz3z2vgA/xStPRWMcm4euOxMW2sGZ7yb0dlc2PFb1
5STtrnLBP9rLpxhMiRi5rRRcddHon7v5NJv8wfWZfGjfcfQamNUivZ6anVbLZh66uVpF/tqRHMhn
zMjMk1My8TPV5uuyXmrfCSojZ9n4bDe2Kxw+79jR53gbqm7dRU1Fuw1WvG6Maq1eDScqb3CknRCe
vJ7YRBmffHhoNnm9MZ9+24tntYUTiRWpULmVOoKx2loNVFuwvDjJwHnIjbL2GKljAD+OYggcbInm
vJ1GZkZaXG7X97rPN3FAw1RnGxrJOC/Xs+8hBqpW+Hi6Zre4wAAImMulMHOSIGh6WJyowrbvO+Cb
GpaBf4FjAlhjyBR50bWWLj0nbCxx1gMtLL+7BM24kXUnPjnilfcgH3Lf6fa2O2zSBIHiTWJVfIgc
GW/E63ZPUJZIZCIsR96+fhNJG7E0V3t814x947RSpISUBdeX1AEvnfyaO7rFBhJH8K/E0GvtoJZD
rKdJWeHZ0iaHa/uI1kw9w/gx9PHZyRrz+HLYlTwICB7uZTWIvoUskrrMuffcJoMGeuDGOTnsO17r
VbaraNvVQj2kcE0ZP+dCqbtPC71m5/xBImEwpjeTkTAwXrhH2rsJTCZMLa39yTkYktXw/hVUL0Lu
e01DU851gmx+DZwu7bckHgq25awHbhqFScZz2YPpFyWacNzr4HFMhYprWmQ29wp8nNfG3TQdvmDs
qmwUfDbBGt6X/jwlBOxb9dIGjZHYP+UrPjSk5v8q+OX5iwIPTOZy66jUv16AB9ZAU78W1sDRP3Ja
Ok/j5f3tjI+AbAr4asU+fAtehoDc5NycFPcwVkFWuCs3LUEfyYiVWJeVy1dl1dAlgdEIhIPS0Onv
ldv7m/TptkfW+3aIoCZszBV2M6Bey+RrVbrxFFGAg/VJ845+RKISOw5YVgJc58HXdsne7w2G34uG
8UxnsuspFa33/UT/z5yLPDX10ApqFJyhASRg+ScpdOrg+CfIr7jaxOy84k5ny73o+zTiwyVqO45i
1pqUZxXkcPzMnw4wLyovvsszyGLrRmxioROH7lLz3VreWyHmm0SUHc3BahJAp0GnIEyMRL5WeR3m
czhg+ebujOhoE+h4FsLYJAnu2n5xJvOc8WgO/ox8I6SBrK/AUdFzy5gBAAIPIpesMFOw4fIArYG7
qSw/hWF+KJ6ne8KytUbEuPq8FHMPPVPPYIEWLh3rGplELuKqiSEFx5No4desk9rqxZIozhn8LtAv
nKaFbGJbtCXHE4jNlMwf2H4n3uiCjvrgw0KO3bD0Wpd4EEGq++XrDVDbltjNX09ljGJ20mwKSKFG
dURTupkfRczsnu2VnF4JessN3/3Pqo9elGvt8Ce08BmUySi2wwXHtwJz70+2tAXLd6oi89riFHzn
enpwNrNDf6CeyV75L6jaxsTNLroiYFkY5EkYqxpVbd0ArYn0t91zpGQqew0fyJf9o/xdnt2gOM6Q
9B3cc6/QAOakj8Z19RLl5lgvGSDsjoUPfA/xYi0eozlf+YH81BWu89M6qtp4i1xboBURqY2TFUD+
Lffx5gNKIiIGqFEKwSK7tcBTGpDy9wZvQXUXrr1gZXSEh2rW0xHqdVGVrU54mNAkKY7gKliaOT8z
bOa3rVH16INU/COfA3BqMnTQqRtzQ31G9d059kv2/J+qC9hNp7OISQdq2uGduoA8nZG+35SdJcxV
MPglKqgFM6vI3KMMsWTTROX5HTD2t1C9aJu7Jkh4C9ILYviX7cZs2kaITwwe3Lr3qtusGFsNPxRi
eRGywHrReXbNt04DkifI+Jrcg5E2FqIy/ay3CWgQYpAAH35gysZIX/vuS1EFT3GLoqUX5QEjmoVX
E0aNCDCw816z5lq6JY5I9HnG9nJ8a7hjHABXgeGcl9KSHzGT9whtbUMqsplkjecNKQq01mK3OcCT
71SmiK4NK/MbKqcon5Fky3qR0Bp3cRaHXr9j49NHQVQdjQuPYGTcHfoq/RpivAUFg2nPHk9qc3Ph
P6gCEG8eTjlAPwuQngnsEX3KhzPWKwMQP1kPfPJonCWjnU7MYDlSVZ/hGLoQU2tWdMJZbvJ636qE
xTTMcIVICjx2iiflstwWr/wk9dPYjs1MJv6JJqhsIweLixMIR+OF5NJvBQAfgv+iPVmaE/ZwN/8u
OyfUTKWtd9OJDHAQxx8R5TBg1akWgYPvEcCzBusTHqlsSI0Jl7XPTrkl4JflpB1yN9JcwpqUM5bC
NS63LV7spBBsdzrSQuMb+z3oaAS6ehLzZaa2Qptla7WGBrFHl0uJTXlf33jlo5yITItn3R1SZ6v7
JiOYbrJKx0mHfDUjUXI/j7Xb5oyaJ4UBDH7jHkPTUlJ1VZX56Aw5kGlwUxM91dqBZTeGzCatNojv
xc4JFlFrjx1qPUWUsJOMAHTRQFelOKtWqv+09qdU0RebKV5Ol27iZGECsXnfBfky2V7Zj6rAUBF7
/JR5OetAz4wQ1k25EOIQYZy6/JxEN/v716fzEcdQ+HXUxr/NiDgea6bc5uKcMnaxFlaxVOOxP61l
DjpUMe+PuryjouxOhaVCUxaBqi19KngJGHvWUd6/YSX6QUJEPFpUyxyLDw7Sgumwjh1o20UxveO3
53wJJOX/oz7JT5qUwHHsOfSnp9YfoVDf2PFZqOIJYzyOjnMZuR4wPUel0/8vlkELPXluFe78GQGd
Oh81UuzrI4P6w8MwbdB2yXexyBHziMoNIiQFkFnIjPOSHhqaNtiziRYU/wGrZKshvx8NDW+0WlSI
I2BxFUO6puGiXgMDQwvzomTBoGE0jOlgd8Hwu6ypH+yjR4revmfMEm0OxH2e/5etPYu6LRHb1QUF
ZzSK4a+QgfLozJpX5ERnbm+RGnHJcwjW/v9DwpgKqTzxyfM4Bhv+odqR3sAkzcGnMqprgkm2CmbI
1QlofrTB9HfpHQK4mDTCfIKbdDZ3KFLHTRRK62hcnTJLWC5AJph5EDCZwmljDrPmbgRuTMBSJJ3p
O8U+tIclmQ4gv9p5vgDlj8351CfJd/AlIxzqiSdmoYHd4dhgAJjLJT+NrMHNfqGKWSTgua/sPUi6
g7Tj1abt9CiGfym1gqMheJ5NtzubqMFI64oL0KPReYCPFtTt0y8LIL1FILUUpCTW/qKuq5aqpWvn
27IwO5oRSA+rDj+bT2OmB1I3FN01wPJPkGySyAWSMMmC87O6ZaPGwwjkz4bupbYpVuduWeSgCfPM
q2j8zyck2OzqJcoOYQn6UKiyXPu4mdfVbQ2hz1hHg6koeITOJBro5L+WesGn0kUX3WXtUdb0qgWm
Vd5PeWT9Ti8okiW6erYDUFPa+FkYgk0oFXh6KbovA8Hl6sHjn5S1ZG0OHZuPhOQtdxdYbQb+Rd14
jLQejq8cCiAmI1tbpwvvnVFxtKfxDBdlf5uQ7GvcL7RG1rktkJvDsMwVvoY8ENpXFRbJ4yKTm/Q1
hL++rI49gLP+bEpQFIBTFJHHU6qkWKcSn+BKuEtsjphczk+irCk8RAIfz8JocVwKG3AeOKnBxNSI
n6ZlwJvljRg1cNKgZDJQ7oroOKiQX4ehjOzh2Qrg6P0kIGxRQtgr8DKri/HAWso0rjTgOjaM5/FC
8UPf1t87u+4Dh2c4t5zvE+3M3Oqn9W/E5skdilHeoGEjuiMjQX++xZMd38gTyGOeYLzUpeiFc7SW
n2OvH/NnVkdzYOQHhAUNrcTKIQXWxROmGbYCPMDBZ39c6CvGnd2mUPGIGvEQjWs0mYMs1ybVaBnF
PJI6CDyi1Caqtu0oxgIRGqUp/DVdveFYA95ta5OE4Feaebcr0q5bIgK5rMaF/tb+fELohKqfXPAa
2zDYuv6FUX9h2IGcfr8IHmApWC3lBC+baYFYWG2PV38gYz5j90Hu0mRjo/eUQgOo4tftHOJ7P/Br
I6RrvrE5RT06Z0qDZkgDqJP/vgIRbOzFeLyL+Dbj7b22PJbmDZUGY0xRAKPsi84kNu3BINlAp14p
uGpL+8mJFYnTHdoABphmpUe0LMx5oj9mA2VwFIGorb82LMxbK5/IVw6Tb1tU06AR3ylyeCLzyqhk
JljgdzncgQaCghSNnoiaAwzPYUIo+CfiDI9My6CUQbs/CQe1c1P9aezi1koph+sRGoWEh/JqxE1e
L6Z7W6UW3zlAkk7ejKC/X5yORasEnL2DJSFJqc+lmtBRjAUKipIPjLdkNZFlB11b9HoLfXI/NhHq
bTTpL43FSqrSBCXYqYb/3HbEeVaZFA+nWpmEfCXRd+fCTyNiBmtoT2EMx0a6Muu+e1IPTQbvxmcm
siODKht2Rq6rblbh08n3JnG7haBf6wKrLc/4e34bQtpHKIyIREvCdaBaos4fe5Z2rkVTb6J2hhIW
SI+EBMZD5v04B22wFVRKzibAlvVg8SflsmebFXMD6r4tPv/g4JoXLAbXVQH0R3JkBA9oh/cKRKYn
lHFAGKV1uZSuXDWqnUKZER+12yYqv1iggcaI1o63tOgDP8vpbxi6IH11R44M4a4WGYI4t0fIbPWq
ehlS33RfNwOn9L5rcSuVCXQk+5TzC53g7JOWD21xqKkcEGI9lhqOPcq7WEe11jLU+iO/gf1TgYle
NgA4mcAHb4/J8iiabuGfFBVZnvEBSNqmpjHP2mMUe8kGyfey2S91JRUzlIs17ndTzrsJF9cdPOv5
P4lg1508ECNZH5ytxyu9g2H0Amtx5BhSameBeCfrQbfp9AmSGol072CSugrYbj2tpfAJ2XgEawi9
aN0vdEXz65HpkjW8WnL8WkkPREcX4MmZKoJ4LVfObar/94TGi4fibGiaUvqKBpVHZAQVHqVQmhWV
nmH9uBVjci7RWxdlQpNkdDtv0ht+eky8HtI9f6GUITM0tQpgPEf8YputDju5V1sCO9t23CIwRfed
hnu46ZqP/Zt/B5d6DeKn7MayqXTLDavdsOw/E6YI0N2rFBmqpC3LkmTx5YeyEomkbo9laCTgUyNw
A1zOTfHb0L1XdHW0/CRzrKnFDFNfG9QkIb+5l/YFX6AAXxatpBH0umnrso7PZIBnpdXrrfHn+JVo
eoz6R3PIZgTZc26bl8vAsH2B3T1J0yt+g5nt8xPgg1Q3+1gjqgqKs6aRtbigksfmNw1nGSfTL/Gx
FG8Ux5ygWo4O0/S1NTB8ipsFErRvMD7SHvcn+XuorRyp2+2d3UZJJMu7l6leQ/93o+OLJs9nMJb5
NEgGuVRw8dVSqOTRrrlJuH8FxTPBQ5/g4wpzgdO4AtXqwS6vnEipW/+pabnFrw2JHAjStFRx48Wn
xvDZTnKShTOGz+G8aBzE7+hnKPUrc68+WZTlh4lLvIr8yIC6rNysFY5G8c2P1wY4MZ39dqIDJO4e
KB193uBWVjm8aw0L2iZlWKpbznAe38AQ+xn3Uk9pLeSWDVCOclryw6b9+nanrJ1D14m16rRA9E4C
dnMvyeSoXXoRlJsojnC0+Qutao3lYzfalOtzZHLbLnTAyStwh9La+pkyaor5rFy9KyDiSlnYiu3w
qXq7YyEJYZzxinJlYbn51tBAJBmKhFhUYVHmRJCnUYLUca5Ywmc868s9Ide/+G68oVvmNFtb4T6g
8b+oS6fXZq1ugZmKLkKSL8Tm9HpLh3sKqFYfV8xMu6zTWEeLo4xma/fvYkEk8Q4CfYjpA5UxyXDU
xtmU8yK8DyhTGFQ4mARTD0m1QJnX0fIHWvWfn9YyyzCqNS/6zFQBZ1hOTU2iMigkGLnxExcgBz5W
ohmQHi0/i43mULuh5pXqiT7EIR6AhezsTuGmZXz78N1mb3ZB9xJYk83Axc3huBK73TxsAqS0Tqgr
gUFnjt+G7+/RGxAWjIsti4gV/2JTYzM/xZFOLdCcchwMXbPMtLrtvlL7NpYv7xQUiVtLr8sUbF2H
RInlPgxruEsKsymlRrdbHPinqj2k7NckW9tH+nGZsIbFM9v+bX45tSkkd4IYWOFQ2A2SrGxbcsLZ
iJep/9JArIEZb/em9lc+5cyoRUSbLzVaG3P3Stz2PpTPHXElC5CeGVWJxraNi38+zuahODqCSZBg
NKwW4ChdEU9wQCSQ93Z8+3AasqRmY3n4D2C8E8tiOcT6K8ikqBY80NaDCZv0tlxEsDfalpKvZ4cE
uYVCDI9sVC6aCZ3eTEZVRlcu14SEJlxwEl3XtVS8OA6GPQM4FTV5FizN/VUMkCYWIxq6subE/QZJ
BzPGoS4Rn+W/YG+oP2d6wpbUfbvHFzOrg4gsqxWsU/WuR2onFm4zEWa5bBB+L8lcfty/yUhsSxvV
tUMTO8vM1JKx5ZTeTAC3DPxVsz5CNLzmW4XALFToRvgo15LiFpkqRqBK5O+SjOaF/btOAX0VcijO
MTVtCdgFaSyXxxMOlZUoZVPbjCnGyFROAI8crzjKzX8k5RL/FPsyCWZT3HjWWV2tEOjqj8uow5Og
ZW8jWhc4kLlPtbz5lW0BCPlqLONBI7SgE+/xN8dLsVU+g4hDRUNR1VVuZHNVvAPGhOKQlPcqUIxl
/5slXNiSItO88eOWVxgvDw5ITeJB+3mlBsZf1t+I1tI8uP4ZxQ4bvfsnjQDSMl3XoxbaWzQEUch/
WvGmiDGlfctLhM2bqZikRwtLISV/NnkGG1OEV7A9nyStK+0pU6ufeDK6Weut8seTFA0IHLi5Q0Hs
2g24r0sW7YTFrcHqGM6cEXdo9o3M7Nzd7Bs9vNy9tAwrsyjViwJRb35hJYd4Qx2thSTcoHwwZqZ1
8vre4zuIWnE0UIJWlrTKUN4HC4p2a1MNNjgxGBk7CuINaLtB4WKdjHn3B40DqjSo3Gz6wobfBlFA
7mIaKvIZJ9FNmr7WdxRYOOozX6LDZGbXGTNc87Olo2+M7CyMgKRkwTkZI6mhAWgOyKukfphzo5Nb
IQPibXR5reCZW/L7QLyUe/P0ofiHpUqa/enz6geOr/MAMYDUw8+Oqn/kZae1XWqMLODxl/h8d3lr
8AOCiLrpwPZ8VJj+xeTS9m11dhmeKT7ob9nQwUBpER+40hSIZeJXKkezuMjDEIHG5cKwV/2E0qDo
TIFSLI27LUg5c2eGBmu6IKL4OwN6ElciV+lNgKCGodvOYLkDAe/tYkiYV0SrHe5xYFZe9PP/v2OM
0sC8sSisNoVPxx+L+hKhjmciVIuzSrLkgFcXSbt1HDcPvcGla/BwgmpddFNnFQ5T41C+rNB18nyD
uuKNHNQBUEr5nURIrxp42ZVoSrZVBn/b6Mb/Cy9Nc3p0tqw8S2twZeBeQpWllwDr+VFAVoMgpUw/
N2cYhTrwpKU8uErM/0NZJ9PF7u1YKVmMoZZj6XGdjaSYw2B0SC5OnhHJ43o1I0D3A0wPbu3W7+xj
E0rofZzBsBDwv6G4/FPHi1t5KchNJF5GWvRUAoERNRfIF4HYBIVQYqUD/lNu4YXoIx2UjyuOW8if
pmgZuv+ClOGnOPYnGGoo4yrjK7nxurrpo92pekf4Y4vnhysEKotKL5eef9B10XYRAVemRNapqU7O
n7eDpleJV8kTTV1y1ijGiNtshrQEDZFFswLYC3orckxxtpuxKdgYiie7JUjQLuAhJ9ZPa43G6AUk
asv9tubJIIFrSwivn1RiNwPCWxQZD1KVGvkDnETHhKJyqQuTch0anOI3YL9gAQAVym6yd5P0wt8t
LihPkp2O+Vm5rkvZ+5bhzFXeljzKkYYHclBTU/WETdnJbYDL/krHCG08JZon8V4mqE3YtkCKAzsb
MGIG9uVthyRaPlhpdX1toOemXU8qrMZXEQ1Zt8y61e6QinXOOGufKPjVUpf3/hHYHAP+4XjZ3L/H
L+q7sNq/tbSiedCCOv0Hj3zZlfppP6oYCXczYLegk6xAqCemXxpFousreraj0OzcJ570IQYFlVqh
QzRUfDzD8JAoeL3gPIBxckcNpZ4fzgGgEofXYB+/eSfRUd7jPVACYeij2OrQ6AvoVkFBS3Ni6six
8fjP78gvNn+NqwRT8xgX6gcYhNAQBtEj4Atatlv0L9EI6LnENGkSYehTZsUKUSPDRLHBWb6uv6d3
YtAHg4GPg9xEJcQg027zmuLXh2W6MiI3D+Q5AHWGlzOi/Gu7FDK/sQCJuMQEMlwQx1nQJbAVlTNW
ttAUiuoRBikDQ9kRbCeVRfkgOMbXqLuWs7drqyWQYoMQUokpDacyrdoJNgu6utR6yjWGauRzHhAw
yEqh57KVvfGWnbvYIWV+3MeCqIeqgE+1ErB/7CWT10STPbatkSVafvJ/YQrJIL8wCH9ExsEz6BjF
JYhpQa/cH1bZWkFC5U16pJiCXiF5s9MgbwhmB+q15iIpB2F+0Y+qMqS9sMJ8TG2o4TauQmtBEILW
5CHdYj10v7W/dhlXfk001UArDuub8FshBqPHE0fivU05JM3PAeztFVbDVhCh+5r7WNrzfkp30as3
Q7/8+wE3WzWCEyVT4N9qSJmjA2rZis9bayGfLtc8FSCPU4EagbCY+GH3Tmtx5En59RFUlF9BUHiE
5o/epoHySSG4JvklSC3pAPdxFOU6+oITO3c54y/qrzdCfwKCNweR7Xm9e+2ybn9tajjzdvbxj/2s
UXzstxfVDuWm5PtEVScbzeJGC6vqSEL5m+8NKrDX61gAEEqAJBpcYzBf9A4VkbFaCC+pbusd3v2K
tPqVpYJovZ/FYW45UJKJN1VP6hBb73U/MTybIGUYr1sxdDLQ3OxWdA+38at67ayUqjEkhjxpTKxi
2HbtzUGh2NAjzOpcfus8EVNb2x2yhalsNFMwAGdWArP4l7C++dJO5GvjWUMpoXBqCs2pialOwlts
HQHA+I63X7KLFVF7Rg/19cFMZ+k199gdIlAIwwzg6nohhVxrIB4/5+4iu2i8a4QcpM0SDFqi6pm1
KPmlJrQmpRAICijf8LRpn1JYhWjCDR/pCNvTflICJjbFiZMTvtXPIXpAuW2r4Xkqdkwovqan/8fl
IUmokW1Ud5obZvelZeXIGti/xjgTWG2L+V4M6D51hs0yBMY56JUFZq2x7GzRqLWU+p0Jv/DLWBpe
ZnU+MGelAQ41sAUZsIz89h44AIVHalzHpNI2ZMjE2LGq3AIYzwg0g9y6Fdi/NoEPMzrcbTMnD9Jm
WuY0rO7UT76QX0dKFyUkWeUuSUqzfoutbkDE3fIqzdU7TYaP37K61P8327LpBtOHBdozhJ5U179J
7Qih31F8Hqlph3qFnEtede8O5amk+nQKlu5XjjlXwbcIHQ4Yj57UWqGYuJqGsus+UWWD1GlZTc9K
qL/Ym2W+DSN4HZARPotyMuQ0eMFr4HLcYI93mt4UB57l981WOJTmnagtt74brRMAJe9jnISc7v5+
CMqc9/rg/D3Z5V51ACaDlQ27O20Wti2j30+e9h1BGqQ8stuVoxhYMDM3tewHC8ezp/gnrUyLuVEc
8FqlKQsjpJVUfllQFL3C1bXj0C3cXVMJ8P4YTZ4ZdS41Leo0Z8w8FVTdve1/c2tYF6yUsWE/xjrg
Ct3X6DKbKqBrlL1W52WF7WZEhuedQNbFnC51QgysRB0ThI7Nw4S9uDP8f59MICBHkUbgDX2u4R42
Uau+FRsguIu5tqJB0DBcB9D6otDn6ohorO0NVmLcMHetcAppbje2y6dmRXS0guGe1IyhQxLnRj5r
xuBLsMJEdPfta1JtGlY8p+Gxscpmz3+c2umgZgXFlLGaOk/w3OVQ+j9lbqQIGoW2IejVKLwg12T4
UbKFCZQ+9IBCCuSb+G4+2DaubUNiOK9+e7VbB5E5fbtVsO9Zl+R5ja9HVpjYlxoFvUFhMqvJSRyx
82f2JdaQpP08NZHJ0nIuoUaVGEPQmoCPRPLewhn6kZOSEP6trnjinwLvCOuyeOGY3woLSxG5qne8
yfYl5Haqf5bXiMPp1BvsQ8FBEQjUJUkuxjHUtmnOtC/+zR6zFeV17uppFkIb3k9KCGdZ333miE5s
zUvoyUOxITAv06LfFeNGHgKGcTyt7slJwJWs1QYLn09ZkMONciymTwqvGf/9yh6eGVCpgE0eL+4E
b7UMfucjsiypjQg0zKk+OYf7fd6q59W89iGvXfVGlxX5zAfoi0jNfjvanjVpnzCESRBhlVYxTLEt
W6lL6AriIxXciRMVbMh1UkXt9VC9GDt1vqyjQeiDBpmEGoTrwaOa0LOZLSBe8xLNq+UhULjflD5F
UzEVV/2RhzUoQhCbrcPcxvosie2wXWF0hP9rxPtFcEouy1cYMpwC++zWwxU8Ksx1biWUg1ehVJpc
MQQYJx7DJVKx8WRyZrYxbdjT8dfI1wiYn6LBpeBypBt1xNLBJ68Tx5oRqGaPCyb10AV6Yc0Mr6nE
Q61JU/2jpFqqAcxnJZE/oYZAropwlbwU3Om6rK3Mf1OtZRstCzNBvxSJnynk54vQteTFvpUuLxmI
9mCpq3sEylzlAnNYDwJvSbZ/Acd48tfp3KGlNkGy2r4Vv5yaCtK5Q6t+syq5YS0/SZseOC4KwvtE
+nnrUsn0glgIwJJ90sf7Yk8V+p5t+rYIvcgjyrAH+4uMynZfZqmB6x1hD4j3FDhIb/ryvswNe6dE
CiwWvKNW+Ao6RDNcINcIoOxXbwIxds8dQxWFactCxxi9LmzlrUsWJO1cy6jLRIPvGHWAGzFHspOr
m+ufWj3SzOncJyKKX2J2HVRf/wlVP+Vgv7efaIy4I5TXXEMKw06KInHxoOO7hZbrhE66L4sd/i3b
BR/1O37LYqcvZZzbsKW14XTj91w/3bzJstHgmZmlJYkHqagoHGg9tPHuvhx8dAoJGYWfNX71Vf0W
+INbyvcEP/tF3FIGlVJAitLNMCRYsDU36lFPGrU8fFPMcGEJRzmAoXNXwqaCqWzffHdZHYkii0OQ
sjWCeOO7rdZQKupFCCvAD0R7UlNL1P06hJ9VKzbuRGWmEXl7ey+d7kL67pPtCqZr2HT9ig/afjXN
0Gwxhgde8qqsuFqMwG0R4Y/p9qQXZ8kv4tQa6QmcHWB7zV1ZLXLFK0+Jjukfeteb4XvvssuwkyIX
GpaUlsEE/o59SjrqtsRgle22i2mC2sLr5WwZZIjhnGZUYeg/iu6f5xVNPjvGAzsYBMd5QPfCRlbn
nDrCpSsHZYIuV0gHlCkXCwuWBr411Q0Gm/axL0Na34At+htcurT7aXeWLxx3uQ1oRrO8/RKYoJLu
o8w6JUCnKNVlKH+2Lb/QzxD59q7MfhdLg7aZl4mOwetVh057J30dPmA/Q43o1KgOe3KeC7RXTmqd
tgyp10qoByfwIjLaAgGO9Ea3VHBrHeFXWZ3dCcbW2Fjpc3HA7UUiTRFADt/6bB3TMuJIrnn46qxD
8iuJr3PmN8/xGMP9DiodLbUoMowJ8675q/UPCSJ0EEa1DAHZFG45hn4OYWZuoSmnUbsmW/Fa+b2s
DNa0z9iu3pdffd7rymGUBjjbqcm0A9uHkRj1s9Sv73C5huQfA8lHlvvU0XibXfGtaIzSowi5+oau
TLoUB5OJ6MVOjOTWS33jZw57lsypz492o9moGsAzwrkCUPcSf4v1fp1I9wrFnttclwMma7JIm4nD
ICDSL+1L7yayMvQ3npRC3cf5UQLBih0Hnl/118H+yjIhe3d/9P3aeFcIYAWIAFbK6SWqQ86/+e8c
/VOS05BhzwqNUO+VuMbTgedYdsFOK6qaIHH4MzoxY2bQ2BHICgYcBD7rZYqhyEqLNv5MfElHKlCd
cNbb/a2wVsNK/ERVV7ecDdNpisNS5xDPdO8XEpy7GR1wreDmzKr7V5IJuxYAnNr363326ITNx4Vr
2x+RQ5emYGtu2t8wiBOjAsy00APZkKVKMOUHuabH/3KcRl8TvDHb25wydSF1ULykeD2y7ElD0cT0
7M7awFidkkjoJJ0Ehy8HIWZJvXE9lrnPu5YA7esoLkZAisjKY2vFnp4gAiFt3dz3+PeaHrZQaum0
foSCuDCfPc0RweS5D+FsxNwB/BEcWljdPQwKPRUINAiCE0UdvFStw4Tnb+WXOWG7g1Pquc6KmXLK
WYhrPugoXVo1KJjqwi16f5rUS1co6Enj+khIA3BKDNxavdoxA9anV7FeMXA8Y+ohqn2EXfHlz5px
FHMHvyeTherT3S3mPirFfH0fhrW/QlZxhqgz1r1yQ40NKB8dEiEDxwyNMu+QBCBzsGsxwB5M3hdE
FKp/pc5IZx0ilu9dEHEfWQz6CwcSczO1WAaDMiO8/qbQ2Bqvdp/xVLpRmypfV4zdEXi8bYv9U9E2
8gHufCsASwvqlQt8NkzZBdCgC7EQE/MQWfEhIrn1RQQGp/1NnhIxefgNxfe7u4J/qVdnLaGO6Aph
I2mdl1vSmP483FoMIBAoNgwRwL2tfw43jf7mQ6BSp5UG5WBGKnkiE5ceD1EsDsPy7iTagxZ6/EyL
xK8KongBxFsPAL8B7pAAUqGUchFClsbZJOS+ph6Dp5IX6fEe04+zpHdQkTpTr+8bn/hQ45ouudg5
OC+GhpMDXfo+uR8Svi4KQqaiNJQZCM2wIDZyrjVs4ezk/JyDUMF+bKO/RJ/h9lB0pBR1GmfaUQvK
ZKh1RKqGWdzOsX1arPTxXqqhCRhCuCvv/KbaHByUt66AVGV38TbpgJOqkIDxM5mM+XEFom19zeJq
IF/USVAVUgfjEN9ZHe9Ou0SlhD7xWCor8RpdrXVvPH8y1Z0jQ84BC9h+K2E4RF6dvsSueUH2WEuT
CmxbgU/Y029PnF3EbeJefuR2lNdKDFCaM3MDnLHaQL9KZ8NQyPEPlk/wqBOrTAt2+jq2wLcAmDGa
GSDBZwVA1p/0QGJr0u9SCbXkdbTCE4ihG54aaKAvC/j01X2AiWHasm6yxXlHLwxTit7ZNHNpLeGm
/8ze1ED6yOdFEOn1+6nKRqckMBUM95EsOoIsOIpJuLWXnsBtnzGkgaHZORyFzfJiMxHdpuUpQqDM
HDZaCihXvkx4ZBL08FuTGXoFRzzBpKVARY60/UVZShpOi5dPPXKZSuWjp06QlztJ5h8MKHMjxT2S
Zhqo1lAN/xB11m/nE6omLiceQdk9hqVfpj5MvVXDZgpLZcIfqxcjluM+iwjcv5Z6GO8JbntV3OTT
n201uLidVT6QvHpOtY2qfxNQyp9vgk/Of9jQIfEQA5/8Zmuapubcc/TN+5QFD9x8UY9g/lSmkY47
WObRcAW6qogH3kWe9dkO0JiLWbBCrGmaXPy3BvGKzyOVrnpFZO8ZZpBobOwMz+/kei2skJ1viMRp
7iaQ+CGxHN/K4qNnsfElQOfXV5NbeNsMmWK9UsflfyM+bIykEx6mGE9S6gQO8NwKn2SElm/FeGYi
dn68ovRZmeKv8XAOo4jTOxXTboPvTUi/PbU/s3l8klkVAAzrdw5wIFOY8KC5c+levTrYBN2s0lDX
DioUTFeM/S66ch6T9aJ64U+lH4GS1VrLH1dIbbF0NHXcONCVsKrJg9XpwS8MwbJJURo08z7Mv+lS
nVg9r+l06Ip86N9hUvr5WEPfhFfzJufnIwcJdmMkcH8z8OEFbQEct3Fy0BoumnQGvnFzTdLOhESf
Qs5YuDjhOTF9L+SX4za2zZythxYQWeMmSFEweFW2o+YhH61XsdD/MkKopM6aQ9hs1xN9f2iCDurg
W+w08VIFOhDlLscYPRSmLZwK7m3cad60NuY1+1zhixKinxC5GL1HfAKNeD639jsUzb3rvh0pmPeY
12p2eFyBuDIkMgvgCujERzG1nWJIDanEO7ROw40lld0RORC2jTDOCRyaE/M5dRoeqK5UWJXMmkDl
X6vwmWnbpVOduGbB3xpocboFs+QntSP8axau/8mkqiqZwlMxupeGe0dXBWCF+up/cTxJNTgA3ViA
YKkB04M11Sr/wyO2ezF+/oUBSGqa6otXoTresDKoPiYfduoChTN1tKwIlQydlepJfIzVXH0DLyMk
rV5eslLhijwggykQ7cIZwad1lGWwvOaphqPPENgxqnbIkpvm5TkNDtMWLn9W1XHmbXNHTo5dAg3g
ZKO1SYtC8fJU7u+z6ekgrhfTIcVpBHs6YZW+pe+yUSHuT5jI4jD/+uZXmVsD5sVSrQr6CFj0ZkcX
6dWImQ4j/owjFDRH+od5ZQrjcAdalOyL8rnqFBZrGbrjei1pWFCmpvHZqvDlu1UqU6xFcEAqHeVv
TIGhMKljCWSwRUK77T1i6jcv4DdPkeaFe9FGUFZbqfhFughHNPpVKUoJlDYFhE6gyCwqUgW6iwEb
+qiBnEzR+8iFfpqQsyVT9S3duyQ6v4OIAXiShPJOk/NKuKuaDhBkq0VPf6OfelViQyszjwCQby2Q
XfqTny2N/SMk2vE+vRUNOCXg/WJssgTZ2WpPDjuW1jKGXq/gryBR/01Chbtp/rs0VIrEK4809G44
yOw19r4Tj2Quy77uwAZluRrRkFExxbn6F1ENd2LBoQV5v09BH/E8bvLm3Q//uZr0ncsfltwjdOk+
d+aRbc66UfvQ99AoivSbjKClOSqce0VeWlWWePOSYTRTLGdB5SlLqA/aiUPvPt+8a9SyF9wXbrYg
0R3wnvH2who538yuK8cmYHujGftQd/hGehLjApHX9m9FO1PMCsAdebgfxJhkoBYhZfZ934PON1pC
ClJ+J+HS1Yz0j0QvrjrIEVCNXNCguAVnvQDcGvCuQYPaKp5FM4r16TLNtUdD4izG4vJ3KcxlKK4N
KMYFhThaC0/5bLrCLtoDXW2oiKde+G8IcVycdw8e7NJyxClZhbSuthuKnnrRXZ7bndogCfIDzKR8
DR+j4zzs4G3i5cdXtUL7+dKVXTFJFJKb6oBjEAMcev3TuZU7op/t2tgebGBpRsF3rChLoeFY26lG
PA7gP/cgK5Itesjsqh2ewrieAZSG6M20SckwVOk1OlhsA/vJwe3tQ+1lpcHI3UWwxV7VHIcf8t7R
FCTyfhUSX6nVN9aFcdSWrGWTXXUM1WwPneU5x1C0q4F7QFI3f53n6O216aQLZfmjswq1+mNIgxOp
ujBOEjt7oixcomAn1orAknLBD55GrQ7Pr1BLyCDTE/vMuuUgKUMcdJUe6jNTyT7pGy4d075wR6Hu
OUlgEBAT6O/fzBz4lkWLX6gur7dtGLywMau5gtwQ6OQ8aBw0FLm6orc+ZkpjTe51/Q441/iOcKsw
XbCRbI1vZep3DpBFQ4pjowTcp3g1JpIbTqecpESfX4nIaP/EqzKJuPhRA+0LTfGMO4xmIDiC2Y9M
fgx1zH+ELZLeY7ivJwRMbyPc41kUul9F4xS1MsUQ3YEMOwVEZ7Nf9ZPD5Mt86S28e4s1GD4eowJA
BWsBvtZZgq5RRapJT//81PIm2SW92lAEVEaDo7DfqR4SAdytiKRnQgh1WcOO7DUfLi+mWzStt4GP
3dWMgc5CR772k9TunS4RC2mrRMxWkrqdvtVVnMSWl3nenXkw3zbGi2OGc9qJ0xgta5BDkETQMM0B
75LKUZNG+6/vBEHvCfym1y4/J3pVSj9EAooxGTboB+RaPB/UrWnFrfimDRFF+YRe6i7YhCL77jg8
+qLJF1fFQvljDZM4Nm1oHzZ40m3YZp3117rn1fyn84M43XE/xOW3nOjxu2rnd0vnUdmZ4wPg0CBt
+m/MMLWBzDtHiNhScEjHi//A0zSTXROifwd+ekmqO+cCOjierYFds89XAm1iHtuFm50CwZ8GO2iG
rSE0DCTm/hZT2hW1MFKim0Xj6tFcg4nTrjXg+VE0j+nQJx55P+bD00Ummy1tKiLv+Nrd2JWUltM0
CTGIZLE2+MpBb0zY5Xaw/s1qeP3/2+HJxhUMRwqkVOP2SuXgkva/OXuYNd3fNjK2fgO3r9MrQTo5
6BnCqmgQ9FbF+mbrwN7XO/5upzmepBSUdnwzMqtLxzfxCSJmq9axoDULOd7YNTSo5UW/zeNYUe7X
Rq70x+YeLVXLU5N0V+eQvETwlFKWprB2yHoGT8naUIp9aqa2hNuX6sQlLU10qPzNl4pLh9MvT0++
isB+yDNAlSNalbveiLkOFcMObkplcc2rhtspN1ZzciUWznQF5lpoLLSfD50sai9cKBnGI4TcsXJT
4VHcEtQOQyggWES4H/oODP8c0ARPwDWHFk2KtvugZWxLRTiiur0Xv6VBEgkQGJhmc8OXUygh5VkZ
QxzgLvqJZzIDJxQRRQoJjNav9S5aAs5Zfsc/s77OJEAGvBLbQ9ZZrZY0zl4mJbNkGsBvNT3zorKy
OxNtIh/eCexoS9hZPBjk+BiihEWpRV/JSB59WAgFqp2crODlQS0/i0qf2W9bBW5JYXp8tuKU80eD
Zw0zP76WTKYFt8F4YLtvmW66Qgs9cUiKKSOoJk5Rc2JK6GdKm7+ijmQnpuXatv8udGvZ7ocy2IZV
rZxgTKdI1gWt1FMMtd9QU0v17S5ztmBVr4hG2Jr7BPw+hbeEKBKmAJU0T8HTqnsR/P/IaDxXIjJM
4IlLqoFlUS/p4U7/MvgVXYeO9iljGNVq/c5qMoISnWcaPZPMwy03zVsPMeWdBzDiWQjR5qud7DdK
8NOADzqUTl8KKjTl8UgnLuEV0eD8J03YLCvSfafzzZA/DCbh7ERewOhXm79pFGNkwqjAfNaT0JL6
0AASdKypQLSsuoCZNEymnJskIFu4Awxj/makJDXR3fW5OBDxPpRizQcGP/PbWAaCOzK8rJYkPNkA
QdUhVPTmeaCuTpwadWQ/rqRkQmGjkopMPpXrpoRSmRIgkV20Kwm+mEHM4wpt55TAawsMak4xXyJg
QxGYvLmz1bvky9cWiEhsu/zsM0WRnEc/lLYz9dh2M/y2kojwFVfkMH6O+Llp2+yJFHhi94UxYC5/
wVnY6JvOaX3zzzGvGsmWsjptOMH3h4X84b07O6EebaNr1NhWReqv1c1TytFr9d/71mLF/+DKyBKF
XHXM8qUUFt77/YeoRE+uSYC+swWwSYhO1whHfD/HbYNxelfIqiV5n5loR0Q45YxfTQTzi4hN1zvh
iOEqOo7jm3PYQtADSfIt3bhE9arQUshWmVUaQSwDzEDA39s615LxPG3tPmrkkZTnrqriZtFZaghR
MFkh52e6Ff6phFJ3fOUQYNrQphz7yhWrc0J/IIHEOFsKPSmiroX78YzyuQ0gVGlXqhdCLdhVwhpz
A5bD+rW+ZjZxaKjIWbrODDofY/oKJWhqnQci/u2DXkcxhbee0jflpEfA6u76Wih5slVLyb1wzHf2
cYpC4s/J/fp7Oq+JZQ6QAgK+fyvzhVJW9dX+I3KJD3as5To09syAyHyueHzKLCgrHJ2C3dAp1E+u
0JEa9uiHN6xPgUGbNui8vk7UWnukuZ5JJKYJxvRotgYXb/4z/JcIVS4W9blsKOQOhkHBtu1bvai8
szPki/OGseJkAC7+W7PgCm9RiIPKaRBoVJ7OUbjeUHu7M5Tm17sWDQvR5Zynu0NLlMPEr33BegQT
O/smsfw/2m1gjFLimmzVsi6mtDqKhYU2UWVH0yktSz0Mf0tXTsoW1lZVTxekJo2Ya9ioMQavz844
jTeBiThe33HmXTp13lsiM4g0F/0PLg2MVWzqHLPPM1EYBRl7UQ75VKsnxM7tkZ+LpYz8jdjnuyX+
evSJ1w3pdTRr8iuYRPkIwMBA1iZY/kEJU26TqBpiJC/bszzhrJPQv1rVxRxBMZnjzOlUo6bYBdzZ
m/UgMDcC5dJ7JhhtF8tav1YLAwFXahz3wMaxP2CCWakQFNpenWGrLN1zCUJemY3CAFGIUdXHir8e
CKfVvpWKigllQABC4As4SVdKnjvMQ5bl5SSM7ULrwetJpSwFloeCmIPx7AdHjiY6maZh0qpDX8IK
Y3F9YPE6vRfDXAlWTpuCj46L/q7F3sGBEI6LkDCzh+Yv/yYQkDViiXqCPZu19dOCzBNpMiMJ6HTF
2LyxCqTsotYHHiA7gccD2l3Q6aa6PdZzvGx8flihFTmVrE/VOPjYASY1bYlCl+tH+W516LNu0N2t
LY172JdIxRw2ioVEBv8dEceiEzsSMBPrOkHWPws4gQtdJRA5Kvo+cBBUlw+SlfHo30aBVlSre0Dc
1+tBjnuKRDTvYxoBUXGeyoyhshoZG0/aEmjnZiU6TNPSeEqUukLtCtTupa6sUMcOqCOoeFAfhZDe
mmP2z5I+2n8W6ED3nGyL3wwCCQUxGAeHbaMTbBmSEEjlJGZc+xGonhERWR4JIsyJVWw88qHUFxMp
HNXPr/w1uCnFT5gXMlCoew6pYOTFqw4KTdwez+Hu37auuk+Ps1kZwDO2qyE70qSL1MCm76hdCZ0w
Xn6jndymjOeYb2f4vxaXstV7Pl6hlycTROfFMbS8BajUHrWfTj+VpYEmAAdCImSDzXW4JdMo5/Qh
K33fzZHdgV+oeXPQdoMU7h2ynQMi1dXFNiGJc6H9/TOyBi/sIZXPIo8lo32E7z/B3EOPPXg+GjDf
qqGxAMy9OMuCDB+Sefozn0acNjIqNkB219fLPc8A0nbgfC++u0MLxhY2lqRYp9lr4F1/c+2PONOk
+sYPV8sQGE5S2u4d00gNf1izJOOoezxg2f3u5wLLiBG/M+tUZMck6GsS9SVDqe8FsOKTTywFoCI7
47lbT0fIvKuGSHD/VmQLRwkZ+LWaTQOcCxmFjuKau3osWF3gR2FDVWkAANWVSXn5f8ev1CcupB0v
fAjWUdztK/x2e24nsvsbZAATSqU/Q5yEKzbtOHVEZaNPZdyJlCJJrfCNrRvG75e5NDkontojXv6B
eJPDiYpw4dReQLhKWOZTqyTeUG7Rm+lEo4iM4C6n3uGykynjDU28bBnXgW1Tz/aK3PeLkIkr37mQ
UcTZNxP5/1nusxDtI8cBU8DTy1DK1aD1uMV9gUjm05OJWUQ5cWOqKUwV0WQZFWWi48YQeiCDbxr/
Ir4nXTqnWAxh2rVi76Tyj9EUqn2b5MLMNefC9xhmZNVqGmX5Kgo7qdh8C5WKMxVjzD1/5r7H3TH/
06TNLVvfDGGBiPZP8yg7tXCIoF7ervoiChj6YOBrzMZ4XkFvdA5I+MlUQ0D8+w+r4F66XPQJ5AIA
HfaSfEO88MjwuE9j/PtoLx6IT+KZl6LvUzcdmpuChU3gu2VdCBPVX4uOtQqgkgFZMYnNkUaLZbVs
7ypQ7uCW45GrhmATQdv5UHZwwZ7gQycSfRKqA4iHCU3nMLk/H7M2iTEDx5SkjvBsaR1iAflsLBn9
/ZPpESVtZo9YWHJCJLU5xAIJ+c/CKCmp3CBOBr+RE+BuPJWkEvpJcI0rmmXIEphYTnAvg0/IC/rv
Sj+f4CjNdj5vzJO3Z9h6PcHoW+CWnHyyMCFT1XZKbDoLLocGK7ys27e0SWNClFcXNfXUvifzNPS4
igbk6YX4N+rFBPvVvicBeGRk4k9RfCXMt9w/Bp6NqvyYgRq/wQDmja3cL/l3FjbgNLAeAJSP7wVd
A2q2Z5XZlsrLSfeMcaLkWSPOSf7o2taE+Pakxp/WvolwH5FPJL5ZE4MpGWjPHFJTTFvFeimNu66h
a7s/8ub7Nn+GRfW5B14q85GwOs2+1sJ+m/PLtjom6RBvnHsvl6/NprobRd0PcWMM0yiU7wh5FHbA
8zu0EXl9mQZLi9n0vSYvJ0BzqeTX73NEwmWWrFstFvOv2T+A2yhSaS9w3eSFhT/n3XHPmypGnmsX
LBoyQjk8OLgCiEoXykm7GR8xMEHEYXmgisYU26BblreSp42G+DjHewE9qWNbd5DbYSkYExasx95Q
0qgbNE05sRLKA+i2OvFoCZwqUM0WQHmhpVJbSYVjBlxjtWbsJXno4XlXhlabr4rvjnih/ckJidWX
Ar+HPlNcjvJv5WNVaC9EHu5Q6r85C76P3Mx5KpvSfBETJO2w8ocLJmBIHmKzL/jsOZ2qo7RCRAYS
SpROna26BS87QLphxVLeR74Kws+Oilnzs2P6NlGOFtpYrZd/K4EHJbIgU3K5YwWwB1Xegk+tMdh8
Vxtp0lAe6HUvuHJwIAlhfHTeQSc/neL01dYj7f1ut12AWqK4yFcPblhZ5++6tCFdt97d4cQ5y+ut
dIPTuBFxlrj7hLWyzbcGttED3ORgVGLKVrqhN6c/srd3D0ieT0s0OwnigF44bIMjHLphmMFiEMuI
HCICjIKrTAjARwtTG809L+G77kSKYshAczbqNbSBGibBqrbvd1RWxsFg9g0oip48bWZZg8qe1oH0
1KTq1oKllLytaLSJSH63bmdUWYm0FfABiQSuJtOI33KdXHrYOx0qanNAPd3x6OyOQcgsgZarKOM+
dtXt7fwPAIOWuiM0D7SbqFSqsHjep7VGVw538EqpklFTlSNH6v5nQQxJz1MFLRDCu9IOTBSQ2KkG
NAr6JZaneNeNpWl+9infNgsb5bxtu/E8waynJqYyawRekQybKJThIZGMZWV8CK+B00k/PSf0OUIG
rz3Qs+h/8mu5w1PdscRUneNerurcn1Uh8H07QfG5jRok6931iASWEJJST2sohhHMmWTNPRurWNoL
PS8EZF+CswW1wF+DAEhysCqItitCLUgfAE8HuLv5M64HkWhzNwU95HCrht8tgnlefdmBLKjFoRO1
+tSZVAzAzAVcGnE8A88gl9Fr37nhTdOYow8dkkh5KmXS/AfZFgKIRt8Hqlg0xLIfgAhkW1Id6jry
8SWZOPd0KzglU+/bLmdqxSgP2f7W3UohkqNepWUl/Q2yjlLRU+dMJ6rMRYXJv/PfDFpD9uIEKFro
WBWkaaOxm+21hdK3B/BK/a0esOhlT9iyJVb8ZmXc9Q2/YNt0a+tJKqdMo7sIRljKFI/yin0YwN+P
sVHS2ng5vOhgWy60gCivu4rakfzPVwWoNmRCdG6PfPVO6FoYXZQPIbFlswHRQ0kKGD7X8zmaf3Ry
PBokFyR+cXRKwYAvTz/ycDOxzh9ZHA1hLtW1ycV+cBtXrnUJPP/airfhnOMzwpbyJI9+jCshNXSO
IqekSbeLgVrC0cTinmlmQKO7MFJP/ZOrMOktmHfFmD544aoN3hUKNAXObJm5gCpEZFCAWpoRQmzP
9tXj8LLkv30UNvaw3QbCfOaWW35DT2O9BU4gNttA7hq3034Ta+oF58djH85B82AlV3AlN/4Hv3DR
bisxmfeIKLahtupyFAItRynaiMkB+9vb42mBfE0oqTigR5pATPGB9Ih17Q12fVstfDPWTQ/UhZzw
dQZ9Vt+doFORebw0+mZtEs87vT6wIj7yBK775jy87Wv/pINXLGBv6vsF+piNwEBMPNxiiG69tl/2
lj/7u24w9PZzSUWiFOCT8M5QSPqObO1SD43MHR8Nn9LLRJUkwhDBo5CyMnzqRcO8LFEtYsPNAKzN
N6gHu4eeWkAx1JQXCRGSlfOGKyvdFbEL4t+YhQs+AEgW8OUCcrV95g/t5bnckahk4iXScLfWfE71
CB4I3hXkcbaOY9Rg0b0n8iH3nQo6XnEFEK30832mqo6Kvko8bZkHP8Osk9wCBNaHltnV4gixup18
QfvrAwjQHhjacDajDmHOV/KO0yQzBGLeOAOWfXP4ukAleD12t0HiIWULodEYoWes5y1R6X3y3c8Z
z/m63rUCmc0GrfhOkFPNZiSXlj9IyBzffRJo7j081Aw/G31MIpxTHYKAVYancFQdDx7xMp39SN8v
QkA9pBSVdbzBa5/mPacwx8DzenJJ6kZuizw2mM3d+vhtcoy+9OCBiBewDvKgIN3upe8qNG3j5UdF
Gncz0B4wdaiiUVCyMa2SB8oEecY8tPtWRNV7yFcY51WBts/YQwM1NjBX6sICZLOw34YcEXhZKX5F
QkKMpF5GrBvnxBsCa+aA5kjFs6mxcxH+owkhrbNI/0m547RJ1Fyjnxrw36RugHJR7cZd3MTXn7ug
gd8DHY180AqjmBKJDKZRXoCq/w3fNFe9vxsqFvwAY92G/6F8DpAc5k4nSvKdTiQXfy/76IlXV2QX
e/ze1PsDsNnsHPGtm1GQRtiUvaKKSFD+Yj9Y7ZTuC2/O/JrCzero2wvBn8UlBTLyN3VQ9nILYgrB
Ebt2Isjg3I1e1ZxloPjazqSP77VsBaSb1EgylBumh+xCM+mIuqlyUeG/p5NLDfiDyIw6UFC+fFy6
0R65gCdVm6q1O5s6prjvg8rZ1e6Sle0Jpj1fEtkZcJj55W75JqWhu4YfLUBapNwYUVwSNNXTC6na
f+wcFkKY/wmYJ5t+MYfpXpAq87AG3zzJ69bSA5PvCM0R17QWicU15ZAPQZmayymzFaieb0oMag57
PAsD3Wy/6qUvlKdFRXnvU6rr2VUNDg8psirgzhagWgNnaNargBbRmHInjLIjZaOFaBjqo7NXEUWl
6f5a4EgtROpEiI1gIZR0oMDMoKnDJWBsXKMoO6cLodht+PMZ5joMDgP795qHAC3F9i4Ce6Hyi9Xv
h/zcvKq/tXmn5d7KQLzbh4ZMzRthN5BytPeKipvIzaP0LcizQHXaSrfQ2IL8O5lxEq7FlwrMRGx/
i6U1Uu8YmS51vt6Vv6EHK5mlLL12k12QeEeESybAWV4Ub3b5YrVn9jZRkiQyz5DLNgbmPM4ciEb7
ii9lj/a+OOdsVSLWyoSwQZlJWvahXKi/CE83PJ3BZCTmspJdsi5Ddh0+sXjKsfzXxxJ26Yt9oD/7
Sdbal7uTsNMqPAJR0zkBwAyjv+MaetYAQya9BXDjfyXLynNHi2u6RHfLafXOPyjcJUMvwP8tQ4yI
AjUcrYWlWr8C8JBjLQ3dIG96jt4l1zm81YOVhQ3gSUS7jmIZ7sHRQr8nOKYh5pKjmzQWubhBRQKf
z136CaCZ2H0kFGmCEWb7iyyV6XniFdAoDsdtd7WGss2OwyycNci1eqAzfIzOSj93xYlcYqAbxXx2
aPREy0qbIcGCVmVdD5m/r035r0hHgKrJsDsnL91xEIGfFMhkni8VeVO1mf1dAs4LmGcVF9/JYv1F
sQWGirljgp48g2/mU6mfidtHjNH/nord5VMWCeaY6qOver5/KKndN7ObCLjimr8XwiCaQ2/HHzS6
GSqzuVdUC1V0islp4SVVw9zGcccGCYAFbrnEe6c0jA/YlK+McPtXUWg8XyQKey3Ml4rvthKIOg/0
w00xqpYgMFLJY1vCFOMJq99EdLwVYsJiXP9pIAWF5AYQ6kd1AgnCwZl/MnS9DEVOLaFLdZJQRbdf
i5eDEVFCsXuMDKp3cTaIpK61yCbd8tdO3jcPSTV/uYsku+yPawtb5qBAGJOT9C2oSRyXQbusbmDx
kXc3EVYyFQsXq1ASb9/8XG3jtM4eIEv9ne+Sul1TyrRBPnp+uYIeJQbQ7X5/+Om7+j1rV3Pijsuv
26fvg+HeKYUDUvxtxx7XIhiUwydteCrMGnOjzkOn1oiv2PxoIfOhfICYfVTTo/dIg1t4w6vN2YSV
KjHLAmxyADHLLP0NIcHpkaGJIdxXOGP2TraEX0/OlmQ2xwC3ImfScehrjdJidN5pExMD2+CZVAWE
Y1YyM05LUhyepEQ7wrj//SCeTb1ohiVI+VCzvgOq5PQLM7Bm6GrmKdGw49p0/RjlSOh8zik3jdyv
uBuFBaPcWSsvWGrPVaLx35R84CdBg+fBZTjn1d9mV4jfAdmAkeZm1pZNTDqsuOoWW68ujsQv1sNP
sS7sEI+yFQvzhbuU5nBjBrvHUNsPnkTa6BMfJ0k1XOo5gKvE5TiOQ9o24JwQnP2trF5/8ZD9ZAQJ
gduopD7koPwbUr98XfPc2l62Y8ri0BPlAcB8Dr3NqUY3pUDgcLekmA/lroWOXnLTId7YIu+lZlr1
G17Dqj1yxnbshkOJLAFslkK6Lv0LKYUt9tlBkSJsJiQpqnTn7g23MHwlkhsBgnfmJWok0XXqaFRF
JjW9jX0QYiqvMz1UXNneqXEdNKohvwbSbm2TUY3q+kpbEuHQ3I7D8patuGDcFfnn8gLPIUz5BIzC
h+aloP/k3MKCVtKvuJUac2leIRCom+hbxJOS0Pvmv6o1udJ6pqie53CWsJcJLWAU2RsApnY/RZVD
1ZTVxnhPB58Wye7b/IJXTgk1AC3EhdAEUmzCLeQM86sFsIjRtNMqX1CUkysd0j5HDPAh0F5UcYDo
N89L0C1TOy84btC8v4Mu6RspdsO9AEIyfVsh9riVfszU0DMZBuNeLZDDtcaepZUGlqi+3yGtKVhz
/lMZn5e5cX3t+UKItug6qlKHVHWZuvcOZrAAgVCBKlb8qoW7TLSHfFrg1rZUBLRa/LzapnactLiC
6JOmrn+dL1kiEJCVT84Pnhu8HoBtNJS8p7V0n+0LEZOSCDsls96ZcpmY+AChq/1yZIVqM+nNfbvT
PktctgY+0YzJhSi1wMtmBJJD0D7BEAVMlGj4Z9dfI6HWlMSx39h9XrzfZzqOXatqOoJjcPyLk7j1
YvKuYH3VrncIqCwZ93kmFBDEy+ASqnFssiRiY78KgslU1UrDTH9m/l4pzWI+/AQ5kyd+T8ukMz9+
IzeZTEcL0jxkmPzb70RyqeAUY6MwgokYhLg4t7B90gCoiYFVttSpP/FxstrsxL41+lMkgXtpi49j
I0HxW0Ff0udovd+O2WdYlB6vYYPpiXOaMnNQsyjeZzWBP1rDlb3xPVHJbo6GHHjXVRrJjvBbN1tx
LxglJcmQvsLAQYCefXlaWegHpwGpxpv4Wlnml26m7pKaXp1DXaF2bO0OiY/74OvOtF28XRivrGuY
wmf9MaHiZq/N8zCiP9+EdEQjCDXdHw/fFbEMuE1fEEu/B6lYRO1yc7XWSQXfJbOCEp3Vxl4hrWQA
THEbkRarxxOl2qf/nZ0g1fQUvrDD8OtvNw1rMzP6nLe/YU96JGKdHRA4ziVx5U07EXjP0RXkEvTt
cXZHz/O5vhHN7Ou1n1fk3a5c6UrehHvpDC43IelDHQUtXq+nioO6bgS1agyL3Au0BRaqCcWGR3TJ
7vQdqKSGMVEazvhHm7E5bb6hwgnEkFdkFa3zt+7SrwCrMMoKNmybnOXSMlbSLnijpfw60eS/K/E6
JudtsHuO3ibBiEcwzeiPCS09mP+LgAxjvoTnVGBXLRA2PttG9+OWXyO0TWZi0HJVH2V3zrAMMEzT
KzKYfBlITw0y8J8JQnnx5ADsl6pLPx89GDz07vKcuOtsaTbYCfGm/5txmUhstJ/Y+0xOGNdJfbCL
tFMjjmsIM27eoPHuw6sLDK4XQ08Lz0haxmPdYITKH1YLWxRBeDSeUUYnub1HLzYEzNBe4gXNOLCU
M+Ygxqz15/x1Df1McPVCmGk4v1C2/MH/aaX2lXzpWM7ILnlZul0I2yVLsHkTA0wHEFyBwo2X9Y8z
jT0A4WUmjTLMKKgSACZToKC8BtpVr6kbIyE7v8VboAvYgk5M33iA0JgS7vUVOm/rA13hvvzZx/1H
HwrNELvFxfMRrM+x9eq5TdfWaZ5MxXkNYt/KZwyvyTRk1XuoBWFMoJ4g3drycV32aWqIv0i2DkmC
AhpyOAglAomzPXcu+MefFNOqD3RI0pjYWyJ1t5wC3d4QKFs9wc6c+mD+NOg+L8Inud++526kbPpp
By1dXLBy/axy3bFJtlatPfI8fCA75fTiY8USdyF8VXRq0w3h4xCqZaUff+g0c3ZskLlCuJLoNcJ1
WggDkJ0nlrTvKGXi4+Cs1uJiFqq6EfJ8ygmH2tr0+hYEtcPqC1HQFmE6+qzQ0bIJkvo5ZX00UIH+
5jmYu6z41rBqIlZQXTQDmCT6SAsS6jR3zVfoEPRyWPgFWiWDEWgDzamYAVZEH/co3WwagZbNB1gE
VrxG+rmnky5BPZkuV//+Hxyva7BXEmTasKS8oPeeXoYLWw5wWMcB7ILNCK5iIVgAM1GVTMkO/Kaj
wvfQdEyzTg7AI0c/0LNEkJCFI9vOSK6p+YMGdoTDPL25bCNgLFES3H3mcWO6wm6iNMzMNLYtCLcd
piAKnbmoRY0PlXpAcYRZu33kwL/YVqjhngVZZQCPb5VeGmW+5x6ZAJ+bxnRyBd5ykyTaFhkDXnmB
dHSlzG9TQ9bVnmZHiMlOqqczKWXw9gZ6gyDOBT5INHXlNHPch/hmFKg5qbEPSVsofQh7Fsnfyqzk
wuiRSJjiVMJSTtO++tTNoZL6Oi0SfmpCNjGezEPVIr/l+IhZguKQTPgH0mrxpi7nYAzfnHnfbVWB
G2znQ8A0hXwNXu9wrQWH3VzMyj6Movz5gDa+aUZ6qMKFcSIX42o9qH7u21VNpHx1yluVITjCucNO
J83pshYNxg+DSKgKp1FKcfSXa8/Y1m27IEa304EHqxKQC8bcofpo+68I8X7o42En7kgiKVzJlGwO
jvppt/w3D/og8ob9n2dJDDquX5XsVORos1JHCpPLneD2Z+NAJ4j7pfuzC5KyuvNGvP1jWjhx/mKg
/cszdLfzSNITbxlbg/PFp1wwnLLVyoR/jeY/3hKNlUTVpgt1IxTIqYEDTVscbDsmtZb24NWUwGXd
skcrGrU8QR6+ht5KPGJSP93tiy/QqoBemMFQVmKQgY+M/mu9d/HqDSWbifG5oiiRZO2DueB9yut+
0x8ApTw9n/THhXwszbIYLhYNE7cqNELhDGb5AuulJ1gFX/BvKegvzEfmgVM0rWkyOYdbqT1lZGry
hsCeV68RXmbEC/yytWoCLWJViqyeF8oyZunawBztke7o9h4gtPf63nzR5Z6f+hXh1r9aCS1EsSXy
5eVjJsJ5pJ5XOSPoopVEYbp0s+N+b0/X4i/ZLLCoc9qYB6TrzPZq1VsQkYfLMaO8KmdK/snz8eWC
k9rY/qW/jdWQXCDwxQ2wGTQG3SzKZXKZ45A0GIBCXVRO7x4iWBTSvKlUSoTvER2ul3KvMy4t1fhb
P372JCABWT3vRG1qiH/5c8YgmZ/rlVVzXK7Vqhr8fSXSCvtoNGGJWrNQInDVZRTpV2fS/o9b7Iyv
u819YTbYVuHU1cyZTMbWXwwreBG2/VG7m7l4mwkDvXOWSjK1Jb3gBcxwCgUsEEJFPTjdqTgDpbKM
LqBDxqjlgaGzJcCFeIrZ/XsRd4GfqCSQLJJrcFPaEAIknp0bTCIVtQ2iQ1KFE4zEb2FWgUXlIjJ7
Wq1zQzZYDrXo32AVoy8IUtt6L0Uro+cHipgNJkWtIlNLRUAUXZLFVJwt3+eXmyEVsRyO0sVH8qR3
fJo8ypmX0KrR6NWECOy/jvEFE453sPKGUyvp/Cf4UqMBMjBVJw8USlHiiktezXt23GzBeTkhv0gp
L8He3lzBK84pK15am7GHbVs/rlldNFjgnF+MYMnTBtMKequa7EBaQSZbu/Ai5EKNKhyoWOVvw+Sm
Fxew2tjytGSXtch/lMF0yEzl9KWdMgx2SP3h2INTlgmKghrDVMQbYuR4lnnz4ZuEn6nUwFwFNmgw
l4X92oYcoGTSKtT9uNsI/A6OZEJSNnA3GdQ051Pie8F4m91+TUb815GpqCpxJ3fa7leYO6GZqfJV
LYUgQ2nNIf3U/vXHyjCGxtb/RcoltqjcO6+FgKqqHX7xqh3q7QCjqGDYnxnr7h9mR3FqZ4tI+UsV
EQDlIPLEp6zyix+CVC/eU4BZZsKU+kGoD98Utau/T/bBP/fNT26k+iAZD7k5nlb7NOtRVnxnTuzt
k546z9swrENaj0q5nI06eMcmRpD0Jrhpl6OsBZdHPMJ7IGjw3Zv6FJuxdhfabMU2wxqipff3jot4
LpTt4Z2yLHKySERTl6JahPdvZFvOMs3iNmuuR3J3NQW8ofZvdEwAPc/12lHwb9TXoedVpx9IwTQw
mKe0gUXlf9k9DCLbGGarjGKYeeFS9Xq1zop1ckxMkhqjCkJTpeeMbL4f2EzC7wwiLIixd4Wulxmq
axhE1Rd/i7ee9Zcn9G15IghbwI9gNThiSU1DogXiudJiN6PPZyQgNmIqvxD6SZ0AL3y9to1alZ48
Kt9uHt7gA/OfudPE6yHGqSA+J5N1x5DTvHN4qeVD3PxiynCxf6D44eSptueHu7S6qbPRDS8QyYNO
pDnNuRFb7if2CCnYGsSyMDJo12pwQPISjC/kOhhNYDNgnJ1DVsfmW8U1RgVqjl2QlJFLXubck+p5
jpoeEe8OaVdCmoE9vyYRAA2uJJsBYsjoObXqRxUHurBhEbtiuqMDdDl5uocA/315aVcxnIVXvdG3
7cJEWIZDIOUmv5PsCUhOJ/viOiRSY2fO3vLnft7jLpMlKBRvBAZuqRUEXYbMSLkImALytra7RScJ
NerNzBo60nYbHV5V9m2A0lBswILIb6yZtnyvEjXeYnsudfwhzlqedcz6Akq9++v9h/qjcJFkENQg
cISIRB0NK+zpjMcRwlDIusfAUVt91TH/BFr4QNSPrADroKdmA7zsqOccYuEnPL+JCi9HM+vChmhH
gBEGGVmN5nWpefWs8bNQupcGrRx8qb7oYXc6vzjW5d60vTDuV8XBB89MoBb14MGFNV8rcn9rkXEx
IAyWIDSRzZWYZ49Ro/kfbCF2nkFl09iZG7Jm5bm+FpCpIIo2Yyb/qRu5ERYB+TaJ5CkS5iawf58t
Ne7iwLHaVs93cIkzD3nbV5Iy4Z7R38Wzk9ud7WWC08z+1EXfTaViukHjmEDacUBnQ1xWQiuv/kVz
JWPaL/eW7YXE5UHhf++rP3tH1W8CZR6htmTFAQsy0yzlE8a35uvjYgeK8n4GkHjmsKbAvBvnQE1K
4urSv0mAsud2h3KDn07YtmVJRvCLwlITZYOUEMkA+LlwQRTZyaztdskbNYaZlceEvkKbG6O/m/uv
8El5EYG2jfbpLWeHSMc1NjHiI96J829krpeNJL6EYyPm7fSTLGopBr66aaT/9qyGNslL8l/FHouC
sULP7DT6lZ5gU6KMBsENLKxBDPserVEPN0xYzvkCdGIuAgHHGTiG7X+7byUteG39GqyjdUZ6p9fP
NS+Ha1awEkr+dDv8Gqw6z11A0tJkJxYrL63w78+b6MoTu0OpJ3IQFewSv/oovAU9k+GL32dKuX0K
7Q6hFXw4+hXtrf46IawtjHDc/Zj+3EcSpjQ7NR6e53HDUrL/DLnI4lHlzocpd2IqrJLaT0Lyjp7G
a+/JKs9733yzzxAJhmJx4aJ4HO3rRWYB8JnGaZIbkIpWLgjsBDml06hVJoP870Eb8PzemVO73GJX
0QaVheMi1CCK4pq8i3DUKNHT/BVc9AFArPgehKrJyXSYhJN3ULHx6BMYLncZCtGock3JWrJNik0W
IvXr5w5P+/vl1Edp0o97WgrUpYi6VQ6tA3TVxwCoSrJoD+I/yuXdDkY+IrQzKRtwNW8VWzsBAuRL
oQqZex1mvgn8Kn8Ue8TQC5nYshjcx+jyB9rVWCLdrP93s6X+vzDP3GYUL4x1odGxcP2DhvwD/yFO
9qeWVLE/dyENpsccwQoupmkc9n7C2QeRiS34IrTGPTvpD3LVA77pjsttW0+jpJIQiwG4FeK4s+LQ
ftRTfu0kJCZ5QW2kpm04/Xank0hz/5b2gUK1b51Mkh4KRWeMq4GGJOq9m3U+x0U/Udf1ThqPI65m
rf0qG8pz8ORB3B4pispixQy/W3HSTkHTDbwHoNw7KQ1GE5mzoKc8EIP+PVMyvrQT+Ugg0LaiVAyb
+hE9PLirQtcPGDo4k5IVvwEvalQkrYd9o4XJ7EL1lq02192+n13/bgwjkb1fdJorQZDewi26AdH8
IhkNGiVN+hLNrBRM/7ucRJ/O4Fr51CNVeDMGYU9LkiHhftNwUt3Rfe5L3f3nB0I4RZdZ6Klflh98
JRBlEhk+IN35Qqjx3Rzmxd4fE6TwXFjePEpYHZ3YCG3GJSwejy8uozniMP5fosJ+/xW4ICiNATeQ
U4RtnaFqy2GQgMV/z9AEOVuTQ0td129vjvH/AFf9USzixzXzF7/zcYSu1Z9kBV0DFTazbHV2J++E
pSEneSwtOxUXXW2Q0yNDVrO9c7mrK125UVsdxqYnvoN5Ca3p6CxmQRgkDVWUkVL3WT6WnUHNniby
vfhAxlcjhr7e3ip47CBG8MyjwaJ9DUTZXaeD8N6lw2k++r6Bb76vxzTYZz1GKPN+JieeJi1wzCrE
3Wf6Q+htzQk6q4SBbTwl1j4gWeO/slAM7E05O/XoN6qQBP2Zdf60t5BYxuRybO+9CMiNkpS9Skmw
H/sR/vq9v/GzgSMDpiM5JrDTwGizaYVd6xToYzeGS23G6xcB2XLx5nkq+HTLfEu8x0l7WTcWfrvf
PgLr3ykW4m4LCaQ6SgFyxNrM0FU7BXk5oJYdtBkaNAcmCQ5ep+iR+4uNFZgBF+vY7JcV4gB6ig7N
G9Z2sYMc/IZwvAImoGN720Vy/LRP6pIz3LVOProqTv71DXd9Dzi2M51BeJq4+JJtGXTjAgVaAofU
cfq3jUwtOqhkbYxs91dUkJeKassPD05p84mW1tikttgpm2SHsE7MhHI+8HU3UDJqRl2CuqEFVxh1
irWydO/yQ40QUnptsvxiuhTa8g371uRsdTD0cZ8958muba949adRRb+1pA3OcePmP4CkyfDYHRCf
5OtrEi4JfR2ubypJ210ROuyH4aC33O/moWcU42/s/t6Kdljqr42Pij+tgATtzrERqbjrwNwVX+JO
X44c76bGgrZXtS20V1OhOVjp/TSRSHaoTA99xJz+qW0HfLQueCg4wjmx9bsucAwD4R+ZW0z0UjG6
R8SfkXkW/XFcD/NjlsU5D4C1Gsk+pcOsugW9n9QqU2hGi6beRlPxzyAjZ9nfDKPTYDe1iPxGks5q
c3Q0Y/8zwK7EgE5rTDMwTpF1mB1RE8wFR+1wecWJnVej2DZmVKCgVUis7kFLD3H43iGDi4p1kji1
7cGvNtq/B5Htt+Y1g2QL9RQsWBSPJEhl9ODYVkXdytzOWiIdfSD8IWYB6AEWRX/dxtyvARdcvm5f
OXLgsuL1U2QHyETcUawOGSF8FlFR5MHGS1A6OaB0UjguKbLa/7/AWsKsqB01ROyIOp3m0PJOAQVV
lg5lGRBYbmFb9W6IzteKrKLjGX871uu3QtQKVcICFIhmHtGen7FVCXC31mEb/4oUHbZY5oIJM8Zu
1LWETmrwLfR64/WBYZzj8kId6SHCv43v63L751Dow8Dv3CLQ0PZUz/uDasd7sr2OUVkPFJgV2C7g
mI3kM46fP3jbdN9iSdtKOOj2LOH0X/qIa4i75c9gm1DG4SswrJtSy/1z0NlVA/ZrJHnqtPTBhNkZ
pv0Ek/X8yC92S92mnsAFslusVrYovH6LvteTMRVRjaKOv/VmcNLQKeCh2CseF6yS0yNWADWXKHRH
uZ4GcGJIkLcRdDhUjcBkUvX7lrZg4e9QjMMap3L7omf6Alqkf343muNdvUnnv6o7Irbs4WIJtVTX
um3u4M001J/zVCDQ4GfZfM8MD7+prm0xFa7NBgJ0Dzu1Iy+IDLlOKXWdRjkikB64DHPfAMAQ1nCW
Pnpr4aieCOHMcd0sog0F/cZ7eLabeJ5uxe0jKYoeUPLrfMJMoMYAe27JyKBz7TPYq0R85d050ZM0
Oia143CW97sksSU9+oRzGZL13wdIHEVCeXvH6AIAjnFzXzw2r1WrTHdJNHAKTlF8hFTIvt/qp4/n
ZX9W72yY1vBsS6du0srWIAmhg5Gu1KPrpk83PK0bTIlKywfBzPDiDWSqgruw/5CsNCZk9oVUdI5T
UgCuC4IQ8nUV8rzl9TYYjJfwyMaQDA3oVfXUpQCTPIKysaMhSz5uaTXKozEIzvFqa3SVt4bAp3OQ
sNIuL4rVdKqw1dy63DE7YVk59WKxc3gm0adQmVhcVk+X7O2YisPP49Poxo9CSttLW7289qXf8zlr
SvBnoA9JubNTd3vIlYuN7OYlGj0mW/vRwzaxrv14NtJuHBcPdNMOwlHnjT3F0/+OkDyISbK3gFY5
KyQFlL5Uh+xEXwzapFGDRdAebyUP8BAan8ohSyJSxbnG/ZxygDqMmlzDaClOQ7K0P3xyIwPqwyrv
8ZObi05/UKKkWy5C76LZWaafT+vCB3ar9/PoYNxi2jzD4r5j+GPk/+J0oRiIqokJgLS+DaIWF9Yi
ukFuzuW3WmFUZ25Ak7FYYXN+pzGcTwfN+hqQSkNncd3Y2iOC3WYBqGTc7OBQtTrmq9Oatjc6VoRl
ykfIwIwIVRG6bYBVjDenprejeJc2996bpoVLkWRQc4rrUqzmOJwfzYkSbgn5Ei3pZVmLUdRkSs/0
rbjGrtBFvbMIVh9y6AuBukWIO1MQgZ/LDapPBdwyYd/5PL/xBsWNZdRgAN+JC+C0t/YP+Yr7E+/0
wAEyAiyIti4KLwFFC9cSZz4bMCkZAgMhcL5yqD8kfRkLRTfIcrOc8nVIA8Ealc9VDRwkotVsCfD9
NiByIaFPCDhh96c0tli9rP/LDtxu18Xvw6ZMkFzV02boNP/DvuJiAVhZ/dcu5lb/r4XxhtKPTM8T
Jg+kuXJYV5fx2BsZmgTAlBi2EklEXi8kMHq1cf6o3223w96S2Dzl+wQek51Qjl8aoIxIja+Uam57
FE0lZ34NXcDCsdxsWTSxYtFCCk2beitCV954OGBEVqBml1fRYciDuM3XOMNYgohdMvciH/TdPHI+
vxzG/R2KTo6c6W1HciRmmsABO2O/Q4k83R2A7CVYskbY/PFR21u85NZ9q3sCkBYp5NJagfkW6Aaq
5GOtDYnJt7SwjsgJdLZN427Fx0+7Iw5QvzpxkYw+A7zjFcW+dTwqwhwKKDbdB6PWlyvevZ8pLmaR
1t0TlLrzeEEc8Y5yNzf+5UUg+R0H5Ivm5qAxI1TPTGhUO+EotkEOZIMwnykD9PPrSb5o2YFx6Hqr
ovU58PnfOqje3l5jRZaocV6ECoIJNTM97A694bRyh+jQHIXG4dNS7ExiDX87tPDFD8jWdg8oDRQj
j+0bFC+KOYgDLX9yWsl4jdx3eUHMBb3Sl0l0pDm0in9I2o2QvRU4PKkvfr5qHjaEoHhsAJNcp6DU
yNOG9241S62OZYNoGQ5jGH1c4g9tbCvYLaOQMGOiK0fg2OHQAa4FLUiEwuqhYajMRocwta1lVSsv
0v1pFAxr78V0oyZAZrgS1qEGdJ0dxOt90PsrJyP1l48w1lAA+A2dTuWvYhtXlT8okugbbclR8LNc
KzB01Mj8nmh2B15IKMuqICVkNH/elEkn1z80f71Wy36Hq4pPpD1HiiI8ewHulOCLMaIRRHIaD4JT
yKfts5kwBTP69JiIoPlyQhww7DWaUgDZdELhuFM5wLS1WiwxbPMtDbTgfectdy+lZ+8cc/akVksY
HWxDy+CkzxsBwLqjCYMY03JfDFyMQKeMcyDfTgeLgtTjrl2hkhASE+TOG+x0+cYZjoSGpCXBI8Fr
b92iA9ElZ2U+J/CByncQQ32huwnNQWgU+rc4VZhIferRM0DUeRxc9tHxi1QucwVLv9xNfvRy2+vm
v/9Jk7K5yUMPjnae2PeFzVksa4PrmdONltUpd93lMtklMxJtoNYWFUIrGFs2PA7cHApNL1M2Hgxl
cuCOEooHxv7uOP+tnn0a2DOIIeyZd2LtvIo74ajwkTjlWaYlXFCElcN72bBzHxI7dNrR0x3Gabsb
Tt3cP7RHxIDddOtpE1Kj62VWNYsFvDLmO9rs4/R+1CHYIi5ygdXlzLrjKiXQ9GJMrxj2fnPmlJRm
p6mCIRHB2dBe77Y5Y3wCaLPahQCyLgI0o0i8g49b1dYV+6rxfZPSk50pLE3QeE8PVVoczasYr3Ha
7LzL3/k9mHHGGuZTY20jZDtge8oHyro0S1nuLXPnaO9OJO5jXgTj94iJpHl1wFxfK2491hb2DAIM
Uak0x97m5L5Ld2la9tTrFLdrMVQQSo1xR8gxuGKh5f8nqOrUqHiU1qBOgoBLN3BP5CIOTf29Ang8
vuYflj6qJAFNfByWNcsUNCtiqw4mFWcwPlYimcTgKuPBMo+nLFL0V+Ett9A6NB631ChcgHBdXcWI
wHlLHmxrKFHGD2cc3tQf659Dcy4HmHbEvodwSqM78oC8rWDGPfEu+/Zm699lC2qtwz45GnsWWeMm
qpEw9/Qqoq/CAE8K3j20tWk4xjn7AtXR/Sk2J1Hr4+lFk/eUaJ1tPynXoW5s3MMC0AEBb+GRTWgH
kYzctz15JdyICZn5HVzCZpf8nApM+/dCipBZ2VHoQcztz4+a+B2VjdBQgqIXEVJ/jQt3UZmGMgwX
ENKeUBEvgbhamb6B1z19OMI5BNKeTQyGP4xkfbV04KNWaSiP/zlPwg+x5O5ro2o7mxVRVmRe70lm
OwE7QdglV/mtFmSYuUbXqH/Mjq0qttaLtc3EN/bnfTuLZDxvZFysMKTD+VCq1K6J5Hxgo/lpz1J+
Ae179dkd22imhtnjgCjYOnYN+qYvwDjaI3ASJhbQaeuGHEzwNxB73zlgot+6F3+gV4Z8q75IwcWW
GGx7HJ8JiylG96s8RpnqA4OlxqX/5VAvsmwfVVB7Lo5sIFRjdC9TjuROxqg/8mrVKwdAShmAweA4
BU/FxoEAJ2/4z9/PlCK8Ke1dpKBX6pOP54ZAcPkTR5qxETncdtVfo9CPUkgCQV8nbOD2j8Sn8gK0
OspVTEPI8t1yDXAzP5w5J83iYUoDLx8XvZYdMg/tzgoYYAnz9TgJaLwV1i4kBtzMuUXyqv4wD2iC
Frn+GvDsMkmOeW19G37aeK0o9UG/IzJrXP89lyUhuk+VoYdPvO6vaubIxT9EIFZS41KO1reNtXRG
7LNiNt/L/QdjsPe75zvLhWSA0UQxqh0UCTDz67HSPkgpaa5eA42nuPzX5I4BkLDeILi4WbK6bE3x
TMq3We3uDPnBLbFS5BrsHsljBRDIjBLLGMLj3xGPrQAXDKPpGdvJLnqZmU26L6SPLTHgGuFrNFPH
BbhJohXCKIqDqjCuGJZJqRf4eMSjujhrH5W1OqqPcDoxbOStKRSdr9ha8VRCP3vLdoxgZNj2wNIl
HHCbR/6FZijEtsy/1AgIvtddnoxlBX/amtV3ijagd9H1JCrHIcJKV+wC5XgRgZnPyls865hk+yTw
btXrme49GfGyoIZ27gvWAbu/0ZbD5Ry7rRbkcmyf3caJJ3Me5Vd/SUWEVjAde3eUIEIO4y4Igs+V
VgvpXt03hikilyzrr65vG+dEoDR1I7sN4TBInpyllPQvZ86qoletARaZ69JQgt1GfOophS+zsrfO
n2NhbqaQulLMA5Vz5aRpRrdrPJUdCKUfVjrrBgzR5reJbHZxOe96OZ6Ld2SxYuuLKAQmxl5UC8Rt
pv9IgD9civr9as9atf45GNTaprDPd1+AT4MpMgiRm7vILBn1i4e8jF8L0k/LEW3+ZszoH/+gKvTK
jGIUI4nyt3G0i0JrdRe0tTTybdkEZ3Zc3gJ5TUWaEg5RtpjWw+KLk75iNm8Xuai519NlvE/Kbiks
qiaCqxvbS/xmpWM8P6UD11Gy1B9RtLwEowJxJbMm3IqdktqLVwfEquCgHsDiK349TWgK3Xf0+8Bf
jrNGc3lkmPNDOXJmLJ/s2+gEqGpigCuAHbTy/FTdiA4oAO9/2xhFYLYsO1YBYW09lkuDndWrymU/
AXwPig6BT0LQddz2QKbcAnVdpoyXJlk7EqAsDN3VsH+onZ5uTmyBbpRhwBBlc/qU+pkG7Wk0ZiJH
iatVzIQeWEhwEsjKfEaO+H/7u+bHm6nrT2chx9431prIANkXwGhxqzTbW1KMarR8SueaqM2hSFHj
bU+uIHw+0yGmtxT73sJzU4tE1BWDJ1sLnHd6ZuqLFRtuMVxNrDyx2Alhj3HWqPvzrSxVvt0OrZx5
9/1IMD2276jXkmjuZ1/gLRJy7XOENYYqlF59Z2vBxqI13yylgjtLT6x7s6KzSh+ddNCTfOQMFdgS
iWNJ+jKJ+ppYqAM9W9ZQnY68x01/j5xnq6AkvHTd2iukJ5VDAbSxoRoLwz+xe/L9Eoh5fzNSItMa
AsbPMVixs6RyqyE1Rv9qLqYWaTduCl4Bi4JOyzsVWpRJc4KxQVntmZlA1mi8+Xiu6bv2rk0oHvuT
OSyEpsQjCbNwcQ0QKDx98E5ZGf3y3Qr4+0wERyrHsRmBoxvK4Ymia4f8XfgXZJT0M440b8nQm+4A
FahW7w8GiolYArpeo0ERD9tJ3HGZJJqRIXz45Mv2NF2dqqiPCxpT26K7SIkmjvuPzFWc0emlow3T
2PhHUD81WxscinVMUzTkMnhNNiwEHI4g6jFMG2X+GJskBCMVwXOYrJz+AMGF9uAIRmzOFvy1gBHg
yq80geKJh9tZq9nJjquwgMRHXLKEQ7aEWGs9OSwIwt53AWxzWh48QFj4Zjg5u22CrUMYfJtz1cmE
yhBOZ59a2z4s8pF11MJsJKjwziH0+gVt3zVdhAuuuVa/m/UOEawX4i2qzC89ljrby4mTOk7X3hCw
d0XYB22H2K7um2Aqq/vjeTtrzUGVnLppp2WeGcKLuT5kCrsMC2N0lHrBeRCVn6v4/oCSbU8ZTjFq
4q1X17Iqb7mHBkKEabUFPpbKPEBQkcJhBtcHYVATSWjNgDdEYM9jAhrNqUyprOUuRHBxqJtXCXkj
M4h4hJlqFOEV4DZRz2p6lGiAs+/RXni1UVUOrTk3kR6cFb8vx0ZAkvHfjvruVHAFxGO5u6yXhPn1
MTTnFRafhM4ec07maLl8F86EJunYsqE+VIolm6zva6BvU6Lex8nn38fKW1PdYXuXJ/WJREA9MAfY
uXduJOYaVVaCl0SjM5agt47ztUguNpXcjj7ePikD1NR5VXtoGuwujY0BzgEriJEpJ2qPTTavN46c
OhSDkNIJmWNQs7op7+kgLeGWCxnYkW28rZo5f3O+ymite4zu9cXPVN7koTWjV7jpr14lsvJ39PNv
MnJyKOjrEnam0WpA2LK+keaWQjNTOayxbJUbbAjc3gaYFa1s7xJf4nTr+UiCRUHX8eFCrhDMfnIL
PH2c9JOXiWS7c8sK9o7kd7kpCL/Cb/Esl0Itl7dHvGKzMShrgd4H13sLXuVbs7ychGxXHyzD0lDl
JQnUp0gkyo4wTXLCFvgrJGUVfG2kElNkr4GarJfskh/waCS1OTRSu7M2wtoT3dF2vVxup8C5QTos
nSVrI6XMCXPCZzFHbdSjIeFbbSkY88s46ILYWOd/CYd9+syRl9zkPKanI2M0MGz4gwKH6TQXRgjz
kNcct/8HbeIOXJMxQsnqTqfaDVRguNA6MRzXsl0xwns4boyxsSYD/EdXZSBjPk8Bvi/+HUS788rs
O2JcKdjDjheHuXDtQWbMCiAPmK02lZ8ty+HORz6/MfvBkSDd2OPtPGEmfip2/gbKQZ+cPfHYdlfM
DI0aXWcol8v78j5Nhn8UqkcYitJc9R0G7MqWnx3Z0CYyLIf2UPT5+X0ITYnITJz4nhTS09uG6lUT
JotTNzJImKAJvsvI6LHETD6KPrt7Gf7Y5sP32ouTbOgslhBdA6nZaFHpMWaAPkwfKEBD4WAfZF8c
8aLSM0iorSdCK/k3tNdErkzd3b+9VQrmjnlnyp/Dm6Y4pS6FWtvL3XvqxHUz06SsrGSl6Os9RS+n
Sm327SwtxTSkLSIz3G9V3hd4lvN+d8DgbykEPqkfXi/1X5h17VX6UblbRDSZ7lUF4o38Kp5qBEp0
IXxpO+yEzIB2+7122PV2SmDV8m05ZvfW3dxIloahPEq6j3wbOSxP55zQ/t2qjnMHtuE5H2oSx75l
mZ9wXISV7zXRtgWPu5WyyMyM7k3D8Ei6sdKOmTWj90vDlxtdjDbJrrFIq7aQ4eo5RHwhFEMLdQfh
OdvBup8M2LKexWYbu/YXkesLUIxYEB8Y+hNbu8o1RQq+hUI/Q0TDKTYymEA0j6RTQCn79JfLac9e
GL1hm/U/w9VwHzGNwqer4mEyFB3NZKIHvmumfvmYAo6ZYmVkHTaiQaW+l+0hvObdVvFIT/E/wKrK
iiG1Ct4bk7D3vcwpKKF4oEA6yt5ZraaM7jruc1bGQ1AszPABH50GePioP5G/LbWCHloMha7yZDee
cHRaklkvQv1HA1fw2ujeJ6+jMHTCjzRrveMBF3fgrea+TSSgcjkNTnvGFfxjYeNydFzJ6PvJZjfm
Bigx4Jx2tUeiqHYpDnWnfViITK/egZUIB4fFuGSX0D8WTbfFhjWNYbQbhyPQhy47EVJKJIaJMhIh
dNGtMLd0o+fjrWBuaKe0hc1d5F/o2SL9BYlRZR0eOFRbvCrUb3M5kW7s5Fd9IyLEpWOusJil5C9T
LCBlkUTBIyODr/KkkM0o15zcHBZf1oI2KxKfpZXdOMDWaYx0/YCdhL5jP6hp+fd95/8oB+3eLGtS
TiWZ61MCt7ClG3B+KhZUC0X6kBP4xvNQHe/Y7YV2qf5cbb65p8mLmjXKNkSp9GL7hubeYfrnnPAu
L91u4086sZwgMuovy1XvZy1c3/HzIaDbnMYrK96/oy2VQUy/6fIXISf6aMS/Ok6MYpNyJRyCu6oL
mZ/y1JscII+ZBtUQug+g8Neud59Szd2190D6EpVkbjoIDSmHcICgEj0dnid/Wp/Y/gD4bhXRwnQ1
/CM5i1AdB6pHBK7YbrWyzuWDVsJ7Xd4V2d+7FyXle2A5yFUt6jLI/UbmjRlIgwmRz6UcyG/LM/DQ
5h+B+CuGbqNYIZ6Nwvkeka6Nxzr0wv+Qq2QBnXrJqMCCahlTQly5UIEs/Jy146AU0fh32F5Gnov1
XtPaYuhrJo4BnbupznHEa48l6Yu2IX1rtMP/VnTS47S1ILA2O8x6YCg+YgvyW0k4aitOCXMwipqp
m1VEjuyWysTDqp6rcD3KiaMaxSP3P00vuqp6YHIvtgILOV/MoXv2sJsMhFocbv0NMXb4ZsGKVsyG
hvbQFXF14afbk6aP0WZjS1AFaa2ER4dfrR71GmaVLn81mxdug76gHtiwyNtIFtUeiwjxw7jAqOMN
tc7n/evP5K7jezhM0vzJpuNhXXWTdBotIsxfOIWaIXwnKYE/5EW/k/9DrmmVSKUIIIfw8/r31Il0
ow7USPvLWP/xF4K989IdFJhA0xQbaqSUzZdrN+K7MMwhfX6yz6KuXtQCfMvoN1GjksFTgqZKS8ek
mWiw/PWy9+4QuwwEEWnc/2fH0GzIob8fIbzsUmhSaZasU9r++x1FMAcPyHxlG8fB9UV5Cq3FSvnt
remjkKBYclEMpwMAGx1x0YhxU++9uV2oeLy8l204iNY8o9XPDA8xgXOm4tUotdIUJzIly+CMg+6v
wu1thJrbzA8RpSb6Vr4SYRt1cjhQC0WJYHBfhy9dCGsEWwr512zrtKKyIatP8iL3NiQc3V+Nrhpa
pvQWtMvvmpaz/MUQ9bXRx1Gbf66MTcCNN+7cItoPY5wQqmAEevoGxquUJP3g8SbzJeeD2vsr8nVJ
27wRj30il7uKjgAzOrySzpw49cPVcWDZm0/tiFCZcu8khShCaaVNeA6xpPJpfqjljaMNJ9G4lbhd
iXaJvPLh/9w8L95AKN5Qo9vlQafrb3X4hVGV/8rF1UF1dGgVFEPISDFHRtmXMRCJhFFBAreLDpy8
p3kMjgUNkU4yiRt2W5IsA2Q3jvLDPPZvm42PZ4XTJN2xFrEKHC6BH0BVFGrlN5FZvZgGnSNalBWA
dBWRN0A+vbs3WGDDf2S/ya9OptRAVEKbgV8kbkdDBWYQJXRlStiSIponnLw6MeMs1gdTBbu89Dq0
sehflzlyVvElXyH6HIxO+GMyRS+kKs2/opGDK4Ll2mHbnLIdpD9M3mI19sONyxgbURc0r79FGnuS
JLxUeihgodJLJrpXf61I2wn8n5S9FkeTSC0ZxdJhga9cPBaSZguIWYWVkIITOF1E0fMCIZzt53Xv
ZXhXMnX2GmJjZUshatBVHXaMwXc2Xzg/611wmNdITM42xQTGtH/Jmdmp3luIzlZ39sFCechGv4La
Xko7B1G2oC1x7EwSc+a4Q4qTy6bSY/WxObRTAEAsp92nA4TtASYfn/wlDN8XbYCzMlUVMbvZp3Ze
fAd06UJf43pfTiGX37T1D8VHoqKT0/GJ/KdsgU7gaCa5bQlRY1m7nvlDeif8yZI0pxH50XoqfzzZ
j8eqYdPIwcqZlw/3w8zY+a7iUSl/qyZ/ckPtWhuVZb5GsavuGL+7w9SOFVc4zLH6Ast+Du5tmM46
FenZiCCsT+jU0AcbCw8qFMTLjZBkrRNlyaO6xapITxORM/BPa8u6X1ykFt8JRZ3pAxOcgjByC+PG
SQET8nXUVv6zEmLSagHEZqXVo/RkCGvaG5l91g9Emvva7r7pjJGDEBPgJY6Z+u5OY+0+XQa+sPwK
eswh6njH+GHQozgdnEKJbg2ePL/M1ZXEJutLjYBC9sFVyKLJl+Va6fW4pXWHeg7/o+My0bnMk56F
0nbfWnKXmN4Vv6v8iKt6qkVxyHBLwgUvQig+KL/EbyYD/xoSN3GUIN1he6dqklMMk1yfUkVVfyK7
JRtvqbAgHKJfhIZFFTHbNz1Yg0Ji6PyaSm/qXDwP1pJ7dUasDmcHicTDay4E5FTKPBwRTmqLM+kk
CJ5i9wQ9SD9wymNc8jwLGgf2lJ8n71f3gsO8k2ZaL7VuQgwd1nKT5xRNFhcDPR0u4N+v6opzxF0T
GGZAUoP/8ANPMC154TZysZEWFG315n/1YWH2oD1fhLgAdKy2t8eVyuX+/xv6e12rG/IT9x/yV4qk
PZRU/34HXRharAMHBXQQvCH6m3xT1AJGKQqO7xxDYEOt3Ke7aOW8GQP0iePbk4iSaes1fcmpav/N
Q9FN8WW1Bwv/nqQDyaGBY5JneU0LBFgNb93cMfdiW2S674Zu3jcK3Uk6zXg2zDfW3vBgJaLvyll6
9PtzMuISPvo7NuAJhBKje9zHJqPFkfmBp+ke7cQcPMTtv2DvhI1iz4T6WNL3N7H8dlwHzc+zaX2v
cWg5sAKDLhdPqZXaz8ekp8zdPVRb/jg9Dn2SChXqAR39BD4Ikg580Pm11WQAojDGUjR2a8Z4Ff3r
YWAs3bmsy2Sy4lVq9CVfTlbjUi5Wo22Jgb9ifPwteDpm8oGOaEy5tbXyuSMcbUGORqzo1V0O3kkr
W6cd8qJ7maY75fLx5SzallBLNTVSXegSleDQKV+cls+X+BI6dje1jCqKIdeyQ0wGK4mQ61MUcRRf
G/7pt1moBnb6BBa+U9QLZZ88pYa3U3CC5pDVUo4DtgAFWPV0EnJFtlIb8VqKXF6Y4Z+EcMalrzRq
8c3oSkqpVMBqa5Hp2MUl+ZEWZ2adgYPxV5xHSIqbDrCqd8dabP3AepnZy8uMKcDQoVYSdD5NtVXB
nJ1SGxq0eSz19Az/uro5J24MS2pDb6IVSv0ekqhmBeWyS3yGg7lRf7IjRPbReq6TrEEnQmkpvoMR
BkxfdSb8PMVCCW7Sn7RD4fDQlkhzIj9/j6J1BfN+9Y719d6cPZkez8+czLZDwdHXw7EQ6Hot4IDQ
dCdOVDtLdhP+vmtsDkM64drs/QUH1gBfscBK7dY/FgUMO7vx370w1gK5ROCenIu2fUi4T/MTUuxl
hVZU099fJVvtKkHxtMATCSHdUBI+0RQO2+oYlyVQImybg2mn3VLuhvxJj8im76GHvWhq0gbEf1oC
EGpBQCW8EyS6UXepU+XpLBSbASkSSRtFYA4Nsfan+4GyY5uZQzMvsFIwz9FCe+GY0dBmRWZR+MfO
2jgxGR8eZJhYsgzDodEQrYSL5cSzZCfqfTopgckksO3lsFFOvBTV0O+UjFvcW1IyO2nB0lU5uLhg
VuNKLyhA8NKeEVQ53r5NVwe8+PFgAhhYDDYbmjW/2mb/NMrkBCU0jOwB17qcekY/0164jXuLSlaN
B+oNOa0Hebds5iCNtB4VfxvjoPB4s57/Ptx6ztPB93vzsejzOBusFFxShqHcBDTPsYmvrT5syDxh
wfawCE4d/v1ovuCLxUabkY9qYdeR5DPu4L90jSH+P8VEXZxcsRiPoKMfU/jjgYhRm0rHaxnXdvtC
MN7DtCzZ03CeLtvN1uz+FvckaRQzrkZ2ccbmR324KkBBSudwVb4Vuoai16wjDaSf5+nxoboGu7rk
fc//8XV1Ze20TO1cqaigoSGDl+e4hgpkwGNMgTCay8nB2HozTZV9k6NpcGn9zBGTwlhGt45biE3S
59fwUoagxEXkg7AWBZwJ+Jnak7UNElArc9r5GUMv/VvFiwh/zEkehIYQFFxLV7PELwjAN815VqLi
X67499wZI8HVGs8NjY6+lmpwyhRgp08WUtM0DWA4PNa7nY82Ev7F2KSq/7cQb2UHmY2oFwsV6pov
1U2NR7i7PE7I0uNneV/HYXMYmJN7lbWSOgOdh2l/ETflRywlVvgGOBpDJ+YVI6e7qspeAyNcuoo9
6VAy63a11IpWMJzfecymF+BtfnGhGzUOFeFFVHAtQBYiM/+HTU2bYIy4+CPtmkcSGXBhbD6oAupk
kC05UUqb5CBxeN7VRim1+x9D6j5Awqx60uz4opIVaTtJ4X7J1uEykfjrZhnQncPEnM8vVegfmP1l
7Ek88Hw6f8Cp8cTxypoGCKuIp7TYeskM/jTinqbJb9C7aWPaS72BlGu27cBZUcH/fpSnfHBf/C9I
H/2W3SGa4D5n7xKi29KOGXDnJabAqiNK+6fw5TW+rrtIHCT6zzxjL+NeXlqJ6tb2PjSGswdvKH8P
JoHMzF3UbsoQBaojMyzoV5UWR4dzl9WWcwMVh9oBCWfjTySaTgJWdL6s5o9FNawEwVfNzqpvKIzi
5ws8ksMJYSuTe5fpCFHi31S6qbYuXA9+iPR0zw85bVjHezALqiYuPA+79Bv8+z76KG0ED95aWxKA
2hLA03bTX3DPJVqYtHGKPsvKuIWC+Ore5XVEec8oJUBPpWFZk+BKSQ5wC71RW0hpAuGfVBm10qJZ
/kO8BnrV/JkTx2PBCIJsXoy5tHLiwz+0xfD77t+Z/EO9DVRTtQPr7HXemwJcXzh7wpD9PqRwDWF7
JAk69uTgf4O0tVGA8hQqpRJkCh4Z9BNaaXKqlYtaWRy/7Phc2IzFAABI0OdLVz2FiFUBBDdfRdoz
LxXTKF/ujUVQbkgDM2ZGr0S0ZXOFRZ92WYRojMx5IzG0eXHLysiPQcyQt6Js+JVp7Mr2b0uWQzz+
1ivLPUjoDdDaM3RXPNePsNLzyq7B0lHs8A1i76Q7DLBfHMSq1AvHDKqUndNLeuVpmzxiDsP8RFQV
3zP7UF0oY+rYuKVORlJfkokakCawT0aPRVmWsbQfHElImJhSnzrHX1NKJUYoTgb0vMYuJphnbVix
GoVsZSTdcaeNGLXXf2+RP1QRvxr/EUbqVwrR9bXiGU2ZyrzULkUGIWjd08k5lbm423V607YniIgm
rCIyNuRXMc6dGxGe8/tcVMiiTIm+Dew+nVq9StJuhDfME/QujND2KN0hujBizHVCnaGlxbSH5oBQ
8DOG7yFSx1U1dcR9RibK5TfBg2vMR46o63CRlKWzcYtPSk9WsYDET4oLIBwPBpLipFzBOarnkBt2
j5WBjn2iuRBGcNv6nhSW7dqOvblE69J3T7VtASnWQKiq4QzsqGiL65zpFJJHksFfMYgcV4Jb2CoZ
nEN/JC0HLZT0yrDZcL+Wap7QWvmB+hQXaT6N/RozzblRdvhXK36Y8ShteSdnoSyMKRHCBHqUcR/D
aWb2TjTc28JmjKeNKdLdSh6/xy0TwmRAZoPxtRSIbYb3ffIUAwHlvVHV1HkMXSKpYmKVeo+kSyJg
N8HaphP5ao9rysIOzqTykij2JMJWTAiU72tfAMk/1/yyBin9tXUFjCV0J0PDO6KUPwPvZxpar7EE
QShIQ3fdmYLhYhemm1L2uNwXb4MLCH2+uzwc4qtMJxhZWPr5IM6IBHIy1GjArd0y81rS6gN8q4jM
gVEURbA1BPYzDIp3/EyQ1mSfIFDFoQ3pjkz903LPpy1FOi8bgwqEmsRNKa2hW35Y28SLjqwph4wa
03hF7cgHpL3H9dtBfXBJtKSmX3EM6gN5frbzbQcZML/SYUcSiT/q7+LL/5flg0tJpckuy8euXjQl
U7xkA6F5ASyS8qVkgcADHjAugBdW7aKIjSSLhYFAnZUgEYerbhYjUoMWo8wGtibT44RcvvrTYOzG
hDHWqX+9b4hu5BrdiuydHWkukz1bHhvF5toYZAu4LT0zZz+t/BHgntSOZq2dlFDJdf7dq0806sYI
E//5TWZI2QiGN74g/ZgNBWWx8cd1V3jUtjfNTZV8mLV/o9uzL4eHsrw76I2BAlqYaCwSsopyvZly
a/qqfQPQ5rgaPTWXxN1Zyf15Jrcr7bll3RzOPk4B6dfGiTEqO/VJjSFha4VVFWKDfzZUi+MRv8mv
UlR1xhAPMw20NjuUazoDhovc0HEXcu/x/T3EbjVDpfGnK7alfJXi8/9ZawXxp95hNDNmKdNECUh0
2FllflTVY2obNm45WY7BucJ50NR1YQZavjrlTo7DMRqU/7l85KczhYSHYALL8bJyYWDJUY6n2KX2
FoRuip0/8jZHtrnwieu0AbsxvQbgyxDg/el2jU0ogV6/pMpWwBN7N3cDrmNq+wtOqGA/ICq950jf
e9ng1KT7WBpQXsrDmewOXlF6vfbQNJThKRSQqUZupf54kjEEbCaNBmgFp+mKAYbPlnbAr3YpUeHi
d1K15/fGUEYVMC3nXgewJbrmEDmWGlmy9G3DKPWwCuxQFrfseF9PoVa9mnVHpdWl+sJcqKnhnrBj
kX3eIoDWdWAzTAWV/OnnkcGDbCmhqY/gI3GG7LvEErbeD8rBc/pyvS0JY2nKswkcA9Ut+PYoBYVz
S1zXCdFL6126Qlb49xz6cyxmHVyDgChapTT/1jfeCHHdPZ+s943w1Tija97zFeXbqI2OzoNwFFai
tRxrEr19BNKEKe5WJKDhJVIIqLb+3/o+2vBC6fycLH3quppbnTh/Df7D5JACo+8vikDFK2Ic+X4b
Ima4YM6hdgjzx30gaGnKu6yX3Xzo4IZ8wVSVB90xRDDqqkAAcU22NyE14rnaGtDur1Kmo8P9MTrk
p3oE3zU9D6ShRO1IfRuHUJYDnJSLvFpM+Ynus7vxXCKN3+Xee9tqfom+WEOJqb52B8aZo0ffVO50
2tYkaW7q+aDOAom055HsQ6ije09NRJoTEPSdIK1TCgA2QBT7f6v69FrSlX1xTeVlnIdhe0uH+I/g
VmlaM76S4kauyFRG4jVkc5pGfjAlKEg8UUg9jmKWxtT+xjEU55p95K+GHsN4xa5/8MPGITZsDqEb
3BA4Svvb6SpebyAN9OxFKRSPMVYOrkPmxxCc2/pBCBe4Q5zoaLQNbfiUTuvVkHHSH+7mmnCVGs+r
PccNLVXEy1oOpcorHwfOZy4igJUGq0DVbOgRhfGbSESVGCZo9hamJY3BI99A+v/LotZcRwIWAyzp
Z2A2W1UK87qc4XgMPbxItdMS2iKSzJJKkTWyTVPKpdC2niNhHUjKmsQGO/jnHlGAF0BaihOiWIgb
GAZDhVjgjuUfMXLxjdXzMVhmns/7k+wF4zDn7oif5DgH/6RBwdePNXAIK/UjVyMEGp0mMwhIsbAh
M37KZmul7/sMz9vSIwZPztSUyGYOExg5doob716so2y91H0J3RqrOEkFoScuKJ0Pc8OH8IINdjNN
F1Vk8PpFXW9kBCIJC9JD1cOf7tDAhE70dB9kDCHr4nmIf0ZozBBkWx6SKP2UDqmGeqZc5dWWZM2h
zF9kXDpW3Y9b32GiEpDkp7udCQOhCm6zI6zVnfKVhzd11V9JOwNn2grAnZUvHIVg23O8IkKCyQLq
lEuyL2TXpQQlbYanRj7cyMwI+sQUa+n5SPAwQE0tVS9kbJS13DlHtjCtg4ps19oY8mq9XSCgz66G
+qRQh4M4csn0JMZMHfyw9Q0Sw+fiOy76gRhFSd1KQI5XqyiIVhBemjONAy+gUOivGJ75VCSXeL6x
QkOyHw8AtY94hmB0Q1uzDBbnqFWGBVy1lTgGPNyM1GUJLdwLT2/Ke8mpgo+oR98uMJ7si5yje+t1
xQogZi9ZiM8wygDL252qm7DjcdBHFjhGeC+qeENLWJ5LJEhhR1zldzN5607FGlVKeVhEhswxjDP+
AqSACAjCG+U6qgZAYWvAEK/CZvnsDU9UTQ8RVVvjUQQZY0C06plkKq5kht1+ugQMeukOI05q2xDt
RiunMspri8+SQAiGpdzSZxygcsmKL/rq7OJOJl4mvx1stSV6GBvo60Onr8OcfMOH+r5NWDojiw8g
Aj3ZI2e0rUkhnr9vP0ZaKNJnouAyqXBJahtFZIzdiCpXFcoe7nAhYKm1R9qAiRUtA/qIiMWzt9W8
lWJxWsqfc8J0/t1lDJFlBrk7uFZZRHP63WCG3DAzk6wXyoqzctdIp7KMORT4bhLimhVr4zNg8RDK
f00FE+itFrMGsnffxbCB84GnmkyTrNh5Aa1/gN3KnJpo34daocNW+5vtfrN8f6FjmjBxfEn+DLO3
Ut+kQhiwDrNqe5U48TmF/ewe1HD63bH7BWTZvOdvIDrPy4H7RYguWXaIq3szMDKv0AVDXf9ac37t
jfzTKfdx3qxpK0djGT+fcpK2svkEVXRn4m3e/nFhIePurGduswIVYqDkOe4VqM1/gIL8NCSVWtcm
aC4APL8T+cBJjiJR+LpjVYPms6Rqvn1WsPjDEM0gQrcpuAAUHJVIKixkXnrsHAHkG7gGUrwKmgdj
fV+OtirmuIeqvHPHPzQ0P1jsg4r4lLWd2aLeJMkaVViJPoq1nTsdPNQgsP284RlNLRdFXEjOzyQA
xCktukM3lhNGxmE9em8uCLUmO/9R/MKIyAKjZZIh+1YF9/7uls33Jy+nD9QOz5tnULsfpUvseKTE
TpxKTW/+q51URKWx+Kp0uuxlyOGQRjDcsiavL6lu7rruF3RNa7huPJDLpNKOIpOBMpG9bPHWBJxD
+JCEA5/kFzkjfiAXhFZG+/Qx4vM7z1VAgeRLRkbFKp1j0NdIc//up1EVrmdkWpwduKn+TgJ6Vs33
2vGNZU5XkqDny/4CRZIKfJak9pX7Vw3zcyTm2aJmp8u+n6votv6Qs1UrwNjW/dSmmOgGmiQ7/z7R
Q2EdRoWFNuED2PWp1tkVgs+I9IhJ18hNyFiFm45lCNzLzV1nZA12oS4yK4RCVAUAlmpjHx+FrIcZ
3QKQp1Ri78oaN3hqyD/wBLc+uW09XEO5PDwwR11P1mSDJ735JPGTn6hwBBDPjodiLZQGmOr0WOVt
1AlSk4yzlorSaaWjC8B6cdahhAESUxNiyel4EoV/0Yvmg+shciD1wqFWxztkdA8YiFromZeX0IGE
FetpYTpMlBEU31vFmTSJJXp3CmMUBMuiCahkU1fMs6jBMGVqFFM0gyBF8ywz2zjvc3bvRMgChBr/
HcE1cqIU6Ccd7B2spVWVI+A8DpWLUmThlt45AICGdtbR02rPu1xaUF8c6MNUnS5U8rkqi09Mob90
5vpyv4SjF+2xFqEHtkEDAVTPqkRWQFxgNs1ew82XsUd+SpfkQVVWZmWiO0CtQcbAGhBucTM0DWbC
LxG0YnmuZDCA6eEXlEfe3mauJTt0wEfZsboYFWT/JyvJq3wiDFe5Hsvp6WFuwiXUgvoZYpCok1P5
kKqTxe+taTlIhCnpG3JNtpf8sMW4Ucsh3clHvPDY0Wzh77710aWeIOTxCbJSZ7eRH9lftVPwxR5u
gJtYIXxEgvob5YzIH0GfTYseMtJdv8WL6rmJ1hJn8yeXy5+fGLQYTZKZsCrnGv0EIDOAutsvXwuu
Ar6LETPQnhU9VECBKv7OLxHm0v84gbquDbKkWZdr5j5fCy4vsG014ud8mw4CbUNx9PZYOdCZHDzP
2ou+efs7MdzDpkHWaQZAUjrUXQPvdcnjf7/xwIhcNJ+pR5K19kzELv+K80RbF2gAGhGo1BuhrXvg
hjnBrQdmaPdXTYjsvep8ygZAPmjAqBbDSZXnOBF2tznGoLO95gQ1auApgnqibpAMg9AeApwY+Iw2
XAejFPR4Ps5Y1ENJb5TU7opx31APu/w417KH+ewEFZQkUKQk4JUVozM7xR7WOQLzhjRvVXYev30a
Y4WZ4meFHz6Fm8RNQSDQvfktnIpCQK5dgUejeFhZADw1L1Ei1c2Yb9O3/XZxdiJ+hHLtXVtPqyZM
4bMB7CdPp9lEUVjDHunlfL9QhdJ1iI3EQGP03Pw5+E7G5fmzam2ZqnD0u60t+IZ+y6ni4q43gNte
GOm/Jq+AvBHsL4C9kjIG9QOIBSH/TqixcCbeU9JfQbdKY8e67Y2MmaA3O3NuO+eKAEMkV/slfNF5
03B5A5TgsDUqroLVy/MprNn5aeJUscq05pleu85BvD541HKfUelXeRvgSOewy665QGV2wtzUp2Ml
8F9qOAyGdhO6cccvsR+VAO0HKaa5rFgDYkXBU6qJTJNgin976msJdnlNAxMikQCdKWN0zijQlTer
mn6OjZOk6SsfnqBJxPNi34xyd6iyuvauF5RJhpfGYjpaJlr83er8CUTTZ2MY4FYnZKUCL5HcN4xD
bC/r3Nt2ryyPsnr3ZdGfZ+CeyOKKHA2ROnZP5IpMqGZWNpkO8rZzl15znFS/nPcezutA6SwSjvIf
VMTLGB4FpmcSeercMcZkkyRJFab6I6gglstQFJmhAokSv6KUSkaLzM2I0G2xCb0mHcBW7Po9rocs
BaGXkGMYrO4KTi/9nqZ5W4bX6N1spqkK1090E8UJ+0YARZgVVu2P0sLa1VWVSOnOGND3dxSB+T1f
lHRGEkwDekda6rz3aRKMfpYR9FFMUMLBcyJ2WIt6vnrcaWYiVHiBKTg3pXpffgJoR6MFjtel2aa2
8Udos7G9JItEpjALz78t55o2l3ySCr/yPjrGtjypTxGkK+Vc5RIxRJYeSzdLJ4k641MhLO6s9k/S
mfds5JOT3RDGP+AuxUrz6Z2kUCK580gyz+l905gCiHUbODWpnBGYWj6JG1RPMc4YZ63fI0YAX1OI
Z8Uj89l8/O1oRvFJJpcf4h52LjIi1LUTfVXQBr+IgSlqkSCOshho7ho9/KNgZGMB+2dHnI7TL82I
JCv6Ut2CYawo2FCYt09H+nQHWCLcK3lHFP+79S6YjPxVS3fmwr14CGvdjXHeSx2dGmI8FKyFxqsl
H3uya3liweadakupMJmeHDZO6b1KMdpsp72q943Kf2b9zeot1iXViwrnDcfnJoJl1wkZ5FMPBWeQ
ZZXYeeIGzKiNeUraQElv5FaHkIi544yAxUCk8b3ecam3IUBFsm/9zISFR+LgygRwyW4WUmIOatUE
wp51sN8tLvWV9xnvAtQ0PdY/QqhPwfEKfeuHfKUoGQBNgtwaMI9XJeq9R4CxRQgDI/w1t36Wxeh2
j3iQXsxKKFLTLCcK/2c4xTb8QKHL3cWp9hyH/WwLm8VXOdtp5wOTeRXfum5q0VoEVXYV6wKQ8hMp
5dYhhb95YlsdquMXjShncAxu/DF9txshMZ5YypussGPymEFGvVBysX5ZB6mVfzT4tgaBCVgEHhLY
HmfaHRl17wSkoEOuq45RsWapLi7RmR/DJXq7yEKoco56xC94BR9IySjAfL62ycs5nepr9+VGT3j1
sOTCZKJgQU1ziqCFwaCgxNts4FKFfIS5zAayzAT8N4SymMIKPL6ylC4QbYGYcBapak7WE/HJBFFv
JNN9L/2TrsmjOwu+YQca7cfHqLEk2PLA4VklD4P9aQoqMUwrLdPCEFJZxL1FA4AKeWPCH+7+rTbU
Lqn71wf+HeI+zsVJIaQXUCPa0c05u/n284574+XWFyva4JQW89u18/u/5k8GDptFQyENIIOtFG1M
wcPBPLOYO+bzUB8I2YZWiJ84zJ/axBl/Zw6vmtiAlfNhFT0nvgfffgA7oK1w7ci8VHZSxsXU7TAx
VCW9LRZBCmW+BeSUS++ZYPM3QhCDlaKI7J2aeKXeVAKhB6EZ9XQp6dfFH+YbOuW1L8LTcHXhyYB/
U/x4hlXZXh2LWngZxe1MQ50MTq7FuL8zkiokvGckiMxGjH/y7JOgh8At00r5SjC8T2us4awFRuAW
5yMigmg8VZjZNHZrjA8vD0nrDqliyVUpj13pUQtfl/UW/BXTz27psmTxS9WdP0ZDiHmqSOP4r4Zx
TfzTZ+Rbzmtrd2WNj5XNyZou9Chords4Pp0/Dc4Dv4nYmThOIZUL3Mic7BeRXqtI62S4dW4j1ic8
0n14B71AWwk3yAEJvMrevLWacXOEJefAwq/h0YkMypS8A5/JtZmFhJdUPFoOVmKOgYSDzLijaK7s
7K3WZFCt1cwzoptEFIBWyZkh/IPJ6+TfBtcRZ8o1DjjWvkioDPdngmYNw1/w2Zf3XEBbssofaEtC
IsEtB/Tit2NQyf6bc7OHGnOYYNkMfqKGoZGrnh36qxwcM29iUP827FRkwL3YcjzrP4V0MkynSWhO
AhPfiHwTWPQvKFiCEDakzeJQwi6QW59hldRYq6uAf/6OVxKfqczh4OtYILfo0YlEO2LQn831cXqJ
HAOciEcC/h3+6zNoruy4lECJ0diMYDXNwstHxVSBneaYlKxrVDAkwDKqpJFHGVKbP7+gr3EXiywO
gr4IDTbwLNt9ncrQLxs4vFluYxGZ0CJCOjrRsNKSaNxSWQfyRySk3Gq4qy+VG3GkEHCciOX7u4ah
RToSZdsBfIyo/Cyu7a6M+/qd9CJ9IUopXiiebp1aP40Sr1f/HUTfdde9qTheHncqtAq/v8cV0rdA
cXCpghyIGCRkTL0UFiv40r8B4bV2i7XfKFQMaF7H/qTZgrHQjkpSqd8RkLS1Zm7Hg47kPiiRCFdw
asarNqU0oHtjLl5qbzmpecErI3FAgqwOsFwbzGhGGlJBLRNmHsIzEcVt4/XA3Xu9qfQJR3WDlVFl
8vDq7Uczrl04Uja3NYiUn42SPLOzJcVrNh4L/mHwYwj0RzXB4NAgkNdTfQnvasobifRfmYzTUjKN
HBkPcYP8OWC4ZQKtFxhVSRi0wghKkv4zNtYB9GXMdDnEsE++0/WqXrOWnRGfQO6JfES1EUldtYWL
VTIovztOhtUcF76A7s8aXOPLxFa7xi97tXk9+74pYHm95h234U1lEDgiH8+gj1Svftu66w6dGtCj
AzpVvy3PwUzuNZ3jrwnLHxVYF9FElmOoAUpEW1wVW3HrSEMcQiG+2P9D6gFBRm7t+bIv+HMes07t
bRWGepWduR3RanfH3TVY6+oHJKQ+1YZ7UchUj1J7twmX941yAUBBiBDLruU3Nog+Ou5EL6CeK1zi
bgl2Nr2vP7N+V/82YwOxwv0kmHyDmXJJ+oP3z4cQeoe6WXHNtNX4/LK3b7TN2ngGIN9gnUSjqFtW
0zQqUIh5jSy5nRQath68nmEMKma2BjyHQmpN0Cwl9lhbZmPP/i4ADAuOQrHeL/687efcp91gC+FT
4l9lWoD95LYNhiI1+i+jIII3urw4rQjJW14Ib5aXVj3WKUsDQ+Y6RXzVa8B8aQru4qcF4EuUYeRK
eWf7PP+omxoYmDvPt8tiR3EE322JgfzHUMsI5FQ9ppcuCu3BpRxuzksoYwXSdAx+4x32w+TWbvZm
yzYWvhM46OiJWjTjsQsGXdn6yA7OJIIEL6DRaE3aARxSdKtRpBFTYwf8bgQkDF7CV5PlSh/1AfQq
GYKxWGnMbbBEoXmMYIS2Z+GCqJIWzvi8nBeHHVS0j7Ny1AWmMILwqe9TyvzB2jMNsXcLjn9fh2dl
1Os4PNptv0DnadwSiwH7S7MbAdWtDuoekYGa4AXDWd8QTxmR+RCmEYhh5yoRPqOMZVYcwPi34Pd9
GhdcQwKIOHq+sv08HONhdKHl9efBBSalE5IfVdBwNzE3CGnclmFL/gizkIi+xOjFTXyAiNScUfMu
ecS594Qso9ruz+ETDZRXqYs0NuyXsutc2JJj+kz+QW59NbIX5tRGVvURidyOYgeanUL110XMXoD6
VbQoWEXp5+s4lBgYHh6jcKo+mm5bLen9VesMK5CMBQ5Etzm0qSLXiaEndmXkZZCvfEbJKayzydf1
hpOcdrFSKcCzIVeR6MIXcU6b3jzgRw14KrKlvCs/g8BxvFXQ1RDoVq19YfoVwa+7KzqEQquDQFR7
dELQNHgfw3rBbjzH7KSIB4+hu2fdnK2fTgc2/ezY66m/c+fEAzCtDEliaqMSYutD00a+43eDXvii
5RSSvkGS+8GQ9pRFbw+Jk4U20AvznME3ZNwx21DSwy+rMoDhLYM34nxQA9b8YHZZ+eeQS29/Rzcb
uw7YRlUnkvxuV0d2Jwr5yalbeafD7Lr5x55H36m13KJf0nm8+eXcooU4rjEZJhfZ4Y2Y3D2pL+kv
Lqa/OGPCHxkpqhbBkRkMweTs27K7Uef4Mnen9dHg9Yn4a3lHJJJMEpE4fDxAoIWMi2gEQEEH/798
bvOc1nwBJXPvXzguSN35uzvs68G+7EI6UsmzpZOEg9L+YbMbLt1e03hZXX+KkOJw54W+uKGdLQ7U
QXfLyN1DbmIfi7Hg5Se9hHlJnSijjosjbi/Ko0rQR9bDkTuZGO1fm89sBLHB7TkG+2pFrR/nAE3J
y/PZB0FcUZ7dTSoAQCtTX6ueYf2ISAUnFPEsvmQGh4VwuVd8R+Fid+C3dFkFmGMsMj2eXnZhdbLb
LKdT+qP745qtwSGpykICDFjiBQ8jRS3AdOiZzkgufg1XZkkXke73zyzwtfZvS09b6l4xuBoj69Vi
bwV9eVMM5elDYuTUvlSUI94oGWfphcGr2o7udefw5GknZgI/wb33VX4j2Ccc8yT6EnoRoOsSmkKm
yM1j4neAQnKVYQaJkALbjv8VSJ/RUXZfUKTAwHO3UDNGX69/viKtAazC1ibcvxpt2EOPkrg95HVr
WbCxabw2FXw7Ou8u0VdG3I2UxtwJu+3tFpfQ6tgfyXmOrWKKGattPh2rWkXPz6o3Q/pBV/lyqdeY
2yVEqVMxJsDduAry5pkOly/rwYqTYbFYXTbmbHtW9cXUYUFpRXOPaLlp4B1CwcQWYcrUKFNDsn+1
yte7BQTufqU2KKTqwrydXDbl/yuES7LJGt5ZISxxesCHLcsg5eaNvxztZyfZHNl2R48PTHBwIsRo
qlmr5q8hfYjiMiSxoDhS2FLzLbuupDhgDYfAZY0+qiVihoC5SGsWqtFHQRnHdK0Q2mw/xkkZO6tf
YufZvdGItTZgiFqejfNAOhP0X/Yf57fTiUd1fvXhuPaz1IalQaQBVK8IebNlcVQQzKx9snSNznj6
qekB8cVvFG8o8RuxfehSKDeIpFYGidjetBftvZroRYz9Dbg6zw6EXe5WUaitnIRyDSl/NftRd2Ph
HxQHpViCDW+r56k4oLnP0oFcmjpBoK8PHGm4pv674eriZaia759tzEUH06CZBJItUJhc+iBH3udt
9ydZcxcJqK1gUSIn5QM3VoX6HJAYEC7naONeQGZaXO/i28Et1dxWG6Od+CCGlNsEG54lJ3ViP2Gz
e9J0G9fjethfOaQW9NLXQILeo83VpeNX4wQv0eCXOtlqwZ38mCu2GNPaPb9XV7lJgXwSlfWk0gCK
EXtM9gxnbkkoHBUn1P0HzJLTJ0Odc6KHbMgpqH0hhFsWCJoobNiWsKkYI9J1iUpuenxmHzdiD7p8
XJbMQRbjM5MIKveB++ukK4PeMF4Qchfxeu05cL2eIAw1BT2jT5eLyclytFl93ZAcpPmVI+wE8kNg
zb331U0yGnrkuQirSWwzp62HRi2/hDNA+i7m5/tbTmEfdmvzFJVDUkKYu6rMmIRp+4LTpSEWfmz7
X7Z5g/gPHN28oHFIzlkEIUSF7000hWu0Kvra+PO+tw8kLjyB8vusHZoaWADnjbjWnUH9UEitBIVL
9YAn8Ad+tpOF8ZZuTQE1rNH5Lb+nsXsbhtBWgJlY6EckDQs6JPtPwgXfpySDSeLVpbMW1idGHUwR
McddNjtL8g4Htv/DOjat8KS1yh81eK7LvZirOWsD9NqS4SPqdcgcvsioUlmfVxP4+r2Q+37VsB9W
sNtXMMBTjzedBVnBA3L+qajTxjQX/AwB0WXC2n4tjo8nv6y937I1lYQFQDFpoHOSomQ3cOafrDLO
IrOUcFBUGZytRzjpd5iZabo1Njg4kmkcu0W7wxLdZHFEYIZ3zhRoZxm4xtZLx3XnkCdW3tD/DfdF
B1eTmJBAf3qgCrU8aHZ9jvUeogDuwOmpJ7ntcipMih6Fk1IlJHWPgVOdaOkH/nXsfPRz5e2/8VmK
HmCiD3oTI8pTVXgDiIlnbA1VsnhNmSNhdjwKMjFkfe9lGHwU3v3YycIH/z9BsVX5EAfrNXNLAA/G
oUB9uBqFPfe+aulnPU6gW+LZTt/0YzMWCrhmVE9H7e2nh3+tf7FYklMhITQ/8U0why1v9r0RVhLT
Ps63P++4YxY8Cs770DS+5mP86wgodS53Hz2b5Z4p5un705j7VmWGjVvgRQEAYYKD77TqCdH9S1bj
4qGoEogHxM6Iz+4v39lYBZb9SJLj9lep56PExosP2yFuD2lQyK8S5HhHGfWR4uc33YM3EEZu1cTm
z2MoAgGVSePbN0rz8S4sx//NSo5LYPTjBn7UiYN5ciod+/t1DPhwq30Ym81tFT1thfjydQ3SIHip
pfzQaB19SiYetpuwHHLuXoN/VhPleEycDKuyZUkjKGR+dcWFuum+M3zujm7+Y8/louWmRxa8l/mW
8095FaGSO/7Iv6nfG132k7VrYiX23wXMApjY1NNYtlUHcmhUcqRWaWx4JKgVuxw3dbSm/8Jk3aMs
/CVf5T6m/kl1T+yrJ18+G+Um9WzkV6fTKXaFDsHo9/E1/jvzuTWuYuKkjZ6QoAG5nokV+73dPtdi
oYD+VESJj1rEhkPtpD66hvfLAlGKnK/jiQCoI5v0ngJ23Os9qHNpu86J2EvfY9WWA33RTEjltnBb
4Z044LnMGuTwNZGHzdpMDs2HdZyaohAXJ8KoW2udK0XPwgFaFvvoUriHPdOcUrr5kodQjYUU/AsP
WN+V8bB64AVa+937awJH3pOXH9C+tPXB3RbAyT60S2Qdc0nvFTACBeYQMBcc2teyGkTySNGS6Aw3
iLsU0bN+fINZumF8ZiFHc+FYcB+Nsd3bKZGfl1iMFTyNpwDQb3maELRjsGBn5oTqM+NhFeJpHtIa
vmrGCA8T6ACQqox4Ugthl3ttfX6rfduJFClBtLRkotonEBI+ErxR+0sGzGVKa/b8CZUof/3DNMD4
FWI4+sbKjOXoAN25BaCQXtF4sC1KBHA49qxT58j4ccwPLJOnmvWM7t3z0n0hrVEa/8rkT7xOUE2X
YpACkCLmRishkCSWK/eAQyK+y4ELZAP5zLU4gU2S68Hy8xzJHXJWyOyd+O2Y1rsLaxNcnLHebsTx
YrrlUqkxltyIAB8mdoX82t0/l/Eo6ArDTYrzLgPHZvzIMxoeLMZ9nao+E0cICPYwjgcGubDmg5B/
s2+WQRz5DeQzvqNZqxM9SqnWo+jXJbYjHZnwLTUPHza9Y+wH/0/hiMEm1+dzvZT5Qe2kfOKvNQUe
R7wTpH64vaLF3JHnwAFCY0aDmNjIRKnvJ0rHNIxYLnHdyChszwoGuA/+sQ1kMVLWEFCullPnP/oS
3R3OghE04M+wc7JoRAA/9KcutbqXIITE/VNuQ2wlP2FBqr9YbBeVeYbcA/ARUenv8ir9YXg/4lQf
7aogWJ3j2I31aHvpzUiuZ10+X51EHUpaZW17cjXAon9XCrjmOqwvb2Kui1ZNazfQ1nofMM0bCiQB
k8stDav2yDS3BHLy4q0/BLqD6BlzyuyTTL0osQsGi9xrzTlofPBo6645m0qiJl3FyT4PoDbqYAnn
5cKd5SnK7ccTm9Zeyu4mDPFDRg8L6Vi5Npog5u9C45bk0lKp9c4k78ODwZBrfDm7NrJbrqPEP7i+
fpwF7VW+bt9lc7Qxf741CSR5ATfTDPM8gDpAbXpJyjK2CThLwk0iU/s5juK2wA3JeJqPYLGZgZXh
rUO7DUbha040aGhJUqfj5LCkbToo8psttCqrp2AIUnD/9Wl2bjAtkgQ9ugccuP0Vn5X11kFTB9Hv
gC5h96TMqTyXcytElnZtYWyMjat/HP1sXKm169/W1aCR0+GqG29O+ZOg+s2V82znjr5NZ1qkRE3E
6ih+0QjKjyUxAQHufLghlXUbgsb2n+byqCFJfooJFC/KHJzdZr8W6R6yHCS1ckO2C5c9s9ctjTr1
fUSFUeOC7Z7oqOLCzRlYffwPwpIh2KLVfqT1CvTV4inavLWgWShHsS6PQVXCzuF9OKWZBc12nWvA
vYXc9sCFRaQ90ZsafBHtUtEjCJTOD+apD5DUBm+JDuFGcr5K4N038aHYDysuj/44KSzfL/92/2Dn
DORDvHoLxduSaxem3lNJfiV/8bAbtuwc7nB1qaHWODf7mbk37eQYIjzAFJhVA7hshOplU+fKIexk
/SLqrF6EtWPJ1GI1Av7+4GrbtPpKU5WDbRpxTcyZSL5M+dSOnv74IMRjc3sk7PCC+NB/W0A78Oxf
v1B0in8VMHWVDcRGIIe12yw+edo3+k0jpZ9lYCMNhzVdA8lDXg7QfN0mol9POWxCsHKLhiRKLAZi
hqUjlTWbyO+OWHPeHVicWIsv3lZs7KSHq+ijkFnEi2EkUOfGSDYvwYimHDbvP7JkUihOc2DcwSPD
wSLLjT0v2/qDgncDb8lJAnZSmEUu0GmbxHWuqg4SvQNWUolDwo5wW9FKeCwyvaLIJtpjnZO+y2oA
hbgyvZCpiT9ZrwYbgzoYiaunkZSV6RQO04q5nO7NQQcT/1V9CQGwYVn04ewdzk3Fw8U3O3QS3igt
3nn86J2f4RURPUpyQ4vyQBVySvDedgSeJzb1h7dIdCb2hOd6c4QLUxZHGzXOAn9wblWN2/qz3jR0
ZEPXFYR3YqGrV4wjn544ekEQpGE/Il2JC4E0rDJkuOI7Y9+5rRtwtM4jIJ6MZF/8cpGdWllOOWHB
N6MTQoy0icUHog6GdYdYR6Ui80xhwBK0jiNCcAd1g6ydJAPw2/pE00gVYdMYxbjvilHrtOGiuH5a
gYrntXgLpErQzQRriLwtTYRSGvqynP+XPWTYoyVDpFkbYNeDTC/9Q/B+4oDR/smCoyPjzkZxEmKd
bxvMBRKTNpb2txiPAURHCiwQfTYbpd4u+qECvzriJXu5wrmS7OK43mS2MQ5bv1ktb58+zTEvGFgs
3JWXqmCxnavC4AJxJ6SHRDkfj9e+mRo/y94HeOIzpnr3fnkSahF/gz6ycOU5rxCdMrP0yyeHnx6Q
aDYbti7c6vD1IKu5/pCRN88UWXaN4bCJtWlLPJVgfuU0/DlJa+hZk+eoIMKltAQrSN2EBnnMTN8H
d3Si5ihNOKPSQi7nsiguUQMLiYXS2Djr49G+fiUoEO5VkUkNzlhTbtDPXxFujAJeM3PggycKgBjk
K2XJV0qLsUyQIrJFB2bmhfrXsWPleRjY68LNPOGOGBIQgqauewlyxA2NE/EPWvTNI2l2BZF1s/bG
KZZVDhfHjnOtlR6CSd1jsJnRDkJQRoH+OM/dUhWt8UbhQ2VZQMRhooKaepr1c9hcy8w6V1Bf9wzm
DbdVjvjhbuLVLrWc9uNGexrOD+X7FJMIUIQSCliX8Ws/+Zgg3wcDKtAvYXtvTVh9LBYEHAXVV49/
vlnFwQOz71YAbA6ZABpJP4YmP5Cnetnvv33rzDDVK9nSXj89w8c7mBIdszOXBr9sGbxc8Ayq/+z9
DlsLI4go4XSLkly+bI8OCLBOnzYCeHlhvoMC6heMLc/Nb50RcWQc5XUOG8ZSO3vMZ4UtcUPP4mqc
nvfTEIKzGsD6yPH0KBFjIcBL31IaiV7YsKlGqBg+qqar1o/CzVIO9KfHMMOBOJ6Fkgmt/yxl7d8I
160KYwJR/LULf4Yco0vTCiM0A7sAIeZt54nr8skCi+OqXT/m6WtZBkLv5s9W/MW13z2AAc492lYs
6gqAF34/zg1AzoYHvw1iHYHiP3cOSrFgGTAnR65sKqdJQ+QWRey3ccJ2mA/AUCHwrt7fhqUY7wrt
YoQp9dk9ixqB0UufhoJyMWjpOC+7SFkywLyIDDEFWMe/3IkDhXfQO1VQRsVrzTVCDIopB14JKG3S
EDS3SIAP1wzuaTb1yLSaRw298+IkeE46VCpY5yBKJkZtVDL+GoU3qDhQ2TZYbseU+i+I3R5WD28A
2Uc8c5askzifelifDQnTGmdDqqC9QiLG5IengsdLX2eF+R3RRXK6GXskuasydWB0bzW8qEmLnhHG
urHUwvCdf3Emm9auayCCa1CgFA2sUdCC7v0wjxffJ2vKE2LBj6G4v1o2tQdXSwhHFQxU5WHBes8a
eSGYBbLZC5g47BE+1SAvSIudnY1ctAOijU7uB8siATiOQO4RzH0VqQFjtxDhpTFnkN0b1fdKTD+3
3Nw5t3bTn9vleaU36lLnsGmeagxEu810N04fovtan/+LEt262eF6J69o1Zj4fwRiND3Gf1xdZfBG
EDNGR5FW7mx/vjrp8rh9ZaBjO8dqklZ0+i2JwZpaH3zh1FQMUa6fdtQT/6a4JsteKQ/szXstL/jO
jNNvWKMaMZyZGTC0UPB+lVnoD8/rqflu9UTZ3az+IEorxbLCRV3QVfMB8Vcw6i18ztFXgih2ray7
CfCla+n6YUaGcyg4Z1TH9UqjsA9unMBnFv73KDASJoQtQaLQy+Bqak8zi0+Pjx7wl51mS43U9eG5
wIda0va4zjnhlC3A1rA5iCHhngqcZ7eTAIufW66vTG02rx5rPPCJcAQeGeT97rdyekguDKN6k/YA
ubnrs0piMQuTtMxY0jGAyd5xO4CH0Pc7zTDELE3P4tIHgP/aGrbQQNMm/6eH55igYf2nsjVdzQpV
Y0cQtwCSHZGu02zDA4UPSAdUuCHYUAA+0P48BXUs5rmyfDd7Cg+x6NqTgwOfUeq27h3xbUG/XSIX
HxfZKUTNvLY3IkcKG6APUMiX711CJSGeyzahlsGwjUlI40ETX3nz6b8RyKFfAZ6+i0T9nG1voZ+T
ILI9NMf8QfPEuDe6UlSeH5pp3zbUvKt9LCToCDo5FXhPamRJA4pupdxgGRne315NtkB1GeEc5/HG
VOXS2KAtmprELY5RCy8rb+MVGssXs9saOWof26OtUwtjF10Gs1kcrn88yGVD5UtfjiSd7VsZAcgQ
zDYY7S4JJ2hTkr4YHa58FctUH+E6SqFc0wNva+uiDjLUcIoYbPHRkAGXq8OVEzEIWhIwK3Z7Lzif
9LRTffKmYsXHgjZoYRq4kEEyYqxyT5r20jEa8HF3Qs6Kg+Ue9ydSl2BCq5nHC7rDDRjmrqfKtCAs
Kq1ZkGl7U9kqLLz+lnIXXLCy1ZG3SeIn7nxlsbdy7qtR8ynfvLjl/I+tzJ3ihppZvwbaRmQyPSne
ToXiskZTdLdZvZuS62jqki1KQCMJ0no/dGd4ysxyO+YRNcDhzUMul9pW9Xm+o8uGb7mX0RxGYhnq
QFxTLp9sMzgCdi+npJ0PAskll5m1t0VDkx+FtTB0MvKcom7859maBOXjJ7UDpCutG90ADHqkL8ah
5T2BuMOOLIo/VArdDV24pMGHwxw9T6uy+VAA0qgfKDhaJrmubiBtRhIsuJcW9gsMtnjBfbtsYCOr
r/m1D9hkO1vAr9MqUdSdBY66eJSY12tpdu8//w7dAPbNfZbFklI/Ju6cdNxEd3RcNES1ZauARGnd
ZGSM0TJR2AyrHefJoN5mU+BrYYf2+F9iJc4B7IPrPfCZCKfOXDlwWs61YEufht6jcJ1TuQ3+YqOt
c5YSyvdsB3wQbP8Dxh/I1LwPp43sMz3gLR6/JAWzVMq+2DOlPavjKjR4s71uyD+DtHE7rMJDLrWp
RoY9mcQizSVoLf3rpEob4t+f6fbzPIToy9KwZ9JP+e4QKwPjHsFO2CM2hdhob2G4Nkz9WQQWiVOK
wreus80PWIzcn/ttWNNW9mqvXfoLKIa4aCWW0RnRtbqmPVM5eFwmrgdHjQ23BY0A7EH03j3tR5mR
kdyKJaEP1w/soqI7sUThI4UOp1gru7D1CPBSCU1/P+j1rZ8ABS4ZuMU0ZImhETlUkUE0Sdal5Oqf
oCipry2CdEzkT801K5Flq03mRwbZWtHvdjP3Zuk6mZ09Q6b/fyxTw8OFXgq6bGzUV4M5KWa+MN86
oPF8erhjzgHE5idm6dhk0QkvCLP+EDWQZFyh9MqMgKxMXO0gdrlE6Ch20TPi/g7C052fWxuni/pl
femRnnLJJJGQTGB9uuhcpl3zbVQkyETi92wofN7g6ge0cDygW1qcXAiucZrhJP6AzbCB4MF4oG+n
pBuYcvrhMVJgquszErrmg3jHXk+c+Mh3/TIRbnzI9+f3JfBLe1fL+2GaMNyi0ICxa++KX6KDX56t
GSFX10318KjPe7zxS42ZQWymi48vXMTy8EZV8h3drzcNy4G9yCuqX7ewFf7Vflf1iv2c0OKC+UTR
6voOAs0YRcwytpU+aRwcLGIDtYYBPqby/uw18rIkbHw7tsAqgDwf02lTqoo9jqc8uF42VHaKi405
M5ZXT+QjIKrnJZt4RCN6/bnT5E4AYJkwgybkLpYaUAN/U3pYgvDdjWbRpkExHR8HK+q8HJKMGDSL
4bqyK2ibVE8mQB7xJne4UXAHRH4TvWVeiVTFbcVByrsPlMvE9SUICAj+iAPrqOPR7uii2HfLK2tw
g1stg4zALhbD4BdxwuVPsy0Aj4s1/Y1DKuIzUVi4JqUK00lNtF4TR/5aG21YRXwES7jQz/dDbX1o
pIXO4di1zbvREnfgz0bXWIQlHxOoxCt72WwnSPw7Y7FUBYsxIlgiwvsiOqcGH0nLSUWVnHNTXfr3
ddfGkVBZPQHTl1U5usoK5nlSaLJWg7H+VbGX5Ticsng6goyP+SA5gyOITP5kloNcS4YepFDrLoUy
gOXj39qhj7jUXZuvW7tEVDWwHYGkV70rg9ZgJzphIsKQMkZMHyD814ExO8kfhOBiAfqS/HN52ZrC
ufkTlMKn5oHtKVkr5a5cSFIUewanMMtxPc5bnloXhzsmiG9NsCLLRlVUEM31HXZ9KI8fF8TufdGH
Ekycnf4qXiomG0v+U/qAGWsnPvQMiWPmKrfmMMsjT59ZrIBMMPT4dqbA2SzyPneAUKIiklldVFgI
eJodQx1dc+rpCzGazQ0ZaJGD6jLA1agGNRgl6AOpwkMCKxf6cajOaFTTl6k2nilVWRYZoTxVdYh3
5GNDRNi2vRWXt6QcPWW61VEbDpzTobO12LkgFPOKAYJXWbXtZuPkoAvbikc6xpdWRy+3zXnfKlxe
HUnX9KQkv4c/7dWol9XzrRSonvTEQuV80nBDA7aJPAbSNkuB4bN7oOVWwMmcHs6ctx9MVmryHjKJ
U2+yjzXFlJbvsC6OzMNworX8vuzqOoDjgjOKL2Mw03tKtxzlpZOEySk3F3Y8fpBiDBpR72RtJa0X
nEgJmhKu8DRKWDNNPksgYC/aZW0nIYy7YQM+pgILb5oYNCtqcTxjFHCHCioMRy/bTrYySQrDzb8w
z1DOOw2BH36U3ytO4GZYqHT8tvI+c2Jgypt9Im6XqNVV+91wV7//g4g8maM44ARK8Ca5CgwCeooR
3WP4No2KMMZe02V9zKINcBKJTxUw4bKLgLCa2BPAWZb97nTcBrU7UuWRL3OSYztZKRWibB07Csb5
aUDpfPn9U9LHeQ2bIixWil7pg2HSZ40Ua449mdPpfwyBQAgNJ4j5zTyUI/at19/IYaW/adHTL3cv
hM9/bV1abdVV424Hqxc9fD1+V0+Hde8RSkpDen4U7FuKuuvs8aAupvWQPBPFVgNnwSge8xsKUWtN
rMRhYu6e5YkXhP51URZ9jp6KR+EytiEqEeUpz2e4mjbX9h8vBfN3EIK3ggYUQSJ+zKzDgCaAOjMC
KY1RPpVHDai6Wza8RnBRgCdfe5b4w99Gxi54PqsFjmSNSKS/rzHk78cy4txx3H/xAHuTMifx9qJ5
o+6lwfFIN3ZnUesXGY2IdrqGgMl93CSoUdBIxqtoZaWuMm+6RaK8r31TMcM4MSLoo00YDIT05M2N
G6lrqSLVdsWO6LBAl/tyfaWM3/oBmvNxi6U2oDD+oigP84uANvbl+wVVq8xWcjbEaiCPkyTHxlvF
hByJ+6UoSxgBaM3WL5iLfYPXTPZcBRqlUrJ3Ux4x3/bRuhD38RHqZZUWWy7BjkStLLncABLq/WvU
iOGBLbQV3ACz8mTHDXcwV+jakKjouYx8Hqep0ghgq71hNsQicy9DVr5H4ShnMxNNaNH/bzLAjge6
W5P57rpQunfdVn07BLw94QTMLdbbuL4sFGCKJGKfZ/RBsDZIYjreuSD5WrumxBOuUj1JOvaq3Ujy
4rsv+ZEbpeDrRnQ+xa5KtqzAsiTtKA9bEFSAZ3UBicEsQQQFW92bddKdkkSHw72euZ6j3Mw7KFgR
56IHyUNDXioYZOu8kNd1exzVersNv/4iEsnYHMoqlBpIys/MjY1wxl7TnU/5z1LulxzUKoAgnOaG
FAT6tjHfgJ5dtZoSv8zjiYwJWsMvl2HWrVVJCpLXPI/vaIeY545sLmHGePtZzEvuoAgiOHxUWYFO
7DKge3cUzdjUrUXR1Ys5RFMNc4/rEZr8HcpSBUjhWa+AetemjcNG0XGfm0SQRNt+22PgZbcGXxQG
9dAhtyNsz7i/zuS6aP62176hRw/4+PTiAbiWCOjcE65IfBVcn5BXIpnajAHP86qhyA5nnV7aJSFJ
ag6htEmNwEacC0OGttpbQsJcMbPhlCj6xN1d6lcQzDG6OHqXClz3VRw24d6PIHcf3kU5c6o2Vdjy
4cXQQZqt/nsBY7AtwZsRjCoLURMVRUVQqhHpAnfnh+V1vroR1FnYwLwWrwH7y8lVD/vKKjGbXvCC
rfQi+8u+fmfaO5Zs8DWOG9t1R4EHCFFit4AREzWZARFc4QLup5DVTyBi3o6lLJmsXGLt/viXWFCU
orzFeO+2LYYw4peeK/CzTu6waJpg+Ik+dwEBU/n3LRUrzZEb6JCXOku08jc70LlX/yAM1Exy2G4k
+dC1e+cwFssUn5Ndmv24wkblzGSRbIGU4Fz7QGIJQrJkk+/i9E+46H06Gc7Sy9A6jknz/LmP7wXI
L90aiGXSdK6uncPs6fGJ/L78ggr/YnpL0Wj/M48qBqPnNiK0x+zDdBFZ5EZoA2tr3h8tFmzO6DBx
McUqycGE5AgnQ/1tgWsTm+ijBfIxs7tE0Sp4kWDNXAyuikVGdxBp5iyCzTskchvnuKDNcbMTzcdO
5Y6vfPP2s0GJCY5dVSVTbHRT/kx2UybiqBPXOsnB1mCkFNpoY/hsp/eA5QEPBS/3Ux7sllzVHlPc
lua3pmZ0RxNpVhHUNzm6H1pqiv+pN7tC93rNqdK2DqieCOjruR6DKDhAPo3LWdko0PrUEcdY0zG0
2yYMd++D57VPZol17hOcc30rvG3NhaY9hOtFv2SQ9Zutfh8GDo5tlhoQl6+pJt5amL4X+kD3aEdP
Ke2FEC94SmRks7HCeXl7ogy9d0B0bJtv4d4UAVViz03sZ/sVWYG0xdUWgCNUzRBpv/wbMx6QdVtq
rFrEMfDRZacEyN++Jtk3n1PLv2F1iDvdtntWlzDXgStuV63M8bfofzv1ndJRbZMlZiUnDdKHvyHO
GI1rXZ9dfxjDqmkW4mfoHB+FDtfnd6paO3SzOHMJgQW2/7mpWAOWhTEO102lr4KN+111pUNm8SUo
/TtmoVSC0PetTwZ0gMpa6bWB1+y4uf6AXl68/HAQeK97OlZ0PEw2kG0+KcGtg6RYSVVLtKgONfe2
4yqJMi1YDdaTfiJrV/8g/IhKxXduOFAKZ99f0kwfSp25vqU1qeYt2NDwihepNznd0BzfsZJWJu9q
FoQaqTmQQpKcPt/2Q9JBny4qcMtKzSi01rw87Mz+Fil3SkbRM9t7I1K7Pq9iM9QTsEhIUj/8Dhhf
TFBtcOTR7q1pOFNfB4aKiuUom7lvBO4gucGidhrKDXLDNy/wbuIGekm/pNH00ZjGF/T/qtJYJh6t
E3pcx10nB/b0TOW+eKTUY0bV8DD4qh2WcE4x/CWb6NkXy9wQzzt4E+7h5Q65Q2HHfHl8WGPLxAvc
m3PJ5eKQQG48IEG9umsOhP+20udwjPzzgOWgqgD0ZQeJ/Q9kR7lbyDvNfhbYUkKLtyohWsqc4ym7
9e5POjcJP4IDjJ8Ec64AkRjggw58grubHJ6o4hP/5n7HPyCKX+aRXYzlITZM6YpDVAMbdoQ1aBUb
Hoqs9xQQ2ZV5rITB0pXnW3w+pAdkmBF0fshFj6ZPBuPycaBsPoi3PPAuKEgE/l4Ihv9z0Dfl5EIH
SS7b29Eg0L1h5qFlYyojG2jKOFXGYogTOFVVVNM15hqFkAxulBHE6f+RB80m1XkCOetfr5DJ/6M0
Vou5rqvbLbiDCYEX9nQYjocnX7fqV6C7MKhRv7kbnvsxCZosSS4vixUxbRcnbgY7HxW/YV1WJ04l
GrNMZkAXdAeyX/zHgZ6ni5eLDGTvGqBjjmjMh3VrtLEnZqYu0JXY9nZU6JgDjUd3xmB2xj/ag1DW
82W6FEueNdo4vnLuKX8P1QWMlizX88lIHvm/kWcVGsQCI1pHABlcrie5ohDYn2nGxABlNskn5jo9
GeavLB9Lrox1MVGH9LSOBc2EypG5n+pWzZ2VVFYooBmoa0Kw6SHQClRAszhNc+FACxqm39iO2EB0
C2j/gUGXUI4YjeHRKNpDlcI3Gmm6U9nmp1Y0FBD1QXt/SnX3//wwCRTZ3pPfw/9SZU2tvfXSPyAD
hZii+CfKU6r9odVRmW9f0+ZFgxu3dM3tN2+rvel9C+gT4Y8OxjjDosolk6JK3quicTkHCzkqF0Rn
Hkzsu+grwZmwqK6St7UHdJfuzz3USlKvvmFQ/vh8flvYq034BBydnghozaP28pZfzIbcsOsQz1JR
V5HkTgaltAcoPCFSI2kDXEQENCWJ4DpcDD5WM7zb0osAiFerllowG68oal1nWArb/bxFUwdKg/Gx
IpUdGwxKjrH8VdTDjm4YDDJi1trJt8bJIJJw9A6fDaZLUr+LLE3YAfacDr/W7blDK5OtaXy7eV8P
ve1yGEqXu255NfpGGqUrFfGrqMj/h5NIn4HcfKQQyAzaXDKQxX5DiRtu0OVMIp7BhGAgLBVbDEFO
tiA5GQAq8bT88/VhtOZANSHRcdhrffHeZBKIb1dTs17MtZnsY20Lby72uENFpgLhxaBrusP/lOKo
9LkwfvQvRAAjFHdLTG9S5ZTyZoYI7jV8LDNU/lSNLef7QYfHo9+s7cbdFk27Q78gOptjOUB+8dxe
9XBg/7YsVFKyLBnnurpn2j1prsfgQ1w+GVKgi8Ag4BPC9eiLEMTJFeggpY4rS63eDfk0h68KjMox
BQJHMzGsgg7B5e4sxptzhkDzzgm/peN42xVs1xNU43ngmhKmU4yHRy4+Rnws3LbzGQZcXUeA2jiL
VWlloYwZ755utmbTIqGP+G4u2Etd8PzEUs2GeTJNxiaIqQD7uZx7oEj3I0ilNsDAvCGrMa1Vu5kC
1tr2H1eg4IeG9VUUdP3eICNiy3lnFQwOGx7zt9LilVjbysZsqszyAeBE2EStbJbVr86ceeHnby5w
zpXboqK6mer32UV6L8n84HNRJkodWQzW3XLR7fAiaHa2/aODvX7lIGMtNU5BKlSh7Qr9pNRgEm8x
ZTL1pK+6J+hcOgVhknNLyerxBJdgsGRyINa/t6qf2ayqFbNZMPNxhTSJGDPjcA3qy4BbbZy22/Sa
86GJyzuDIgAJKIvfxiiER4RCGGu7/YTxOoxgCu7Jps/TXbsWndl+tICtMQHnG+DP4DkxTNaoxUed
ZQscnoB8lgjZFQ4HOsjN7GY4/mW4Pe4LufwDT9aRdJ5YxLiKVLwZCrHQBxvO+A8Ineyoa8v/oT65
Q0mAN65ulzrzciLUAE2u2dnpT8bUnnEjsCY7EgPVxy55HNR1tYqSY9fk5tGUuQkckgZ3+qZW+rbN
QJmE9B81HnNpBnbRDXT9lLWTshfa0izCfMSSJXsyynjzskwE5JOOjvCeqoVklMbkR9Mt7XkJsXRe
53HUwGMXfAMNR4J8/1tOcW617RA16rRonnM0hCYigoJQjOYIYb+giYxTqSVEwxl1vBFyM8141eal
x9Cd2HiqUS0URp0QYz7mrAMAJVnatO7RugNrKeEmUkRpS2l2LBzrLW160odW8OsW6NXOUyH3y9hy
TYwNMmll7LbyBnAZaTOKAoa4FWUBJAPpso4AjH+UhxjwsfNbtjhr2vz8uWnNa9fdxQVqKKcyqkKd
z6yDhvqqSvVieS84FSOlUKsahWgMzx01x9z8JLaiJoULditiQcS2V5yjK1zV8TAOZS0pG9Lhk7Er
VPLFwDMhDFF3xDPUumErgw9/etNrgFaqpYKa2NX8zes8qkFh+0S2fY8SF3RsmxZVLs9XKETwsXkD
900eg+D3UlpbsqDodGmEKzL2zeWYAeyonnmXBenOWbbv0TK6x4Et5/9yqlYIDVARI8gwM7wVVhrs
oNJ7t3XTnnJ0MDiHvmHguP1s5kGVUrTONiM9cdW+UOutCvoNE6ErpWGDKq7i48PqWYTGKaZpaN00
BPC8wLQ51AqQNRcJRI3HPBqDyzM5WEVa7zlwhtPMo+2Q2lTn2U7UkTpGC2TfLDVUMYlLTlNB2ce8
zp9f3oQupGrAXlV6jqUFpmS0KxJ4PDr9hxWDNqZIFYbEANp82A3C27NbJB5aLfnqBqJ2NO2tmRFy
a1nFQhfTUiUd46zhI/47fBjifIVfafdsqYjNQLCQAn5FddOE5qdTXym7qCsNK5vXJ2uc/VkZW0Gz
+RziYiuB/ACSOczstF7mK1gPLgySC6p/35UbdTa0nNg7Nx0Sx5AZFSLmSoo6RmOoirzQOsjM+2C8
gHLIOYcxQ7s8qH0IBvE5nye5S8FJxTddIxA0QRRTVCVFwmqq0YYCyPdrSVo132PK0Xcqk5fej3uK
fnt0aH+63kNI1ctN79ZrfOSmvk/HoJ7sX1D9TLVD1kWRLtuKM71rXnoOc8BhthUKxkK5eivShfPs
4AGOAZhEdVrxYuL9wijnOeMkf4mU8yJ4nZwA0NLTZWOotFzdaDPeVEvkzxlJQhJt9aRP5TQrIKMB
2Fu78Ugl5I0R3Sn2Z5PBON2FeipRUuCebZefqN8j9jp7WDss8YIgIFpJViNMCmsVPv+TOJCqfCqX
7KcGF9BdFkPKZe3l3Wh/yF9cWSTWT0sjbwJ/5XowCfM/V1yTjjxXZ4vdWzRqkWWASaknllBXlih7
Cn6Vy0DxF2v8J0Q+Fs1KW6+fqpJQNGhuSX+DpBJ378N9YMGlTyIVWnjPQWcjculCb0nx833FqlcU
5l/DWT/7M0lYi07xxlqEQ3OoU11lFnsVOall8Pj9gcLUvCyunFHrAnmp0x3xu0unIiYrZ49WQPr2
ggFvP4dRGZz5VLrjhdd1zFMb+ACyfCFec25DVABZOKRySNhIGzB4ZpenajsVWL6TYZR786dvoFMO
HG3m16DxAzm75MvQ0G9lMtNhOwX5reORX/TTnsrlovu/PAx27oNpyH23HTTNCFiWYIi7Fk+LEel7
/ZkRkLKMA19MvlIkje0BeaaMKFYOVHI7jnZWhVBGIvFiwutEESbrYfjJ0NkNc5c21KPqRNvsJi4B
jnBHo1Kt2TIb7Xk9CsJ+WuRghUAaPI0eZXyWpHLS+4Se8LtjSWWQ9Tfw/CQMdouw6EndSXF5uw0o
1jrM9My0fWXoXAaTFa2cCaG1rE6NyTWPXkb+0yOG4Gy43Jspynx3sRHK135t5hbzTerX/BgzQmkH
nz5p4H8GZCPbJjDdN/jieJnP+93zadga4zKhrVpq6AGcwU1LUNdGR6kc71UDtFtbH2HJsuJeEO8l
c1N57btmKsmYIiMfk18ihBB4HNH5m7oqKMDsqROGkychA/k/zI7eVsFW1WzwSLHtoCpR9CddDxJR
o3avuS6t3J3hOtokKwtqZ9/2rmHZlA6uxJhR+GdhtSwubv5toYvA01WLGWri8lap89+dFtYZd1Ji
H5y6l0oygRXjHHTZPENcsJlyJEX32PHngXW4PVY9mcknMUg60YR6535v5cY8zUDmf1jfBkbeSQnm
Yrdeu42saYFjB78yXH6kbwqmoC48lkC1kLqRQ/7DOv/SlNEYJVG//PQpcziTSN8wVcSw9yh4nBi/
TpML1rdIqJEUQjN8n09PcZT3d8+lel6nT1KwnMrpe05iBbB9G348iMyQLHDl9We1g3VKchq6kQ9H
l3U6cDDbZdrvrwrCZd5hY42RE1QbvWsmK6m2CtOGOsDBC3amjSgCT6bvatgLJdAg3+lNjg/rudOd
BYDJJnw8MCnK+uoqRe8+5pzOjBn257LvrV24ieg7aj8ucu/3Wdn3yviLgISpXddsjdWfCzrlZJjK
D+XJvfayydwpQooxJslNvbfyUZW4zOQqQIRtDtmyXc9Yc/z8d3nSMVemNJCY2QMzIMGNQMxguatI
ycVIl+Kxd25VhTmROO3e7b/cuNRtV4G4sYPRcVCfdD7sPFV6ULvTp6yA4aByhaHw3TksRzbTg2S4
O3xIX9XemXJktcu0pM6fwYUrAy12/4gwugQUwW+HjW4oKf0DwdJHslgFgMijBTBn834I/wolD2nN
9RsDTlo5dQn4jjGobHft3bWX9kSiy/njae/b2foVOJUw9WADejEoh3FujUxkgBAZQJdJhB9aEfPq
3foQHSoKoSFCVK6Ehq28FfUUOr26BeP4d9vvRruZKGjvm3U6WoWv56ARd62TVB5f9SUbbCeyfa2o
WvDbUPOMCVbiCkxBw/PClkNMFTM/U41u9uIFfB+3945oNOvicKMMvM2UEGXOK8NNcLMOTjgoJQiE
PEZx+raHwJs+Dl/RaN6L/NbhKz9jWpvfvZQl8Xnah7cFseFSL5L8Yan2zmcX/ijdVKKuJwBlWpaq
n0dyfE/+y/aKUds3H5xzxg1wfNLJWdDJbrh9maOnW51uXCDovnqvYXu3NSL/cmIklzxs15JBwjGh
pk0ySnjPGNSvZbGLla2mXwW8tF+hKHH5rIe6m1EGHwKc3q3RKneeXHaAoKkVIFSSFvUgH7RhaIxe
RE0aUjXr+aTCmsME6/eucy18SQF1ZoSVzucR8bOm9Jo1tPclE436wSm27WiH0dneuMUDo3yHrLFJ
zUoOS8qy/HvQ3su2BYxcZOhvEHHNfm0d4GwLFS6NINC/GEzdm5xId6IKi1BMu2QkY7RPlAwibbBJ
Wvht4Bcf6Gx7pF3UrL4xVLEDIM3205rQPF7Nd33Ykw2u63iJQID0cd04FOCcYFEsudnMI5wX0Pow
DNiqNeoA3alF7Vxx3v6J02sfXqcv3b1FGfs76CL9vBof5S4zh11T5c+3rIw5IKbZjNmRKda7uXlR
z24Vc4/K3sDhJ1RPFxUqZkxCvwj+w3gj2EoDRKTQwJQw2jmLJg04Vy35heS0JXFdVBRl5egD+f6G
MrYaP9ZcTLJjrbW0UuqWerrxNcGsMWOz9BBwXnIGJncwNgLJAIiw2poslrPy/J3tltjYgLxEFNZ2
Qb79FsgFdIQckWGPdwmn7jnZ2X+VH3/eQncTPWyJqh6ie2D4E8AwEHOrq0SCRKuExiMkCP/Ex/68
Cj2aWs1iQvqH7/h/niG8T8WcrCQUalsqtMdd3aiXYpIkCXpJbcRQ3rlL7LIH1Y9i+bBe8palMrFE
pFBqowdi96uYPK3VzhhTqFTaLizlVrJL8fu2pwRMuT9Yl5CCvADNi3UdGmoNKD2NF7SwZejrELiN
sBA/R5+jlRZR6SHXl/X8f7chZZfaX+mKw/wpKr6PfkJXHJTHM+l65C1orzXWoOgSQ9MFXiHUt1qO
haGXorhmcTKd6GqUgX2EsK6ZT+cmQdp2WC2YSBJtpeqs6tdNVgvjiBGrjOQ9B2udox3V54O5pWDI
m+lXyL0seqF9hsClmSmAh3k+vOa06kq7u4uciinMkBaGHagdUYi7wbF8n63IEoKCLK4TntLxZuke
lsgoVHlIkXjfN39+I3+xHh+aTYHjdO0hOxkuwQkdhtRNP5azEK6ClGCuFrZg021j7EzOiytrTDxK
dz1SUYbLhcCbIP48J2MSEk6+HBJMO9+/0jQIqk7VCMIvh56V8GPhwdywVE5jitqm5IOaRy7MjCGr
1/nlh6vTOxVWJrQs/tY251IO07u4bwZ0J+g/miW9lDn9oFa3NZx418efXJ9HCcuORPHFg3RDVrXB
p+tH8SIWRNKx2/sZMJ6vxt1w5lRkB6QbXYzHLQkEU7v7/TUECKnNfVMQDX1xMio8xHQohml4btDX
JorJERXhgwBViCE0PJgTvcP6nlwAaRDDnAgFuVIk5K7dIiD6nk8d9ZGyKQ5SJ9I9L105VdWHXO6Q
xrk/xndtTqEeZrQjSXEKhe2YBPHkS6OD+g21x0teHmCh2rkn3/2xxJsE1XfxnRbmsjGrsjy3p63w
yCwe4v32vhwNm5dVmmFDDm3Gu7Tc1dCaICK65j2pW9Uc7k5+Vr7KVNemWU0FIl/eDRgpwZSNv8So
+1u55fFp6YmBlNOyiyYPm6lUUo/7e2P6i7h3zNI3D+Vn1C0SaA/Y9hCJI24b8eZysDLFHAj9nPTh
q/lMjMTv6+KCE8wxfHYZKWIcCzWRFbaji/zbeIiPtG7CRC9W1FeettrDMe733nLQnmpmoyYboQr8
4p16JYlaah5ugKQTgmuQcs/u37CANlNSGVap8Cd7OEc9mN1tCifySORkfCBvVfShNG2/aZ/IVF59
NASZvYNSOINeYwq97MjtF5RP0GwwbF+6P/HrwuPfq/WrhwxDcle3GC99kkMRYM4Y5p2SicHClS8j
m3pH2UwMsH2JoRbqZBE9HZ0/DNVVcjO3PvVCPfGyyfTDk62a488Roe78LTtxcZSFToYHn+BEB5eF
DdYhQ4QURnwk3TLpErRauib+PChFV/Cpj6I9XWvGLzHUMlnNYmAc+hes9hIi8QzuPpCHcvZlOdwK
miR4IApMU1sVIIusSfoDLKXVbB5GajcUeNBy2Dp9ucL6UHArnTZQ/Fx3xRcBW4qwooNPJ74Cfvri
f93mLg/nk4NtvhbJ3zWmKNgZCehH93xrOGVCVPPkMpEZ0DIdxDR2LBVEy5dSJn3xalEfEAAIo3QA
13TioYLqnaYKd3JiirP+PaaHX+2+G8SCb1oZ8rkujhqpn//YwOQI/uXcKle2kvBEXp4Nk78kVz7V
qh9MGMowWJ5qn/T73nz5dctJsU6bbRoHdrhYRVwKI4N/yCZ3Z0LTcqIcsly9XJr5BNJumk0+jvdj
ZJU3WVgjHmvHJs4xYuJpu1Lb0ymv4UTmX+5+eK0DH6vqP7k7cgPPytY9U5dbDBDF+1dy0OnaD0/3
z1nix4lcOcqY+uEg/bWbxep405At9hSDX8vrpYrHBBxIvTm1NA9FL2kKKggc6m1wANuwzbRt8e4d
PoCw0w72xf2TZZc0yFFHHZ7NbF47I22HZDplSXBpRQIqT49U3ukMFgM2bbvN6yzsRMhO/FT4zaSw
x3wGzcF3Yf0OJhl3xG2UaNiVpG3SIYiuxsOxwrOBM5g40/Nf1m16ZDPpgzN1uOYsB66FLcfCiaDs
ZK3xDbWdIbd9oj8YNrVe+FRTB4koGrh3ZBJUGpzOG77FZnbpE7c6wyvURV6FNMXp8NeizNV4WqIl
kU8OUtpTjYUIjZ/U+wRR/iZrj33zt7BCYWT4f+7TycrEjhB55yaBvv+XppsmtKtbnebQqBXlxnCF
2oFBImFGXeJMArMnuEk7V9iZ07aup/IJwaHb0BPzFsH00SKI/AzLA3XmpI/oPod0i4m7fbig2puH
5UwxwZNO5iKLWjD0lvMQYikKOsv2Rd6Byz3WifXHzpmj8bWLiuqd5se0fkRdRexBX6gIyQTRKZUN
mpWdoYT3kpqO4Cqe2yWnNWUVpfN/eP9dqCBx01zyRp7CjhP+3y2DTSFam7MdPajBBxv2oouI6E+y
OWd991ur6skykc/hooOInQ21OIhCAZP9C9qqtIwxgI6XYF2JWGKb1fdAmbX6JaJAJz9rehc8L7c5
3AcwnbiziAUoKt+J/F2xhADnWXLQbOuVGwV5nJJmfLUx1Qz0fkB6vHujmtYLB6F5xR/3xRRZ/QiZ
czhx+FUA5Dkp03/45dOvY9nn3ScOw36muh89EL4v28Tp9WSpyOl5wfIYGWAb6kgOifRrA1oXlwN5
LqjRYNw3lfON8qxQDh6PaNsm8pZzSe8AgCFQRH4QWS5HSBym2gaJBb5y0AfT9colisT6E9D41wJP
py8tYol23rkwA4DsoZRWLWHowotBdDiydQZRiHRv3S4JBWoh/B/FIvQIqx/SAqBEuad//bo8uGxE
O8u/FY3S31w9ZVv4X1l7xNhGPS9BylykYv9ECFHEVhlFjCmhEqDTIVdSyh68vrfEPeB0imB53ULS
mgiDkZtJWRQepi2FN5QtDTzqVlNjJgzE8ALjnqAAzZ4rLbJPcCFygCM0NSE6T620J0SQBPkyp5na
41xqrV/rYs3TIUcwUBOyoy53GKO4TvE73RFC+AsZ1iDfb0jDD9ZnnrMx/ik3ivDbU9+irE9N//8A
G/g+Lqa9QiKkPZBBooVolNTV7RLP5pNWEGLdklQYh0HPHrF013ZdLWWJC9Ar2VvFSmTJyYoMf1jq
Y+N+iIm1DPUUmiCBZZDw6hxDyi61cT9R7kRsniJFOiftyvWeLvmD3AJ2e0OeJUifrEBb9umafHaH
Fi3AvxRySLu6Dwxn5PTApX+/SOe2vb2/ppBvhIwFtRjOjHNXzDEzNMIqcjZtpdlYJNu2thZZNE/w
bTwz+7D2eu7KMlXuUX7dx7pT9iDluIXdDYecvcbOOuhJvavGAbe/fSx36gl9z6J4p+pJgEhkp6eG
viAdc8Kx6C8kDlK+bF/NReQtPx+DKtaSL2ei6CDOcQXcJWSw+k11GIYkzry+9OJOTxckIAd75uZb
l2CsMVvMeyia7tx0wJVCMB+Cgd7ZLTuWNOWGJ3/OaQlsXCaQdaYY4Gd5ZHbk0F/JWRHOk1TlxKv9
ZTk/sNCqEt2tRpOnn+5F5/hqy5vuiHwdJzuOrzgbvyfEkbyVwMy6hyVsj9bAUh9sx2w93zNFSu8O
fqNFspZAYokWVG1I1CMKTEOAJHAwYbQI+Ch4Tj+Ub8R3aSMYgyftlGxyp6I6JNbro8hJ2XB3wHUM
IueWzc/52CBL9zYFG/22hrOrIsTiR2275C24rOYOrAejqEksovUxpq15e4QaVANm5l2G7YMmoikP
2yGE1PVZrk1nexR7q3vkYrlWZj/4vaxHVtbTXoOd1T2GNbRDLP8uShgJUoSU9CePDvrz4X9ur+3c
gesRqWLeXCF/utE9kFLSoxPTKecKxneCm76mVuYdtW1Cq7/HYJk662pBOVrGS8u5lhEw+9JxAMXm
tTd6x4MNreqDxxrd4Jdv6pK/EIo9uBHcWosS45uURnxyjVL0jthuDAzj1hRy+gV+4hsdxbV5buiK
G+MctkbtMUpllZfpNvFiMf5tWPacY+iH9oiZwMezezekhs2sUnzLPAYXG3iTJW01BJtFKCkmNsXz
5+KS60LB/uEFU1TP0sqtd676js5XxoQ1wNNR7kyScIWluTHkxEoIzVQtn7as7bbR9AQAwwStm/iF
21lWgxl4HRNxCFr9jJgKs3bkZ45TRJbzSgA4CAgNvkZAzEq/Zyaeq+rXYvU4NBvcwv4qOZ/isDv0
hNu/LVgSV2+yFvwTrw4pTlRVILL+TnZc1TVXTDuQjJfaNTxnSI5ND1FZncHgeLCRJkjJKPgKiQwS
bIy3vPZuKUysHqXrWs0raP1uHzXrO2cS80gV/jHfGZSvI0ET+6XzXW2P5XktpNhL2si53jnkiHgE
/Yh+QJhHxqA61NBKfYwNHwbwQK/snCcKxEooVeWBC4X8fUJH3HmpQIJizTO83RteNSbVVCjbiyLd
2xWKC6noR5j57dc6xMQQ1Lz5q/MhEyrxRV1dL+pLBBEhgE7NzJVMEVE38OWQIX+o7KfrsVflbRPR
jOTU2o90ObjmdUtNDCcOOgkpANFt6D5eoxQPs/+VXJaUPKlYWTOBkPyvJGuR9LWuiO4cpLWjQp0X
xCSDVabHRyD0yqeObC40mbI9W1we89xwazbHj2jCppYlL7HgQ8wvwKdUvh04PagbYJ7DIZ2wwIaT
yTstVfhI12yoH/ciuKs2Z7374TdSv41VM4XGYct5J/qzJcUdo+eCrq78NeBz/mvlJ5KwN0nSIEu3
d66tz9mjCQnq8ROjrzje4KePjfFFWAdcbQk+dH6gesWyTy5j/xwwhp5J/Hz3vC18G4RS1wUYOJVW
eZxd2dKEof5eYYFeJm7DkOVUtyCnum3F59d40T3SW0geJO8vKtzV1E6hKbWlsFIdlNedde4TQw4W
FEloFM52XkTfGJbHDL96z4VKQmjxHw6gzdC55NI1oOew4Km1prU5ssXWsa/grgV3YFCChwIuPC98
COBnngu1Qzl54m+ZgyU4/qQYjjOGe9GsrSSBqACal0cwEVfo1kkM2/o0xkIVR6ML4LXcBTxaGxmw
I2cbk0jZehKACYJ9C+sK4hMT/reLvVz1ohAtCwjM+d6hM2HBNPPt8Xjf+N607Bx8uWodTAI2Y9s5
35BblYOoLko9veZFWHOWlzvqeFG3ihrgnhnNV4IDf7YqPFhe6PxEG+37yomMq+uQQ/bPpUc4j7lm
tIQmAhKTqTq90xOskiJ4FOcWeVaI8Fb4G4K7BZDueTM/NtTm/zGBjPMlOnx1neJQEAK73i5Qclhw
PK6zsBr/xmDDfXc8BGgz63qlcRKu/1BZ0+Z1PtN3zUBzW/EAmedHK6paj2GBL4BgSM3Rg4Ojglvb
tVs+BcXo22Qq5rfbBj7VwMpvNUDqScPzVCOmVbACCQl6XhhD3fS0gYHNukBgNd7O6HaIv7Vd6tEU
3ZFKvtrO++CxSpEDznMh3JWBP6DNgamBIiPpxMUOcUh1sqt3W44U6xOQOtAWp7vWANxqACzpYHxl
EOSkNUg4ceQctsUxIxgf/dT8iXy3uKgEpmy7+bUc4CNM9N0NPz9tctg5GQWVCLw2dKkOlpE2ImUt
1lDDcdOSmyecy85ix1wUrKEaj3O6A6FqJwq9SP218TeerPx4hdNxVWyjAS9FJ9htc6dzadBnbPTs
0iwlp6UjrVwk5+7wZxocmBJIQoOarzsH06BMKfGw1IMSrsQi6aOxBkHgZsnPfdrU/HUzFOf40s3x
bdJo8M+lelUVsT/BrBQ2JuMxzQqQtIVqfwditap376hAwwD5Cv/8E815k6dpuMdJ7Om3szKhW1Hs
r/QTSRQhjlgjqzJhqHonSBgEDSJER3IhdEn8NRovDp4AZIicMNtT/nPAukFPMoqJpgk5AJbZSyqg
Nq/LRHpkmsnffU03BnWjPWh9WpoGRQysURURUrcgaJMJwVu132yQI4+kM/U0T/MonBuk0MvDjQUi
d3PMfyoWoqgOwyJq39ynQSanhr2xctxK8BdHynqgJ2QCn9BE2jU/Ca34ziL+VZk3nG97TQAVLcMx
Yyg7sZM2p6cB6Ehfj4UT7L4ZcVK5UvE5SXMNXZ+HLbiyt5gNJZPlr2ouoRi8OQ10Lz3hUSPBV1nR
PcgBr8cgWQebJFqAyS4Fn9AcNdExokyOP5KYAIoBvH1b/+uWUgsnLqpxpuu+X2H8cwjnk8yUVAjC
23q9C+ns8nKn2NjjWok3m9PIkkF926dkNvQcprjGivk7tzbYeMSVaDm71UAxNE0R2MO2jGhoQ1ax
XX8uEwHv3m/HeHx/3B/KjIRQrDG4QNertKdkz/IPG2IG2AzSO457EmNNE2cQ1RJpVGAWSE0OyMI6
eRrzLzb6JSYrDNORUq5xqTx5iE7TDHcMtLTyMBh71amt1ViTLDm6GC5VZnEI5jLMEJWMZB3p4Ug3
v7/ZFq8hCIiSegIPgVHYJEOL4OAaZhmL2clsnFlnc3GiZ1aoHSo7szssjznb5EaJZ8FWrUDcr1mo
cpjj8iLxqfFimaObPX/Wkn+rugLMNlk7KY7xoxUNSJPdP7GuwOrUF1tQQJFTp1CSOlAcaPUjHPoB
5CctEIjiXArjAI5mNOMvzJ4EU/3vPKlrSfnIMevgj3o8dLtBYtaCASbW7fht5jElrq8+PYnmsVLN
XmvWO73G70W7GEW8HFnur9bFI4OxV7mb4pTb0YWyQBNj/g5wrnCRfaB2uq9ysahN6EU8KyVEsqKJ
xvLnpRwQaJAo0LhT+cJEEKawv+yBBPymm776VtiwtdexIx6FsnrA03adATY3oJwNumGc4yR/jx3Z
IX8NjLZxKvpLvvxDl9vwybuwlFarncrl9LmADd3mr44RWVXFBH/5tuYQzNohFg0qnPNbyqncADTp
nNXz4SAmpjy/JhEuXVrgpKnTNaaOkyZGXxT2mrpABF1OS0n6kkFp+/HssOV7C+urU0IFHzEhs08G
l8wZzndRXZMMYXXMIfm4rOjdwHn7Ewm/rr9wJEsCeW2cYOSuklw6kLbE4Fe0QVUppxKADFli6NtO
35MtqFWBq8wMeuJfdTytdXCORG6K24LbHDZq7HYrm04VT1mymIOL8LlRvhGmCh4G8FviMbvlwiHu
eRXJuijTKyVWl1UMte/Yu1gCaTonSpe3EXVbYLd6zYcEejI6PTxLLYkycyuc41qKTXsTWjBKD7na
1XUKquX4rPinaHsM8wtlafSyJfbcdtSY9TkDqBFrPpddeL7DtlC9IjpkgWf22g/4lcd+w7UJM569
MoLrFTfSvCB8KrEu2DoAQkFI7NdoeTQqxTd+BfKZMNT+ENx0F7Tcrk4FGQ57832JNRzIM5e2cU1B
HZhji0VmtJvGNkpzf/UL5CQADMGS4RKOGbdgbxNbf/sjeB8PriUSA0dVfoeTdTWa1oq1XtSAtJrF
mcuCKyKPgPnzBcqoSv0nrnQ2zMff7e1wt/Is6RBigWIofi/Q0MwI/Ki/kpRw5acE3gIxtdpngE2n
S8Hr/j1+RdJpemKofr3AUe34z+RyfH1KNMXXBmqvYTiCZwyutfDmc6uRo+1ivaqtFQXgB74uqJ/s
Et9cFGczkyTrFsqSYsVDnoqeFg/9uimzS1RWldenbxrItGXhinBmK2D7Jvd3mgNF9FXxNQv8rWxw
LtntaeXHmwaVkjtiRpkWjXBXm917WN5F0AWm0+ya6l7E+228aKLKJ62GAKckxyt5Ng/JAL2NQZO2
D2kdIq3MOG2UoHI8SBxM9h1nmIB2Z2yJm4MXwG0dfcpqOPQhCLouW2uSDzXjh0eKil3/sOwAFI8O
qRR/Twy5lIS+bOOE3vddj7stjetJI+Svz16E8GcUWEy0fP0XkIkvwGSgvaUy7RSJV1azQpT6RfDy
WZinzdgFKp1RR8SEV725qpYkOAC//ur9tauzGTCiN62U+YXhK8MgcHbH50DbEszEjZXhU5DiKXLv
uvVdLuUME8a/wE03QmOGUyoPm1Phcrkv7bs3r7thiYy9LPRw0F0LhD6dKWCSaeNgx1a0rDrsvSf8
EK7xjNUkEdubNYHhOIowSFKRU/Yt8XLY+RGQLa5PoyoTnA2OGsiOgf0biCOpQHgYaSa2kwLnB7ny
DVupWqIrki+/yw+ymvLLdU7TJrHfIQRWroVR8rXeh5+ul5XapJ5yo9xJqKGhAZnTVoDiux1naSat
FDK2ThNE4dioQOq/p/vQm7ql6whfil6uB9bqHfgG+c9znss7z1wfm6w65N6go2g9VN6iISTmKYeB
6Fil/anhxVAsL8KXJq5dLp3YjDjFPosXT2d/qgZ1enzlmXdhcnTck3IZI2poR5QI469k8KHltFsA
1fXjQYqRceCfnFju1/Isvag8W1k5EobhD1jA/lcn7m5nyL5sJKf0jv74WYso8bSBceIsO3/UEDR8
w7l3tNPTtf1G6tcfQ2QvmORFZWD+sMeNMY3iyjcv+nMpwtT0kEB7CcoJnIxpElUMp+skCv+BeTF1
tUmMhnswKZ9anYUIDZ8Kbop3CCSZ53vkeCEJLclhhKYnRabJGvobuLZ0sAryTDzZwivqaOSAx+VR
byZc0b4r4lgty3w0VWvjr1WYzoDDzU6FgE08ICDyJ2SrkzhVjul/lfsIx6CnoXkKkZdmduqVohOW
55IuJUmypqa9+VT4RT89km1thbiUnJRhWGNoqCDe7VaI4zJlovgi4nSmSds2nrfuXLDYttsEYKSW
noqv6y2AX4nl9fY0yYUz9wkI0kynoCIfLgjjsm2IuzxgNMt3GcUMHLbxlVoV9/J2TLjlvRKI6zPe
umJrGG05H++vxsQfuWIXEmRJ5goiWgLh1A5QDkChC5P55jvYRaBEtGCTpSb+vRPapzV2UuxvAuQx
Wnwy5KjqGoX/eeuaMghI2wyRy029PooDEPRBzj9OUGP+EYY/5JcoQXNh2KMthbEYW9yC/3LRvmIA
GStwiagpjbaYen1oVGkcLtTZ43fMmWSwYES2sE7m8IFJfELCkr6joUHth4bqQvO+a8aKEQptvJYF
zSCpxroUvx1bpJ4Xf5Q19oIzTxfm2rqtkDtR7FDPo4U+JDqwlwhxRvp0VSU+

`protect end_protected
