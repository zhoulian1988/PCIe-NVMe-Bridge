`protect begin_protected
`protect version=1
`protect encrypt_agent="FMSH Encrypt Tool"
`protect encrypt_agent_info="FMSH Encrypt Version 1.0"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2017_05", key_method="rsa"
`protect key_block
u8UbeCdmNCeva/tApe0aKx/Q2fUL8oiA50PzgNF0iH4e2CZsOQXfJEakqQYwQ2ZsrZmBKgwx2OTk
xFHcxHHWANMpbN3StBrNoifSJ+e95fOZXCTCkg+UwCF4KVCUrVnTB7exTmzpUURd/wcq0CX3XNVR
LD98vnyJ8zRoayyl/wh1gw8MGxmjkfVwtyOZlsOTBcfIFxjv6/7/mLvaMeCmoz9h3SymEqP3h1L5
sFZotTik1fj/BLiHSvEXYbn4GhJo8V3yuUhN4ieG4uUM6KtGoaGqHm05WDM2WNKw/77Wg5UzHtO6
v0oe5+rbjMtHd5/hGzhsaqo5SBLLRBIKxI2ulw==

`protect data_method="aes256-cbc"
`protect encoding=(enctype="base64", line_length=76, bytes=26688)
`protect data_block
psEHpTuVKibKqhbkrbNFim+/KOnFVD/0gR4kJV6Nz4sjtr4Hm+Pt8LjAKYZ+PZ2ZCpONT7HyqOpN
6+AlRPV1ZhZEt9hWa+0DUPdPVMOMQBStbWjxq07y3ea+23gzaIOJqjUBHw3y2GlHIx+A8TuWFQ1O
xtceQ7xU8kGy4hpr9CEB5N5Lgu7wUFlwZSzTDAFfMk744PZLGrW+wFp3nZHcLxHhU/WRsztb2dgM
r+ZbK3Cj22akY5BrSuM3yRWYG5kLJkzLKqn7v4PZwkYy7TEBYfRpfkYOFlUe58LOFUG1gKH4qI8o
IZaZiEqReI17Zasbhy7NEp6qJWhpeOM+v2s9jvqCCR2bfgDPa5bkSuQ2vv2aRPyrkd8UY6XypLcH
msd7xexP5MUNdfWsHiDlYXChslpVaaZ6+csn02q5DnSRuO+2HRMYxWhMpsM5VyEGsdvkPQZPOAkw
ILAIOgB1VGpri1yRyTht724V29SU84v39LoBQmHNIbLNXaPxUM2OFwOdOTdo1LQqz78HQM4j7/EG
geyLMZib6rNjDZ6FxKFcc9G1L2pgQO7xnc0vDsHx5LVM11zU4sSAVptXSnKqQYGfdCS04okj30XK
sDXfz5ZnXU9d1DMaS4Uwhs+0yiNs8ONky6xKteabupIPRidETgpShFkF8c5ihHU9n66E4TJwbQZ8
lY1GVMeiT/ZyW4CVcqKh++yFYJgyvddbWpNnJQrv/bOVK+qvwn+XoMxKGlCvrl45RdNXmJVgIocK
PEMtpXXbAX8OotdNrXc6jsKKu7icZwLSe47NBer5uvuzEFG+CBRrrb7qwM9DroDoH6g5UmFUCeW1
9l5z+bf2y68aSB69KGNlmP2slCmmu46GNxKOPCFYPdjAVlXAgptFCDgtjrXjjyV6UeQG4eSBvceY
ZvAUs9gKyfl7SvH/Vc98WIxfFgjH04WlTwm4pHPy6xzd9hQGc5PtAJ/pvj7bleXKQWRAOrsSwidU
cwE0XXryXwgASdXSijrPfRMTsyfpU61kKFbWWxv1Cy1wYAI35V8g4IabJbMgjUOw6tE901WnH2+g
Tpy9DxmGzR3VsZG16CIRV6qnmZZzp6gb5JmJ+LCm62Hlonrqm8DdjQz8KxKXaXHziTvF40RK3HHn
2mAuQoB+1+wyQxQ2JnsekJRZ1Fr7CO6Y0spO78wzryAhkpUPCZxo6kogusnSi0uTkUHyKHrSnDSy
zpoVYdb817bnCqlD3TxVJkO8gbbdmfe5eajxCnnh1Q4vs3aSD4+/K3ynfWafPjR31lD10Y0l8OTC
wGaKy3Iz15sH+WstV5yCb801XdGFod+tb7TMu88FTdFZKcd5o6QsDg3N/caGgAJHXMQV8O9IwM5A
WodrtiAmCcYsN7U5LAOUXwqXGGmKAcvh+OFV6UY6T4EJs9PEkrPayTzV40wQuEXm9TiUVrP2LujU
7Za+reQXOmjShq2vk41vudUl3aBfXVhoz4U65nabRPX9HEXb4DCaQY8RQ5k37Yi9vuibD1TXKdci
ERXvBdVwSdju91vDGIw5PveKFSNuE79+klfoboSKuI2yjxlphgoZts1gBLEMtAxVJIDoyXiNIm93
LXcSNJjfZWZdUPfbQ5R3ADnrS6+pjESsjuCE7ZWIuRzHQNwywLVQ1z/jhyFjAHUe/DHp+jqYAxsX
OuQj0RMVBw8mrdi791Fsuw/1N0HGvaAE6BnDE6fG63V2WfcaEfijO6lCmNShsermdrHGq2r8Vr4a
RuH53+49NQAL3jWKXmm5Gih/3yiWvuo0c0eWlM5ijilHEmBWQiqH7kRlqPN+yjj1lAY+0KwD36V1
JANCLr1c81Cm0bxsDDgOImx5hAXhVqyqQks2KrfuSUHmuHtNCl/oxXn437ed3i0GbIkd1IZIQQR9
KTz//Zb0COZpiRpZF3vWUhiCrq2yHHbb0jRLNCUH5kzXbJioemMG5L8z0r6iJ70Wqzx5/GixsATl
hIy+3dZFuB5MOwxYyTnBfzgMNbMak1Y84Ke5+GaUam8SmMCb5LjOCaLfdw3uGs6nTUxX/oNUMuIu
py5mrvFgb7khPDkAYB7C9Meh+Yp5YYYEjuWZaO/OBXgBDUVd+pgu/w9KtZEgYtgIpl/tdD6SGhyG
+039cM5gT/VtNE/e/hR+3WoiNa1YIgQyYRYuIVTb5w3+QbrJOWEGiccJKpfP3FbmtRdTsgy5qnel
jGXQnB7B/hZykaYTTfpwNaxeCGOb3K/6JfTD8WljrPLMPhT2IVWJ+RjkVJkxoB2Re1ObkT3STgek
zH4GmVefUP/5/qLbT/FYe4S98bkWYIm47j/ner4k8BRkTCaT4De6dbi0KZQgKeggrBJrsK3FL37m
/2HMVxR8Q1b5uXsDvQdmEyQG1Uu2rfHY4NVd8nVfRPpxZ55ijJhEiRCuIjGs1g9K0d3JcbfCtxvA
ufIM/fvDBBigXOTYbq6WYZom9grMJwHOzBtLLcIcf0nEpDQHoieF0G2SoHDOJLIe4cIG8DnQI1cW
H/QxrV9g8p2p1JWTSKlC/Fbo2+0hGN3G8uBW7L0+iqo21Wd80D/qCB3ViqLR6tAEdCLr/83cKc/d
uk/zB8Ge1bmlpcIT1oEDTAngukJNpKKFznCqBSNTzid8VDNEiyU46u1L8iTZnXu5flbZxi0zxxTE
/OoPseMz6EgfQh7DtrdvXx4HbTWonKNpX1aGqwECugyaOmJ0/+wIox7opiR0f1yZlRtQeMDRN0uy
0Z1b1tMBnv4l59587Sx1/3fz75UH6MkSIHZTS4OOKiG/ZGhzS85oe1pr4Adb7hhOeKlN4tZHBq7D
/4PiQYp/WKNMVFToRyFqZ/iC+KJITASYlDM73APNBy5CtJEhtU4jbboSFegOZgRI9dj+bmksTL1v
vxr8VFjVT1jA4xlJjY2HDK0TIGyzkn9dvQkhI++iG/bG5b99D9cWSNXNRQBYBOZf6vgrRqaeF4ej
ZzHs/RKtaTci1q+mpnjnGXckZS8E868FplmZFzxjOUK8NFaxGBdhYw3hQZ0Jk4uoFkxpJgxHeNmI
YLP7E4KojlHaQ13vDk7aix0Td9y/yzEDPNBkKEEdXlpR0Gnrzo25/d/fgI9K1KH5Mcfu430IzwIi
kqBjk2PYCxcp93hs4diAv3AcNeBJSjgPdDpfwY5gDOiGo+hUxsXv4STzasRkU1mMQdoArB54WhNi
590H51V7I9Ee0CHhnajVDUpCS4fjW5vOzCNoPR4rSrbtxf+ZGG0IkYC3FnCP/HXyyznQ/GUBE7hQ
dPMBWmHZLoXJ5kTB027hg08C/DjBDD1YnUAItEGMw1N8vtYv7VNrF9k/OPmHRZkWeB4gcqyHEjaA
g+f7CU6mKwB5iusOC4pOypHdFlFbeB5oy0VZ6TB0//vnhoVPQEETcaEIkWeeSYZGBzQBD1XfJnTi
Lao47vlDu8BUL3tLnkqQpXmy1miKMOJbTHUQ98Qa4GM0CASmzpy1AuiEe6Q0ETqug7UiMuoo3bKf
GPWhjwAYk5TAyKs894x4NemNnIkwd7Hvvpj18xbB4+JQK28BPrMxzX9EVm61KyI/KBpbPT15wDaN
HlqURDqjQ0gahtxNmyhktGKxZqVLaHs3rVFbu52Wc5qjjLVEymA9POzA2ej+u6DClK7TQmINbHmR
tq1W3GnxdETlq0O0UyBCgP83HrqfJv0DkZ97CzPE5SEE1rMMjYQylNWtUn9Brx8q1Hdmf/3WKK9L
WJJPUcpye3+BWwq+cU68Sto6r/g1Z+BJTg+oSdJAmgDSoljdzqJb6rX16E/rWjYKcmjK00+IO3Yr
5XOS93HOY3i/PXgVAcwIf0Ll1mCDtD2VgGD2W2ioarr6+GKEAdnAdZN3pOAtwpmzKGhZ3Y1mpnhO
zoZuaWkURG9/620Nw9uGdTg8/roAzM0Cdy5TmV2otdQJAmgJbV7Jf5u9vGgPxqAwa7xB0MvPQa6A
CBzfa7qyRcBbNZayNHpHoNubl+qmAyChBe1LJ9CYGvLyl6ybSUdtVE/e+Y4w9Pk6RmE56/a0sxpc
Ffv3DA2KC8Fa8J/xzWlqCnS58JTTWKKxPNKjbQHjWyUuu9Q+OO2dwFDN6xpBIJKvYFnEWmAg4Urv
eflGWv+C4QDwg6lnXJYBF6rIt3yfTHB/q/U/TWOhMMts9Nw64Jx+k1F46LMpbaOzCQaLeMEGy/qt
JdZ52ZGDARXY0EwaiS+tQEcLrQgXLuLry/wEMTNWu3vgbm90Obo1e/xSd4uPYjymIItTQLMz8FtJ
digjvb36McU1+CMflebWdhQwJhK2m2bO4B36JYKq72SDkOfMN2/igtOmqQ6JfjzhWYS5hcVrMRkY
Jr55Sq4G5JR330WA9SphcTlDX1D9sNC7fiRfODS5krvbmHUNflz3xnzRoMnbKgLEG2hmCaTV0X30
XEpFKGct9CT3gaq7ll52obZbgVD/CXcCp6PQo7hvFDMO5R+Y0fPUkNgM/H/yZBazvoAjvMI9xlCu
fgQXYk+gQwtap99nVUrt0JvTawLNsLfriFPxVkUiylRnVA7EzLjIHjxIMUa/WmJzVM8wX6L1Nr4h
LxNNvRiRPcBMgvGCD9U1MQTnf+DyWZPJidFIE6U9piv4AzdRW2+YN3hm1szbKaJJU00orTzXAJ18
0cbLd5g7KxTHRRul60qcTR29GEOoiDV9c2daS76In9UrUPODYTv/RAumLWoJClwdv+KMvNGWQp64
BnVyIYTEfCYeLwisq6RG8AkiRFMsToj+UjXlHNoUF120wahX/ao3RAn9X4cgyVQydFMolf9qJcxv
dUUOVcG/93Tq8tWQeuEsJ89DmIzpL2Mv1z7h6dHnqiD8lMucpc+27LE4NuEgMWBB43J2isjBPqZn
r57YQAm/OAekDxyFN+xpPctWaF3zppLFuvu+n4YiA/Dwd7YejhlulrWCPTHaK3mhp+OSLHmS5MnE
xsl5vWiVflNYLDeCLQe6fgrRKcfojRa+z3IcLM0avruAwjC6Rv4KNCBuGsOelNTv8steY0QXQAcs
bl3YsuMebYc+u7fprWFFCSnftkuSMC6LZWC8iH+oFq9KMacJGfsXptLEtju/xVz4ECaSr4VO9uUt
1SxGiurLaZuFJqhDHr0XTz4kBmsArgczWrdll7LfEq8JAQccfzVl2cpKar8BmX1LYsXI2QQ/2VH7
IGbIBCi3iX0rNNDH7AM51BMGZjDtROn9SzI+ygrlucEA1wuvVkYlj1U5bpSYB+oHwzpFqFH9dKnr
4cD6bFzZn+gWKrTvvAvsrPPFZQPsbKo6Jaf1cV/4tqvaQEVumKJqwdRrZPS6Ej8d+K29U5A5mEOc
SL0D9r19ric9eGumrdB3154O5NDrcQ3/hUJj7CKFig9w6BxnROanvMvqnUvxcg8hWJJHrl3mwKO2
i0bIat5sa+WSkoWYRAIMpczDahfXgUtoU145vjY3vaCGOhtZ38EynCrjH+yFistLGnB8ZxGaz9W3
WBxJiGNiswjK0cL6yPCZG3RQfX+OR1pZUScE4J/+2Mt2ftpJYZSxEOZ13gFDc4vzbTRElQtuyUDN
Ss1ou1tmS8Z7v/M8DTc6RMqs3qSoM7xrIFZl1GFGTZ8DgZfIArdIbAszM6ZBaVAcip0WHjsC6ZM8
ht9HFOe4xuuTJ7PBPogEtUs/yNDKufUrht1QgN6ZHXeW5SNYfxPB9LoMGPlX+/RQIRCKkaFr3jkE
hYMTZJrSdZUKfLeV9ZZk7jeIiC1z8vPlerW1f57Ip4jETmsCGqnl7CHIXXG+4C8CUcfItmUPEdtI
lzLEqY0j7q9azMQug494T19+aRq6tg2EWBJzmSDQ/og7uU9zaMSqAxxrVdWLrc3VK97Thm1KdrEb
n0m30MURadCb+YX19Cc+ZO67yR2pWGvIc0wkB3OlCNVZQKSCWsyWGO99xgA9XyIUjchAduDu2FLw
bTtLwQugAgUJg5K90TEM4AlpBMZBFxG7QZNrlKWF02zA9nB+d88Xu61zZb0u9J9xkNgcsB6n5lAq
IWHIsHgFlCEca7geGQM05gjfU6nwyWVGJ+rXVaKtDJlPEdlIGf7Ai5ZN3lkM8huuGWbtyPKMUl8/
cXTuIKiYU8EDH7+ofTPa8uOraxiWsFcFC+OfuDEIUqvvX0M8VcmLEV2MQxi47vTgcnlj22v9ePbo
wE+F3ornCjgCBETNdGfG1UqOduuSdpFRdgmjcF/uX8Rt2HZAL6ljnaMV67H7Cn1SQCvTVJdTQbxB
eL2KiCuaPISa4bUUpMquTGM6xEHgc2rDKYYErormWy+s7IlTcOlgnVy1I6nGvMr3ZiGtUjsTAOCC
XZOhaIxGCgcp71x3T/FuEG0ZZFKFiHDYCyWBbxslCJnJx09ygzarchsUxQ12KlxP/oOQvyZsfzYx
fcOVLvWlVSVKKHjRmyvNqfYfI7XuRoojs289Gp7P3SE/ebo1kK3pdw5fZCnWIbmgTBYZvHjPlwoZ
VFTRifx5jJdqalwLse0MGRLnp2oCjDQddid7dDEH1mT1iCESRrsT5Ztgb3xECSXZOai/7R7IyxmY
ZGJGnFUGjIWYuVaGksHCWouD7UhiR5ZIq5OoabrWhe6OnrAfP+A/V8d7DA1pqj50Cv6kzPrk228P
c2sQDYZIKLWQ5VLdClybgoxVrcuZxEOkJoVDSpliW2cAGUmNzJz9NAFxdFu70NF89jkzPnpIxpPl
otvw+0Dc5kqRr8BPxQRKQRbAnGEjtIcPIFW5m9+J0Dtin374G7flMCTfNAPJANyVNs5wbui/wHbQ
6Y+6Qwp3K3fRIHiuoHbOXuiR5qbJKnMxrDWgWwIULuBwi2UbmUBAWaYeJtys7tddzL9Tv5fWEM4q
qLSysec3ZZ0KYy2EBSyQ4AAfCYaLsWVFWLvoPBng755hLtBKfQDAYLrAA11wb8rCpTSc7ehUa7dm
1wKMFDAo9ohV/nbKsN3FbhsFueu2e57V+XBGld+cz0FbTjh5rHxWXwRS2lYoLoFGwFa9JFxmCPOe
rXwRP3rXmUtlZwaI3zvgCq0H8DwvlooBj3GYqaYRlENKAcaGJ8yoovVt7Lmh5LHZg9oSwfBPFFD/
XwL9yqt5ffqBjwpSg0kMKhwbP4pf1m/uRnp/HgKPrMWXHIcGIzTZ7IrUDhMz/2cFF8FKbj39RIU/
ysBI7HRiAjWEmgsih07bx7KzuTkDT7aMOfqn0i9K71uiO9p8C+eZJ9OVBR+oRzDrrj/21kjTcfWI
x2boxW8cKF862EyUd5y4Rau6V0y859inuMrQwzBKe8BReEt3OTxZcSVOeeKvEZF1m60gxeWls5Xw
PgyvZh5RajpkbcShx4KuhGO24xEPirTNIZsmdPB4RBAM0Sh6owZZ/09YvRD8V/hiTqIdk0uUXucV
H+PCT1fuW/dfS3fw3FYnhfmjtnEp8QGLMKdszNTmQILNiSgvh4JUt4uGneUtANd//yByTirG1KAF
rlgZtMChFvknpOmkEZemFzfCNU0OA9wf1jEkyttYs0Yfve64N1zdoSZz0d+OTfXJnZB93JeZv7eE
vdQajbpkTOdiWz8YI4czeWQ89XSOP4//CzCf4fz6BO3ZT31l6MTHzGyEZAcnGMkXSOCL21TFbhDW
V1fbDueiNClUQhsz3Y3xaOXkzVGX/w70vp7zTbJt6RKD1ldzdfJXf5YrewA5ZNsy44U+1IyTGALq
cKFC/N0Drj7/DOIayZAcNWQzkGrWDAYRP0l5X4zWbxHmMaau4WLAkymYLDU0DBCOFNb4+H1QhPZ/
0M96CwQVrsBAObwjUZpvMhJwIBaH1dniH2j09F2I33HK7JGUfuISlrGqkFdt9AcUCE2goe7MfvX6
keptfbJD2zExv7U4Z9a9Om+xtOmdLWZjjTOXiD0F5T9gXWrgBc4GPIxA16ZrefvMZ/dtKQ6N6hZb
4o9Mhdjf2QcMnmUADTnyHuAarEgXN3m8NosNkbPPloMQLVMTejDp9WVIqhnAmtDzoPk7Mnz19ZiS
nKrubiBVUUEGWk/soPcUrAbJ8S6cDFplgrGAzuytYk8f3AZAEskbFu/eTjn9PW8ByzihiNW44K5b
eITSZDKCQpODo7+b0aRpLARhTOs/zcdd8slpB4HLH98g/kaMy1gL93n4YjSfPH+NaawqjOQNBKTu
cRCD9e2RtB4HkYaGcteF92ci48Q+x77XABV29IEI0vKFFFOJW66X4XxoLsRebV6MIGlkI2mewuXi
avNIKv5BMnWI6D89yDnnqDWl/5Mn+iGlx+i23ypQMSdo8nDSESVxvNUMYv35eRxPT+vShKK6Asfy
Blxo9fLbBSWAe1ev0om31eqzlCtcTJElGmxR7cEgEadF9vy+FWQtQUR7ojR3dRHGAJhjHXX5MRIV
Uv2BCeyHmOce60AsiqAvTd5yXCTg636lwu1EO42+5zcXFsTtWVY5uiMvb8YMBfSz3zwRd04S75I2
qVFVLIWBbrrIJD/y02kgez0dIVSmvW+J7DC32VAfYD2ihjnlIZlTdW0Lh8DOViBjqqHNZXOctn+I
5m7i7Wuagsch8FnkWUuBBu+8K2BFOIrP+Srrc/ygOl/J+YMOjeRWQfA8/cz8x1FoADNKVRetSsYW
8nLOPXDLnpzlr5b2OC2v0DZAxz7EakZO2IFu63qwEMR1B7fxQ/I3JT0kg+Cixo2hdGB7Xjw1UsDs
lLc6ESPF1Is3Um5RQEF5O/W2z4WvMNf+gw0HNUG1S6yoS+jW/6f1Ijgs3xNv4f2AVynILbjsxeiy
HMOG/ZinD+LlCIuB4/sjQ+Mx8Q9VPYVS2CmcL6lyY0UWMHEK7DhrZjLW7VwFsepKImTncwcQMpWM
zSvCV5PcNGKFAuuP0CsS8ks+A6nshW72zBiLrHQqsXAOg+tn/i0z/Bf/B6iLGsoyJypVCkVtIvy4
rWYOj+MtxUwp0MxyEvEn/gQsLFJPzMMY8qGylTmeyFcobkLfPBJ+iK6IVVuHHZhk2QICHokb4x4E
m/ZTJbVDYIRkO5313pnNSkrMIv/ZqZPoie13hQ10I7djN84YRWtbRHkYVAMteXzAXCuLyvpGs5pl
GLcKggRjr07MhA7PIZUsikoOfMxhEHxMHUJbEqKZnm7y3wVtEXOE49rl/gq4jojcaghOSC7yMxib
5TGzM47/1p01NxQgCmBhe7ki/pMSSABVlrN9VO1/B/oNGYcbpg1XtLhXIbJKma+Moz5UycAcMFMu
apr/YsE4YehHbpe6q0o3CCZyU9bWzj1zXM2rXD+2gjx5lhHz7ZTfz8hgg+CvVippV5QqbKg9Clj/
0BcRp2b8wnYmuZCsUD0ozLM1E0g5Lp7hL7O+QfID/uWab7MzYJl821/5NsDTLN7W6Kkgo9/J6/r8
8cL44VuLw576aNxTRWCCfbA8TzZAQ7PiAgpMA2xL7TsBBywM5mtLUcBcu8rdGO/FA2QO4eyrmNCJ
/I1BiIA9nuRZfsZnn31Q48D+m33kjA1Yh0fIYPhA/YA6dBm+8AAvAu8Qoib3boAfC9ExxSEHRQBs
+aUjD6yoROyF5NxlW2o9RsU5XxQyhFbRNI47UzCPx+dIM0pfgdkxX43VpVswH7prqE4sEOGa2MkZ
2Bj4se5iNc3x1CLSfuK9AJd1ygMbWRqh6au062rofQAFF4EFxELc24tUz+EooTaLI9mQFED6Alc2
RE4YJDA60mzcNXf6ngVI74LgRlLQqkrKk+Im1H64brmyzEmODFGLIr9/2P146M88DHRJZtvBssf3
uK1WBnNZaH59a4pCoYa8CJq1CXx5SgjLAH4eEcuuBbISIWwmJnt/20/xumMh1kBVH/ST16sNAnCJ
NEPgBoC+I08OBvUu2FESZcgIa2FpFXBErmsAknfzfB7ERC7tUcXzrJO8u0chKXT0jofFc4jnLc9z
qGHUfAGrMAo06fW0q8Am4BHnveq6dgKeXuA8B3b9O0DS6FyXLLa7HDyspWTG9QFn66qlMZOALyYm
rHjedla9cDbNU5tC7hyRvTlPRm/iJX97FAsBfoDtzQvSaleOsgR7z99CXeSnQuDN5ChK+hmTQSxX
UthsX1S3nOtBbOFUqZem+fvT/MZBVYcVMUhxxi6cH6L6MCbiXuAUkWz9dXkadXaJskFS1yi6nApw
VwMsOuo1NWHB1aMEQIeq8jw/qVgtOa7su2v2+aCbcfHGvvKEOY2g+qGSVdML6PfsveaYsIx3RUct
bCAely5dgZXjKIDlQO7nj5Jspc4FLoWkTkutH08hrWT8NTbRUALLXU6SR9k0FjjXoG5S4xYwTMBr
iY5vA7JBGxNdOP1/xlhWW41pmWYdpw3hmpDDF1e3sKPrm0HqgNvfZuY1Xv3P057FHw2hJwoyx7Kf
JmoAqUZXIGP5tnv0u8GOHAiTS+qgdd4vbu3ekoW0/SKiSTPQbAtit5GjbuT9mXkAgNivB2UKMejg
0Z3yFpPg2nrC11vlpeCsjNb6kY5AGnYwWPA8H8OP56der7djuIfnnaeeajsGqthtbrS899LO90at
8pqxUy/ssUJvanbODK8ukFiFr6ooaDOSIH5TLrd6tOEeNflnFw5wwxwroM+yOLMX1mNG+lcAPCj/
XokhaRMpOpbUTf215N2X4DmlCkYM6MSsTrZCG7hPTbO9znYy27DhQgphRXSGFsYMrz1sAGEsq28N
MMTnbzXEx4G/OVrJQMyoVZ07B0aYQ4bzC9W1vnIqPk4enZktaCe2KqcH/8O7wYn5vg+E2KlX6sm6
GTx6hYHzpqWZzkDl9lkAwEnuZEaOecTR3cZataXK094my5dNTkfxjo9YG2avJEyESGetNDDo+CEt
EEYctW5EmuDsMZTHmdF/qcKA8G5Q0Jr8RmoGcRVA1ChSBBt1u7iZ+v5Vnr8cwYG23WR0XVnvOUIt
JpcPBo+kZPePvb05vjCg5puN157rhROSt5rkPB5ooj+wsPoswukrUR2REjQFkg+SAknF63fSdimx
9tFz6X8yZe0zNmLLpvo3VS/tJU3wqU+wdfRazYpYo0dG1om9l6Maxn3yAtkgLI7bzIQfgZzwGJkw
7FwAxFV6+3X0JLy1RD5mkYhYgjcVFEjksVih90Lydyc6q8BQ63EabtGkw2f9cDI5laKuQoEgR5V0
6BXO0vrYc+Cbxeoxid7VS0oz7rSJwxlhwNniMpmp8enVSx5C2WdncSJ2YS9kkDhRGt8o6Wt0FU2C
rpczzSNnaSQE44WJfN26TnA7yresBLWCYzMbiZJebUQ2FEJEf5N4qpSveL2Nn4/Ia6wfXZPi3pEe
p7jnGtGRs63A9Ryd9i9fUsaPTZWYldzsFMSOLyT8Qzf6PIePKsgo9MqakGgNMa+P7PRB6XYCnX6a
ILNybZSijdzlyvaOAioxCHSMKNPO7ZhKGMelhFnq6YSmcZIBGKoD1wQJCUSSmW4eXNYxZ2kd/hyz
RuM5ZbeO8+HuOtBsb4m3K3V5JfHPDH9C1JkQ+9BL/BqkBu/anytd1mLc9rdGhM/HHPSetVFDNTby
P/vZ9wQV48HIk0LNHoWvcJnGxB+t1CKsGST0u3hfe6kqjRUl4EeQU5lYk4xVMYhZ6FL8KmoaFDfc
Lm8l2agByMzUbluCGJlAlbr2DgeR4dgxHNmUzJRxbtlhmGEYwqC7dgcEVFyHRd97LecKTj6Dzr+y
phnIcA3Z5SCZ9Ffvf0sfI2MtpMz+bm/8aYlYCof++ZgyqFuy8kXoQdwqEhT7dpYI/gK1ncmSBU8Z
WV6IXsXrssV03NEyxw2Oop9fkdZE+zx0QZAuxaQpO8L5+6RPF76NB6TwG7kF39oJ171R839IyeRD
2hcDPA+5cf/9RnnMxtDeUEts0BGkS7jW9p1EBSpTp+v5wjac/Gz5Cv4GQOlX4iBW2MHREZ6DoJgR
brgZa4JCw/SR5rIF+j1dMhKNQOf7c9HuWqkouMUPJqNYtLfVYZ7xksM9Ifyu0DXNRCdTDSUJdOfc
DwAeP4HvclBpKV3y/TyK5upw4iHJAnODkTWQl0p/iA/tlAHHQDpzK2hDs7H/p1Y1awMJeGz5PHIZ
aGcLRNg+NvBNwr13PgrOb204JoCglylk59eW894+7sKnGyk0zAeK93oQSg4i5VnAGbLZA37UezlE
pjEPJPMm349eoFEVfhqnME9zFYIRUoaXCyOsL3h4eZMo9YeCvoNV2qek13F29ASNZa8if9Ic4hR4
p5TdnUFH/ETlXjtAhad+wI9dEmVUV/pOK/3Qzv8byl/EjdF/6biIlL3unVj8uoyRg99Ds+1lqiWM
pxCAV9YavHhQeDtD+P7E+UJLnKgSwbkG4PlAyjL4jWSIKdTyj86HuBjeZLq6U8cQ/the10FU9cpA
0DSrkgbPceQw8w9ELNUpCw2nSRsuALMnR/yjHPFBaUkA5T7f7tlk3HMqaNbllAZQB70icNrwcgf5
q1CAkogzPPf4YkJTkKpNvB1VyMLc/wiEcs/Qo9iEUhkMshYeEBMUUoPPhp2LnrRDfoLLKEWW7Rgv
WGsmj2Tbbu3zX0LYcl3XUgWYdMuCHm8NO28rrGqyuuBPjXAoC1XW/taPzeDzpxYQlpgnI7EWntCJ
MGMBMLm1F6i6qNcNwrv2FLE/rMGNGdyjtlZg3DAFT5k8Jro6yvVuWVhpLV/1djWFccWeFBTlbfih
4x54dOLzix2lBFO7+AwUQoh5Mw2kFCgWQdcyHFb4wlaN+saXcY9LhU/tZsWFlZtJbaB+WngJBoWw
/LOPBPbEb3+n2m4QyuDcCcsP6FhP3HVCJGLM5pxvP1JiP95ZHbaxR4Hp/a7qAULVxpPOnel60yKw
tX1j1PjX8RH7QnQzckl4xY98xmM/q4TaXfOU+WbZZVlP+OTe/he7pIJ0nOJrIzEauWIV9Aa6DXPd
lTAbndemhAh0JK2TxetkwpDmvo01OEDcOh8MYdUoU3njYns855fFpS72kiTXTfLTOW7SST3T68xK
JWmnOd1O0K4t/PJXs11X8hUbr4l96mqX4DOxmi7AovmrrLuKYfJUnrUTmJ1n1vzg401SlxVxnnM2
ZoLCUo3WRQdadlYyhhMN2nlsi39LG0Tp8naMs/fMSeoNXStmQ3/h/hhrzIkRVUutfXpN9fE8yVqQ
zdqU8hsL6+FzW2gsseGSknHpvQ5kZAPNaRRbnfvafeyYN+1J0igbSXl4STtnswCJ7yrbhQcmkv8w
mabQ3EkJuqwp7UNw39DGaqNPw3U/6kwk2ayarvbNLAWaWor7cZ4H1YyooVwikbtqzx/UpnELYrm4
Zv6oRixp0mGX9g0z+sjUpGHKBn7/+oHyh2a9Jw4K8olN+EZFCH+rqfoKIE5rXrt+yCwbVtS3dnZ2
/7Z8v9jmGtBvLXhYmywqqs3Kc9m7RolBKQ9uGl96eZ3RrynUVsfDAK7ecil+7GDcVQsVuM1sVNA4
Tj6FDlqmLlhDApwjRMpjFxRp3XArNNerOWZbs9Rz+9DTKvYrhR1+44C+S10QlYj1or+IdiwORA2k
s7OZcG4Yj/IaCDK27y+qtJ76Ct6ZHsXrM6uURHCWPmK+xLqazWxRXFumma8Yo5sJxMhZAbTyvKnl
yOp7OzvkpIQyDVIByo1QnXt+zhnbY7VacSuVVO8UiH0HJN3iK+1JAq7r6Cw4VAyqJgvBKAFL9Zrb
1e7BUdoLh0ghEoevMycR65WrmgOglSy54zKy9hRuFiGXb+cELwmxM7TEeznm4PHYcWvcXY2EDUaT
vsdJ08RxzA7+9giySVrTFt/wY/RnjbrpYI/u02yE2dkJOYy/4Bq5mPRItJSsPF/QHUFdQ8hjDzZl
sLDJ4zC62/d/wbWJS5+JQQ5pB0O0LhW72ZOeWPa+2q6BtzeAb/kSkNv8qy4jGT8fsx6OpnPQmpK6
Fp0NxVBbTONQGFh9Aqc9SfkvHghBKn+FGLVbMqHXG3lWps31EFmVvv+SaIU2+soP8Cqsgj7U2oHY
wy2F98VBJR0+/wUID6rwGy5iGZMoW0l5YAkeH9PAVRHnawp/1uwGkVSAKWtii2MH1s16lvVseequ
ZcDZXVEABuwDr3Vlm3i5cLGzgk/3Nf+djg2B9x44XWmyLadaSoIzauXrWcBWnWYkef+nITlSeUj2
4EFZMDkn+3CY36ngTE2T5ANYOwLHp21EuVCwz28s+W4eBzcwhyfakpmHRMzNNj7vGa8+L6cT+u/e
3B6yLQDajxGbHHiRSLKtZiG6BwFes+9CYNUMCLdTWSzz3bvarkDIJjUARt5mP0eCxpuf9+PN68oj
MXWKF0wAdxo/3ce0tMzpYyqDHfFqO/6Sr3NXMhc7BDd4Vqfjm/OcQ8hkPl+OimRPtW95IS3TyDo8
GH64I7duunNe3OCkub97NO65tzKGA8eWdGtu9O6aAVYl9ykX9N5kvrWm1pcNsAAwk0TPiR6oPON6
um0mtoR28sIV57XkJwz9dB+wPB3ui6gj2aLaW7k/T/AgREsPdpbidKtVoTQdrJdHFAiEF1YrknOq
4UKGJY8vgUNGSkNUHN+1Y4TdME3Q/kDOoEeLAULfBrjoD1mQwgie1fVSD3jzrsPwcvGShahzYxUj
s3Yqf7vEuby94MlC4Q6zBTSOgI2+HUgdUfr0Cy5z2XbYfx6/HnBJgxv4V27eJgcyKX7MNvrFHNxp
zLqZNe3apoYzKwtgnCMW4IDBZQCReOW6mMdtjea1jI4NdjkxJQMQQWFfpNv8C0UWx4x2Lmw13quI
Y275jZ+ZZ6cyTtAVLlO6I9TR1EyblvX3I5WIIpOC0jHJ4PZmXMqTKc3oq4H3gHrOJM4Hz533oPem
CItO4S2DyAcOY442IP8tpB7Ha4Cj0wOZqdwBOxp/UMYgGfb5rSAlxijgEBw5fFEXq7OTWCtLJoNM
tdy7zTFj1JJAlrnfYUEEiXH9sz4r+0LwXNLmtxxbkIrYFeDioBCzs9s/y3K6WoXR+ef63zP8t9RO
hSfLA4+WjXYQfXlEWY8BNuRwPbQuWquPz/lZTHCne+qRqZrZOSQcgRDvH8uwKBL68AoIGR+fdHpg
VCVZLnz5uK8bzWKbJJ5/r2sTStfz3NP6PUcsf+m48Zi3+AbGHUnKslEiMEHKQ9qmI70jyu1n8JT+
czvb63cavQXhWMJC4O1oERC404NvWnEfvrvj+uVexyVItuH5Ux/xDfcPGO0Zp7u/atwjVQkVzOH1
qtXwcCK0r6eAclzlGAPIe6JoSPLhz4wkvaLWRsr+8dYB849IOCCZaSMtQ2P7blcvMCfFJTZQZ4Or
IpumeCko+rnD8Wxl5kN7NnB1Jz0dk6UV+QbwGSxw3/bgZDOx4ycGfjxxYQZABIk6uP0sSGopmNv3
vellwpWa9LGr1Qk36BX4Tc2jO56+iHLrDRaeVT71NzFfrPfd93JYX+mf0rPitQ3p+FeCWWO6YfGD
UfahcqBlO9ih1y5/0eIrWPMy6KjWGLffGNCNG1BiJ6hyuPlSKHu6EUUz6aK3nIViSj8STPuvCpUF
kxbG7oyLAwS8XzHRTI33BxOtE11kAkYYw6k8hltdKdB9Q/wRMbLiAkniHzU5qjd6v63ETULduNxq
HR01JmoniskN8wkxytnfuyjFeb/L+RiMLb8/iapJLmxWbp+bnSU6agndC4QqLWj6EaO1cf87mD12
ptThDsLBnocUpQ1rZkMLVb7yNsIFrrdn3DoyR4uLye03SVJID1QZO1tgRqcH4lkar/pMeOqjNoVK
6l687B3CB0qRobBtyX2EwsqffWldf8AFCYj4FlTTiPx6DRovl5Ps0hS8N5CkgFb29Zk6hormyWHM
m1DtGxmkEfd28tIMFD8bi1YL64OI7jad/dxppZWMvJp1QEs7jP01PM7BuBo+Xd6Tbg4ZxOXj7ULs
aqMqzAdR/kO6KTW29dwlXt/BfuqdTvNGJ+vHOj4+NXPFRWvQZmmNOEI+6VEv+HFSqMVX2ESnzSBR
ORN+9abLfm1NKYam5A1bXUBs7PHof0vXm2xGI2SwDTIZoN3V80mVQfWHBril+w1/PUDQO/GwXT4E
CrZtygPcNMJs2LpayFnm4N0stBLjufMTK78pZlQXyrbEAfOh32fvdAGmH9M3Nyg7cnWHXb/qHaK7
OnE24d71ZPm1LsE+4443AEyAt7NkqpaVrRMfiPZIGE+pjPWSyG6UXT17okomaw8uIQX+RqeJXxx5
83fDS7UenpvUZzXEzBdBcKr1aDx5Yu5WUORYhjvXnYHlytM6j0g0hufky++u9dL+NImBtoOXySjX
CwlEUOtJkwSt4+kQcbT+5CCRPuWRbjsDqpw+TlVcWRk1l5M/ueOZlckgjH9UbyIvdUEWR4vWmh0D
pq7JK0DN/v2CcovTbb99HqH3omPMwEzPF94YDVNmSfbQN+cNWSpHRccHYcIidsZ1v3SbfM03m66F
LjiS35pf0Bom41nPmdHEIjmEE9+rW9hkcNI9HXVVLeLYITBA5qbdKMPFz/NoP8CJ5Sbm+pyqfG1S
vhmaAZCXrsJZR1QJltZPNRrgmNyJg+gyEuG+pr6+qIB2fubEAvAO7zL5CsdkojapeIzfTey11/1l
rtg7rDi2eOMglCfR9hzvio/VmkTI5tES4zPL+rOlp9OT06oJxtAi5ELRE9aJlPXbUI3zAWdDUO5l
F3rYb++4lx2SQQvMzRzGE8AgiN3zEdvboUZHUMzW6IV9PC59x7B+YCZwtClaJRC2CD/+pQ67SSBZ
8YeelkVK+R9DXKChIEEBBw0Jn6bUt8/HGndsohPWlSAn+fm0mV/I4KVnGgf3kUT4+Bm5BXiF17KM
JPaz4pIU0UkMITgdyDuITf6CQNST26CB+997lX9FMjUP0LSZn1n8onUbioyk78/gC5a8WEzdVl73
+pCT6T+opQty92aPyVXlaArjKM/bQwMkxc82qKQ6E80SPUXFfXrZD7P6iov8bliDxb9q6WDuSi8/
Y2Mj+wEKHj6Y04xXSdrlEJemMv2bTkG2/cjaHFOkVzqbnpNpiR7OPWr1HU0nSpT8aZTooGKgYGhg
08mo9cleDOSofbtn1EPts9wKbA2xEF0Xiz7GnjyciiDzMbZQGW9Mbte7Otl8tXUBcPj8XigXIoYU
TkOW1KCP2EqLdT6RhZpdl6/6tar2Xqe+i69CPjGVC3E0GLFpTPwEg9/h0DjaVmQv8RUr18faPcS6
bpIa65BAytVImdgVWCMifyTJkrYHVfFAjeLYAM2jXHOz1HY3w9ms1B1z6lyaCdPaeNiw/4dnG2rO
FLr+iZb0WaihTps3YNQPcyKxYmewRd574sJnWgijoZp9OQLMbMey3Ze+Szaa8jLpuonpZxbOU9OB
MKLnItelF3MofUgjrpPd01nELe0hVZ9laZIy63yZRakDsSoY5c7BYCmcm4zyZjixleFQJzjirXyq
SQCKn+OrkP8a8c0okoyqWMhBEsnWfhQdITxZTKN3IM+nIEv1k9EiXzy9hpXYXtJAFPkBT2xXS/B2
11BHXI0H9j7bsUNgQO7yoKKd6d0V27x+Ieq25LB0UBYzk3VCcViWU+HG4rOeclpJGuDWpPvfFtbf
f7HH7ovCTIv842vGjiR8tSrxkbKRuUJFOF7LEJVceKONQTJOmiTncWlMmqEGtnY0wkLlBxu1RYVY
4xYiBujCumOpb756ebfj5CYj0THy/22MJDV5qAebxPQ3gVDi1Wjf0ePvvBgj9vlzdKDIZlLGpO9Q
WGW+H78wiXeVHUfD9VWIHfxP//VJ+ij/KjUz4+KQfYu+6rPdrqjqqBfEK956OZ5CdW7vkuozhJyv
opPUIqjg+tr4HxcbLmN9GSzLFNNElYH9fIaVt5Z2JkKi9nyFxc/5K8uD7MKO/SurCn+cOUuBTMbh
+PrderXVQE3b/jRB/44ea0wXpctASN6xgjjkErPi3FVFRhk92RVfZzIzIej130FocuAItiJjYlG9
lIX+OeslFIbqpxSPCOp5GaBLrMfjkBhh70+LfHlNXMkvRl/ocy5yN2M11G/TRAR5Et5DBqBCjm2J
+GnlN1+glhAXiZi3um8dQ1pdWywC05BdnRhhNqp+xN/x6aZCYHrNi0ZEzn6TH3eD6lI6YpmpPtVP
bD1ZUj3l5Dvpd3GWg0exCBDqypJZ7kKHb+svrD1NIJ4A+EEsmWg65CCl+XigdlBdTQLenwCM+6KY
q4Scy9Qio8e8RPFf8MLhVMnx/VpyGiO1sslq20uqnDQeLHXjJCaHmM9otP7QXt59wnrD1Ekppzpt
Mr+wWyR7bDm4YJzt7oLdrEsLTy5tyZF+XPPHltGybTf6Cpb8IVFmYIaypNkrONKU16G0dvmxqQXx
wywhFRnc1V/bTC6Q9c76hS7HzxrThmqyoMM/twpcSNa2FcVq2X0yQRtmBrlFWHTVARdcD43ppD6/
62BH4mmGU15rk07HpvPIxJN8fkxitj7EdVALGaG2/QgFiE4Kv0BnWr9hY7fAkbQgvmFzG6rLXaNZ
8s9jZe6ngfV7Yqw+H+VYZnCY9GSbbY83YQyyrdYj6c0QS/9hCQk8XxTZPX07kF7ezL2zOTfDwjPN
7IcL1sFUMoizpXhHgmoa+Aa9SCxZb2D3ToMjgHDKb/cWr9A1gc8XMQUH62q7b6pwCo+FGdh1sZA+
ZlTse8BEsXPSDzjUZR8+LEnb0VCLLKWSFih/kaOJcpPo2cVqoEuGdOi1Q23+jduzxC9mtMVz8Oai
dmIaOtSZwHn8LGH0rEPingARBdVyetPrZXS6CFaKrA5dQP0Nx2IuKDRTkinaOwq9adAyQNYLUtBX
uP82wSblg+d4HdpyW7FrCUjn4q44HJv9S+aEwSh2OISaVMlAN7KRRFDOn9xNtkGdbpRgPADD8UWq
R3ByTl+/EIx3mV3HMH+4TWEyKWglnwvnB5YwpubFueZIEOTB92JyZ5CufL2/iEaP2SvJn/QCZPL+
5J8649jexOAyNd2Cxc7lu8GfzU2zAk3XZj79o60WqvFPZemp3BHtkTFJ/EKs1NwqzlOELVmmuNj3
22WzZyYeGBv4D3riV1nZ8p1hCrJ8wp+T9v2rBzjKHixOSqNlwGjfCp/VpiTaxs8DdDuP/hTjBQOZ
w/FaxNbxpNy0d5n9cqjDvrADsEo5w2t1uJwPAq1K2gP0o/sjSiBnxLg3WCXhY7Q9vxMaAlytGDjG
kWxkGxRz6sTv43x9PhScpNogJdxuU+wCVAAykpxYNTvyPTqN67OS/f9JismMoRscRSVYYxBVMWG2
ECepw6J9LqlK0bk3INwsXdjQsY6hHI3D5o2Ed4vHSNI451rrE0fPoRQbQVEHeCL7PowkXIJJp1Yj
KaJqXMcydYK/SfY5/S0L0/cYLHXaZaDoHY5EVZVrXmZZxdJwxB58CAA4GJIkfcthaV2P45W/69Df
6132dlGzNK/j62keSmjUNcYg8bYJHR5K4saN0cETBHFZou0/QKhD5zs6qc9ua94PFMRxkVN7RFmd
In0KgFkFBRtRFjoAT8U+PDjeTBEsujmxm1KAPhkpfxme9Q7Fs1ARxLzHDIFrIT1Rvqcx9WGFrhen
dR/u+TTz9DFMFz8ZMZbbFf2yo7JzHf4qqmDv12xyL0bVNE3tv5WdfSUGFKukBUgdvlOXOZSS+Xry
o/wLXYfj7K/v0cfOfqA7NtDuI8OTn631ctCBybVF0vvOUGrcuBALkFG4QdXiYP7ip1LjmR8z/oGT
FO2oykREJjSy2fz4G6PEzPDYrjUrjaBULhzTcqXlBfC8W3m4nHwsCLIDZap18FCWUlzYVujQs+7W
8O0X7j7UF5EngzC894Mc0wYZKNV83mLRCxgJePWIMw4oTh8/gAIj+kGG7baecR8fIaeArIfdQsO+
m2og4I+7LbnJDRIm31m5vxYBPxEkGyWNYYtW8WjIHm1kd9wuHob8obdspPIjCtB1tcWjFAPB5vf0
nP7ZsIyQyITLUfivsSl6ACI/QJHfauB7x76z54ftyN5zCAGinWaVphdgZ0R3kbUGAhrWVbvX0spO
d/KKJEpa3DGG5LB7DA0+d2boOwKSilDOQytyE83ATuZFPllMK+E+RM+DQCGnlTIzG+YqP/40VuhG
BEWsOxEOUJ592MNEM2RDs8tZFJUSRCyVo63K1NoGT+BU07WmviCi5gjj+h0U+3qOzp9I7+aLnqy7
0wjqOoi/MO+64SStbMpyV+apJWDEnBcgZZiJALhTmx7jV2KQ6hUG+CDXyPwVLa9CmfYm2XuI0j6k
UkR2IEYZSf5DKyjGN6sOsGd1biR5iboVU0idpvY+3pXrtv91dKRqaJ5vQuOXaQ68qU40H+M8osB/
YROAZ/NG0f4py9jv3t2LcF01feG/l8l6Zes7UvAO3Cv7zv57GIQTfLKV5IPKusgRb9MNVg3Rw4AW
/m8IfIsmjNKJDtnGKke9ILth/MNApxnWz4ad0XYydHevdXlCBg/XpMk0/dboEjsETwsGbjyvmg56
fzEl6bH7cLhxb8eMNmdbDUGwmboNQ29zhDyhnEsZHggIseaFUUCyY801z/ESrBr68knYJstj7bDd
Lhy+fiuHSiL+bcDbmaG/sV7jtk5AffvF9FGo0f25lNrE9D4k985rTCFe9V3wU/aZO1nFaaWG7F1c
x3Mqmhsc8sKFs0wlRz3sZUPt8Et1h1mAQeg8yHH2Y2URyucl63kM3Oion5hpGpq0yJ2f+xOUgKej
LatlV1KFVXgagrXDskvn6/2NWqZ52S1rkJzV2ViRknPbwG7p1YKVfxG3eJPy96y2e90pWntI2Qtn
TL1WsGJh1F8FnD0bbCev+P0/MoECJGh6Wy4mndIWGn0cgdHNeB9cSHs2gIzG45UJN8FaWGm4Lz3r
HIVyTwoRk+iJGLsYRqzbqYLUsE6t1PV25lxdbD81u+ljTnWBwcWk/1vevUAtU1BNxWJrNu5RJhxy
F2Q8zJNwLU06/Lxrq99eLhX+LZ/IhXvf0EH9LD2UNJVFrMB8IpBHjJ6ndn0U3NnS+lxwcisoV9eG
mIpu3XHSirJi+gCM2eFs7qDTAScskMGhzgWHaGskyR6awgErJOUeQnnxqMmTk6LfBaZip9XdS2Gz
BD7hWBzgj5p9Yzhm7GthxRB1g+mrelzWEly82Qe8sNx/JjIT9CHG+eRCo/qkWh7i4cykGLlY+9y7
7BUolkCu9bgI31Z/yCD4wIqvseXN4VXIxNpAFMkgR4eTRPAKyQf0TYyTd050Zhi9z1P48+4LGTba
LcRdJgdzsBBHvnckwy/FyAFio029koh/XjfWwIDluAObwlPJPMNyvF4UbDPBjLeFFgm4/SyEDwxr
j9SdJiRCI/OmWhGRNci2taDb82gdHkmLP0C+QCmplmqcH0RNARlPRLVqC9fioS40yPZKMasP8qUl
jlSU3YxkAhVNrBmXOrEkfbUw6o8C82QQflUp7yJDw6jIFnCFk6mxPQ9Y4YWAnFQpj5MHUlbU4gUa
Ef6LXScu866iJ5ATJElEHbVADFaeiH4KujHdosz8ksfeJE3bHi9ulkAsRXjXGYW11j70iu7rrOO6
SO8WZkmFQlgw2sLJmSUj/oqm9QsVuDfLk6tKCkaT3+VbiwplkfUaNKBbkOC50EQYH85GhBm1vpRP
64ZIWZ3TWOOUyJEI/i1v83wGIY8Nw/vXZZn6FzjaCKqE/BTv7MOKR7G1eW2ryeUnHxf+Z7notD6k
FMZnBKXQ06wDot9135RVRZFiFPGSn/1VckxaihIZwLUyJQoT7ihwaDFDLnGljyeohZ0jM3zR6dTu
No21YkXcpYie++7CnQrrzwuXL10p3G6kBjtLcLL1e462i4JAjfiUOER6lTaQbFLnHxN3mdly3/KF
dvZqRvBSYmI9SpVuzXH/Qn9Y1X4rXczwdsSX1Ti01Fuv8rAwN9+pSBatRozn9wMUSC6PLY0f8Rv9
dy+Nbk8AJBMGgs/OefY2GW+KMlxHSIsA3C9xYdgrY7W4VCMyQ2zasBu3EBlH4EeUytsuV1cULIKb
3Y8NMM5mcs6scYBQqdB+15ri6mFYMZ8Jjay4Rj2zOqApkGDmAsgmOIdIrYJB/KiGKyuDsbcoO+gA
gaIZ+woo0flmI6mnInVhpSqMnTqkMKj0ZZJV1fxFGsKqj50LKZ9b9zt6gT5guD9pVIckpWwXl0LA
HqDK0RN4MPRJ7rGBEVjVGa0KS2j8U7lJXnCXdbHjGUlTu9RGpPun/VGgf4mzVXZ+iVzWe+XFaMdQ
YXzuNDXlOMYskeEyo+CU6g01/wB6sBinNvFPyzMNgLqI3K4/CTTg80FvNu9pl7ysS8nrpuxdaKT4
mKFfOVX8vQQbCaQEe+24T2q+pDelZnrQf30zTZcCUCVd1mOHGWO+hAWKk2Cj2d8POg7d7jhyaboI
puzLMo+M1Avx5wXeVteriGhTFvPBO0TBa+8yC5d3KNyZKDR0v4oVGqm83kRYIc9yCCrcjb6R4s0m
hZOC9DXdnMALa+W8R32gRnuTudZIYy++UDJPFof0Ari1evK4Ain5olFp8XKUf94hGGud76RsOevp
twGV7U/103/WD9LB6AXbmHz4reKaQFEsUwN9+ztpwtXgDKXhNndtU4O6XJ4gyu29IjPdVubfScd2
Q/7hkv2KCR4ltnDUP78pYrpY/4LwOJFL8T2JrmozlwIJSuVlL36QkYPNokpv9qb/jhkGn+h9FOfH
RACvIwJUSLyr2ZJODAl8QDUPaFIbJjfIb20c6UaqY0+HPn16y2o6lI4Xf9EFURIAgFscuT4YR/wU
JpprhQg8UnHtc/3dU7G9H0bt8fWSu2ijT4xqv3/KrC3XC6mD6KYPupp/OKmHPxyE7NxCWQvtczk9
VGXNZ+39OA1ED8Ed9FyjQ9R70oxiQMiOx9tVdvtdfiHsB3QnTsqwGJc+7SuV+Q3I3jwdPs/diT/o
eu6JeQmq/qw050GeIj9XhtDqOlp5PPfx+LP08uHaWJCz+ZQRKEFBrxTsQW6nf5ds5cvParN2vXTn
BUWl4s/+zNBzLdd36EW/HfINfCSh3BkKDOja6LybX5p+P80jMNu+JqdPLA8TI2pYawij92ahOOJw
81MABho/As4uMHjfSir5JefhfH+s8AV3ZLcdqHRrF0C6O3cOC/HG17KkRPA/U3lndxmd+I3ijpOv
rrkzL3fmO6ec76HlHiW9fc7z8ySFLtHRAcC1YJInfoKNGr23fa+dGQ0FQ7s5QTijGaraR61Eyd68
MVtj7SW5ckLlX/m3y6ZUGme85/ot5qbi7elXuin9A/vRx6IvUHH4QWvdpPQ1KTQQZRlv7ab4ChEn
xvPpQBIpPDB/TSXqXnaaysg5/mQv0I3Zq5kgMkZjjOef50cdWfECbdJ95hYozOvfaDYyr0rhQVE+
vbO51hb/H6SXcL2tU8sKyaUdUgfGEIOGZ4uLDl1QhJcPdR3C2vRlkqMwKCUDZsNHySbnN02kR3xM
3ShcXUEboawtzN0YJDGojCdP+Wf3O3UWKR0Cpexa2b2kx/3IBLl5GQlkQVYgAj5lW4mK3n8hxDhF
lKeVK+95hYAdN28O8gSYo4yiSoapFeT41gZBJrgKV2BKRImW2khhYkZK7eXs/jBK6OpQOn0USDI4
Af0UqudYhyAJq/UB5WuPAIFhvCdMq8rnPay71q7ddvjhUzsdzL78IfRa/JDoU65VSobElZRdWotZ
sWX82YuTELUXtTT9x/KiO2b5DFBsyE9u3eoFsJ3DWPKpRGxtj9eNNl5d1kpqEI3qQcRHLV5xvYwl
m6kX2XzJ2RK5YnoABERrL+nS+2D1611jiyIFF3+6lLAfl0bNQkjljTRSnK2VaXefuipptrN86Egs
lz8dxMUiudpOpza22dX0wesk//qr0adkH5HmtqKf0pJHVTlAQ852VtWRI8m6wO8yH3fHw5KsMbuM
Fn9mag64uDI8JgmsYHxeO7OKYeBjCfwMwYaPVSAp8DOqlC2DX9Ef2LSNd9n6YnZuEd3CxowLxgWG
C1PoM5se+OIL9OAxbaZu0Ngf/hGj/Dk606+cf34D2zxhf2msK7+O8cADRJenlbaumFSv7Ccn+fl7
9TyPnRpqc/Y7zcT5ULDAcR2a1Ga3l/LhFhZGFRV2VNc9P2I5xKPtk10joGuCGJBDcd6CNMvjM7nR
jQi6nuaMjsaJ2Tcwh+AzC5iFOputARGWx0RbCzy+0zk4Q2mXkpWP4Qz4npTzdYHnabdSr7blEnza
ljTGldRqlX800vkPFKK/8xkgb80ZjQtqjXyZODaj977NkRzqjXzAvduLol2gi2eejbXpnIU7+6AO
8VWGC2wdxzNq5F0kriIhfcHrVTaHnsqTF4dPpyP1NbLWcioCx9vFUPbnXz5UNuNMLG1o36X3ZOda
FVk4CfaA6flMmV0aydEwqDk0DA22RRqtM/cBFz39xUM6ZT8WjzevlNV1ryNDg6jHfYPS2g+7pj1d
7ldI5d5L63hJMoJaC0oFcEcM8NicAnh93f7TH5kRe1r7RHiChF6n18uOAUAfWjREiWe2T37fxN31
ujuduyRi0GU93WR2tZI2CVQ6i1il6NnX/m3CdwtWM+pcX2W/1XJci1Hhx53cKrOv5/e2yFA1N844
ZewKkkuf5B7yU/nRCRE0ZjK2hAcnJvhGkUUjLLgki8zVxCNmvI6sLpWVE/ulLf8y2X3IVomQsBS5
WuSw+yySz/6hu10NHFnwuFtdzYI0CSUCM/RUa8UhuWFGXIKlqhsQTkE8DAjBaoxBZKcD4HMNWRSp
k2ti9gTvRHAvplgFxhluPvmN0MVAyHxpqbzpjAgPOOvcDnNkRjDnJCF4kL3IYbZJngyqyI7rSSkF
6NzFEn7ui4GUXVj266sU3bqqU9UAk5KRnZnnLwMxmNQvgqgqDUFYIMj3j+n1jmaaYXnpT2abf52V
i8lNuA1WR8XylCWwKeTp/NJ2cOs5GrplWtgpo4fa80JGbUwwPW4w6fyamHiO3AWUyrLWXX3NBR5a
lbLxnnbp4bscrPe4FCao1/lKidACS8wN8hzz95jf5jwWM9vr9RAudt7rJ+l1RlyeTiT1s8mQ4L9K
IEoH8h3TBMTyhAjItqBhCfmueTA7RltclxJpRIQUqSI0cCovzam4pOR0E3RVkwbvAeMpGAAvbQa6
kEDit+ykWqeFS2FPySpe5JcElS17mHjfFGz99j66gpAcOT4O7ky2ssaXv8QDUsDkXiwoho0hZABs
6XbZzgISeb/tQ4sj08wUmlArzQxdGYxQXPQBNSnCL6CnDnPXP0tCRWWjUuOJYWPa2GC4016gj3IJ
WLWtVEMivmBqNMH6LVq6mKxiuUrHRECuOY+mS12i9gUTeNCRYE7rEGHVs3L33HMtPDAad4vMx+nU
jYp+ZXL9R9WSUkZWGTsfqDC7ZeC4POw7s1qKdUHPBF+3Zes3cTAx9N+8q379c6D5rOYGNPYdQMIW
Ia8jdoxqDbscQR1M1+l1aCnujRzg64YfQZbCub4YTFiqsNrY9wQYOLVzUmfe5LX+kuPIfAiOu7k2
8+DFicMUABnS+zUO/123+9bKf4tIvCZoOeHMttkigmpMe7euD4876OWnHrj3n3oRky5mlVONd4pR
3tu5CGhdBjVjDYmkwxtg5XZ9xifhxqfM/9gXLWl3AbPYLtmIO4GNhUEFH61GODl/3PZeDB3f8KPG
MDwobXPhwPRKLwos8hdufLO9m+sW7ls/PZx4YsZgPbod/WLtcfamdB7uiJ1WzUPI8KODHUxlKZMa
jnBZeC+EXbnMrY51p0US23i0fLzdF2ZYJ+ViZucmVmMST6rONhsmyUmRusoIl40waCPrUk8DSPe6
6wr71huBJvCsxiJxVW1CNbUHTX/rplr46NRmTAEaD29RRRrY3Gg2ROMkYdtieQegQEHXflJDVBd3
L/D7qXOISRexaGb3nSC3nArpJMjW3q5syyLfe3LhKrXynhlMABk0wSgzjKC3J2hAhS9TBgB6ElzO
WcMFBOMM6Wuz38g2pp34YvbjU7wYRA096HTKFszcUcQbj1DTwojjKukt7Y13cPquOKtCieoN3K7T
uxbYvd8zmJ1AmZjswsq0+QtUSVDKkzc9XBmtlDQiQWhUQYzWX9T9BxmU/nu9XxIeFjFXbvI9I6SM
9aECOM7rQTVAOQv341iLkTHbNBbsUAaYt8//A/i4yBVb0S6ojaI+Gxho1i2YZCSKekYDXDyJLHTl
EnMG7mZV6jorUmVuEq66kzv5w5uw+S77xYunrzX/4pCWzwyRx9FigAzS6hiZTn+ofLOOWj8E+7UJ
q4d0000eqBwGfP3O/6CHZE9r0AJ5iVnz+K21qLrADX6EeI0RuP7nk4B9r09EDKSskx3We2cfkhiw
NoPYTuXRZf1NU6sIVHzj1CW+gIC2MgX8/LkXgH3r09D1rf/wRU2D4DTdnLd3c8OfXz7Xee6B3rXH
9qd1QOQwZJbsgDaWMZXG0mF0cnsRFYA0pMgARic00l0QmiRMdOlk+nWjKyW+czJzzSpvxPYFArVI
W8H508RzUZzUFinmX5XKCXIRi3rR99+4NFfE8TVfojlJ+4ln05/bbVpBrJF7E1DpLHsHbLgjs8HC
f+uBVstENtBlAw9LQs//NA/3Effn6AfuO5940bfhW/Pkjb7/j33+jxB+ERFM3cGPI/qr7JwCVurl
WwalG1KrKmZYRdMlbKpYGo4KL3WB02FBO+G2RHJZjV26FgXVuY9srKHwAfVJbWCsRYyFOkJnBzn9
JIDaP5RFBsd7YNwXX+yXGsGLxyjlf9R+GHTI/aNkyfamn9qlLNmc6IaJEp9a702ay6fWneKfd3xI
PfxDPbMbURS8l5JTPyhZpCthDQc//enQyIliXMzf0ZM4kXzIMhwq96hiaxjnoClZsusnxKmus2mp
DPr10Ck7UPBQW67hJxiZs+Ep4zzJYibhWzXtG9SA1Zx+AV10B4civGRq1XD7q5zdH7pujZjQRPKx
wxhQW2JllFCWK213Uqt7WKPxQbh8jOn2Jb2HePqepcslbjMmzDnyQbdMj0LOlXtbtqMSiIC/vtPg
ulnRYmgrfi46f1rFSkdoYKiSLLu2ioe9/ZuSon5lc6FChWhuiUhm5eTQ/Jj7ud9owoAHgPx2R3GC
hjldhFcUB+mE6QbLG/oP3tGxNsQzR+xnhCwrqh6tHe/9jFgh/3b7LbZGfDCTaKTxZ2cbyKGwtZDM
/szzo74whb4eeer/+YEswc74QyeUuKBH85eeKfZrnw37e0ckJXw3mN2ZpZfWvUbSbyxoXisDOIfg
YyzgWG9SxbOYZdqtPK/kNxT183zvxsGDthDLxEaOsnIyvDZO3ys1AVPsPnfWafJ1m0Ynp/aXUQ3R
RP8hPb8VJz99H+VNwAImFJ6OnqhqpbmFTBHtE2ZtOMPTkN2EdPCDbJBGiHTemu+MTkCeEWB8BGY5
zccUBr6aqoY2NpfuRa7ADuCTf/5knMOrgptd2YFHa8j38oqOGt6HTx9M8V1h6rI69n/5N8Hn44bj
kXUmKzunbPXrKVtX3k88tGNSdVsnuJlFMw1MlA9sE5sAQpOptljeBhqkA8Av1wCX6sl5jk2Bn0aX
ZXM3eXeID7qXiwPjDFoRRSF8P2VTPA/3Ahvj4pRH1OeB/4ooV8k2FgHIjzOep8eRh5KQZjkn/+66
a53D9jgtOW+FZ1RggRSG6wDn9TAbLAMTsgxWm7Ki+ZUNIlIyaOHJ2QuuqgzVVby5XVZEDYZq4i5x
X1Oq9Ly8LJwG006Ylp9YXxRHN8npTtGM2aRlXdh7pTCGmcwmNLDHFHG21xvRViiANzCkLKAIb7ww
uSO2SpSsrIXlWSkQvCLbUs8heV8UCNUSFLXWJ8CR2ob9Zvpt0mDUaXBKZ/o3wcfXInllF4FPYHuw
Wjz0BqrR0LRGkPKgZbMszm179ANt7nTJMxscChaRdF1/G0+6oHFegG2tGCKLhH3mP4FbPRgiyKV8
VSrnf/k9ppGL3qrtUPEvfq9ySZZgoTY/1u3j8mpXCN08q3awpMF60drdknWmWSnJE8OV3DfCVw6M
wt6Tzl9e8dyJ2eohQbb42lluTWCd7mw0G0TVLeN8dtsAPgpQ9FsKmZw6vc7Vyo2x5cTKUGf4Jwjo
99vD8/3XuDMo/ZTft1VhUrvFqaEWLNPzhHvCFRnE2lKl3dHtubuABiVKnvj7wxxLsIT8/lJaAgKb
uahyaTHTq5uk1sDUBUMtszTM2HynYjXJfzUjtsU6vg9xGIkUPUVLsUlOuvK7P9ZXVPptU7bGwNir
UvZvg7PvHIQ03IEnjhscbBlOhOvN22omDDWyMNiJgdS/OLJ6ChP+szHCHZPM5Btso0N6YYhn7lWf
b1Fy3hhaWLREmSQ1TlZC0fdBOf0qE5VkkQs3FfFmpDSPNiFqzpm0XHGeoUuw/2fFp3IT3M01Penx
FROBFhXDlfhQbTeYKaBRJpm/KTt3DnV5uS80BsSDVHxxxFBhW9b0t+x+XA/vOZdYFc+UFpw6RJtU
sRNIjiXBgTQ3bQfLHuKDlL9bJFASboJP7kQizG+e/354JkVVs8TLPVjOGvRFL0usUY8MnHVwg3hc
U7b7wcKsjkyaSkW+4DDGvhPAL901FLl+eqo9yLf4P94CY/0de4AtJa1So5sQZrYpxXZEdtHjTPN8
7gl5Yi5UYMRUdy1e7YfFOI+/LavL+Z8/oTGLfoOHE0r0R9lFvuwn1E4BBAXCzVXiVuVcl7Hiopka
4POFMDaZ9AhsvB8mlmwcSRyaDxgQZpWHH9ewBsUOEp+0OKwkGwjUhe8S5lGctvRXy6AIlEhJOb/T
x4dyuV2hc5FOKZlE7VWX8mJk61ve/ZnyNZirlLZEV7LB+JG7h+1yLzLvtGmYqbGQyUsAhhrGMSKa
0lM005yGRMI9RVCJc89/nlF+AK5vY38PFuKOxUwbNdwFUx84DEK9KjkluxRLqlOR2XkECotMI2Ee
VqJVq1WA/tHs8ExY9bBTTFNlQlm2b7jm7s5Hp5t3k+GLOmcgIUX4RxKuwLcrIApAApMIfEDEjUwI
Xi7U4daF1hc0Ap+4E4XLGHMzGJwzp1fwjyxhy+7XlXQyre3H0tyDlb3HoBQaFbRhChN8O7NRZPqb
0WjbdxrL+mp3qlDWCwCmbvyWS7BGe9N7pFn6Y5q7fZUtxesc9suxYEErLg0c1LTxafnu5gX1Mstt
VONYDjnhAEWNCJoVBifQVTm65C1gc8lsUzCiW0IyGplzTbDxpt0EG9biyiPXP88qoe9srQZYcbXB
HRqebz+B88xMCC71zY41iE6YlnJK+SaiVQXhg4f5dVn/quPzMtDIawxj/pFqnEbHwstgL5k9dgxF
rn8re7/MdcWNv7irGiYa/fOWwHlNXaCkPpStx2QzqUjNQewaRfcu6EWOKDyAaJ7/vlAWZDUVhtmL
K30yCxgbTGIKQz0+yzOXSrq5wJqS2yO34/yXOeWPjT6Wd4HpgqgNGjPS606N9SO/UzZ7RMyL9inE
BQduL3fdmY9Jt+DWygEkF4Ddv3Q5APbJUoPhIfd0f+goYXXRK9pTmsBnuUBg8ZHkwL4PuBDxC2Z3
NKINHUlcZe1k87foGjZDk01A3sE0eu5LwQlgTIPDjdzb+gbVfj2duySlWDmJKz2ufcAlSur3fePS
mResvIw3pUUIpL0JHWJ5VWXfa8BOYQkCDvTCM8G6OxElI+ffOrS9WZP38TzhHwvQMpH0ZPRYLOUg
vbD+K5BwsbnFrNuxMZolFZvXbmYbii2rBSGAOxwgVneNGueeTyN4qAhsLsZOwiCx9utJ6z5HzqQM
htYqfeUxubP09uRniLQ2sV2Yjl6VE1Jt650qVIvM3YNPKF41AuQTI0EqalbyQC+oKVk7pKiv05uD
jKtNZ3t9wvVaAoXsm9g7KvLAwuAyOKpnVCy9StB0fOTwffz3Zs7doEkbuAuWSCC3wqyPf1YXDsfd
wY/l4GrUgXeKlvrneqF4Dr168pvZMadOmotpxgkRyDQKif2uHAEIBH1enZQrll6x7ASO6p3nvsk3
TA6YI9HsSSeIevZGQoHsBaZAES8kRCUCwwTUBWAY2+1YYMXefIoe30JLLV/6vvjXpbLokWdFjSsc
61PL4c6GfRlhcjGS53lH9UCtojlgfpxlvHBAxs7iBQkGqJSqOBKmjxiGnJ2RudAcxFxsRvENA/fC
kVXVTXJ3VthJEQU37X5z1DMdkSYP1739p23DzhhjchF4O/TdIysrGNnZa+c8c0jHpDw6H1W774yt
LzejPl0TyQr7a6j2biQPJ51JudAUM/b+C93H6183nsKK6Ge5AgSecs488sXLSF5pIPVbmYEL0+ZB
/ht3qNwgP5GYdaxrSyUfX0fHr+W/XTYe/7iGt7j0O0SUGJl/6MK0xMRwVr7N64tzz54C9mCFIUvq
tpKxtP8VO25YwCYPgI/mt7SjdWX+zLtI1HKGHX35h7Ad/Eb2C25oSSPt1po2LV24v6cCiMKqG/FJ
tdBvTI6ue6osXUq4P8Y6BnLsdQjafESHnP8KXFpWzldeOBQ+X63Psk8W0/YWpOp0KOUHosfDL17c
CLcJYdX6LxQZyn4c8btIV7VvwYaZ/jlcNdlOfNcfnySXldjB77q38QHfeLncwpYBK2fOEeo/4Itg
iuyacQHz89fHVJnzX7CFtvMmI2g5I6Zoe7bHAZgK4cl9e1G7VyXzDG2kWq1MHH+T7dHC4ncTG2pC
WodTF4lQwOfYwLrRvgF9kLI9lfjerl9s9iv9S2zSjEXN8Xz3ArJfJusqQa3RD84LI1LRBRkh28cq
QIXaPYPSZdZrHof1LkELZBVk9k7+IRd9hyDS+HmCTrj1T3G/sbTfeUvjgWLgR2CNIfndBwrQa0Bf
JHhwMdjJ1psF5yQSwouzQ8jaME8WazowOL5TGb+u6rA4Obu+udeOMU0dKvLy1ZTWxQVEElysO25Z
gpor3r9ag242tQ3ZZVV17mneSrmTfSrrL5aL23oFsL8k4Ek8V5PdT17DwJqZKpcIGFpo9aENKiXq
MJIFvR5OQmoTqdQrXI53Ri3kcMnre9qtly0l7sMgNxVRzO6OZ62AcDLg7F1iqqM/gffSyAbSq9of
Wnu+N5E4seVmit3iyF69lCNfrte89ITHgpvk4QvEKIRNc1Vk+pdHE/70xVlGS2YngZt8msBG7pJE
zEmLwWhUWkGRlgwyF5nxX5JFmkFjofLYpZGZU2WeS0vzANxgPkjQAYR85HiW6JT6Bo63k5FWdrh7
Y0UKwNIubfcT1pH9IZwNoG401h4UlzvxIMviCDcnx3RiSxsDEfKJyH/Zhr7gq8EzBgFOLDZzG4xo
ltBb6MeTM/nekgWpi/ix2Nrke+EB9NJXCJ14bxGCrVap6CdpBVhLFbk3ismvEXIsaeikGw+9jx34
IUnoq33aTHu8mN1RRSUCBRfm/6dN0MXC4rqhiYiYVrZT4+WHvzi9+boFh1lO6UFpYYgD3+Mapiyw
9sQSSnWh25mOkRjGXckEQmrjFxx+tUBYU+b4WWPRdtT9H3sMA307TyFdDaleTJCChVSCasWJxHrt
m8TiMwrEcJEUpXFE41BhQaVQX85OnxFBghDufhvinPnvZqrgZCowlUiNIeK5F11r6FbYYnr30wXL
1xk1Fi85gHVE2h5qcGRPCqPVzt4LXjuY6iDHkdKaRrQ0dvGgq3Fmoa092bcBwqyw0KGl0JVV4iS6
wO2AQ5J9Ua8YAgolGPC807V3jG3PXmqaz6slVSgUaZGYa1jVszan6wfJ9h+ETLLREobxQqd59vma
h4miJAtfxAYw04Y/WUAfOnAIBmDQyEFpC6zV1qBHwiNcDQkn7y+BNkjpa4Fbf5+t7ZFeJoMlYaWN
0KOFKy7v/8qsMB47+K+Kq28KuP4rT47dE3WFbJIn+sFDB1gLPYUBwg6s2TroFfzbtWVDWJ+mtCcd
c0NFBoJFSesRqCV0seYtj7lMfNBXX1s5VpaAENQLvh7V4KB+JE1WV3Ma06FMGfM84xZpKb5kkxI7
9kYdZTYVh7P2cfdervcOhdV+vUfmdsPA9B+LXkh7OKWNW+4HYqeFjAZZ/6mf5gmOJI5b6XhisVoj
BZLUv0AeYDQS0Y9eBzw7mHSQJngDowTma95LrBE+cHQukR/XDrG9erP09ftBjIuc+rydHT2K/tK4
q6ITz/C93mfxNpMH0p2VgGAotV6DNCPKH3kzZICsy6kWm2s+p+004VcE4e+P+m30kq19wmk4MfBC
l4j2LOrZ0X7HgOemoABedHeMmtYveKBjecKnDYmYIdpaGzBCKuGykGab4Du5GFO5mRCKsAexao5g
NVfOCiWF7Eopd7W5MNiSWyMlYUD4J2yevndGnsdbB/VWZ5k5pX4tu1xs5ZxgiV5CM8ZrtxkNSQMl
8Xrd5rVI7MJ2hBTYDqZRvhkgtD0itWqldrqWDzrIOvMt4mi3OzQ23otmXSb1K4t0/HUBtPTv3HQl
jlgaUPrjux2pmMONXuMGCqafpGf9QG8lH/HVlEgi2tRkzm9yoMkNwIY0wX0JEmWkghHMRQkkw8n8
SseYkhHX0WeTiXEHikrh9XmwKc9NP5jF5UIXLQfa3hgEPYqOHTTK73wlutoXqZl6qiSGWO4wrmyr
A6EUt8JUfesc7v4w1/jAjD/NFZDuWVSr+pHrokN3sPFvdvd0SAA+ttTiGvx3KX2H1lQPhbPLBJXX
V/9lxEKWJDKs2EVgQvwSspWbqqxyRaORc6Ke7L81qArQlG3uGGgzrBcM2heKoyC1+N/hz/f2D1P2
lcVQ7Hwo2svdnkC26LmqDXabfsW3UYDcKsxqfiNj0+nUK03rUJ2qzQdKYlYADeTuMg+KOYld8Cfe
YTsOnBE0LVHRsgoGL7H5BuLzXr36X0Pc0Gb9igP4wqtOO7YRLZ1lmxgPCBBZjzdX5WFwqrKB6shy
V7HuiuwA06yq1qMuDdLchmjHMJgbNKyhh0RFcXQNB0BCBQQQ+yKlBIaNq8TZ5N/eIFyssve2w5k9
JyT3CsEDDt6UTxP2n5wcWRIFH8JmDozB1oSJtaYddugkNAuhkpsVduW7V0QQNvKEgG7ptypbqHnU
zEDJ1I/0Xg6qhFs3wuXFhDm5+xAVNyafMM0iWqd09Uqics5raUwanlPKK1QU8dHLp/oVVM0SKy/l
OzIPLYRAM3eTDMzDWJcX6tXr8VCNkfo80R4cRSsY5W/VOeCpemFIe/SlNazq5Fqb4SDDHWRqBYHD
RGYdY2rRxwhLPG6KyBL/G5QxIq2KyM0eJzwPRhphDI7PQ2d5YfgNa21/R2zeeukjzO1n1qHWqIJg
uP5KCtXAiGfO48Vfs3qi4PNSZEZrLbsDr5Eu8Qw05VScSWkFTztTw+lX2RgRv99DbPimtIuWZWDj
Ldhj4FMyPPscEn4gNGOxuGQzt3Z/R7msQWHLDVkmzwna4znDk5AaktzEbaEoq42jE0hkWKuW4fzs
ahfCT53usXVgYp2F1+onRm+FsK1XayLskHb56J04GkRbwG3oKBFOFdNslEuVEApmtlbWiSiYwZ+g
nweYqbvlx4+715Vj8nqdJIt9FtKNfnCaPhRYBnD8bL01gkLQ2+rjkngfGeAedvfIClZULEe/igoy
x0TMva7YME2YeHCBvWWTSeRvZ5u7Yzy+FPqETmC3cir7ie+ZK4gPLRGOAzYukZ5vsSnmbPPld9TX
Tq23q+FuLhKM7MV5Ac2wUXMvP0l71FFg0BNezvAb90c+VYqusQwpms/73F2luQPlqdoLv79BHw5p
guRDJwvPMjW5DNBSxEUKCwlT8Y3jDoJ13dMd7cuTdxFAU+AXn3Apb0FUpDPSxlkPPi+aFRT0bz45
jdwQ2TEOC7rf+i/Ew9sLXj9Z4hIHePopkYla6oT0oy+9aCPdc28QXO8caij4imwL8GjbMobucF0y
b2HCLVrt5cjS4ueo4RCMr+gJFkcvvFSFoqXgnirAnRH1s8D2JbazejUAPB+ZerfdeDNKIsb9Iln9
DYdxVa1HPSvkVGUh/8jebIov7gXXJxmt44M4LYprl4F9gjBTn6Eiqsw5ck5/2a0rSkE5HAEawuZr
6gg+viFIOf3Tm+VXVRIKE2CKmHnGY7oAt+C81u79+VAYybRHXDzjAoy5Pu3dFFgt8POQHArkMpuK
DotBl4Kt790MrNfkCpFONugY8WaAUP/psB6OnCVtNvJfkcgtcyMINos6eDpIKZh8RCdo4jWkpLcc
MPs3aQQFpcr8W712lx8t1161LLkXQzMkOzDzCBjDO5h8Cs0KQENlkAZAnaiVruuOqE/+eqcew8uv
7VAgQYJwRWgCetLRORGYTk+NpZfKlEy2c9qhvMO25sQHyK3QOZVzYeaweO5xfjeTbg6+y75hhJ9v
DTMTpiCOiCY5h5ZYMCWmKEty3XWCgmADbmUyLGfRhgXL4Px0tmBx+2won4BISTCnQZR8vufKkfPE
AQYFtD5fCDyIRwrsY/lOS8DPvGmIQRYNle1hyXEtLW8XTEzHcQ3fLYTOUXuofvSHj4ojF7civvci
AhT+VM3AxZAwUAgeBJIUQxQai3IZKtt6HPv/1h4NuGg4+JCc+/yraaylX38UdoNhOgkTIRlfS2Y0
1+k9eD3MMqEHWsZdeDSPS1uoNuQiN0Ir+SGEPDlbC9oCiMRcIXjfsHNDyDWmzCAYrna8KY5dd1jS
SPzww4ZtRsEDaFcjrJK86A9LHVnAE7u+XWOKxqnP0Q+4Wdq88qmheetZBlQVV713wyLFNkng9gfx
ogcHc7MeiJt3ZwvetRRZJChR4biYnKiJEJv9OIlv/KBcHVEgR88SukBMDTxcg8kDtWcal+NnNrzV
akAVB73WYryhwO4eiJger0BoD8Pqz1bxRMPr7uJfGhRqGSDF3J+1NoHI1o7rzSU7Zhu+E/vc6KoN
p+h2EKtIH0k10QI2Chls0rTjUpHpjCpTFgb8TTApk4VLrG/eMWsI3OlZmgQMda+/2yZahDzyUtba
x7kLVU6ekswn6FycHMCFeRBHOExGBW9XwfHJpc4ldq21MWoiH8N1caKbPyrzwAwI1+nsRyrn7a3V
74iIqf/XKlaWl+Pb2FkDDZIN6bNhzSOT9mFZmVZee7ZDHsG6+xzk1rtE/nSOUTYpAmoNLXgIqQYV
B5budrX76lU/R2ovLLVd2d+pRZnv6xWyDl6TcRsUWHmgfmvNHIn/nv1wcQ1eC4aSYFMhFxBX6aCK
/FzV/22ZKXoHdWq7X3zS2ldyIvzJFPTO7dEu6DGX+ZuZ0G6xt3kwdtBxUJvMIW5PQPCfMh0QPXJj
Q9INrMBKTsNQxPhQ2JWMzhMCsJmefnHvLkNIGQeNQD2THCEcLzugki+kbzOOLEgKfMMzxr5RMhDj
dtn+ZPGJ7QSQariC9A8rkin6qFvSjfMz0hwxq/yx5/LmfCd1zLiNqthCXqpztN0rf2P2oESWQYUV
GpCFnETZcD7MGIftD1Mxeyg8ILCqbn+wuoPWKpN89po4Zbgc/RhNezUDpImMCGHii2fJh1UloXB1
mlojAutzNjE9I2U8+iiCVMocR8DgwgNIG6T8CD484qkdFoQ90w/roj++2EnkiIkJTFIN1RIkcdnV
k+mnXxwlB/T7lPEvUS2v1PB6DmUB9Dghw4G1Px+efdf0My0ywwjMUbXsboMPMDHDfnaRQji9DKFD
suYr+QrJ3SxwhjzFbbrEXfn88YF67feYoIIsZTmGKJXyi9hLBF38JdDw01JqRnmqtPc68KZpM6EB
EBrAObLdpDtY8nEX

`protect end_protected
