`protect begin_protected
`protect version=1
`protect encrypt_agent="FMSH Encrypt Tool"
`protect encrypt_agent_info="FMSH Encrypt Version 1.0"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="Xilinx", key_keyname="xilinxt_2017_05", key_method="rsa"
`protect key_block
Ryf0eQyEz5q0PHiHud72Pf2moQtUUOhZ6riqmlBrmM44cxriCmqsFC8aDwpFzQIRVMGv4JOhmM62
TerN/FwkAD3r2+IGYdTHf8K8H5XGRMpLWkcQfHcqEm5ARGrYXo2AjUPbtErNtBTT5qYiLzxlJof2
nldp2kyMH0cAl6bbATk+W/nRIDGNPUlDwdDODUzCZeBzQYe2q4XMq7hv/9U0GDjHd80omKF0uDnJ
jutGPn481O2Ld979FFDva38mOWKTjBiih0UMzpU3aZAvxrv2415XkFWGuXp2nrpieHuqB4zgu34L
IZdsSo1Fb3ZgLoT+mNA/uISMA582uYnEx/CqpA==

`protect data_method="aes256-cbc"
`protect encoding=(enctype="base64", line_length=76, bytes=125104)
`protect data_block
fJnvBbEWPJ1o5PiJWI3nsHHu93QsuuicTSloKSQH0iTZ1aXJhgu6jmwMBwzWt6jx4iB3zORktM1t
5GyJXahx6DEX2LnFYgu2gkB9gO4MWN6hHOs9xo6IeWDsFxwGMP1VSoyPTwD5EVSePYgJh5i+MFTZ
lh3upsXAUG7EbReWMOUlHUdwvDFV2vYzFnELhk1UoN9TT7h5nF6iCorS+H0yv27i9jpNacx8b46P
wHhIs4KTQXDNUhr7DJrL4fPrJzK6lx51KnqPVl7NX4xz+Jj/PQ9Lq4DKX56IHnzqqsyb0AJw8pfx
Lf34f8+w47RIM3/m6ENapjGwPO9XIz1dmv16zieIvWQyslZL7+U4gZyHUkmhmopSv9O7mQJwf3ex
gdCVEFTxxzkZ2MiSnwjeY+UyWHOacRFRXd4JmAyVN1vKaiEg/KERK2A7aGriwkHkAH5rK4Ef1HGc
/Js/aL5jdlSCCJgOA3EzPUOyAnB1JBCY/SM5xhlXygcIv/HL5T7cvwRrqlr6ukwSYYMmahmhj7Zt
sCVfeSY4uwiM+XN1GBqSAL2Ix7MXG4HAjPS8fT/yTCXbqKluz1KhVv2hnlYDS9Xyxjbzk4zeW1Sy
s86PM35xYHY3W5cTVKG4toEeNKBBXGcSJx+xU4fj/7d1vzXLoxE8YcEUqVbl2rlrqottLyRmBHXT
N0a8LpB8BGtgXvhmauCKEo6tQYGbQhIrwsKq83rAbi/idkl/wqA+X70h6k6z0E1d24uNTix+AW3V
iPVXCQ28Ip/q1z5xkcRS3DJE6CPKk1g1lbt5pRZeXW06+3zL5qDNtydj/rh63YY74VEwBFcVYQ9j
PeLt/AS6tmtMWEvgVJ9mzi4R7O8N0bS2exQXNVU8kLUHy0R1yIJ5ydvgOQIpyqs7B/TbEQPDuPUv
Q5hkDFng1NCWAJ5HviXI2iTAWA0m9V55NFiJtUdIW7V37UIjBJUfqXQa5Wh8P5ogQ30hTUsGysC1
LCCnWgIFBsJjvacixYhXZ4G5bjXHXsOygXLQT6CQF//CrGAreVTPGwCj3SdUdGdarUxHnnkUy4dz
Gqf9qASmxgpkzrAmWN/sWwAj0Un8uSstXGeZsyFV9rYTeN5t6KC5qmi5lD18UXE8Ze1Ij4F8YFxy
xHyP4AZBFwzzObaMR/giBlRpd4QTsnSwtmKkiqw4cCj5pU9gS0efAcU3bGsRMPTM9szU7xld1OMc
qp/CVFvK4T7mRnWM9X3EamgQkL/t6C7SVkn1MixyAATZbRd/shPTcimQV0V5F11njf3mkYOoAVth
WCFUp0dg3/ZGbAxTFuqYktrr3yrr40OrlUE8ch+JPWZhIUOd4byCC22j0YKK9VuiNx8OzW95iPRS
w68v0DlhsHAOl/fT9GSsqLK1SJ5cns7zHsVH/L51Cw0fxr9gm7eos4Q6nTMsLOIsY13oDbyBq5pB
Irb6oXRNzasyOyNPVbCaxYzLa1Oojj0I2zLYIRIGcTUrGuGmT0xSI986sGmpGf3Yg92QnngNE0GV
cEfUMhRpS9kbwRsokFsDyIzIwyy4QfwueBl37uoKDiU2dCCAEZ4ZEXYsBqM4Apy4qKA6nEgA7rje
zbBelV+Ekt5CMK2s7ESqX7BctcyIambVgU6gW6tfrfmweVRquO2yrghcCvc6wi+li5zxdoHQziYA
RqYghxcoSdcWz9pEC8ir4HCAJmA1TUXX4MoImorFoYZAPLol2hz3ZghxbW4BrPMbM2iTi96mQj+C
CcqHkZaOBqaZ18qFzJhJ0xcPrPtcRNEiOqY8nGPC+w/HV6Rwf/lEuNhIrsY+QNocloP0M0FsqUFk
bYwyyH0f+vFfh6hVIgj9wxyVS1oRLeRSt/xCV0Dvq+qOx4zTTqhn0Ap7tLEsM2TABDSGD+oOeJsu
yWv6Lx1B1p2xFAhqKr7sQD8UxzaUZT1DIykTBOsdekCiCFtGcjIsWofFq2FVJCJeKw4RQ21iK/yx
J5Tcie02uGoLEfn8Lxi0th25r2G7T95mRXNfTnCR5qqKiiKgJdgKRzsvSrtLJfIk77LMVZNNR4d0
JpB0JHL7sLh6eYVGonrDz1IOYelSL06n07oRiyipbKBpNW2/sQDx8cu1bVtScsL0VvoR9QlxyXN6
ofJgU8cahRMesxc8u+ZrHX+6oHUcuGAG1EPaZm9wVP7iySnz3Z8U9oDDREOyy+V9kzJEyul9p2H1
0IyYYzCbqw3tiTy40ZwdvXz6qFBDQo74CkUrhD6FtimN1FKJcPFT4mMQuMu7y8G65y3S03fkDUxr
P7uQ4Lu/9bN9JoHBOelZYszQ/FfgqUVxkAiR5DBhkZ5IW+PQPW+VH8fI4a8RPoo+M68qROlpE8Vx
bzIVzCreXSIIXIAzKMbKGg7bvNt/FcdJ9lCY5aF1pXO3981Z55hsXXPsITluYAWeq7UtdZ8uMNiK
bFQN11Dt6GiQb0PLuQLxKN+cPiQgAWBUEqfzxm4PHASWtrdwEo+PHz4GH4eyJzzsDBvM8UQP9aKj
NBa1tOfdavBGZ84kSWPXuzf/IFr8Y6mx0H2cMoHVW8iTkFxwOdg6U0NagOFGECdkH75dE2g/SDDl
Wb2vMFsb0HN9DmGlEjk+8+GPUmDhahIQrw2HlBHtCY7dBISoIp5uvbyr7CQtZ7/bimjDUfkVukBH
c/X551jH0jDiyYT5Q3NzyMfAz+QZDYO9SUSRoo94B3noZKFSntSOHh6mUX7A/iZ36hN84zhCm3Ps
BgUmsuFy+pJaH7E7m9ddWdLQ8HUuEVGVzi/jzlb9Wad8zVqbmu7zQBYEMcg/3IeK9RIYymvLuA8L
5TWPpexXF/dLV2YvD4VsOdOwc6qpq6Yk8ctIac1NNxVSfc8ijiLjNBCrLXtnFwU0MD9rDpcEERlu
AsrNPmkTyK8V/am0UmP3CfqJs0BuIudcrxDFrW8V5yWiNAxXDaZzudmATz/Hrxi2H1UBZ+CwwXk+
x8+JderusOtMFJzxjqbbpNHaofcqXfDNoX3YXrxzdxvnQ8NdnMIObBlZEjfIplDvr+z1MUo1a6iB
X32QLSzohm1UfsL6VM3/gOMioXbe2GRCMO2C0qQpD3NAu9HHisuGDoAhgBzPMY8UHozkYQthoiTu
xZxsOR6TNlCWh3B9PS5iGDI4+SE6PATo4XFuNUqgefMYCxWQp7AbgOtGqTna+/STk17B73PgD8t6
zbCt5HtqIQ7oLMW04yZkL3drGg7NcyfxtvjpKasYoJwbkDoT0onTN17P+r5Rlf3kBUwJO7Bdupa6
G6H38wVI/F/7dqUXU9bLq40e5g7TH/q9ouWBAKJK6Y0Q6lOwfzqj8TXFKPISaNhbgu/a4ZkacnDw
auI2vO6+PryIl7ig2dMZUNOn/T5DljVOKTj06M4d/OPN6+AfF4t9LM1XC5CJOqXO3w9n8p1uRPrU
V2Bx0mRIY8TSwKDcSUtLJTAGCKCKySKokB/HvmvGMvtiE8oARYBqjrJNtyhYp0XYIsvJkQlL2+Un
+m7+p23hR2yy5VqDVziLtb2BSM84oL2mYZNReeVm5SZv73Pg/RWVqRLNWZbNJ2gSthJkED4C2Kn2
efvkIEzS37w9NmcCYUR4e5O8NOYjTEr744WMlS2HjfMt42Q/Jkxx9c8y0LsXkRaOQcw3lUTUd5o3
0zDXy4XXzIcl9DvI6F0utLeaK7IHtgyR0RGDEMZ4lnvRSGBibsseN6KN71ourSBsIOZoIFVXynRb
nL5WbVa+vxx/SyC1w0oGoGVblybYS6pPa5k1rYHXma7Y3JIZwb1Rxw2sVNyKBazXDp0ozChK1jJi
/y11321RXoSNw8CBh4KTNx+eyeGDuKc7jtbwpfYYac5ig/spEUQ7laUNGRH2f3lxSj6UEMXW8Un6
fVfs4nIVeE26DvYX4sa++Yqs8+Wfy/DEkoqqZDuRL3i467vrBCt6/9CP9zAoK17wVm25MulTsMkX
DWkkdKqbgVUkmiRCygiI9Cnut+BfgCAITQ7aZvfq101g3IzRTPMGDmjc3THuFyxeTsTL7MpHLVX6
/Zhnc0Zlqpd9B5x+ByRPmQfg/0YUxqw3iCbrs0q7TQsorbEP7/WhWVqsfne6CoZvuFDtFEQ3CGll
g4HvfgYOeWrbUEXdmMiQ7P+KX4OWtNjB0T3shf7kAt72FZsae7JSndtRqbVmQcT+CXoogm0QJ//f
BCH1gLY4UU9CJiYxvEIkqSB2TJU9+mueCPWWQSZ9dwxR94kCCUsnPDRZNtK6msgxX0me+zybG3yJ
O9/xPzgMbMiz9ShhQKHnHpIl5AayADh1sAWqJqESnhIreiw6MwJw5jX18pzsX5Jxo93Jwt+7bDjg
XJR+fcAYTAeDshHRUyzM8Svd8qhSCrkrVaK20Rwp6+jz0VF/CcXSm4QWswhgHXzJkRrxeIgZxsPW
L3zt2PVb7E+8HsBZ7wHXTNTJc/RErUDlIFoo/d8DdowXA3IS+9C/yjAcHGgN5bfg4nWVUxQDdRXy
zj8zGUiIvXG1fXCdDDSSJMOZjAEUsidK895NP+BPIkNfqAp4vJbPgebOvJDDBuJzQ7fNGoS3luHI
tNt4ImgqFBcM4g1ejrAUcHPDKg+U5NMriRel2nP9dMTzxbTTpC/BX7T9PilCb4AkNTmTiiLNaDpY
ooPf3MdRQJO7U+2Wep//3iZDD7ZPPBt6xAbctpCOUkYcJvBCH7tzdme+/Qscjf67TW50t0eUw3YE
Ups2OlL/gZ61AthL6Q9iYaeaswSQdRSkONQJVp5wXOzx6nwYdITWUcR+jmQvlcc24n2DuM3D27el
N48Qh+kSDHO4eXGLO5yLiZD/dB8D07fLxX8yRLmdIvOok/+Az6G7tCAa+ZS56LA4izce5k0+9HxE
Kl2N5vIt/FxyePXYJRlQVs9piwLzaaqjWlmtFLqrio5xefUYNbMmCGk6vFaE8ykMOf6MsC744IZ5
ISI9BvRO9yKsLEtd9GhwKY3i7o3d5cF5sWVw+n/OdSGELvh047yykS64UwnxqmVr4/G4Wc7GKHm4
Nmja3Pa5SD9ex8l9AtMUU+bMLEzGGTCs3AqDAZwITBjVUBODuI2nrFQfAq+DmedeS7NAvUs7RVfH
vn98pxF8tPqqzIIuBFk+WALUGjD2mo+F7zGFHd16yLdLhUjqvRGeYpN4EzKwKxmUsWAsS3a4Y8qT
4yTWlz7tVCKx+8vxPpX61AFGqrGBrw9hW0UBjmoDZd8kiF4omLx73cpj+EEJLFleKxjd7sGd7yvy
E/p/0rpuhN91uU5uasOR0GGWFYcPJdWoeib4daF6uQ8hNNN8MH6eFTtUKcOCF3aAq7XU0YUPrqwg
OSF7/zd0PvOlgoQsCR84QFMMImhSstotlRYI8esNXxnOtnp0/1FOPpLs0PZGPPTF0a80RQ3Nfnw/
Qr+b04NGx3xGmaQ3V305hACKfNa7rdi+4AhrzMN9krnBeGejWLJ0xhr9kyADpzn3w6Dx9YCnGdjA
OXrhIKhUz20P6WhaVprMzmotX0ntJufMohYY47fItMP5/wgwQin1EpLTKFiZAfiV7VsLBY6IOK1C
Sm444ePtwsyDjfQZRODQaF39honcgLQevMTN2IyMeICi/CPFb33CzjZ5SU5IVVC08li0pa+Jm27V
J1mDMe9YeH/uts+pNDIsk7k0CgASWZ08SjfvQtjLTnK5AEzVTjG+3iF3acc3CGxzv7/IqWvLPXpu
IfB2qxauKv+psos41fT0Q52bBG0+xmwk1JtrywhmNzuK3iZ9crIHFOSh5FPHftJIZO/PKiqDw3+D
0IiJa/IgciN8V6fefJy19d3nUm/icKVlOwtPPB9lT/NLpsKiQCkkQu7CUHZ01hozduhTusTwKccA
nClaMICT5wSBEZkeRo178HlHV2lgZcLSgqcf6oi57DbYZErm77iOlSYZzCLV1vO+s/g9H0tFkY0m
irgqWP66y68xt2b+PyAjWQCgMooqDnoCOe0dShTatw8QSoD2ruLIvxdgoOnaOfo8ILw1baJ7TAmv
ueROyXvjsaudiVjb1+CDs1i65kYFbUwIyxpzQXioW5tw0NkVr8yKhg06KTS1GjcKzy9hwNCvCM6I
lT8kTUEasYufhcSj2SrF4Bv5a1a7gCj2Nuk2TSgbzKsib97KCQt32o3jTBy5gPCu4OT97UwHmPFG
vWQEUj/pPeEOqLScPGZUQcaCl3burRFfEGI/E2qwBpXmU4K5nE2NyAKJ5B1ZubfnGsv+peOWptyN
ysF6STwd6FUC5RwPy0vvQF8bpD3km4c4sgr7HdnzBEq4WfIu0izT+JTlrJiYGxCyLtQKG/48qrjz
txOmaBe7KRPAEhFtvMIt0kCl+91yUFmDjP0/f90Ia2lo6zWt2Y+0w53QPaUfmeczJhElIcVe5L/M
ipXYzXNYzPG2SClm+mKms8VcC9z5sEEl57m8/lGu6xGm5CcZ6PPI3SZ9YHd5nKi93F0xvRearWNh
WR37+y+YOhCMiN41BVKNd0hQ8pGa1h/9fefpzaJBCzmEnULL8Y81BLSGm7Ggi+AqrAXObVaKMWa8
wmMaEOlefXruz1aEvUIAFzg0QTvdnKvafQDN6XO7eqhGIjiCUkVPZCF2xklb8snJStCRhJ/lMN/E
7RRmXr0T+9G6JwiIYKZBXKTEbT9Ip+D1zVogZsZnrR/DSlTagpIpoqNBG5YHQRIDw214g4x2ddH8
Jjp2b3sBn6ennMGSK1O6XHM6H7JyNEpvJ5WckTob4YFYugk3fwEqe8iDrRlQtYHoSJg2f52lf2eH
+Vwpv2D8A1Hzf6RGXM+42MYrBuhFHztbYxITNRxTVErXFQMv9I+2xTQflrD/ZfFUmXcrBAxaoXNo
N1B4kuny9Jh6TwAL8Oj9cV+f67i9xYnMMJfYY5h8PZvRA7cEQ6Xbgpff6I1+TeoV0SnJwyr/O1qO
jLmUmZ8O3MccBq+BXAxFz+/C/GhGQ1+l9O3ee/WNqo6Cys4vNXqRPUSPDa+9DWMZfsJr73sCPv02
HSgfarSsDxStgSlINwnNCnpJqa/cD1guJUejPYR7usW0cz5wIAe8lK5SrjK/U7accan2QLPkUj+a
xKYTJK4GAdYbOD4Zfqlv+VUCLulJXRjSCkxHO3aiaAVbTS6XFujKMuoW3fK94BtQe5Z+0DO2fiBv
QsjcBQsLhkuajMz5+zU9e6YEaUh0OOHMY138tE+Hm1pQwaFDV3AOi3tvEhFjIK22aFO3qo8iSB8q
fqEG8PZnzQDRRR8A1McXM6Eh62Kej5lYl/WQOGxCG6AZDDX+HoKcWUvZmkFRYSjwMXEw9+lQg8zC
wVm7Nv1s06Mxh5jWFo0GJWhkCBx54nUVsODsEyowpLTeNfIbFXS43hhTAcQ5xyUqJ2AfgJ0x0P66
Y2XUbHcZCp/RDHQO4N/MRtPUjD8Tt7C3LK0dtVNozrErllVAY4lYe5eJupgqrDt9LJ2Df7pg6nXk
axBmjt0TkXnQpjbATZRIvv8WuehSx24VLPaIBVhPEDye5abiUijtQ+htXbWzGB+g8uhvy2pW0oF7
V/DwcApeCfqZr5akWlC4BL4S3Ca5pN5Fkd2NhZT+OdJn4vnvwm5ZhHolBm+qgZMMssZBclUxiUiF
uVTbTsGpQaHJl+Ck25iZyyUizL+i7P9mCOFKycRHWFWOKxJ+92abCILBB76dDZ2mKxb3gHP2CAbs
71ZWa5Uemefk5k38drM6QFh/J3OxpHP+vzdydakGBZS2kjGZi1QbO/xnbGAVbpQyVjTI2coMPA9b
D6MdGajhUOLGTPZgWmFLsL5TO7KxDetjaAENhXkhpbsSbFzDyoSNkNnVFaZ0RYaXc2ODN1CKb7A7
GZKSVSkZM2hTEkn9Z+c5R3FBfhhsFvwbrSKWLrxaTc7DE35rhvmV5rG3uSy4spanxa0jQC9nKkqg
2+GjrLtoTh+wDCM87yAbDpC1zCZ/EUbHk18dmMNqz4lFAZLdc2OfRLbPJ7e1wYdgsi2DTRxsStqS
o8/mYyK7KHt5KdRlvLn+YSRuiwKVIPgJ9vE4dNryJe4dOSgRXbxqZl89SyMbowg7iVTM97RJelgT
3/VD75t2lNo8hC35eOOPk9X9GVoYJbTcum/C//KXW9lv9pI/paCesL0tJQUHljlNv209pBy1h9q+
dKJWkdhg/lY490nBv595JRg9qweO/Pg9eX9BvSXVLAjaE4Qd6DulMX5sJuAgJnStY3/kRHBWOO7G
V8sc01F5YtyA9W7ejCbN2kCU0PnMshZfI6s6NQ1QgtSXFGE5LIpJFR9qOGe3314qe8yE1ZZM4jXY
sTp8c0bB6cdNS/Flpk0tik/TB+JYjTowCh1rzdZSDMVpXcPXl/w/YNjGJ6MadVOb/0diYO2IrsTa
OcTmYQLC/aoZqBORC9FTYwQqpeMce1rzHKaej04oo+JOrAFYRVKsy2NTpm5m/cRvGdUKIkk22Yfy
UUe2GbIK1E/iP9dPYv2S884nt3l5BBROn/M18kshbD/2zTIaqFdgxZwiq8tgYWxDa7F6SjWSY49N
+asCMw7/h3/0qIZUg5DfIHPD5H5QfgkhDkWs17kuI8eOaxYqgxyzsgzRJycHv3CGRv22Lbl0WO3b
96MRKuzhRzr6pDy5KiCY36uGYdum80+2Unzt3yXNp2JTQnvk0h4FPAm/W5gFdK/PC0+6MKbMzJYt
yAnGvFE00tvkpiMQmZCN62EjAGTqt4sp1MqBbf570o2UidNZHxFzgYkRtF8v7FRD2dAP4WIimJ+f
Z7zIWbiaUSA/2T6x9ZRMYpTBhzyFXhNasNw2imIv59xOxmrymMuDhT9whDR2MSwOH2gLW+ZtzrD4
MOamebdP8D0+pxWp296Yj1LSeQN0sSaf/o6s8kWl10FIsMw/r9Hj3fQ4K0Hq3u2YXS9RT3YsZF4S
Wm6OU2MJS2OoK2lEWTtWc1V/tjH3jTONaav1fvlDyEjlGeuV/TJ6lDbA0AUrqwa5lMHu9vMLaklb
/QoS4twjqqiQ7LWoB37TGMVCafX3geARwejgbIq6EErmxNE30Bfpbx9gH87o1tfyVCBOJy+Sdunw
D5mxVtBP9Zyxodxw5rbIgAQvG9tq7In10FtNnJDsCkp1f4UHofb4m80zzKCCTQ2omKLC3/qNYnKA
y5RC1JVXiMC7gcJOoUVL8OypqH3PFue1BYU6IjlBwa6O+57BqNP35IcME5kSjC6kLAutHgLXrwaE
gzYOVjTiZab49SGTcrLYpPYzvYlUqo2ssuchI5cl/6D3yae5P8K7fKkE7G3uH5Assu4l3OV4OpbR
HCwKVJLoArlA88KtigR59jbPkIdnzX3w0E8SNrQybLFu/rvp25Nk27o/F5yv+i6q2cqrKUbVqplK
WjIgmM5xVwydxaa46fvffz7veoMTJrmdroPobJZfeoCMYjBjL4a1LVfCBduFhixmOiqc0+aIv9wW
9NZa02GTvpGiGxH2VuwB/8BnyyDeG/5ZmFyn00XM51rtEMXGsoxcyvne0P93IjdcmGnFfWoo1yi3
7Bbr5dC8hGvQYpNKcW+34SRAo4oECJnAyxR6faRdnObh656RP5ewK67y3zHvqlOVsmnfhfGWyKCp
gRMBkv+8S8I+REtAuGptb8iUxzJbKFocxclyxp0i17kh4yJCfRTbahBbr9pXy8dneJFY6bjW4Grh
kBZFwRbRHsLQ0cJEnxn1JtRI2GJDvqV21U9+yyNitVig8gDGL3105dMU4E+JyZ6MELfk987uXksO
FAxxoa2nqeRaBzRKRxgkEh4xz7uhXTcn264ou10O1TnLeMRiuxW0jb98Ti41DFpbuB8ilY9ZvXtX
3k7zA44GdGXU/uPQ4idY9Ayszefv+kFmYtt/fOVZJBYZSO6Ba4pWlZ7Ea4Kib1iy/TvyIkd1DKw9
1sMx7ZaXAJ4T5FE8bVjp3UQmhgd21V5A0h4wh8a7vFxKWBT2TQbFRWmr5T18LfHjEKFlsOp809kn
sXpTj4whzxuJbTx1ZDV9QojUJ6harDdNm0zY5uchAGB+k/2aQHEArnnv7acfNBxflmEi5FNBiKGy
2/dgqUsFPk78Jyuk013dOKTzosvU/RY9Xm9ZqW0JjADxK9Rt/qOolfo8JXehXx7sFrmk6W1enRpD
cEgDnNlXrk9UEMCHsN8aS5RqTDF+aEnhXOtIH6u4mh3bULLsdf/R2CVojCHXwMVqDYqtAVAxJ9T/
76u5UZD5/d8l5zjyp8cajUXJNILXwD5fpnWii03IRtZ0qwy+FBapHQmSwEoJROZ6EmacpbZELspR
rO3Q8lrpt+vv/zPJJriZfxCUiNj5/49hO6sr5AMDCpWzfbAs8wzjnT1w6/PKVkwINIWk3mBZ+tdh
lPjEcQj1Cggvj1Qhkw/DuduUZe3wTW8NKESdtEVK3f9yhAaEQbp/c9/WKLL6OPAufb9cOtrWQ6JE
rwYkqi2WmzYTsdrI4BRhDhllqrPmEyPE4cJylAw+5mJw85q6AmM43e52oPD2nLa0xEWSwr56LsGA
LkY7CjEUV5nDwjLIX+LImarpZWtJR1dDxtU9q2vS+xqLQG/N0JYaC0tD90CvVTmavuIDD/cm4Y8Q
1mmEKd87OBGLarqWaNrgwCoZyqzkd8WSZFZU3tuIawGa8SP2tVYfUV1xjVMdv+EiFfX5eskx2VoK
eu3cALVN2ugk+4umCrt9hB/ekxHf9UdwayEHI1diel3z/OehGX/ogyYJIHUAGYZWzrdispPLoikE
L8z2Tn/wSl0f6NA0W83NgtV4ZJdILIAcrQ9Su9pd5ngt9L0P5Y+bWWOQ+XxxIxPzMKq06q5Dr1U1
hyn/FUr6lzS62JssVh5JheAYgu93ZC16bQphruZNJ/OxnFFOXPes1cGkLe8oJOALRAM6Vqkkt+Au
6ih/Mkivx32mvjT29N1DdrpsoKrJ2KTgaM4YUNV3gbOvAVZRa3+ctYXXZ/QMQG52276wGzIN3OzZ
j/Ydh+oukPC3AxAb14wwiiXjcRtI+roKEWonFfXsfZGH/xdtmSfC5ZtnK4PUFKOIrBAu0QBsV/pK
G6/83mk+pimh+km/hhNz5YJQj8wTRvm8F3RBrkcdApZEv6HrJxA4fgBl7IpiXoqqABjS22Zg/A+H
RYZKgvWGeGlxmxaU4JvHiEDXHYmgqj+p1iT1AihGHsjsDtkM6K0e88G6+wsUIE9YZOzYPuxbQYFa
APtj3gGtghHJG3ONSgBgvXhfGurzli+33yPvBMvCKWtRlH/Wirl1aG1hkxWw9bitf6N6JWH2w1hl
B0u3I5U+KTCGR+iSFDNiWCQuL3qKIWozYQuZlNR4hHSNutYrZ5YrrcQv9MfyOPQjEj1bdZdPmDgY
9RBiAxty+5cMOqyJVioCEwY8gezJQkGioNnZVkgAoT+JZdmOA/9yIOz5W5mI3BB/EQjtQSOWmDhH
H6bEMT+8hWXqiKzELh8LVcUVEpHjDWm5+5HlvaYvqKGnTjy6P3eTVlhTtTx0PUwm36B530WcfKZW
M9AAhL6doA+z/YUf9sjiexxlI7qt5dP5f4I30WxAYeJ00rWxiiJCHSCnF/L8Ew+qB/6xvawiWgaY
uTYfN+zHBrOcwHNCM9Rxux423ZSxNZk1LWzqmw4lq0G0wSmQq/BhEv9xL7TkWdiZM9qplvIwgpwl
VDfUTLEm60ImlnJfPhu5WLhLEJ4DfFAGGlmKBpqqsy2ooYdH19O7vy8ccoMFmFt3AdR6/BrgUN6U
IZDKdVGP2vylPmNES6XRWKpB8SXDFKnOOANuMbhoSLWiQuDm1dz9FIccGg4fgRVy5MsiFZERP6tU
2lIw93l5XaTxGrkGvy4bJ/+frCoXZB4YOZGyUPSu7C/DLzo71dGvv/YA/1UGbjkO+Zhd4pOGZvHU
nitLMC02ke8yMqoNAJHDL9tJbAD1pI4Nbp2BdNXxL3eccs+g0HVe9GlAEmNO25E/hHcUyiwjGyUY
LIPQeIvf1XMb/4JMzrnbCSuptZPhtq0hGO16ybOGZveE6WqPX0wtGs/0UCxSkKzYEN4JrbraPePb
RxZnbNs4vRWZaRnBfQqsJ4heRBtpSeCz1J0mytWn7MgXrvON9tG61b7uvAZH1FFncQO0mSWAeKgx
POYieT5pwrPjbZG/6GofVrTScx6jlhndzwRirpshWuu+LiZaVh5/VuUlONIU4zo1ZMk0BTjQGCs7
5LPPjlmF5trU7M8AhB0gCvCngGXDZFO1pqgy2TCgxS5fcOBKwRzKjWeU34u+7Y0nvqhq1spmN090
GsH9eTCgIV7eRp5RiUPUDXguEjjGq6oj/eXC8gf18qG5CMkI1jg+qUdSSUwiwsT/JZn10p1SWFgm
Dk/wq34yl6CZSeOOAX3MAf14IRsPuPMN0pWCdT/m+I7Pm/FVPODHKM5b7al+mZoSEbwCB662a4sK
SYms03AlpBetfgAw59vJ10mGaPSy5aVG0DXV7DkqAe0KJX+MC98MBFboSQYzU5A1uC0JQbMno2cj
PgN0Wo53YoV3IIxYw1TafjDoZZ5pZSowhKEzSGzT/G3xx3PHOwXKm+mO6AiLaTPKWVoRaVgVwRjz
c9i3/rljF9zKngqskToan9hF2i7FwDtkFbDBbT5hy7lVrtNARu9Tsv+g4evRzufqIDPGk12+E3mS
oEU3DiJ6i7p37y4/+F831ecllf0tPAiVp+MhLCrEWZxpRKjdq8uJBS20OqqksjdUQ8C865gqxsif
h/AjbmVmrWaPU2MVdyahV1oBszT+1gs8TpsK5wXHUYN6qi3eUCwk+fKIAcp1jeH8j2flQUR3tYfa
jmwT3YIBQmz2H/vtv5AjebVAnZad6lTfu6pPaFq4RyXj6WXbTGzdTGqHru1KkCG0CZO4eH2oAIOL
wY+I3LmgL378dL1OxewJrsbqUsv4P71yINgZw6Ms3tNJGb/Y9vAiG0qY0fp9BxVYZjrQRWPUWRvq
/g1JHDzuo0G0cDdk5NZMUEdd0cXVej1gSOUmdU1a9O9ETjVf7DbcCYpRTIwIFVU5hT6ox9AjShZ4
56s9Oijnph1oDnNAkqP+1pAaCgVeN2yGWXLgzGVGT//ra7ctPj14WOR2Gz2YAiqtBHkEO8pXpWxG
o/nk0n/RSc/yq7YV5aDO+TTPv1StkBUUwd1uoLKnF1wWozSyXhCpjI8JlxODknQIR2V5LJKlsZFj
Ud/cYAqcByzSPtX9NAT0niwxLUyAcCfYxp3TcGa3+rCrhY8KLOe1XyswBGGPapCv0/5KJKDaJm4O
Gts9nHKWGK0/7h92CPpygPfsW9Br+7Cnd8p7VVOWxpn780ugF3paHzHfNkW40AKWOyMHnNrFE0uY
ZZRKu8uMa5x2Mpzcah+0YiOL4ka5Rywx7Lv9YaySa/b31gS74GxM8EIgx+C3KDidZb71JwUBnYkj
hjwxfZKGP+9KatoU0lXx+FxmKDdo2H6Looiuq4wBqLywaTkL+6Muv8wvo2yfGQgMY0TUY4Ri1gZi
S8cOGsZPgUTNaYqaSKTFT/8JiUkTkewVf93eWnbvWttLhkt2rEIlHcaodwZTSvVIgZM8iPjQa7Kh
efkr91bnVFL5LWowt73OMsz8HcBQPPLQd3ESefaku34fZAs45i0H9yVYRONeabWOFcin6PkoVj/o
1Ld5vkUoQ7dq5q6FYpYg2BUneM48b9tnF5jmC8zEed8oBqmXJ6hrSv/kXAxS4TELQg+2NMy8X46e
0KHdo2j6e7My5vjAZrRs19ui5l+M6+8Q7nSMk0CpLyxAXqtC9E9CbY5OKwTOx7STTc9Fv1Hv+J2G
3G+9vDiazWp9QwGNWXprvxT7cR5ZC8xTF37L8zxAh0f+iPKrn+pSC7Fq7/7zS2DanAjrW89mf7/h
jwfsLqZAmtsZtkBCPr2dKvLLcjdEjueM1DKxt2pLlgz4q7ke+djW1OTcfabEnCg9DKs8K8DZs4Ab
pk+xxmr9d2YkXEHdv+3xtNxLXNNMCRp8Y9perVSSin55yMAPS2uihn2eI1GCGRsUS8Rv9jkPG1KQ
RIk6Chc9unVlwyMacvJHcd2JRE0NWan72TKv1pVqkGHH6AkupkKUPEgVeXAWLzK6qa0FX8+/JUEw
CAxfcWelMET0dd4qmW/oX5kVWaDTqihySwDZkxhkuu6emKiJJ4t+AlVQaBN/huxdaQLIRJ/QreQi
6GKY5AZedBCM5se/xa19Jis5Yt8lSJH8PzzR/5krBH9ldRJUTcUQbo2omSIhQeXg8M2lbvqFYT6D
I2DAiSGuKhbTl/8RlsbvekkUUed7MPHO1Vu6fBgF6PvW4uBT8HsRN5wZ71EtAchUHxy3Gw5wgGe3
b7Gt58S4u8i00Z29qNbWUVmDa5vnyCVyLltvQErkXKZ9Ic54Yt60fWgkN1lXlRjT4z7JTvyDYhC3
YK4RTnhkXQRdiLWp9lXjumXHAXBhhATcq8yZ0ns8hHG6F4e3RO9c4VH6n4UuvdIgoSeVpKozyXh6
8hD65OWXNU4mA+WYMwGx1lF+scyNVP0gwciUayzckBYbEAyB7vjKKZ0QtLfSh0RNagdGxw6nSgbM
rfoBUdM1FQPwwcXzwe3oM5zMdixI9pvqoXVKB1b92uYOCUzTjiumRFMajHGbd7THvHQ6XqdAvPPK
3RoD7HcP4f4ICtay4syDraONDYx5Epbr+bqImCW9vR9NeCu4fl/eP9//jxZvebbFkkusolkwwmE8
+FKOWEIkOP58SFCPy1HdRFdhzy5rvotu69U4+AvvP401ukQSMexD+ZSoYzV2SLq13BwyephXl76t
E3fXJDOzlNCjYHaS8OgsGLvNHBDtEbrLBj0iwpbDZcO0XwNyxo5Tvx3paESNgv0XI6w/UgZh3eap
AD36e1MlA0Zgz7cHGcQYd1SoGLvc8FEFqnVV6QPC5BD1f+6KbffELUlEgZi980CK69EKCVHJ+GK6
xeq/qkwTf+T/AqcjZoLNvuoQFLV8RKmrxksPzQIrnFQ5H2b0HYXZpIItojO+x3MJIydDW/hBRRdg
Chnd0uP8vY8Ch3ZakVs3X2jq0j1so50wN5Y2vN+SEUgzpICbUFtL7Qr61WSLm6lzPJWBxotP7dot
Edos/f9gh71vySxcAsMBvQqaaQLnxoXxeEuv6Lt0e1JFGGayoDDrzrq474teTUBcdyjsPackoETn
qri2ac6hyOz8PkYQuhD80AneePbDxKHVQB4Krnf8sKbMwtZqIlJLS1u3AgFLnMohYXML+tBYpxT1
Q1I81997X8PrJ4bQBhtjITyFqZW5AQ5/pa+ugMhFBoftPVL5bJYcmudrqa08//B5/9Ark/G3k6+M
QLqceseJ8JJ0uOSi9+7bExCO5a9rGWIO5fd31TUQbFv3QHssS8FGESNyd7BIQ9HMiNiOgEtrpX2P
tekzaa7kmcptDcowLJEP3EmNrhPPwKwmis6hx7SM/TA+jTaq1Xqz2qKQKNZQI7pKHrKjFXiUGiwE
lfjDtNSk3bVzfNSaG3qEYWEShIagNNk6nx+wTmoy6LKQQ4SjbuZWy+m+rt35usZw/4GSawqQ4Cn8
/bjaPnLbw9Gvx+iD8NXkxTXBAT4h/zjSFsOndF4xzCQhi510tEoAm+Pl+Y4iNyFDxmPchJGg8Rcj
Y273uomo7sTymIiL344T/pqojwQkt+BDJyOc5dOqz0TSpLHnfF/wTnu4yq/Btyqp0oD/q4rWRSdi
IYfnluhh2Swlac1dXtHd0beVftE84qD46Rl6q9ZMUGtYSRfx1jfCtI7M0V/txCF4Fb57yG9woo3K
FnNVpOj00dOJpIAaJPz0sm/6shkt3DbSZe55lCQOBbsc3nG1/zGQDRWBcdPs0atNZ4NrKG44nw02
r7E6IFZrGnz85mbukL9C/gDgts20BZ7XqfvTt05fVCkey/iIJvOob3MUOkjxPRg04bCsKxDXggtc
C3fTAgwwvvt/ZgqUdDsXgMvidNV2txhY6VUBVGWidtpUk3xRRp9k3NxgzmgRVjECyu6IhcgX6wii
HDhjlx69ETV62mm1oqN5ZJQA27VPK6z4FbR/JDDY+bmnYFiQrFQOPWDAIXv/verXTmNipC2rHxv3
ykBTGzBn2XYJ4vDvDqhVMElQxQ8MYMAn8YoQV9KAi7/yPMSNMhA+JMtT0wpuDlRLHlX/5sPAE81I
OZLXsG8ZpVK38C/MuPrnYzgXOhnWv8kYpYJjRBpVdCWXhFkNtlB+/LDqRm4TRiZtq6pgOaRLUNcc
SjAHRzncxSANRU+vBPSHyPkf01qaGNjio78yCD5kmIA7In5Gw3YrzTdxoDOguYJvMddh/JoMW79g
t6j4clAtAJRGK2ymRkq64OOkksL6H2kvh8j+1YW1APWGOlfQ0GGaCEbEQbeZ/dcZkeURXt3eMMiN
G85Pq75LTJqcfP9KBn9k2I3AwPWpeKY3Y/1epygT8oPzCOMeC0X/eiS9SwENznXciC77ulnxKYy+
tUb1AG2y3sJnBS9gM1cmkywzql/KWOLjUNfWWG+HFy/lfG/zBQUJ6vcfjbNLOk+pm025T/3FCPBA
fhZHEdHOg7Wv+mCMfjA3Dgw0mXXTo8pt+4y+j+BQWlhdXGAncbJOoyrr9LIEmsf0bk++pnDXHH0b
5L6zU88Y5fI11p817RmSF6X5lbYUH+dCDfasz/bcFbgrsiJzdljT7QQNHZL1MEwGmyNQ30Saly/Y
kQIwngfXgYQe0K5Gn5dzg3pwVo4TWV/US/PNB2hDZfKSJTpJ8Ua8wlXVDs4W6JfBN9P/VRFimXMa
BwO3gP9m8fwK6wCuU+J/Z74coDju6cabuMJRAqcsAB2w0azES6qDn7ZqMr8Dc2ujyQj2hQdNo6oX
//Z8bryE1Cby1jZNVvvvUXnj2+x7vbfD9Z+vhERgTyMAY2BmxfZlYaoeo/qTFEXkacGBs0+qbFxm
7S9J2COgv8butDNzbhNSONxNOoiE0zPc+srsrp/3Z+yTVV/n5imS1pbPHMpsG9CA2EPQK/Zs6MF2
SiP2bkHd/MFPweAx/A5ePFR67pxjBQ9EfvyFHIpyXb6Y2m0I2H0JuaJwS/Vu9ixVuFpkpoLm3G4q
h3iro02QEC932ArCCE+jMClvY+ogrMF8BhrcM/cuZTHq8Uy15Py4fBlBFNLxJFiXjJLx/aSezlhL
IE4pzrRwGw69IE3eFVL27VgEjpZ3xnK2O6RHu2AJm7k1/POVAMxuW/fz0llp/D1/IvjoX33yebKx
k4tRfdetlVtU8meYQ5kDEJjhT8gPOTXjPbO8tytoUZQ38aDMp6y0+suuF0TLtrkDafSaPrnYd9N3
UJJL9VDeImZSMcnxQQmUkTYHg//6hpWXck0n2ceOqUTJJZkgRSrUWT9ryovJIBmBgkwDOgk+20Pl
PJH3zCpPPhgac1qlKcArxX063YqQA070IIie4d46ClFmdPnJJkn6j8tRPiXJuGyru10G7DzHn0Nx
ROCCW6UQqkr6A/8+FYqrCDvSaWq0pNlSCr8m3fU/Ftz349kuZqZKjAAknMPhVjV02+OtwJ+FdWpv
r7Rv9FchKUmY+dWZZWuTs+NMfwaP+48jSGPbHGY2JjMaOcmj0t7ShN4WwDL49U2d34jgB66UtBy1
bQHhhDIAlQ7O5j207Ih3c/PsGW77yb9bupic2cf07EgFA5fUiCHPtD/qvnU9QIqKYZtCLrt+aoe0
3vT/9PdITeSnxBcrfO8rVONzC+7IcL800B3X9YKv5Lft0l41y+kmSUWC75tDQI3PgltuvULXAKb3
6TMFX7QU17UZdH+whj6oWTNQ9QvwO9mnrYu9ZETpziYbzHJ1dDM0qP6mPqyO9o5dmqEq4zZglKcd
Ht8dXOuwSdqa+XVVRVoUL+UfgEQqRZ3cYTmIBV4R+whir5ofQqTxlB5RnuwvhpT1sA6Ul9Olyc5I
7j8DFefCBEOc5EVZ1RB9zYNjPLXHDuszDo6EMi+q/a5y3YYAj5z+73cPMtVRVOVIZeD5fcMs5gHO
XISkBIEP1Z8ZpnQUcUKKTDRDgwqgb5yTLEGvZiVKa8cV+zgaeriUBuAfVR7TV/kPkDO1jVCeOYDH
1qhkZUJdmlqWfQRDPRQjK4rxT8wwpW7mjcgbw7MiMIL7hE9SEp1KlTthSjiE2UDhyayogUgnWYyA
ZSe6tHuJFtmm4jDktFWMJd2IVAqK5aRHoLpH1x3cuAPG1PtLOimEOB+IxQHZ1FfqKqxczlc+jfco
QgPvXOEyF2SAu7iLzce0DhvTpZdS945dEzjoTOHDmUGVsbjVpOTEHIMStHgVzfT6+3MYp83Wplf/
k+t2kJfEdVbZH3Q4u7B2Osm28E4JTe13Wv3SwIKTMkhCOdE/8pw3TZrR2uCpPa36d5+bulp1k4Qe
TjZfs2jWaPE3DR4gcbD6VDEEC5jngYJ+7BG0DNlG/zYORQEWiFoMgZIe4HGZ9Z+HyZntgE73eyoP
wMoQ8Su3oevggDPpphMOWYG8MxRBZqEGc3FGCEZFOODqK8AyAJXhGGcT7GjoaABaoHuCo8icnpIG
tpDyoGyUgA/Ao4pRiQ7e7egzWIWmOeYQUAq8+9vEu4hs4gwXLnXGzOAjEk1oe3LeO3Y79R19EPi4
i6AiixKWHDo9dtoutNJAmm525HXgEpu67/7vGrGc9aE/1u+wtjgXHmqX6I0Ti65C/HR8aPOPuk0N
bECatsOfh3+uLwRctO7acl10MNc4YY4LLSdYWgm1q9XlkDPW4az72Y2MRG6BFEQTiemeE1A5Cc44
Sgif7l3/uFjd6geCI6Oww5aNf6QxGmfGiQ9OIbGlvWtq6Giq5bL2/NGhyxCjYUX/aRWu8nr6x1kj
5H5jgkahlo0R8WhPReGSQQRLZvObmScIZ0AFOvrTWQF0wDbj5GD66IOT2o7Xo0usk7pvLocMlUAE
tcTWppZYPlQPTGZTiy+0/w1Bf2IFfaz0d14xcOVT/41cYVwcLk7s4J2IO8oTcVxKlaxyG9u7AFLT
G2sbLloz8foqj2G6kWtBfOw85S1lF1ZjXJ7ZghRmoAy7epsvEmab5dHbMUiYvIOgn6ZAfDB2lW/7
ASy5MlOpstrJ3b8kErtxaScxxScDu52KPDQHotxi/VDjEsW/yXnIWQCAR6WLsPCppGRLPxfuzyL9
w9osMaVAkQFlOMJnIi9qcM3cvdU+EC8xGiIM/OCgabmRGsc9T8gfkIHyZc1pHrDIcFcoshrfn+av
QPneiqimr2cScwP8IzmqEmm8wfPyLB9nPbIFdL8BEA3I7/LYjpf79Rfm/Px3uuPTPmbfYhyf3h7U
+DJoOPiock9jQVgM94OdphCoVGMfsZ/1673Dpff5XhBeHRoar7Lx4Ncydx0JkouY4w0JKqYIxtXr
Ux2gDUMvWw9bwnLWPAtepEz2Z0jxaCcyxRI9npP2KmJgVfv8S37I1eGRqaFigVIrdXY4utK+o+N4
9XuTIQr/K/RycCL1VQzDK0jI5jI2rrHq9LF27k+nrpng9JIgfq4BAjw5ULH4825SX7HTwb3q9n1c
IVIYNRo4w2x3h1zLyjNkv/zoxk/2p+BmWTJ7uLPsIH0zFDCSHQTFT8N8yZPQ0KhSfQb9zQ7nLOTy
1Yj1S8rjBSow0YylR6r3vnxoTTXEIREsOkB2nmaDfNzAfSwHFRtPOMa6kZz7UGS06hAcE0vf3uBo
u9akxyiKnrTcZ3saXgqBiyBXirg1OWHwGivHGLYNRGVgkfiNe/t/U9DsZ3qP8ouDTQBJfq29DySE
xxEjcRQ8xHdeiZr6jteVv8kF25sRHeCoYD/RwB3telAAaoPtDvc1wez1pUWY+PiilL/TiDTh9CTN
lTK47LIL1j8lerFuMRZqOQwhZLpe93BVqlNyvbRi5Cqcgy4F8jnaPXsMKw+k/tJtFqMfQsQMTvKu
xcOMLDtvu89HC3FqbQw1uS6bnmZPhDhVQrUw5Rs+ecVRoBXgyTVxsJxqpA/VdFzPi60Gc2rMJJqB
0gHfo6IUHB4JeJPZp14gN2JjvddYRA3VKdbdjJWbpt3hHdY5f/efmTNz3MqJdPxJwEb1YAb2Zykh
mb6eVNHjYXiDGLO79ibH9pCDC6lFES6ps5Qoqs1gjK/bmjayEqqf62Sqg0SfLKqlpzGmOpmY0kFD
Kaw0j4WlBhUso6gbdq9xRfRfAnlR3ZHSzRA9TAJOiS00vyTfJgjayhtG68dtTQcf8wDUkohlbOJR
cBgEvDsxsXFFSjHcokw3L3o/GPnfG4pTLo9FuF4NvwQgMhR2CejA4OoEXve2itfJWUdDLdqrJta4
CaNj+x00owuwwIaRZIH5smkCllTRAEIqqWjd5JilXY6yGPjh8Rr7VpG6c/CCvbatevdF1rKbSxnf
ZHHzNfZ8nWl2Z+ynW2LgJ/DORCaIs1oiSW5Jhmrr+sYMFgTHSAyqtyLXu1zh9EFQP92327WFYAi2
3cJXcjE8PGXph9zI3b3kTqCI2I1odpbZHJpz3ZKWynIMGGS5gRRFtRCy2GpbIuexEc01xuNuo1Iw
/bqS2nwJh/HNKalvReBQDueqRvb1t9pZmAUj3EInNPERcjslKmLj/K+R1JabYKkTiaK71QBepFHX
J6nNpFyybKd+VpnOn/vy/3NRKk03VQQqcE3JJ3d5KgDnJ2CL146bjRGkWfMvLeUg8zrNxwy6edos
ciyb9wJLv/VAKFr5PPrAOa1ZzXADuCPHeh6/t+hE2aeKMrsaQUrUT5UsT701658uf5y30H4q2H8f
+GWwPrFJH0oNqHCKr7UipfbVDNskiA7M6kMKRlO4a0cVKaaRNQrHDP/fIIPrrsAy/9ohebPSkd8E
QfTyajXo7EfBMI0sRIQp3VTSRf5xptHLxRB7761w2PSmk0GZhuQ5h3xElLEr1/3ogfa++7Hf8wqu
xgXk3sLHT1sflsXRtS72TiAyTMpy9eM4oWTRHXg91iIjnfDSB+irHszxr6IvJwPUxjgy0zxslSst
e0FS4imb/EoAp7Y3mFf7MtjvDEojUMMa5fcRc/JNiS7lVFCobQIY5eCmlo32DeO90GzM6hSHC9TE
youszDarmjByXCHCtL50amlv9YhBfgflVagn6JvryPBqwceCrg7dzg4YQehsbopy/4HT+ryTThZC
pdTrlqLsa1QmuIaxK7U5JaFytL7zABrOy+E7wTTmeRwTJimgg7WyE7nnaXqmXBiNsEz/j25QaaWm
MCnqPVRtcSAaHaoWC1TZY33kqMHj7blbGrcAHmADj7pUBbGS9rK6HInbIgNOmgmuaGgA7sqI8NEQ
rQBp8OlgpGbYq+Xd46aQe3796m7XViIsON9SL04tHLgXq2k/hYVJRfaxsHmRtxXEXCmJ7fxNEkS3
D5msVO1DZuVadLMKYoBXAql1LgWYyyp960fkLdhb1wrBup6tPBxEZrh7dgCcKOxmjTzQFhP//Vh4
YCFLCGKbJeFd2AdRJEFgjPD5qsg4fuFq8fUn9KLMDVoQpNjgANf/AA5zXo4El018M0iBjSKGUu8t
ZTjkTHVD72P2dyuATP4VtK4Qt0ERS3Fi0jh5WMchzX2nlHlNDtGAKvjCxvo5H7z+VRQfxG79jPAS
+J33r+n+yeKLJ0te27s/j8ey7qGegHEVEyOZS47QRLrGkFyXaUHXUWM02yReZ/OX6GxGNzXlS18D
jk2V64gMW+eJ1XSMcPQT9Q9COingMReRcfzsG3PPKtwpSwwS3pzjROyxr9ZOZC/fXOUIXM5s0+sI
50IRZ/ovYM1+s1GW0NFqnn0FCaGHMNwAageTdg3dnXR3MUlP2OrhatycI1V4SMl2GV9obNfh8cJq
hvFDrSUtpUpAmyVtDd9+DPHYfuvahwG52Nz6WvibnBqPY3X7IzoehzFbjQT4Uk9Y0YBAlQ0U2fBy
Lg9ub1HHytk0hAV7E/oWC0c8w0f0QOiR/7CFAHbdozRrLX8nubVp6ogQHk1As92Klp2iWMD2cfz8
sVpt7Y922BGWg9U9Y7DeafT/bTQbEnZx5r35ya17rxttTQPi0YCfiHrrmPBEs6O9gMJwgCWcgDIe
3Q4ZYZtzu9lSLk70flc0qH3CrJ4g8yW+v5MhYVvz7Lin7D9FwY86CnRYi2/RxuPfNU2+OczhXPNG
/svPrXgXtyWBME6MyYk0fGrYeUyo9eFncqSduet7j07ptblJpKckyKCbeftEPz9GzkoXNVoWNK5F
/3IunMb9IzjIaJQKmeGv5Yr2NC37PWK9eH6ui7cag9K40TsBbtxwY64w62kLgmoxG0xlxB6HEPI1
uQEBQ2Om0bhvofN8tCaBV5Cn4S0b9doPqbtgavb6+YYGMHtf6v9A81NVFaiNa1z31JnOJizaSmtG
Uh+i6pZsY0rzZh2FCepMaTIsxUYbKPmjIM37y+Hv+zc3a+K3q8KXS3p90foMin8owFGdwmJ+NVRb
dwxFhfJFLfxBaQr7mg3KnrGTYyd4GMAaUsoc38aTEgNi3bYj3DL8IZZI3tRiHujjZRtT+9hlHU4g
MGT4IM2eGHFpkqve1mEQVOmHJdjfv6yiA8dRfd4T/2AFHVVOwKdNzd+21km/0Ni248qlJ2AnM2SJ
xq7iaxzcR0at562J6ce05o8STUmA7X5O2WmgfglnrtfA0lF52T9FX8Rf4gWx8lQdkcAXOoxhfJUu
CtWj50Rv5Izj/rv6VGSMBQREWMZ43TfDlC5HvDMa6oGVIBsmZ53IYayUFvQ1UBvM+sZQqJRI3du7
J22Ow0FjX2HYYRRRSpDvN9wMKnw4BFiQbKWCzmXwVM1fwg/CBO0lLFcWYGXtGx1ZTj6NUGxoHw4y
L7sVq5KeHcawkINDHQ5ZJqvhe1ehJiVvqvkoCx33Yk4dZxaQ6dJ3gHf3hs7HYgP2F+3ysCOhXuHJ
qomTH1SgOTjq40ce7qkvgDff3PPD8lX0cg4xumvHMJ6c3jcKVwLbxuhEW6XtJA7Taaki5I/WP4Oz
Ms3LNC2yo54xufaLub57hvLFmvJnsgMNrwHJ7TC9c5m9TUnnw05Ouj8WO1K1wKEE778kcwnLJHIg
z5ZFcpDWb6+jYJ6Q4JTgW878m8TeFWJieqqU1gN+uXwmCYSY3ow5Mz5w/0ML1VCaSGZo2sETAEKI
Reql/g+w1rvFT7jUy+yJeSycFrLaCcEJGdTBmF79rCfE8+n+d2Cs98ALA9lZJPLOISiKtqRXEhCT
/gs4jh8Xi4LMdxdbIx4Cf5a8TePI4JOaDhr4HpPYoDAadZMXvmDY/Cj80K8BWP4T/bA6EVSJrujB
LGh0ZOZI6lKqMEF88MFvynrnvm5UTTeLCyKUMDDp1pJp43U1igZE8/GQMqjZ0jbZ5VI9zFB6vkv4
9RDljhtevC/llUSLH2BmfVMj0RrLxF4mrnl4HL/f4jAUkYdtO7Zpgto+sdN1/agMBZafwXVETWu5
GHegediwhflNO2mBKfcpSH+H1JUv3h6423JyKDLH16C2XmJ/PlyBFdsH/hbqr1xWROzrG/B/P0bU
8MBVP4WG8A5/q1snel+24B1w2CPHYfOUUGFgmtBgKx385H+rDtzNhh2/5dR5wNp5x6JAieBvym0X
DYYZbfCokQ3h3lauaFhUkZj9rM5vkgfrVtRMRu7SI9qkAbUF38ysB8dUhFQrIk/ZiU+OO/wRgPLT
OxBxO69EUcrGbZDqamSbAlkRffQPsCYoNf4S3xcHHCw4GbjZYfhVNB60+SVvViLIqg4SXRmWCF1O
HDNig4/X09qyBrsuu/5vli7/DL0jduWqFNu6MgQgMLB0GnkDKRqiMxRFj9hIY0VgBn3uD7Kf69nI
hCy7Dl6HREhG6p8MysEpYmfxFpCDrgDcXnc2PSGivtztSIjEZFASBxsMWoXU7IwTgILfopdZgJk5
k32EcudvrR8pAQvOli2MGwwngWBnMAL2c3+wiTAPe5x3ENjpKhwyHqEiXxt6Eq4NIgsc9V2tSSST
b5hWHEYYjMATZ94ChU/hCj1XdJdN5cCf5LFnovk9J+AQUPONAPfSAa1HDNSQ8fzKaXwCaQbrr+fN
2ed/4g2mMBfp0KtAK1Vm+maC1EH9wnYcHAMp35CmOhEsKt8OdIupesXvA6hT8sekPYEQXEedPum6
T95nbXoOfzHV5/U26sMOdJC6G7x/r3BR/iVx0TPH6NP+JLiyI8VY+A2PfKufTaVEDXSNjQjdwSk6
NMYGz4wxerYzNR5GP8ylYHmA5TPbKpHuBkhLB8yJdg95gSyd1KkWgKUh3Q0HpTYbL7x6H26j658T
xi0XEFfXbMksds/dBckB4k8hmooNxq/swcVLExc1cw23FGmua/nxCCZ/BYcxE06dqG8Mautif04A
kz1oOvskKNBqXmC9kYlkeSYymOPc+Kk9SnMSemNy4qMUIeKv0YruKQqGb1MY+AfrVBG24eBjgXql
bqUofp96Ec966LnScdhvFgE1YUx97lQ6/7ZFJDyE75fjkYqmxP0gIwA6YSKZ4cWEJ4Vy42PU0Gpr
sbKqGyQaOQrYff3GUMGsIGvtJlYg2BiIXMz3+S1pjN0+zUY4ZT//MJyyCUpOh6bqKH/nzl80QEjw
pFeRm//mgaAx5Y+PUbn0Gn6RQIAiRb09eZC9YMEiaKVMRrIOU558yuZnYPQBRIMtKzmFvhE4LzAq
HrxS60PFzhsneMbJFisbpWGPCuo80lcNGfOfipv6XdbIeTIQbyI8dxEvN1XAKMweW4BVZS6APWF4
7Q78glZvSH/uM3uO7xmIs7xX90fcgw4EVFPInESOnIpms1Vqu2V98dCxriGW8W5CXqdXBrK1MU6a
xuPjSNqOeT4RFhJdM65Y7sfrirG6XPLRxRIO6bjHZNY2HNMT0LJJfN+F3bKLH/EGXm+EvQ0iXhge
jB8VmHdwTjH6jtZ6WBmXAa7HPeAShWuT4DmMytIdSUbPtYHLzspMh5QSbz62HbcH0yd0rcZJcwjA
3UCO+RkreTMEGcw8ujbY7E/Jg4reUq8HE6XTCVvHcUcc6APlQvbnYnKnVIaDWR+87gUTDjac/DuL
ZrOB4Mgu/RDf+Cg+vcrCHKWiJsit4eZ2Qn2Z+HC8ThPRlngcKxFFE/Ei3elvCjH5qWGgWYsCOVLy
PwVrdfRe+ihbp0MOgr8JqUlF4N7qH3GsZiMv5lxfaDR236fFhVqiZPZqXxHrUc/SMnaE/IXjb0KN
NwAgb2ZNM5EXykay89Q7KQmYodsVWy2i+p5tx8yyWn6DNPk1QOki84KZ4b9NRY5Uh8nDFBPzdnDQ
AUpVJJXBY/Cz1iJakR9kkuy6CDAKSD0JTx+kvJIWd0BI1OPh+HKqr0mXYNrAgUr7TXlWiXU2fRLY
JEoh7RcvgPubvHSIucZCOZos/1cFEfCU6508dk62L+BSSUSzOemkLgD0FF8QSnSBDRhMGrPL8a/W
9GmuKBoG9ic4ZcAvR3OJU984BXAV5MLJh4cQ+0d6VDUJn1IGBB+sBYlFgHdgfzr4XLW8oT5tWjZ4
X/Cm3vLqKF0GHfNx2Ibh/svEiqcFHwWwgm65IgoWol3WaeaZPKTTeZdhL49C5Yu17rfQ7yFsX+Ve
4n+Ya8p4JkeD3vse+hZ7nOGX+CWt1kLxwX4oB7YQwJKpr8GyeS59zenB6gsJ9iCAghnyJGchOez8
Ap+ogUbr+6VCz3kLr06z/51qEP0F9Wstnc8NcOVdMuY4/iY2S/XFs+wIwkUNkLzHMPlhqBnTs7vV
lHvM2n4wjSOD0TleIxlpUWcYsodnnS05fya9L0ElMpZmGfix/sE3MqCNQKLyMcRwJ7D8a2bta8zM
VcU1eBYqY02ELj+k6CfudW0PMF5tzriekDlkiogDiNtzPELbgIBkWUOT5qL8Vt2KjpXne3VQWSAc
3NNtokF7uChv7VaTkorvnvfNesHRMLcQHl3tSNFeHoPFpefSmOcMoyz4+pQ88D2Ec11Wn908IY4U
+byGjH+RyqhuiiJsylvgmT0+/nc9V9JEmdwY6fRaaNu1n6vBpQFI8UnbiFELf2ps9quWiJ/qjVrg
CSiBQLvcnEq0EsY5q+Lnoz+G9zGQJT/JCSN+yPVubDA6Y+ppzn8fcDcCd2rQZaQO5XPHP/OBTQxY
YkxL81uGcLFgZAH6uHPl+cY77HgPyJBuPYiMd/YX3alSBjixr/WoFOebZw/Sr3V/mNj8qzBugcKP
LiIJuLoZvUkSY3MnW1TRF18MngZAZNfzImmo5xaw5GN4r5tNLttgj5ZPKpIU3aIHPUSLn7UNHUnA
cTVkLwaNahnCBTKGVM8fiJBmxIvjOy1C6nSA2tIJEEGwcF6uB6UYX4QWqXRwiEXPBWUQJM8XATd5
Ir1vPZSIOrItm6BawwljhQdWz76es0RCOjcHTw8vQlRwPApAcH8SZGvHsFagzqZDsETCaPOSqreY
+SvenPZ2jImWGY4mU5x+ZtbBrx838ATf2+OoOTK1eHHzGMNe3Bs9vzGnLB0v/aTcmGIBniL57f1A
mmbCrSSgpZmW8kH4JRa439O0LVGDXYvn978TLXdjYRMRXz5RfmwHZ9hx+cpu9D+o8iQQWR/mzsGU
j+CwIAMe2bNGfktxkSTbb7qoDE+jZu5sgDcqMOQtzuP8Mw30ag1/GLYHJSb8VmIDWbV9JxA8D3BP
R7eZ+gX8pfhzVq0DofyF4H30app+a+p1cA4YUnODYqmPubqNwn6Ll76eqzJ4AKhMzqX3NoAVD1eN
ZuAVcSRZ8mnRmisA3S80iVLwhlGvY0GT4tqolF2Qd4hisitkpoW+baoFE6BzHWgsY5g8N6SyczN2
STBmn7C0DmaqwVtdvCKKuNJk5CSMArLxihyE3Sswc01wRK2BTgfp2T2uZKuM0tuXwNUWiYkrBO7Q
iF1e+KnusETWJFqnt7gagLhEiuv0RLt9dUfafq8VFC7ccpdMjphqNwpu1QmVhfmFQUFPwqzi+Emu
SAdOaK9yIUD7CJYcAdDihRFXu+SAzwtkca8XDlRpQbrpg4ZfFf3kqhwZJla5D8hVQZF8IYsP2wVx
UqA+8KPBIo0Dtz2T/43y0Je+MTjRJMt79ZIQaBoHF+4HnlgS6nLJ9RzE9RCN9CF5XWiU9OC2tX8l
H+YpbcGpkqbdZVF739qBB5lfWx7766ij+ZQhZHzRR9kZvms6KChRD9ZQDuE2XNmtx2XuS/yrvEIz
nwIyCJCc7E1X0mh21TsR9IKU/PQBIjF/1KxeHHsKTmtrlxcrGQS2UX/qJlyQYIqksazTZ0HwoLw6
JKI1T4wINYjpB3uuBE3mJKJY5XFfAdX+AliYnn8zfbGQ/qf2+4EsXaOa8B+T+tZ03T+Z74pup/GQ
/PVLjiJCSzWWmvVi+B4mLs+ouGQeg5EOmruZiRTPuG9I8egMAW1qffvVOVmDx01y2emOW/dE0yNB
eNn2q/AeZKHhg9XCLLrEVZ1MLWXeZT0sQmzMa+uP56UTUvojSYgVaCCR9PhAtoB+m+7pdzs/TmLN
3I83sQkmBSNZxH4EaW/PBcMZlpLa8HayCyvVFmEg3xO41/FjjB0q/p2tmyqwT2QYDiar1eMyQUsW
1fmzdIbpZcbmu4v3JyWRosijNM/eCvA2gOHKaZVWh2Z1dLKnWiVdxcb6UHMnjfBEIvgIDVhU3Tyw
p/aZhEV8KZx/ZmAzCBPCtzBJGvuHxsdqlBtZUz7JUinEFJQvP55bUECTZ1oq14QshyBi+EJAvN+B
N9DeJ1ZIS9gzHWBzffkIirh8tCkn0rE9EJToubnrmTcQYohigKTGQVFWLfpz4BzSAsQs2uGdXUbH
U3aeQzpP8QDL/QFAjoSMCHgQ05rgpLW/iYVH5mWbwHVjlJZ8QW+7PHfBIsDicBT7Dxfk9hIWsdHu
5ao/IN4OQc6wz85K6nUiCMLQMIv21szeFXcukrHfAofLrv6POZt2/6U2cz4uSw9Tz2ZcGdmEPasq
1k1ORhW/yszhkhRZ9JH9vNkcz5jKycCtQGYRWaHRD4uFxs5BsJ1k+gC629EpGZKJb4qBpCjsLCSH
+uF/acFLL51PTWZwFjA9qoIiZrCc+9Eqv0oD1+v7KqPlh3I82L7J4SIQC+ixgpNvCcwoizLZSpdm
EhsGKDLo28FbU1HgEzaaXCLVvWj0EY04rPm9BKKndjpDsygAce8TMexNehBs/1hpmQX6m4MqLlFp
eoVoIHOXD1LPl1pGPhOwUATKweNnf8NftKAyg+uqY3NzFbSCdbgA6zHzRJciqteSAG46OuSNWfhH
g63ov7iNIREhMiSWXK4YFnvrdUyrDYVO1pDbzAaEzhnXNi/90hC8vkyNKme8gm2fm9J4XNDJ79Cm
W7/K74EpfgwUpfBjVgET99qJBmEWYo1/Q/FFSPpJGKcTS9/xWfk3oehptzLUypFxMaeLfM43o8tw
fF4c2nck2iK2VVxW9EZ++o6EDWspm4Y4eTv8ZgfN5A5WBvWgiWrjEhtD7NE6gMHD5NZqylGfCI7M
PgaNVCtTg6gO5cEUkHqd1bcArfgctAZPcw1I0ZAW29slnvsQEUtg3wX0aa3ArW+WFFzRxCdYqoKw
M9Pl3PUteUhoVepW6WlMuRPql3K+dnjaPWz4ZEKr+QW7uvMLXPcUQhUv6gEOdlPwNFLWHRFDW5Hy
cplB+VV7MFx0j6N9UQlWyFygarWy4krhcMmN9y7snk6JPBOwDyczgmLgoqfQGLevPKaUxMYivxBR
5TJAE+OI2MDcwdczL/GqE5F72f0QR4I0hO7l5HPSwbiV/tcjTytTcY7dGfUPmM+R4ixOV/BcBFH2
PI7Vim7o3JJIQ4jb584UxJ8+HJeDyiilQ9d9AggDBy/Uv9PYjmpew7uWSgT02rJrst4J2Wa/qsqZ
UnSNITZYbVTVx6RS+loff8/x5zVANoEaUoXG69Eb9WWNDZ4T803oFASu0MpnjPJBINbvwRecATXV
hp4k9cCwcX8SAGYBLTTOg7lkV+pD1m8Vr5T0XNUFvmhe9jr/0IpcoNYBF48Po0IynHc428marMil
LNlitMWtzQGCpAMlt5lWMOT0PtFOSDO78F/R1uY23wPQorB6ylYl69wS0+rnDoYy7qZcGnSyPnf+
8n1cGR+0ovryrJGG9XNMMjqTABJHcv9e+glsaVmVZsPkaxfLJ5WriYrUKIzvcV+sbdIDOt2dEPmq
OXR1dFu4WnejmD/xWHmmXSxFKDymFQ1ZMR+fAFStzu2I7TE9T0YZE4xCuWHPE1cPDDu1vEeR1uCt
qQOfXnBJX25nkwPGKfauGTwMJEsesia44gLRkNtGgRf6KgV6IEKBsa24FxgRrNULU/uNvHF3iX+e
y6TamkxlvQ6ICTUNvmTzkugpUtJJK+d2OZdETRKHMmkWC6D1vy0+DMblsPvVWgsXZbBcTKoAKZ17
a8yb0A8RbMObB0yNn+cu4k7R9IphY/ZEO4qCquAjcGzF9bZFnDDIA+k12VEJX0c30EsN91djZgor
gvZeMrwQjJI25eI3KLU6w23D6n6iI68ov85tPdamPA5k0L12URpRC9Oa/q9UxXZujGdnmEvo8s7a
NrjUi6hC/BEky3qiLUUVYBsUy0b1S453q2pjVMFzJkUnqVA/pk+BOfeINGOLK+KR9q+Wt33CZzsx
4IKiGeIRQPAZBTiy5lwdjBMophKFDGsReMFJN8QxfCGaX9xJcPW6lCi4UsGAjnaJ8BX9c9a9eie4
NEPh7QaYwwVw6j9o7SgWPOB3LivqtHv+BErwSCd9/bGy97loeCfG6tIwsHErAHWmGQwirdTia2Jm
lvUq2NDC+qnULkmnxZczZIc1J9BXQb+yVyvv2EM5YrA5GxluL9z+LOCibt0fl7jNkYtkMseTW0nG
iDG1kXeP+zH/DapvoRiRPMZdPq2EkeR1YBC44rXjEYUkpj9nLqBV/iU2adMhaCXgaJL1xefLdG/+
QYJXPjIgSmCuJsHvnNhh3fbZmZWJcnGgtBbYCvQu36tt+kFXZDwChxqyBVGaLSx2xe/bBY/1P6m2
qfllAShYt0qYItfGtzwp8X9eTRyCN/9uMNrPiRf73MreOkzxzIqnB359nE5Ld+fND0CvQExcT9li
kjpmkDJmEEjkIQHHZlBVEwaZtvfsqAN4caDxgM/5Fz1dnCnxMUBT76E/bPkAfkZpDMxR6wXPpWaq
pw5hHNzICb5UpkZ/GcUuKhnqpJAw1yIb5IhbMX/aH5sShuqKK4b9pc3iS/h9Z4pn0h4ZLBo90Eyd
FgirAOPK/1dQGms6cjPCjOn0rNk9Gf0ZKbvEZaljUzQ1FsRPgUR0Sd2mY20t2EjWhYoTS+v77MeX
4m0kJIhF8gVeRfMO/NwrIZ+dlKdLSHaFFQAJQqfiaPlPkqzq2Ylb2ZlWlZufL0wGDGNt6Zpd3eWT
nI+8wdLT3mR2PxjoBwiOMsABd61/Ma3/v77LEiSL9h6OoBvwl/muzD4oaXbqEkXZSDz5rY0u0SxY
t6xKIZPI7TfGCV7pXOCHp1IXPtdUEHgJKfDTn9s/1DLzN41ovQlRcCXWzKOQXf2jzBdwxIBMiQTo
i14Pm/qbTUGf/W7oIQCthPu6Xuyks+wkhfqxUgguZO04AUe4XRb+Aif6+fOxrADOB7C0pX/JuDDi
D8yzABpz5ZhcgHWPnOCVaClmW0RaVxQdDfmtA6cE93heSF4p5zcLegvb28tMIoS4nAnuEGCzozI8
9AU/22LkmnRForjkRTd07LxmMlDFR6P/y3G3Z5sbZEF8FMjaVJG9EUn5gBzsW7+6ffV5w1GR5CWr
cv9wtkLV0+IIzd4kQ29CmUkfdhkkwpwjKog6vhYauUAhRgj9WXSErZn4mNRA/5B9ook7DR1uX0d3
jU4vFNSbzdQVl0cIVEwPeFOzMQX2WMqwPyttlXoDwouTWDVNdGCxt5Z0QhqJaSBbTphnXkI9J0H8
pcmil8bmg3QSdlucq4M+NfX2fKiPYvSwjTndhYTqJESl2Fs0fAn71B5TSF7gEIzy9Y+MyHOJax7u
ToDH2XbPuF4NykKC/LkzYePBGpiJ3dgIBxG+7RGQpB8CyKQbQriiX/m10eyEXnHsWzp/dixZ0G8h
y5l8n+CDHsnoIhclnVFXgu9pgRfp6XYQ6b2d7lqz0sFUA8elJAC+EeszH23H3hfZNicfBsoLN0vp
vFbBGvg4TPeZ8osvts+RGPo89/JEDnQWTQhWnihXhsIuupwY9Gyn2NwE/dgiqZwGN58Bc48JEXPw
A2J5xjYVJJOt9nscocct7YRh8ZaUHphLB+wmhV1x8K4cBrow9Tq7MGiDN5tsg2LlE3mIPQTpBw4G
lxc/o7UIwvmqdgdBhxgV7lkABd+BitEivnDN3mFovNJr8OYect2oCzGgBYcxw2X9DyrniYxPzper
O/RhV8A7369JQK/Y1/1qTDrKJg3QkJUBGC7jcO+JvW8GJYhVx4A/oZLnnmQ8UNyyzpE9b/RUkoS6
f+mvrDWh+WaWGUgdC0wddw4N4N8k5rIyxTx9se41QmaBuOUAUZumPgifw3tdnA/i/lZO2m7SUn1M
ZErayZzNjQbdCa37utysrRr4sCDZElOTpUi/hZ4vRK3aQiUYm1KK1a03+UJQ33877ptyeu4I8hLc
QvJsXKqp8lNDzd4Ftz1E237UjyX/02vdGF51gZxa4a56gdiuDOrm+jPIHl3U7GaVmy93E68u4Yhx
PoizxiKpKRs/fPKPMVnEL283fuoFuwNBm9/K2rApkTiPPgd0g2UzDf/SxkPuLCSuipJTRQ3uuPK2
2WBTTK6vPLOdoa6e4XoiUgemJg7GqV0HRSXZkw0LpdLGHpbxzrtKl2LGvrdd0rXD2ibyComWYF88
GQZgr1dtlzURxUMB5BOZgkzOkIugUdZmoHwrLXiXXvb7O+WaOq4iFjuNVKpkQlV3Obz9RnQI5QVa
ImyGueNRjZiyKiJ0frz9KdjoAsj4FB9wcjV6EEuUzRDEXLC4TEGqIedJixz/YqZjPJDslbeJyt8X
ZIqJJwLJQ78+0h9i9UGa2sBbvsOZXpSWCTMtWLe4L9zVXhq8gQlNOtMvLo/dnhHr02RylCKV/NNk
ySIIOxEE+VdKHvHsvVGfR422167d+r9EmiveiHqxINm2+Bmd1hBC09kAjE20fdelOyJUjpekkzr9
1OJJ7n+UNi1KyRSb8eMOGUpQYBpy2RtYCW+A/chT0+VQS4AulZiTodtCICqhNi2HYCyquioffzqQ
DJBdQoZSFJzON839QEnPBbkF43MlnHaZE1Ud2s7uxbYV5BMAD6haudcSAL8saA05gk2WlYwjWiLY
qWQZNjcjsJEs1ngcpOpzx1MrHqvAT6oblcZUcRJru8WA0Sjx0Aamt1GM2aa/26xFtrhP0/Nlcce7
3FtaI4pNXbUWQi6Pd4awQeUjb2ZO/W5Yly9Jg8P8VxSnM4IJVD5DlbSXJ9tErqMSCvLSAEiiu3gH
whGzact1k5lCxr6fje7sVP+fWgvSeq4JJugRKWlPDWsxd8Vpl0EP2xuA/5G2nyIMePDy2QMpxxxd
zeERAp5UPSrLlaQsqHb5sMR6YWnkWtTZz+ONdr9Vt7FI8/qYqbN7V1hDxP/pAcBu9L+Anq3Hnlgy
HUchg+aqTyFdSWUMuGIbGX681p7sNWjbaXafL+yiEhrUlm0KhSy24ZHE9XKjNMkUPkBfAksDVnR5
kJKcXPOJ7PPzrbOLsEOLqLcjd/hrKwTvtTPBc5cY1+4S6FwD3Zcl0UwazozfxaYakjZbSw+AiAHQ
p4z2aOaTPTvYK+FAfPy8sKiObgvbz9aSJ85DGbl7NQQpHs9gtnPA90epsHl+UOSQoYRLq/HRixkm
xdMKEr6t3BP6kQE3sGxvjiT/0ukerV/khpKfMjwWOzzG6B5uEMcrVM7fN+Mtyoy0dABdCFitSVUT
qG86AehLjMc/U638EcIT5dOWjiVcRGa1Exoj8perFQbl1k/wJRNiZYWmi/KAa/yAkkgGNxlvD2qB
WVR12VFJqJD8hjZzDr8cFMca75sARln3WwLYTvHlc7pcaM+q7rSUR7aDoolzAsNtWZTovGTePy+X
FUVYkzmdkMwdriA1DqYjO35JEbxbAfdUg+/6WWGRpgB6citZ4E/JMa1L+eJ2GZhDSxo/xdil4NHS
8m3o6LNaolvIB0qbqXiR+0jYNmqOjoQeR/0hW61VF7by1YYFaLZtuwTcMlfQ5GSiZHbAJvwazYWP
dhjd5mquG+PCxXlBTIHWkz863B7cgcmxxHAANqLAOAZmO9IyE0sUA5oEM6wYMyhgnUkProVR2LRh
A9u7U7+W/IEj7yutQl887LILew5a/uY3zd2kerUwaPjukPgvJd+wCggw8w2fXDYVcR7Vqvuq1bgO
UDBRpc+OLWXlwB8iBdl9OKFo8fehK0GEapOQxPv2iBSXK6hXl/yyfnx2YXSpCmXrb/3HCLvE4VOl
fFi2ggupsPujW+IV/CaR7hjEMx/vgccNyehLZN59t8u+vMozCtUb/4qpRXeZStn9xfBbF+Z8u7Y4
mKd2Ccdexh1QtwZma0m0uXTDKnuKHfh8iFfogCYgckHNaL2pzkOBQvehliLDELtnxsU4eDHendNx
CCVYaaCVsk5i9KtUxSjMJwNIkUvSTFFYPrWRU06/lp5RdcJMCTWJsaMMZaLuUt67kIn9YK5+e/Ow
pqF81wJzWb4hWFyk6mDe4ucy0wuyKp3Uh46gbhiPFkMRJ7QGHLLKoPmqmZXsNh+t6kKPE4kdRky7
V9Prk8MGwhYy6M48kyQ5IU2/5md5+cjR9IFO5HVszWjlfjqceq55/wEpHr95c9F4jSLPtutDyKuH
8YNQW2so+dl3aIcs48Af+H1igmuajSkMm1uWLgS/MzQY1NXvs8FYe/q4QNQcACpIUi4v3X7JbSqG
NR9Jd00+IGh2VdGDke6B45323FibAcebKDFvUBPyZzQdeRg389udpiSJmlNjwLMDLu3x7Pxnsc9f
ReOa3/9qATyu7DtLzyuBH663fwe/K8XSmRVwKSsp3or5cvcCJ6r2KWBvjoV5ICmCX+vrTk9QdR3n
H1pYRVcTrtCLVZlm5mdeKrxy6TXJeTl3DNokvuzy0Tg/ZPp9OOr8xidilaUxPFch0VpM+TOeAAs4
RtXLbullGSboeX0WuEmMWsv1xL0vD8/kSwNvgjP2FalJZe9pz6PbNErd/E0b9vTAHmS4rrsBYWmu
wsn0uzdnATfF1ewIJ7GjGVUCEyPX/Lw160JetguE6/n7hWWp1JSlHuLrz+nU0wsAq+0YcyG8CAN0
8AQLA3nHV9/lWnkJJckPs/M6343gpqPb8LuAxuzQ46UUD/P+EYoUCmwn5L7at1h2TDqKFDQBEUBn
F8Z1Xvxpe/ndvoeSB6yHTOq5VvuAnDTwCjKhk0bTPIG/pOTC3gD7NLi1PAGxBNsCoUGkZTDToRBU
9WzAQukIH5ELcX3IqPsg88JnC2WvG06QHbCFNZgJvCLz98fpP/nb7kgzZ+2Zkpiucf6jCeZtfM6H
saU5qI7WQ019B0uFpEwnjZCuqJ5+GbaqShZKozTbJCq2IFRQ0gdCN8HX8xUFx0EpvzqM5MbggPRa
BV4FN5MZjFiro73Air+LbxQ67SX9DVIYPk1eDF7dfUGUUAdd6uMr/CdlecovuroCdSRq3dCx9JZQ
nsRPFu4dXHTuSiMCghXypcnNrdVd9sUUx3T+qBEzPNMXRBbOYY6IcnlQcAT+kr2kQokTw/xIiCcE
jHTLHZdSLpE5wmrUzZdAdOaQge0RsR/KMuXEp69ZbXXpYPZMB9OPCcV29vj79CaqlECwpoVBXDrI
0GsWEbxBzBIudPFdBYreKuSx8K1NwLi0JQwGwlB/IE4JMeapigCu0/qFhyXFjxIeoOjmsIY1OzB+
ewjkH7QCkPEGTA7QimkFRwWagS+ChpmTAzWLsPNegh0csMFYrMxHUbZDkNNMr3qRsD3B6FSMd9am
zEVM+wDNFs7j6wh3uBegOrZFbEWiK2B4xRTcZpU0aVWbWzu0xTmYJMRvBR17HGWXirGL6LWtyP8n
/C+5JRrQZd9b52EDPEmXiMfmYj8dXahUMFwIXXsVOiKiuAqi5cP27gfmgg2PRN9qKEi3VDZPxEni
3hCsoJtZEyd/yFZM1FUyZ0cPUu4UsqP5JkBjJQ3wu5N/96nBzJcGGmRwc1a846Dh+FyDX4Bp1tTr
eUzUZNo+No38SV63oF1ISDBuR+OYrcvyh7F8eQVNEIIxZUdcTPp3mCeB4MMgLFuzGC71nCxZaqpw
19rt8VlGDnT6JVg4Dcc3ygE3Un0TvR7I2JqAJzfghH4kt9/l4HxHiEWnjDQ9TllZYyuKzFgbX/SR
2jdt0jJUASHOU4U/SHI8rEcN0eR3GPNTkIjlh5mufxTYPTPcatb1SBqBvhstCIzRJYWKClFv98yU
7MzZ0zTUi1epSOnoe25U+A4elmJ4tSgpUmOTmogaK8vy+dEtc5INnDjrMrxUkC4+nPROs2VlMtSi
5sLZHjqk4+xckRvj+o6SszuPK4Y9tGcdt2alqtm5fBe4nn8JsOR6v+9apZBSMKtwi6z221hWF8pP
WkSF4H46IVERxJvJTWV1Z8MBv44oktZk8+9ZpC9aHBaIQLtkDK46F3/Jsn2+Y+ohE9KOiUbEHKNX
GPq06Qw2zCCfHqe5Ki+Vdw9hf2JCDS254h1Hp0yzp/ngzQRolwHvxLIv6ybEIZ1FeL1O6z9YAmm6
IhdUbIzP2YWooIuYU66YQ6Mcfot0WVEkRsrnbpdv3CYnaw3uwa+BFHXNcnPNQo298kzSWcpTBX9M
sbRhJF5mICj75eWx4RHHurdCDA+QIA4oPK6v++0ReyrzK9AM3xNR2e/diQ3VH89yTnKxkWlv0Hhy
AkZaGboMEjxiW3hFnZFVewfQa16vEmW1bcMg1+qGCopw5Hht4ZwY/crMLHfBAHW+Yfcv1r/cKxJf
oh8PYQgfUUTNASMnyHQNWMHIKhhO4Km+pLZCUgWE52aUJ4SZhTAW9P0R+Ky3uD5DY1lBtzGSANDH
rw5Zx2ILoUU126qKSkv0I58dc1jVLBRTlV0YAEda1jDVRt3gcPwRZ3QVMQu9uMnUxL+sNH+MLV1T
9Pl2zqIz/Qt4J/wsYwrZlfOWDzsE2nS0z3ftBkVmAOR/BKGLWoyEhtYDETEozuylNYyy1JNiXPdo
3oWwj0vBpmy1UkvEmje2uYw1VQFRap94kFnpcBwXmpzUdm9CydxmSGBHUdbH77CsUkCAAuhmJ3aJ
XNzkRoaLgBH75mt/SgtbMKYkPaSw+cdP1n/eqiycholHMm0g6Hry5OL+a0+/MjkfLave7yPNxH2e
XK/Hz6DVQBNjLu1Dm+5nF4j99jhDP0FnpdLlWQYYT6hvIJwBi2CtuxGLdOtxrSEzkNmnRC/tTcnI
VluwAKNqeQmsu/t7aQttINOppl46452VlwYzDstNZ2WhzKU7uPYJD+ZGXG7aA9DOYn5bmlKgWAg4
shK2ELpSthoFVMsMB3jJq8EW6Gg5ZYqnd0P8CFwRbojxcIe7C15XDLDb2fGSgqRK05qLSkOFmhqC
4qXggguBXg8AUR8gqcMoZJpK1l60F4D+AcpNZFDrrTkfAmwEuZ2wdQ7ZG0gRcVLMIr0KiuBa5sC2
ZNOK1vK22KjYtWewm4JTKu3aYpFaxkTuineM6/sC1ZG5CpOvQeV3NLEOrdxH2Dh0T039dq90u45A
H3waOGRfX+hx/zObNj8TaNQ25dsA1Mb/6wOg4bpTJhx0jhMZWgHRNTZUIXhPqeM8pFSNfo7HMzWS
Afua9Vn5yI9WWE4GkhYgSoYYrus9IkGj1oU8gKi9jcihN1ZC1iDQgPFRF6n5Fy6x1gIO+KJ2TqUV
a/wY/J1OKjyIKNJkwweZGQX+W5aDHXlHWhuOD/djukIA4njgWHR8vjFItxcNvS+s10DVdQE9Lh6j
NV0v89t9sD4BkoXo0iuD26+nAbnp/FGD2u9Jei5PVEwN/PIv/ESnPyjw/4e1s3u59ZzNrnNvpbEm
RqQUlFXznGuVFClMIfTRCTpteZHjGEaPnOSklZIo06siijorpu5rcj9JbDLMqSij59693lifpned
VriVAmWqmlhqsz2nNeCS4OOVujLKRWx2VmC6fkKEdxoOm0nzT1XIsqEWYUI57LNRAO2e0E05h3wZ
0HuGPh258VMdmWtNiitZMis6B9zPmGlgi+CBpFWVQ/+2ssSsXoQVEEovN5jk/R47sJWcrU9TVMw/
v24WJ55zKdoS2+K2CAabKyb4mrOVE0K2y8LWGDICNvgGz7VTK7SRS1AvJuQ1FcrVKADTrCaJCVJf
2TMEz26/LRZ+foQQTiCmjXA6GiUDoyxAo3bAJM/pRNTOFv1m0XeewxRIcZlz57qsWPWjEQHnIach
eyl1OJxQVhzNgmog6MM7yECyW5wykYqpFo3MIy/94cJkTgSKGU5ynWZXRBh83NdK5iapKAvEafiU
8vt0sQG0onO/SBuZPzuSbMNxlt2V5qlVKMSVYFMOooZUaKYFbGg3z0bRIkGmvQYT1N8KWdAvDJU5
iUV0IIiUbJwh9ibgX/m69q65bpmmPG1JE5moFBaJPSzj210nNIjpOemtRCOZJyA/wAflCA5+LKom
AgcFnV4JIupTmgH3X4OkoyZAjNFVPjQPPrT4dkvv5QWXdVF07aSgomAPYQHjD0B1qGsKFMAC9cHN
oZ+wW5RarJepgNH420MZoyJbosZGCNqYo2N8uFq3vArLBOl/aywERNnqHwJw0ham2H5xUe0xSRxy
1iIsx54jCA+VxPH9nECq9a7WfMBAyAF/Td/pq2QzIE/d1yaRVmUL/0VlilIWxC+tAy39iBAGKAfP
WJHfrXjNmJxaJbQNTRlqyIDqC5km3m7gw79TKel/Dbu0SrK4KGaXrpAaAM1U+mZhqjnw7o271kZ3
Wyn3N9DbTEqr6rZrLFeFwi/iEDdRYacOr7lGQYSDNzmi9tLdC1X4vrl71GPYSfyvECzwPANhumsq
RI0oM4eJf+yQlbCDkpHnKJ4H4nFI8PQixlKFIUEjiBT0gAVQjLbMBKdeS63Sp/UgccNa8oc8QFx8
GQ1Mg4HrIWhpnQhH84s2b7crhlGYwEXBPGaKMS723rs9euZ7HKL1PNcrDH00EUC0xIm8BE0WzssL
4+I+VzlUfh45yiWQPrOZ0hG8RVgXLGQMIxlPN7l//DX4hGc2agTtnC0CMbcCj1PCshBj5DWmgmgx
KL5XwsG3kCkH2KM30D6I0qVF6ga3yC9EZxtAdRjPY+0J5dawOIw01FHeVbPo3ShizX4Az2VIvKWT
/TQ4txGJF6cAUNo7VDyv7YD8xhSiIZlS3D/gVkVsU0vgXLj7eS/h8uXFkkIeQC2P+PPvvjrxccle
1WNYF7cWsextVrYQvy/oqFMfCKyzOyG9kD0JzQDHN/D6hy8WAY+S8f+J6zf53rJ6ZTW1n9M1iNbr
kB4SpOOPYCr6KQkrXyJimBVQur9orptNyBD1Tp0q24nX2z/ywOPKvvNBime1gd2TvYajqAfwu58l
ccHMLl8yO6oJGjVsYkJyqVthyhuxvdQGZM9lckjNd+cRaLanNTykkxlLC5ENZDkvAh0lL8fMpzuM
MfQTYzja/TIKlMuPVAncavNTV/45C3p/0rC0eCuy90pn34dvuxDKdQLRwt+IcCSc/sjrKYlLdhFl
SWlXKeOk1LeiSr5/rKf73akMkRHfOKCX4yWbnRmHewfxOlxj9tKj8cMWDzP7DIShSxwLuBWEVNvc
kIQ8TvRavcl+K+mUHsdzSx0WvCHNcnGiZdG7l2MJ3PIIxmxKTp0HJ+NCBI4SuE53Bxh31//2EzuS
I++xrlutCevVML/aMLG0e4kyr8878nzLlJJw6Gd8PgY4l2m3zSzX8XVRFYuONzRNcMuwQJfF4elk
Db4SHYyuPXlX0Y+mFtLg6G9forYAQF4lKENVGZrOfZ2Nd9IfOtAkTuu7eXZ8P+y3gWDxnXD7yEuu
zDuVwVAa7h7AylIYm8p1dqz/JIbBZv92nlzmNoaSNFHoUG8PScKY0PMqellny5lDvEhTRx3FQ+vB
jcR0pibx1ONYotbQ0a9NumkOCd6KcFm4vN028bkBfNG4/SjHv7nQjSDlSAZ5wvg+Hz+MDx+0rrtx
dwOqFzVzyiL4Z7U6QszRPJF4w22HVu1l638/zplXnVEEASaeH2wK3YxccEX9M9Hl0uNmxBrxE9l5
qPUcuRnM7qbjwccxysG5B+8t+ZvtgzQpqxsnLQdli+fYWJY13ggAbUTtnCnSrYDVzTVbme32ILuu
zt0aqkl9uPBJy1wxxbTkn95xuoBUvx+YfJEgBYrpeksZlE83SJnLXcVuw5Cm/nOW66/ADso6ZE+p
bPXMr7sjBPZ19usMvCqphQU9OAcz0+yuHajmQbCyB5P/y1g0IvFV1a3aACvusZMaT9Hm4s8TX80O
3oCukifYzzMuAl+DBj8MSBpKX9Uk29kQuah470Zu0sT7Q0hId1m9CRSHDL6ARjUeDOZ2tu9r0t5O
AbjTh1mJxU1C4fGKd1z+SdTAEp/Np6r3mOP26A+9lf+fIEKIbiuXKsxXyhWYqml5jn8XpCEu2EjH
chn5N5mu4/7LuzJWTBqGqu2iFiJQYiFG+OB/WlW+/HmErPEtcfIZCxoREQ1ddYXHseTOukVV0o6q
yAzGSu9qdyFOhBB3ZMEBXOIn5u+ELrjFGkfJ/lgqTbv6twS8FGdi4ODoFO1Hz9SyUtOtTVYjdpKZ
gJXzZ+Pi9NiLTE3TwlZeoqBaHCaoIrtxOEAWfAHdHiXQ7GMf2Mc6CIv3T7HpkzHtfZljULjSPbD2
2UQh2/KnKJASp2QgrUZg9+S0hV/FX1PrQTKsiPkmfp+6FhO1RJsCBNxUkp7BbHtU9Xq98581OUlI
UefvjNG+fal+dqNBR9tEhXXuokuFztP0CUzOgLgkP1vtjxyOVbtO7SRSUBl439lRAIqP8dpSe15J
yonh84YGwcQePtZDdfH9RP2iR5alOTs3Ta6k6FvG6WY3pq3TFcmccv6InElx23IB4JA4f61L5gBh
zYjxjOKLe5PC+sQg7TRhW27i1CaER6+OpeNBOkOOGn4FtWqn0JePXQ+jRI8HFzVJBJEOwROSKOsc
hJgDACiCndoDs6QO7ywPqQfYImqGtjvL9/8JRNmzfbiD31bbSBFJW+4WCQ8+L4hFp1ZoIqLpwXmG
U2rjC0PHkvgPk2YLTIrTCyUYlCPIMeD6o3UzSF47grsEm0rMxXxHtzMIifEBvo6haJIZmNvuFv/a
LlFG5QQhx36S1ltbcesaRFcrVCslo4APMZeUQZVVM2JoQuY//F1i6bN+2cA3TlsMDYKq6WgugwPa
1yJa7X85DiShsOUHQhhTdVJZyIKptUUclBSOfdER6TVlstAgv8jJY5qnv0wyPA2NazH+7I9jTmTq
zENX31SWdSeT/UifFqKAkPJFc/eywAlvUuRiLFYxKyvW4032UL+rY7gfWcYEW/kgllu6p0sLC34K
ZyZ7VlUIN5XaK3JMpswPh49gek2bEi9eZlULiOdz70n052jYsmXzKIVyDzywDs4ER8s+hkzZxGyk
k8qiPPP86yl2847V6OSpdbXQ9YF11dJDKkHLAEGF8acMDdBQFv1ZL99Unln0fc7M6bVDDDlTxVxH
7qb/J7ij1yzbhGzhJVFLc6VgIzheBi8gdXVgGYe8fZd1DT5ikkt3nPlgdMQ3lOPf3IPpuuAE3VHe
YKZLm2iMufNMpKflAsvuqWiMDoe2xHl5sDSHM1lN/qXwogaUMs68hfizw/mzn9XCNoYtx4N1Bqoa
Zh2yqTnDil1YXGl+oYS3KfDR51R2zxcOM9BQoVXHUdBGg/W553d7ZUKN6JwkBK2pHALkBLMZQ6za
e6xdwfJbXUmgYsg26PoU7ys6YXod0Y4BZ6kbdvP8HjbIdMb4628jrMHfk3N3HepPjkH7FCAa/yon
UICGNoQfsQTA9AIX5yCni0Uz/sZr/OiS+PCzVUWHKafJoMrZPYIMPeG2tCeT+cUOGlvshIOkJw+N
POOZvM3ql8qtH5PA4vRgRKwvYDMB5BbcFSDQH8G+Vr2gmVb17l+bz25/z4A5HGEfJLS/9jhT/Xct
ST97BfDDvPsGKTOFkTl5rHPnUiNYwrxeDfwPQQT6i4GRTGE7xAiXDxqSVe+zR4e2dzb4lWyTfkFn
mS2ooFg6TXZ+DREP1q3xBN6PD0l5vrO85UNoatwXZdmeU0cJ7OyjRizpRcKo+0Fwx7hhfYYwQUNY
6K6+WwC2JY45S8wsqAgWcddMynCC5Mr9UQn7hfqas9uL0IBdXMhPaJHpQMnThdcPCE6baz9RIoZP
8rnRF7NIZYinjnj24EqMCujV+cZaxlI2nYniyPbXCXv2wjsE+t7AgixOcrRGCwvPKGVECd4nmNde
AuUO9ST1tSHD3P/nV1O2KHIiEmfN1aDL8AW/VMwOlMJFj1RUott5ivZ7TTmcmd/JuSGzd0A6ySnE
cyLLE/EdXFnuPIwQCcCzOrtHFNbY17dQ8uFcF1xRZPgopIcHwLUvAXp+ojccxAaOsplrgVX1FuSR
9kuO5u3SLseqP7Ed1ePfJDDNP2qpBLp65bo+m84ev5x1kZkg3mqmIdsUBHaMx5zQXeFnn/1/aWZ7
7PNrkq6lqavVG0Ao5sc73o5d/pOr20A5O32SVFYXNT6GJ0gjffTFsc7egJNbTYmBmxE0B1ptCx7y
Rg+cMJEc8RYjrC3dQAjms2Vow3QqWtaKrV5gvYZCdZBRg2lwyGYyFJym2GDkkCMG4Bo6jFqkf8Qp
UoXfEbqjX3Vzc/IaKvAeEIJu0NGdmezo1j8lPIkTND5d2SLyCR5px2ECQpC3tlLCsb7inoF35JQv
3ANHJy4tE3EF+FfLay7DR8llYnYaIGMGfOJJtZwhtrG3qKrO3yNWvvdp6VBHl1aImXb5bxKa7D4R
xO7Bm1F2Xpae753Od7qZEEnhIJdOzcVSJl2AadlM43KsN5o8BtmwkA3RrEY2tFzHtTQPqbD6Go+n
fxhkuE4b955JVSQuN2qkyOmv1alFA3B9ZflDHs3pOySMk7NqgZXKvm3xiuqHQwbOj7XDbt0pYveH
GfPPwZZHCSjtredi8nfr0m8KTCyK1FrgtXfaZad8qkVelD73U2VyJJuiRv70+KB4aTt9JWT0AP4z
xwmbGOz3I3djtn1rZ/8DPqpViWo2H+Z30TBqVBTlNo/CgzCHjXWSPXYviPdyo89FDgbjB0UUldiQ
yKKIvC/rlkOGPW76QUfdV468BDM2OIeDNdM0IcDJ3h6AHkoY/rBKkvkzjrQC7WX6XMoBZ0dz3Fb9
ie/VLQwlJMbonk7tE3EYKz8vaWfyauyHvrr+wVItYypXPEwER8xFIS4/GH7b7O+/TSAci+r//Zlo
gCMgiBgQuYTFgUmqepHpMqJxaqcDMCYLhjnYhOrF+6h8cFAkAOH0nXN5EGSHAw7dOJx+KdZ/MD8P
uf9BDpCbTQFCuwzZwc+u43Tb3wx7ex9zpYsinYiT80vgOMSwwEV6Naen9MGShQs8kYYVsWMbize3
TUPpOEjWJKZ554K2+WWKq3VDYwjOeBrrQ3ps7baBzzzwv2hp820/Eay4a2rzfWGjvP9bRLmrhNnI
ALpS8DdEq0VQj0liGY3+QRgLKPWxKVbxg8FhDlJutoU5qi3EyukM80QgMr62DrmEJlgrqq7jq5rT
fXIz+EIpPtnrRuDhR7VZIFRzICzUcmiKgKNyRSpZ9GAFbrMnSLPfKW+hJhhZ2E+wV/295NuV39pN
enXHhkTjtH7VLcQTrP9l/6+C3FKTwwTCiTFUTH+mqA8/YuUvAwmzcjHeTyn6+ioUvQROsERHQ7pR
1Mn0r3XtSNVFJefOcGbVagxQaQNDjCNd+V9kfT+g4Jdu/frFzd1IbqSYTARg0YdsRz4ZqR9cGSmz
Md4bLD7lduFmqBgbQy4+Ppn3U7GMGTGZ3IGKFsUbfFBf3jVJlQELhxeyUFchXOHvdEKWLeUvc/2E
GoZf0IOhwCNwcGlU0x4AgfRLeQWHt+QoWshTfPA+qwKXbdwB8STT2o/vJ0vhXH6t1rY8xyURCSpC
SyMs2y0lUrLvZmW4YlkRfwFKP4iwZWpSn5el67V6PC2mmDOgzh8tW2vYRsEu3bGpwk2dPqRt2jhT
FjJOiiLPDB1Q12woHSEJkDa2grUV405oSER0EMt4P86OITRBFmdG1KWjo488c8qqMCGT2wJD46Wq
qWs/JgLOIXlQ518jmFAvc+CpS5q6dBBHIYO2ODjDOynIn8Lf4n5SV2f4hyTk4tEgDdulDlLQFHGY
nu/UMDlihSXCmfLd1om7aXFauURJG6PYz2OILpD5R/K6Mr8OPYBL1NViZpOj6K7oEDrGak/iEUCe
CvlwZ61AaE8tOsvEGzhAUEiWHeVim2HJLGXxzU0LjQc6JPSZM/CgkdxX1Dtqnw2GLGqDM1OSSQl5
DgFkRWUTWmC5N0xGtgZrEvl1MaNEBsD2pvIWi+06Ed7D8yyNzHIpr9iSHathAaoPYusQKkfT6Gmi
nfb6xmI5kKjbxVuVhjGjsffOYlwBWUJJKe82yTxeTVKLzmaqrXx3BL2wy/O0Xrjv7ZzClmC+XKCi
Ukiasr55uH8LS/DfWcylGD52WGpzICFomelV8gg/l+AvR7pRhouTL0asq0h5ZrJnkGpVvovp2UPH
TaVzt7SHU229TBUehk8aokdbXZVc4dBat4S01nYlDOQvY+5Jtm5R3wOQrA5g/ERLbl8Ig1sCJuQo
GcNMWRRcVKa23mMU6XZt2JmbZdCBqo6O2ETxqBPvYsU/UHTT4NWuz4/NHhp4kABiIkkgbQuQo8rd
VGw8UUk9GaNtqXgKfTSc23JE8WYxIILWuq3px5qtUqWnGqOHGPJPf/AeAupcGauPrr1AuV7yDzL8
dhcMxe7wLDRM+6vaLMwF92Fr1r+2wRcdxlDDxPsTy0IIrBcyESaPivJcamgdunjqPjvOOx8TMfzF
r+zHMD0Rc6Yt4rMIoQZ9NAoRx155YwO77HCF0btFQ/InD99/EsDTJpB5rpgi8i54FKRDcXq4LscG
LV6P/4fIPrlkzpkc2/yM3SBOfhxwaXXWNq5Wc6+XRdE8mLnvrurRWhEYFbqQRk2rKsn1Sg5OlZly
2zwlCpj49a+QTpOIKdR1Hjt6tcRr1f9OY0sfyW7FH1OBLmgBH7OccFuUtzzn/usLwLoZjZYAuxh4
golKdLwdm2yykOlvle6SpcA6rUfjwjsLlq8IvjkCdOOZIq3V0ORfw3YXYbq2In1J5CtE0cAndSyN
WsyXOS/oORRGD5BRJzTagWlZpDwtnLwYskbD7Qt6rioiXGBBCBFW8WiX+HpYBRFlzjFRGboozaed
Kf7M0LH064gvxA6CQeKiLuSPEeiVvP3ITGp6+eOEpDNpQ+Aespit264GaJP+PZuEAoHQuOM/febH
j5bJCNXfQqXZcyZRH+qdi6G/1xqunlmetcz8wlEqxFMJPeGCP3c92ZoBnJno631wLlUfH5V/e2pd
5l6ThFQ+zWmLipbmKJYrl1aDIh5dA6o5+/4lEGJCnZeXdg8tN1ei9Pf4ln7t+AgkGP2X6i3WUw8k
kmBrKBcNgPanBu9lxHNIngT73xBK74hN+LnYMzAiW0WS0ZZXP68SC0otB+Zhl3KCGtQXbfA6UlH8
vxkHWqc9BCYw2s3yKexFzhmWJrmM3A1G9wOzxNp+sPlbYrmXpY6JTyHDYshuD3nf7ztIodRW6WKO
pLt3UnMVYrYwl8zDlKWhG5zzOd7hvXE4PB0/ClyYJVBfYeNG4SAiRATz8jpIyqLU4e01DTqQj6aV
hQKBas8D1wmYPy2KpeNkWFIwix16T+4yBLper4zbY25ZBaUy2VGEZHZ+zaf5WkKww5nt6dqm2SWs
9P8DSN6yYxA0N9oWHXdzJEtaPx1rPHbn72ElQAucQlI4V1Y/XWNadVWL6fYEnYQ0CIEGff6/3f6B
32pxmFS3tifEmz7Cf4fSdwVz9te+GVPO6wuJvTsaSU92M7v4QimcgGXhkoy8tMYy929rxxU/SMW2
3c6zhpj8XElvB9BXAHTSlKtsnx7RSwoFI0xSf3kaLoRqJBznhqUGF4NZ2OeZNGc/Lth876OKls0y
2vhuKv3ZT4H69gZI72D0YJuXJ+uKDndKLk6Nro2/qitDyQa7d/KXj1sedDTSqHDurUEh7bVAXsIb
nyCe7zQckerminl8PG1rU7tGGZURNcjqKyr+s1mBX+V0apMu/bF+F0tkQqTuCrIaew2ZuziyMxbU
HP/BgPtSbd7fpyzUivdaf1QFTjLbnfYN1CyjCti3KOiW47i7e61Qzob3jEa+rkghKjhZ1croD3DR
iGsltN9QyaU+klrbmffV0I4dLHPpC+nt4TNkp2N1cLlD8HJdG+N+mUgUF08+0VLtUCg8NiATcGxu
qx4FUEakYMHWStOCZJ9qTskxyXbKPgit7ULopLMH+5ZFTwYZByjf2Zq+8VwISApKOlfJ4NO6VMKe
b67Ks3brqtack2WpfTP5NwJbFuxJNXBTgTpPnWjl9IvnZWIT7yeKxBGysOH+LedWcVvD7zE7Cq62
KDzJ8+t6c6le7xu775IYjlbG8P2xk0vjtfV3p82krnPPDB5/8C0rAPoeBvm/7ftYrqY3SOL7tvf3
nDwh7Lnslk+YDMbD89o7njF2Mg9ouaMItnVm7sRG4p/Z4XQVRNN6AvWxqwGXvjDsyl8zwGAL/C82
t8HsK+48pwh5Q5U7e3aNYnlZqVYzlzXHAmsonBZD9HSb71iUhMF98fuL7/W64r9V1aRjnS8TffDZ
AvuijnJ2mMK05yNcNbXMYc9m680yJjheuL/DQ1d/y+RDqX9Bvhkhbn1NY2FAhWSbrzYBPcf4jDqA
3vwKwgytfB0MOrW935MDlIp42QKJiVVFYy6sSngxIu+9vRFGS/0k1PM9VrTXRzsiStDmypZXN6Zb
9SXN+vrRZ9OjBzCCRi8oXj464YmXJMg45Epmpb+NUFSj/WBVJezYURUcDUCi4WuSEZ5sDHtv3lOL
2qYWCbMTQeg9wJjA4Z8kG0of2/m5In7gDNYHGpHcL1RMNhjL7DAtu1BiUHyQ8fwGghzpYDgpnZdA
oSZGu/9qfDuzaO9H71gCE/0YbAgLHMoATJh+PtKloWXx3NEMprkBdUxqgOWifw4vNnwKzg6Dcd9V
vCZ3ZBVo2UFp4JBPXpIFN7csMTm/suzkRDclpwF0EoG0SKh5WtVLLc1yCqW5KmUlztX20zBJM/6S
RC7s0Gv95as4Ohpz1tdAvxh7yD50emYapMm/8pDJmvg4sxIY8q3ukYWsNo1g413QBlC5ee7sk1fH
MWXfWKisXwXE9jcm3pb7W9300BjvqYGjyuLNbir71FpIWVZOtiaP2qDE5ZI6l6wlww94yjccd+NJ
Omzqvw5jxmMQcNqwL/mV4xDDE1h+eCfWpjgLNT8hw0i1JndwCbpIF0sITb14yVjI3+KyA3Ur9zJc
O/9xx8kHu4KY5IR3HaaAk4uiuEki3r7jVnWg/D40XCyXOBV1sYlni3kwOo35kRWpvNpOYvmmmD+k
hnfDj5M56kZSfeLS5KV9ErqZPLY/UrS27VteQbCWUXgN+xiPqDS6sEatQZASc22A1ApBGMWCgfLr
vdKyni4Fj1BE1NY9kFHGLs6fTmMenP93RdSjhb6ejyOOZRNMxyVJ2nicf/CLybF2ng31lERB9Osr
jmVGo6iHf56p9zYnq+CezNRamGl3gSnGthVRbQj9Yy/SXyOTAWXw+iQ7ZMwGhLxOjnbrSJGB9X35
XC36BuSFDqkLL5WCfIZSGxP3j3Tg6Vw9GRH7sMd0w8QzINgXniE7jzeuVTRm+1tEL7551m8fCAZV
TnE4cCbE8Q76CeJHJbh/TtbAXHtZrVmeOL3fS3DEX7xWsGJabxtAktpNBOGRrpcMth9ER1H3Bnsu
1nxKCUOBRPQKVcEczvBMDGBfNQGs3Zwylwi9EL8B5lWCMUK0bzb430mYoROcdVUR1LKR57bgSvPb
xuwqwHwypSE56AckIpqdUsQWfK22yIniYVjwxrjMTZksSk4iMhctRyD9pwPbav+0KtkqDEGVZ3uF
QcGe0KGoOBvKt2CGaI3hVHtfWBVu5rEpGXk+EbaRMIJhUj5JjAZqu8fcixjZT+xI8HaRd27gdNLM
uR+hp5rL5BQo883ERQdc6SdBMmE2zbA/8IroSbfO2tRKkHp4FqfbPNlZK19G4GxnXVWXjq2qui0w
0G4NU+T7+9Z6ov9cygS2gukv612J0iYW+5MvsrV+o4LI1bkB6MnfcszCl7t9Uzhah9ac8eOoBBbI
Vpx9v8LB3lkoHhE5tygDs+81MQk/LmKttrmuW/ooFjvZq7MUGW5CSUeD6xYQYZqS/XAbj6XcYhTe
QBJ8CV0c/73Frh21CpG64k/6DfToTVgsi3cJ0/dhopzKUUKWzsNs7aok5K+7bt6KvtMfUckiPnPt
/QqUXmgSpg7YhRvs5vm4esM+J5ag4KDG4p2LpBRMneJMqr25ZCpmnxmpnaxmXdwY99IFpymjHmQU
YCkvNlmyTGufCDXO+5y42E+xnEi7/oQFhLEcIAa9FGMTQQ+l256y4lxr8c54U3eLRsdWehjTKK+O
MevliW8GUbYXkIWMet7wcMrij7ryZ5BGw/WPEf2hAKMOMl6t7LnAng5UKIJApm2PBC5JmM8jGGaO
33GF6j7VzROLEbkFPEJX49XL7zMu+yfCltLfbd3+/e7c1Sv/4MOZefXcC7J9GK/dVfiUaF8kzAE/
axrFk9FBUoe3ao3ebLJAKZ4QJcLxhEEKJ34Zt6THqwJSkwxMAkZY+pa7wtwsY5ZkNL3iPdLvU1PD
ewvGjH6DtyQN1Po7vqMWrBrGh6Et0gI0F4Bn5EqIJtDD/r3foTzLKb5kkwynKzgE0uiHKv5N7nNx
s+Pr+lZ+ZAakk48m7W8uQiqKLTslR5rseoTjgBQmkPH1ZF9JH5YCmqkzJknAcxhBYy9LXJkiZfHZ
g9NFrEbbknOh8S+bsxfbkwdIBpiwAISbtCIeyREp3rT6vuA99MFfRqZz8WeSLKpHwGDoB+fBVPCi
fKNgYVoeSUkSeVsTPYhG+ANav/Vn0oKsKXthCiGRxQEHaFCcANadcdd3hwd799gGATPbPMrbbnnC
TKYqNSJklBNS7O/uzeHQpsuvRBzOVQ11j0KCWXYn6aFaUQzzuHbveXtuJZU8MeuAkSN/+EEfIRmw
+PRFc+T/GmD2SmApGolDX7FP8d8khx03PaN3vDHqNLKbTdAhr0wZSoIhD3h54pPpHtV1QksdZHgU
pWRZIrxuK4h8lzZuNvGy4yF3ZdlDkF0ymp2+kZKp7rZb5gaK+Uq60rlZaMSgfX+8IQeLI2H+noeP
sZbrN7lEGRanhdRZ8eu1xmXGKS2BFOtWCbExy0S89Oq3RU54MjEVzLGOZar8x6Petj9nIjSSBb73
skLU/IiaEQIMG+8LHZJqvAUyTMTtPX5wu/QPOIaPdG+l0POV81lZJ2P70bP96QO2UpQt5GTCVmAg
KrXqVAYwp2zdlUNcX2ecY1ZEpudTsM3mFwNtm6Hp6DeRNt/JE82Lvd/oQ4j3Z6AuNw8Ft5Iz5zHH
H2T3f+nXOO0qKBQfOAGB5k3H3QJAhDt5Au7MPrB4BVYBcvneddsRAG0WIbKECCEm+r4D1sK+M2qT
HKykmcxF70MetO+peecjNTd0QLep6TxsEPXdOagTRt7L0L2Bu7y/U3KUQHeJtNftXMUU2JKPxgPN
jY8TsOv4+p8YpmNSTqaoxH/ECLmwyOXJQkf7DStntfbZ8M9zjE+QCw2SPbQbkZpLGD3OhwgQRG4F
4Jr7X70g+a+86MQZgDEgsxekbxsouM1k3XjAw+++fzl14h+9x85Mp4DJzJpSHQfaia28skv4qsiJ
sR7Iu6HWerabTUh29lB+emtKVDGoSW4PbwhussV//PhvZAQi9fT2Oob7oMhGCFdsCYpl1CQfZOPw
zutNrA8BLe8TYrlKpYD7Vzr4jB+9Gsr0yuIBRPzqIY73rFn8ocpNVLf6kihkz6jPjTb6PlSEVR+8
LFF1leLEw20Ht0cLx667HCVoT1Qjc0Y7wIxBrmkxin5jWNZy2Hh/NXhPB96/ZkE2Hj6ByByOUf/A
crFre3DOQs2GcxNGjqSRzNToMKT08u+C5rPsI+3OBCpxC237vTWRy8yA+vDBZcOl6a2BXbzPmZ85
wX9mIyMNsCJJnN8ho8KP0Rg/0fFYz5P5dkRMFalXYus3YLZjeW8C/a+ZBDgQ1nJKAUYV2NRW1Hbi
koXq/uRSnC8LrnclvNQaBRkLbg+dt9eti6MT0ncsRUV/PCZS2xbj+gQxXWoXw8b6w04kbsEGBH2+
LRRHBwmt6bsbuAUStFGBTtulli2DpNf+jV2qfSdnbIYj4DkmcgZIX/S2nALzp9lDk9L6yBOq124M
NH93U4JXJLu7Pon5Xsk6YLdyHEz0xoBUGme65UE9GD7DIptKUSMKvP6MmeLOdeWh4zWKSCqlpjwM
E/gT3LfhzO6bMHcsqWmLaIWHgsCcY88BhY20uhyOoVX5HEi0F8u4g5bSnqejZwDFBGwc5lLCBbz4
ZYgM7hCBm/6W1OALdwY3E02MJXztE+mIOd9SevYdv7irlzVC5bnQJF1HIL8SMnehz5YVKaVciLN2
0XPP2w84y6ZGbetoFvLtii2xDttjsrHc0+fd/6Ae4TpWiFfn66rRThBmXBhwOPbv0qYEIrDMubpa
oNI6GiXF9Awnjzi4uEjN+ykX6TCSBLRNfNz5qzOxO3lVnFL/aKISSLnCk+Sv7pbgDfusveg1S+lR
6RxgrJYV+PJ5PXcNaHP1xZecE++VSOb2+wsOHr3lAR3Fw8x4Z58hCGtqR32JtI15Nwx7uSErQ4xU
zrXvcF8zawJY/lH2625qa+9FlI5Q2o7L8IylnI0x8OpqQ86I39ZEogoS9qBYF+ZGl6Rpq9waAfb1
dJuk9ob5kjkKZOgaxazwWaTXcXGPs3mD1JGKbDPs+YSISvZEk4+6/eMG2Yztd75MVwkjrYkyYNbU
IIYLRqJdmybupzP+c/MXdBC9etLMUEYl1wZVcn5uJtD7ntqTEhmO9vTkPodgoM5tTQIYgTf+BNpG
pNEJ9t4ZPJ5NVyw9Eci7O1Shof5kEH+NdVtTWDIBzOcpAgZDf8i86/czLEmpDfSqXVtGOgktMPYM
L9X6/HN2/XNfdBZdhRS1Qzwjx3HaPIlusg4gGuBgZpVA00t2ru4+CyhpfXTHRvEb+ITXOR2nnxPT
MM8kX8lWF1GlvP9V9x9NPr26YOYYILC7bccfMqXpPDhjL4eTbrCJSgAiBBHEi6mvKvd0/wswYio0
l54yOLliLCbXdHDdh224orwW/JkG8d0Fr9YnNtdo4Xqjogl248adYeyB7tckhRkxq3FJF+IshjCg
c1eMMxHCaQiGJauNyG5dmWDxundaSOnucFkwJBS9KdAxdDrC8AxMTKvEy6xv6HAobtyrpYheyOzS
rgn9OlpkKQY75bJ5F5vqQGgGLVyVduiDHHqef5Q1UJMTJAQZMplGViPs/cMR8qRjLP5HXhIt3csA
FRBFx7GMRJ588i3PzRqdGzoHFrutSyocqsIZyl/WqcFmYxTns76Jyl9qzHuRhDJcS/Gvtgjly8il
udg9IaWc9vVQ5Sq8Zk5sSRed6zDkGdQJCoGAwMluJTTfI11WfVXk8Q7QL26iScGsnOc4uuiwUP/v
4v1fpeNaHTsg2lFnI0pccvFWD7FH2AKI5lOuvSLcv7oUiBl3z9QqTWcQ1r47cgzLw0PhfdtVlC2p
Iw0s9vW44vdFiRJsjM/vz+VuYjutmOk6MaUTc0TJqC2n8tWOEKBGiQSexLjz6W7FDMOnXBJ5SU7V
g0yeSx7wonSvcV/dhPt9jEYRYfcTdk72ZoBoDOBdxszaUKhGOljXmK3rfLwaMa1PG/kWFm1kgi/g
ekCfTg+RnxQBRHoHr+hHs4Qrk0ntZ6volCJ2NxqHuCr+VKEsQX0/xdZN89Lk1Jpwobw1+RI5qhCt
fDHhC+q9gqTZMEIo8KQPrjkSlv+u3T0I6zl3AM7bCZskI3fhOC32LZ0JSvHUMIKQGLQtgapU97fO
KH0QI4c+Al8olA9e1aAFpKbM8+ip1ewG7nL7FZTznfGomxhhh6H48UGItrm6BrqnfjsmFofwKBS7
lU9iH5d7LVu87GtT55Ne9jJui3M3rxSEw5iNi+/FKT/FTqGG5pNv1z+3HrQ1qNx7E3lDnEJ5iWin
GoxCS/eIfLfAzKAAFb1sLeU2n5keNeTm+VjtgHsVcKSHbcDo6UpNgHy9AJRHO8xZe1rX7ya43xR0
LnqYs5oGEGkkAQA++Be/aazkY2sAZNQDDlAu1mgUrTa+++heEr4nd1bkYXJO3zEcAafyaHrtLImQ
rKLfT4qlVbxMKyfsqF8u59RpweZ/mYSKZbLHflv9R7pTaGqN3Q8B5j3xd9A1FCMd7i+c0PkwtAZU
3refdLh3IEQXpxs5d+c7PIB7CeKMBI6BRtUNYB2EPGumj1fxetIxSKYeJx0EkClxBm5XYKdoIqWQ
wNDOiUEfj8BI1LqEC6R7Lxfg3m5nE9vYNtY8kFwVfwK4d89yKTfwEGuxxi6m/vUsEoVM2BCIemdq
5viv20Qvk/zKayxSks2Cn2a4hDFfb2255RQ7DeqmgGrt6fujWnvuZOt9ZC/f71rin8jmazqwtDa5
VrHvp48+IEH8lqHQLaDQvLfeoR76NGEK3D8hkWmREZu7+f0x9Zv3UrQ7gdlkxF6YFiBa1cgvZcF5
ctRPIm1j916ZbPtKwuw7uhZ+NrUFk3PLQJzpS9IrSfKyWUVzeNXIjRkZAXTybhahICwiWL3Laybe
kkmYLxJWTpI9SOOvM/s9ROodWXrCPoycBW4FZUOCHKN7feK0nr3fDhtRPkQ0kTQvOloSBTUWlpmu
KbYUB2HQoFQ+M/+uaEZzHrl79mPeEmqskpctnyuSXEM5YQ6i6PmHOjogH/ojDOEV3qH/v6F5PBPA
P7KY6INqNa5YXDbEfDjA7QcxXJIz7hb78xGWp8x15FilRUxOPBo9coPv4TDWSVHNQ0JRpMVIQgsx
CCqD/UimtgcZxiiut+Tjn04+xGIeHr7rDFoW35/fMDJeux4rQG4nbdqVk9OzNUjzNbh4iiPlTepd
5VlUYkVQw1/Oa6x+vRWzXYrVFvDSWF9DP09SBddQ4N3Av4WSrrnfSTg9pTsrKvfclX7j9/iPfP8o
Qj12gdZxRwOkJo+zxvSHW2TSEnftsRJjJ/wrUKyMskLKukKBdJIGRH5IP4HIRKoOuYUtQxdr2bpm
BN1VZgXifovGSc7AUQ7T/glj5q/4/qhM+3Ht6nab3BAUiNuix7QJOJAYnH9fy8hoCN5tygm/npfe
Z9DdansXyAZC+1DxDvGVmpYYxAzYR5V/UR9SOFHyPEMsTv2gyFvLXHWsEborGJBRTQf+GLbZL4Jo
qfBD5PzMOK30vFD2yPfMhxiaXXmn2UKcmCnk9dSxQndt+pf0DOJPjVA4aRIBrW5U7go4KrRn2rmm
kmxMJU0+dHfXCyW22KKjgA4CzvJSz3xN/D490ulBBAIvOGKh22CO08WMH3CrVyUnUb/j4wyz8frH
VW7BKfV0i7yyiHsakqxfefL5rvYCSGUcp5vHsspMQ2HSOicf6R8nVre5TMQ9d8Xt2jpDVB1oiEa+
q9OTaFpj0Zu/3G1zEb6ktzwmJAAxfL72/ASefSX865KKUlKOMlBIaKV4/Ylpj23P5rC/mJ/V5+ni
ezZMMZVh0WogC4BNpCbiSu1d4S3cChySkOLtoay/cQ1MUdhhj73JTaah9ARKNHZlXamGOLtzuYqG
JxrGX3nytR4GfdChvND73ERQxX3MfDwN1bDRHos17tlnO+/hd/V41PAYQeVX39YjrvO/xTR6O0IS
Uzauw1OKGNP3P8rz2oo0WgwXtEi8v2Tlg4G2aNW2GNgcTVk2GtRRA29HBWyTirGaNnLCBatjcem7
ygy9gI2qVTCeODgNwmz7xFCfp9H5X0eQXU94a5IHzb8HAeGkPblTVPD30T0KbfaUEOV2Pe3o9CHi
8ep2xQhTPem4HzTg+gewXQ9RpnAT+Le8pXyjeLVtTpC1P79Zr0asFL9Yr4W8hWbees8Ek3FDmEWa
vs580kwn2OQEM15NIH9R1EPvPHXnB+EFnGcUu9ltP0GbwmGs5mGqlrD9iTLOHNDGLoj96c3LTUVP
n3RQjIdzvxaNWLasCDUgVJNXZSYqSrIhNyvcz9W+juy7BYn7HjG5y7zxUZDAGColjjAL9qQTVvog
Vi+TD4XTNsNXr9WqXlFIV23ig63JdvJplRtJ4kWPxS0jPehauq/eqSNqtYxg8RLUFpcZFxaMaOE+
nz0Gm2hWmdFFkoOQMc/ZZaYWIyOLLy1HABvuuR6+C67EyfSPJDwkcaTTZRlF48ITOnZkq2GtOzm9
qNS5cabVSoS0L9kVXmNBrkjXBkWc9+8AHDY3AiOllhRZ+B7IIqF2H86nxhIaqSWl7hHvvOVKBqBX
gkLhp/K8zC8xz/8rDneZ9mpSB6eiGcflssfBtTYBhZQ3HeC/+N4Cn+lDr+cwVV9GMhN3HCb9I1Si
wEWeoy/DwU9saILx7LQmKeAJTeYdMVnJLLb4Aingp/mkwLWMV3Ng4jNBPLyNdkVXj8DniH1jmiXh
N6gbSi0UQeVYufpTgRwZR1kvTMr2yCz1On6vwubhQg7rYXiazufeXyeZJ9VWOHaGMIOR0ETpCnio
jG4Gy3Pr26703zgFGzwRMTRtUrC8RatL22VptPiXVb79P+JEe5mZahPaaX6KJYVOeaC7vnQCHHJZ
AQFWA34RBvoV5k0eR6DqelK/GM+YC3HRHUMXpjhQG3dFAy7ooMDpOZDrgHzP61FrGf3PPvCXs/iC
yGgaTMcYZ/BaktspoO7hzlvHQq4RHrbYcyViB9ZXhP2MqVbc2RITi1GYnkEHb2NQZnHH6m3zhXK2
ySgR9+5bSMxoFUNBcBQI439LE/6bGZ4vd0E5dMCdzFjtXrz/xaDI7qcjiuY+ZAE1ezTsk7HkHAov
Wn8Srx7cxcfM+9pDb0SuNTrQeP++IKO9oLE6Y/int0OyPWPYs84SjpAueZeO/ND2w/xXbTikovcg
vj2C1MGFBarNCh7C5BvbSPBwi0t/d9dZ62R2Kgefsjb/5dnYSDvCtmbChf2jFE3zcU2CdVCoWsoD
3R5tW25HnE8dv/0mq99/ps4rnE63WoLjPlX89pAJ4VnDpO+lPq9aVaLLn3uIr1OncSnQpQS8okHu
8S2wk5EsbmJU7Lit4DUAlWCT4iZ5pYC0yVNDp2rUWuwv6ZXD6/1dsD/0yk2h9v0M8VmTNRpKsLXm
7NCkKWzs3h+I9TpgJwkO1WuOAdHtanHqy2zQpnlNhdcqGhpHRN1w2San5eL3wKPVFsIv9EvW+mNp
JcMc+e39uJq7s//h9AGdSBrTStI5ZiyJk5GdzWvb7xAhiQFqpxigyR9c27pHJpGLAZkYW3k6Ghxv
K0xa/xrKZoatPfalVOW8lkdFfUbSEM3DBsahXonbpDS7SOalnSUZVohbVeUiHQhApVliyKhqCshO
hhIbzjLyHaAf8CJecynMapiK9SqIDHn3BsCk0Nbx7OlIjj545nqTMJcjVozgG12J40VRf9PYumsQ
bV+W6nKUmDWKcLlmIx+CM0KxZMN8dw37TlU3jZCSL7SFaPOyYhQBaP4F3FXveJj+hw7E8Xx229zu
bgpG1E2pJY+z4D7cj4AJngegBLaSZPwWRgwx9Ib3BfEAb8ZTQ8ebC+MrZBQXesmXdiWd5mBH/C8/
Td9NMtCzuDdNx4N8WwydOKNJuQuy+xFH+UE6SKJsLLpuBZB6qSO7ayShz/gd9OnxEVWSpYmkozeZ
GUWDoN+21vCAPGFBZ8FNjC5oP48HGcUA5M64SRL10Zoxgvuxi0pD3YMqIpRPXzSzqAwAxryMRW4H
Yp7bo/U2qAs4Z5K7EQOP4nCXZcKEW85Bz/PwVRSlb6TbrHuO9uN6E5Uwjyt/1jiRhM3QXakyE+hR
xZ7y9+sAfqhXjKvUgdubjh4dMa3OE7x86DGZwuAF4xSqIWMIyZl517VX39KBxwcgFcMhvx0ehvZq
kO1B4Ii1fHTOjSWW2zgLAXULPZPp0+TjqgfcmzY0xTJa6MLquUOZik0LW5SYO+rnroOKV0mTyUQ0
lgSmOabiJziqtwztAnpBikHEouO15/jYowdHyCThtR1sY20oHRmCA42OBht6NgRrGQR576KQpuBN
wz5IA0iX39+ljFTcxnbhnA0X/trqRx00IqAwwvFmOWquaQXxWBZLw/KzuTSD5bkiK2AKp0ri/IP3
14OdowPuM5KKB2Mwk75cNswAcCpzohIQbeEMUv+77JOEL5bYxl45aeHuzmgZTX381rcfWQEnU7fz
IRsq7YGT7X7Refa4F/AlPvk3krxEhR1ZJXM6ZMCpttnuBWPqZtV4M/1GsmZ3F5mXBqkrScxKZGrA
CC01QOlixCzC8SckLj/lgrVgIssrVB/7gNmYmXxoP04O5p8VdUVhTa6ZQ6Swrji9E/pDXxUN+plB
ZMmFCXE0og0hpwBSKYjuGXd8P56LRNKy+ghEn3jPCjndqGXxsys8mKWBvhVSp2B93vELwDWeiYDA
IxnjIo2SAOrC0w41GeKsxtC9wu9Ib9briEysZ2SB4INJ38VoDO4BL0R7ry+Hrf2warLadT5RJMdQ
Zag+h3aLKIdrm0MIKHu3mkr1XujhMWII4JT06VM/KWwIWSy4lJB5HJRfF83YhSB29eIIiI5Iu/QB
Gg9y7bgumQooJtkqNQeEI3I2HEfiNm8vs8EH4w3fbvWSXpn+EDBbzDZGZQ5P8qZr3iTO97RF2Ptf
juKbuljbIzijKy+F9wu9B4wV3k6KrqDrzkUNaNEgubAqBFuXRshxBsP5JrkSORg65qMFLkWMXcrc
VNHfDssU9nRr3sE77y4fP6tcKpFrI+LCNrLbekmPdnamL0LFEuopsghCK/Gs9z0Q+HiMNeyGU3GE
HyuDxD1qiwDMeymuBxKNfkh4dsyE78ylNKUfPSGirDZR/wOhgrLAzqJS53x6Demycqk8qcp1ze6L
nRNc62N63Cq/h0HOnn3/fC3rdQ8xtCacI9auEa3MukiJSmCCSm6PR/X2UlT6a6+PWF04Hya367fN
G/9FXtloyQzpFUqn6jDsbYL8AG55Eyh0cxmLVXiniAVPayJx4kLBEw6NSu2T7TtT3lA0jgcpPw0I
ZLXgVktKVerf5Pntfjjj+2Tg/cwzETGDURg4jmryfGr7w1acUF9JS59bQ5SE7QO/4dy03CJ+iKEs
JmPlp/2z6lnwyshceAVJbziyJ4K6b/Twve6fvh48eomWBxfyaAGWM1/HCkRXT73GTE8sqxmElQi2
6/N94tsV4hD1CrfacOO22jrhR40LhAf3UJIUkDafiTCly1G7/PESzR7y8Nlna4kOn7BQgZVs/Ohx
g5so1y0veBwUBNx5tUtl6qlK4Fw6gEVtQFjpEk3mZMnwG65VlV5K/gwYdXnnerdKJgt8YZbJ/LnI
cp+/H65bZ367w6m0IAdLnK7xsDnyJmahu4KWcaMQ60zjbZpvaH/hlm6Mvcd3vR/HqfbnHPyDt4td
PWcKp4W1rCMPJ/1FTzOCVyh5biZU49IALcXs/v0J6Eae1LQFsucx3g9KMUA4QQf0eUNtHksTKqml
1Qx4v/cmYBSGIsl4UWZiA5GYmEBbcFKyn2889neW9Ez6VsSxEvn2brPYTIJm8eLF2zagAjh0y4TP
Ks6s2sihMdEjqVhUmz7tx4iU2OAybThiZPaG7eXTGgY+esBFPirdiuhGXyEarAYZjSsU0iA/EKAw
UifrlXdV+SwRhm088fmKiWIgjOcTwMrNKTPR/TT09SguYSaCdKUbzvkneQVPg6K0pjP6yaC61nVt
Fh7VIqn0IthSfTy66e4IfxLCbqTwrXask+IU7MKcmUnuPfPX8U/r6B6joCet4z4HjNmbn1ze/Xwq
0dXaagZb6DvdAAX/yJS4w02NzD2d15xrYwNjJHHffAPuA6FbN1dYJm88+9q9HH8KbH1p/wUC+2M4
qfYjFp4GvOUWnwIBpDruvCixDOXXgt/gucQw+eC9BzrnKDhQA2NFl2/CDoHhM5TtKN5qTzowA/uq
Mu79gizctOkcIUbUltMdhPLCFaX2mOtB0t/0di+VZYuPkG7B9ucy512/ldY0v8LnqqAqFi5PF65t
7mOe2I1xsgaTwSCd+j4v7WfgTFRrbz/9iE3birMxtCkJfdamqkJw7I1f4KHC6nDXlBahDK0aQmvE
jyD7ZHxN9ic3kdUM8DygfNFeIG+NWeR55h6dOR5SCak/Gli05nyxkgNUV1dcuf0g/VhrYn3H4EYq
bRwQitrV1RfMVmWAosjGCWPaYLQGW6tjx95+fuLtTwXZ9xgGanCkPeqIvnRdNpG6M6W+wmLEP8/2
f/FfwmdW+ecU3JXqZqga3UP5nIIK4zKLuKubMDaJaIDfR2z4ryuO6+D6ChUkGOpb+NnBadVqTegB
ZYuBHU7LFzwaQ/Pk2Ii934NzUde5+nDhWiac5Vlt12a6x1EY/n0sMD4A6je2QxDIFqPq4DvPD7CR
tCP/O1RP4sDbutVm+na4GEGDnZPZKv3z7Lbu9wZSMazwYp3jSyEvAYih44TrcUemeGfp47NOeq7+
wzhDr9xls5VEuOIuYVcU4YGtcXWeFO0mMWlPLaJsaJNSjxJVgDoLHCDEF2yfuQwSrQe7loyub/Gt
MVh1+AJyvEqRFNp4mqlLSg8tEvLX+iJHwBuvWThCGijmSaB/lYfcyMoaKNCp4xoBorkZaZBw1rZW
wnzgl37gN5X/TJRhd3p2m6+f0PM2JHjpFqhtozZd86W8jP62K/l6cdY9ELkUf0cp8f7NvAXm0Kqk
barJkQdoyB+lAYytuCbPqFcqajUm+ESthho5B33hLq2w/GO3cfePL4QhjVpa94nyErfEa6F3IPmz
nEpSec8WUaAKIH9+NJ7PWctekVsA/j9H76XsKYOrYReGx6FTkq4Yh5MmUg7vALUdTnxLCAWxe0ha
GO1xBBYPNjQHyT2u29oLNTUT1VUVAGw2EUnNGoECZ82m1zYhoafo6dhpnDHl7cZfdKWSGNPV6Lrc
jA3yC49wewun7ILo9QwnIb7jIP81ruyYYGT7XQKlF6a2E9OmeKDa7CV3uD25TXm5CCitz6CKGiLy
htzpWr4r4gQyYL4yNnJzQacF9xDqTqC6kYOvLVSv+m6sh1z2ZLGDKSB98FWvO4dyGSjiQViu56JV
jFcN1aA9VYpoqwmk2I8bOzI2JsB5oG4q6tZD4N7Sl/Zkc2kICF0btbEyTwz6va0TGrGy+aHEgD87
N44hZzO3mHyzkEg6kc608wjAikVCGlrBvC1/wRd0LFEOKJMUcd4+zhtTjOUwFjDhih3vTRWPs2z9
Bv4v4irOM/0Kv78rx4tsORHzf1StPql884lu0Kpbo4qTJTxTDX85+edVoOV5WzYoQkXfXIrIClst
hN02/sMLEJmt9nqYscY7A9P3f88qdhLZSBE/oas2NcbN8h5tdlS8qhN1d48cAK2XAQlGTMZJjVRy
nhgn7BE69ezJM0VEWyrYPv9brel/84aWoOMKgYTK+ALPKaSFJMA9QSHPN9mg39wZMBzMqXiRHdw6
Na5miDN5Ss/axfi5NUZdrxyUBz6xdKxu5ymTS0/zkQHlLKhHpP8nQkMWBuzaeyfRUbLCqHpR3zik
M7BXlFFio/l5YOt08NTYFFIcAu1Y4oQKscQVmlcvFdYGCbg2Fov2FMhU6rKZXSJ9/pDf7Or962jT
uG5zKoor8wmU1MjqBSse2i/ThGZUQxSSpzrt9APENy5/GL5kZhPtdbASXVSvrvFZbn+IIkfpZIXk
iD4OMbjIzeVoge+X8802Yjcl9ceUk7uOfSjP9nKihAyRdDxQmyAtVWy57b+hYLpTsWafSBbwBe1M
745Ixnc8IWUoaRKqQfrFuRF12NzEU9A1mB0ep0V8oUMHpD/DvvzXMGgLleakB1sXrO1oUOCM5l9i
oVptlmkBz0qeFKlQp8r3FSAzFGAvY38Dnm8aB0WUmUvTbR2WKxKplrxV+6cXUUiCGI/OGl6bChVx
pcViWzr7bPo5gMceIfQMriJpItLyc0jPTYsPdbN9WQDPhy3FPagJahNAm9gUu+whzcRI2nTNJovR
D7ATJN9ZADLqVfKi65jcTBOGGYzXr8WgY/aT4u9tZhiuOQckGs2P9ABDmjI4WIcbpMYMUwyg/8/q
MJNhgdKS3cv3KGTT8jBnf2npuPf7YthrBzoJ4DKPp4NBnKPOvopuGgTiGp0QRhDoGucOT/KdZkQK
1NU4I6E00L/X5QwAmbUKgR22R7xJrhm2T3EOSNXv2R/ETfEuVpH4fNSiwYJl0hvBGJmCQUoEgO8W
Dk8jI7eozt/Yo6uYyCnR04+D5LEacNkT/ijaD+z8TcvZo+/ROXsv/YpFEwB/nU5aEsy26vINZ/rS
FzLyP//fYSrheroK2nPQLfkoQUZyxXqRYtYaNSBDEdWn7z3UE4T5I8yo+lvQaxgIo0e/T3Wj+gIn
MfDaf70QxE4LodU5f+KIH9IRn3V3x6gjC7LtajHck1jJAuRLJUH+QpPsbBXgEVpsZLIUvoAID7Op
3g6+kQSwnVvM5apz7Q6gKJeM/rdGacKmpV+lZuBjdAQpbFg3bpMe2VmYF560CYq6vwJggpPM07LG
W4A1ZZNt2t37W21wwemBTs1pjuQjH4K1p/T2kpqYjwsQAz6Cx/Ip4YU81n11C/Pi6BPw1gijA6TB
ol427kEdlZlEWllGuInUGnUrLwNxF52i9TpUFQ3ZI28T6tNqs8+eOXyvLbugKcgTVjjyGWi4E7xd
+ArQsDmH25KIt6fRHXgNk3HcNDGSgnbHak09Y7ddy2YlLCcK4PS5blge1pfvWPgn++8xpLslfNpP
MgsxJJ/sFxAvb3OMhh8ft9E0DVjoY5ZNTj/hndYnCsqkN+xn43/62a7YgwupBkw5Td7e3hQIC/vQ
NkZb6MjqkAekZSa4raQ7voBJ0Buh00MYziwyluiWrFF20tmJZH4az4r8d0mC/ERoy9QPzK4XF0x0
Kjo++fTCM/8SWbeQTiy9f1HjsHFtx4B6zloh4EzlWyClaflHscteuPLH4kt2lOukSdyRyVQ/m1aL
ac+ynfIc5vW/XsGT+mT5LN0dnPwZZW+SQpzjKW3UwENyKZeoPT394QWT/4Mb96OHPvZfaLDrZCL0
Sk/BvaKvFRvxLM6wFVxNanLIO6hfNiQ8GCelUNUwq/ur719KKZTXSCypjnwyDpqySH2dwz146++w
cAK2rRHLsz9vEzJKqlHCmLF+rq4rK+CTxGcX3te9gr0xUEsDShayqjxutBkvAIaXAJz3hMoYxV73
1vall/rMrjTYk0qIb8FKyScDmtu+VZ6RgVFpAdj6HZ/3ijjBz08TA8rKJfGnNGY+zbaaLEyr+e3X
VqD8DR50ujQehBPSL+diSrcaVzKl4lxh+gvhQnmrCbqpYNya8xV6JVdzH0zC4lCwH0WL1/X5SXlJ
bGEtHBRRDB46qnUtm4JAoo78Opkd6I2J14s1MJY4t0QsLvxrF7uGWUbKVbg/yxKJbHOhQgc8pBEm
YjIHJTERkbrDAu3THD4mhfhP286CLkbsrG17XPSM+6YLFnmgO4xoYwK4k/1/coIdv1XOX6EOI8+F
5wpJ81LmiDF9l0rg6AhwImZ9GsBIy8g5eKPUoa58hz9XYr8PXrJLOmwbZE6355n2flJtvd6iIJwX
VmDNdfyhUS43f1jh9oEqquugFDa+yrjD++4r1wcnVmJdBBReoR7Q9iL5IGjtDNUsA1DnIBERSupG
COBckxzFcW62u7sNB3+yshNdae/HzVXRi6HX2iNpY5qQ0irCUlHgvFFHgEF6CDkJIJCcW+Nhg24G
bcjxggWPaNFoE9dxeC2JBa0nbQN3JjM6i+4GapFj64eyPjl+tKO7G0YAPD3D4JZQnvclzAy8oxfr
bC70w1HMP0uBLDZKe1qjfq9xjh5ncMHwBBiaC6qpAlwUVK0vPBRLD/1E1QlPjX8vHJmRXFa/+RuF
zxU7wJHkrXh1yrs7NZrwQ9TZ6G+r5fusQG0OZtOvynY2RjrpJ/McuT2LbqB6INXQIFCYDeUpXh3s
vP3XSSw1K8oYVtctpdFsY/gpVnueCzparN8lYsuqL2Bq29EdgXWkv2rnG8vVjgpteL1tudpQ/ZFP
mp1Epjww5MXI5PVO/nGfgGAfNzVMaN2dwuekQ7cIASlm1eBR9NakJLqJ/VEaZMqrgND5jVxd0YsC
uHmTcTvoTiKA7+N8rjdjVXvnc6kHztH6lzHCGiE6AthGPVrn6vTqdOCnpKKlsv8yx54GpJpPK9Ut
UgQjV9JzXv2gy8IXBdl9pdNjYvDzkzOJtlc7q0IV8Y4GfKXF7JsSdjJJVZGHiEK45O8FPjXOR4QH
GyQ6Pq6u8EXo1Vn3LUcdbWy5N7Vc944X1zFnEXPFJbnuuk8jq0q+YVnz4hTPL8YrBGRXa0ZGGoQo
FjCDoCRuAmp9nB48tUc8Fe+ibDM+sGVYg3pUToluL5COCONtcSQARvG7+BAEoCucQyySNaIN6msl
xlazHoNoBjwmzok+J9F4yfrAor4pNHUshx8dwuPZDkTZ74b7bV3ROm7sXPZ+2rbNl7hw9XXPEXFX
6Ppn1R7GTw6Us1fCJ84uBP8XJ/vSVS9agoknVkCcvsWLxKyJ2/Cw8ob9dvZxmTse9vfMAJgLe0Be
g/9FpzBdExes0OaWd1OMXwFSx+nXLyI0yd4hKbH4DLt+H4YRN640BSE4Y1AgmABymyxNd/PFexGu
yBFIQP/PNsVCUpkCYghdXZ4vv4frSLVFhcRddPIQdJiqzqu2HWBqQfUbsU+A9Tt4koBxVwo6ABui
47OOkltZUni7ebAvFoNWWf7QHGiq40j6YnyeC1aTVH/jKNJlPMMS03qFslCvFzNnOU6gmf5jMfDO
x3RH8TCGQMuc0PaXsiJAi7TIPZqmrz+Z+04TSC2l8hOXitnftitBLJpwCgsXarm5bWk8MF4BS4DC
qQLFelDQ4IiC3tv2OHPhyH5xK2SzZLWv0fgjVxlUibLbQhLcoG2pkitqDn7kOgQYveWGR0CAoqBp
9DRIEoM0xYrT7aV/592s6wFKseK4i+65XnF50yiiH4zd5+1L7f2s0S/kAGHO6K/WsuVDS1So0JQW
g3VjjO4ynDTdBYaH59INkOeGrFRoF0RVlOGr15CJ40FAChYpIwItEPczN719wG62+8rB0WmAULRe
MCmmU+NXWl4XTLIPIBuvXKT35C6TP+1nbNJugT49848z23A3JU35LuS7yG4nK+CH3tmH8GX+MPiR
wL+RUMSTdtqI5pp8eSlHmjN30OUrltA7D4bvgVrC+b62PCvzj+Avz3dMiNHF6t3EGIdms8GNSwr1
TptPzoIrrWfZXVq+6ajAmX8+eN1iaPibr1YrY6B/HJci/+fHnFjVjYFKB8WygNpYjj7vH4f6Io2a
li1ZHfVmNXdWksHPtXsTnlIk1fYGMmw/d6GntzNyNsQtoXrFm35MsYcC6eltP6tpYlrKR+WZxd3f
ddyV7uKabEUt8aRyqopa1BJ+aGhvOqipHx4HArzRoqTKx87TZec0zqoNCCmeXTqVSLtaYaitjGsw
Y7jzwCChGhrwNvRh1qpbLy+NLvRJyeh890HAJ5YNg/orZMiJG0Yr+NBNsg42NuADReDIlNvpfQaq
SWdibqq10RSpMaesXhfNKLVUB61ZpZQ9fDJz4C4ZeEoFaAE8Nx+ZSw0/UdgmRuE+FVwuwXOrMmyy
kYcdgDuitGn/qW7b8oQ6WEX35gUwhC0W74VFM32xlpJ//toRH2ipQdwunYbgBfZm360cEqeNaRhb
2tITJzCOY/KvE9vBYNtFTyWnrWq+YoWwNt6KeytymrMU7eEwcR9t90zdnqb54aEupr2XKPnOyhTI
5/xbXea8eXT99OH7tf4gvoQeoce2eBCgPjmqjH653U9fSauWmMN9LRI6NYxgC71GPTGKRSlS4h8M
rCcxgf6fNtDRUFCEXl1Lf9OLSju4vFv3ZZ4lzOmqJgb3h7DYLsxT3+QsdRXSCr7PsbRjTvIf+o9T
EAXr1TUYcDSazoJYPQ71S+flD34ynUiXB+Bb2T//jB9hkFFiMA2hmPLNynAl0wHzX0TTTF0pJ1NU
Mfg1I5Z5Gnnqo8Ci8/OlWOW0GBaimPWHXi3SVpR6OWRE814XaXpGCDtHEnDSnO+zItp/taew0q/U
Jcyh9FVwpTt6PVYLePCKGB5+1U45M9weM0TJwZTX/9EBQi+BshjUxAsAVHY7oB2/kn1I+zzMbeug
zSk5uE53unme5GAG3KZw5CwXx+5nqqBs5xOdcfy5jyAk10oqwue4bim/+Ay/pItXzYZWzn1nKFuT
ftm+JrIHWB/emuFa9EDDmiHL1bSNVjYvVgJ/q1e5pKaIZP8u6vLgqM74fnr6qEo0cSRK5BdtfkF8
w7IaLbscxvx0YasYbMEktKQicyqXmEpoUmn35OzQp/NMNl6HjT+zV6jZh4YrsVpwagMImcaEPUbx
BN6xF3kt+Zf1YczsMdIeNq/ywO45FXTaHyCygw+n027y+uKIXZ3j0p79kRqFvv3fmc4iY72iuJ2e
HX4AApwdJ25BbDBRIZYlltaGYZePVjXiS9Fmdz6BhsGHXtocZMn6wA3qV1UELMCFaiKFfvPHMYWB
Jbbx7A4Kr6G53Dj4WxWw8P5czR80266tynrwCFIcBTjB5/Bu/lmYQvHzqnqplX5W49bGXt+gG6Si
pOzh2n2WEGJCZcV/pQD83R+25pwyBTrgXpYe5t2PYWYrXU4u4RX4Gu37cvmNXT2/5W/R8iolBT9W
kixGcvVAq3sutQ5Km5+QuKR9y8cHsicD+k557cb1W4gTrcnfHaH/7QGYnV8O3nqF0XyrbUEDr1DR
q0qzPNX2tYhSUBZxEibFqdlP2YHowfGME14ag5KdiedWuNRGw0gewRybfuh9FzjSE+1O8BcG7rTr
/DiYdDKjLQ1Yeo/ugPcJJSMJ8nk3HJdZAuJAw9cDetViNJPj0SsmsOPlR+eL94rEuRBhLv/s5R4a
w0nGWyiVMJvNrjuWv/DT/Pi+ZWQ5wi7tGn7SNwM2DQSBhsYaC4069OZE2skVFvXwbcQqdpRARXZp
1nqb+i6WZOh5fJSiuhJj0WmB1rIquY0fynOnCQiKavoZw9Awe//Uo1zm9S7u+Vq1DJZRvCYLsNUq
U3fO6VNzl2HySwamE2FZzqKcs/ObZUVyQXPB8UnNTaq4HFSgYscuZyo50Eh48PkAbaCtj0+5ajSq
6giwQObuH3Rfn+vIFNelh1Xu4rpgv/dMTzfvIL9kTu3ZDf8m6qxkfmV7lUb8buTTsqL3MluYJ54v
Xes4F4v8a4D40yG/Q1gm3OrfBeV9pJC5uqoRGf0sl394iB7peq6agea2/ldqfGHiaR/YssBpyYin
SUkoo4TJCFqug34h0jzItKoev0+wckSpHhH3yhm7RvHCmfsYcZuAftLE9iC1ONbf8UIup8xbC1dG
1TdS8D33odywyawhSXN/yiJJlLezYXNVCDQulBiVrsMvOjkdmPA0A4cC7nrcXInTUWx5AMOHyGNA
0j/9ooI/9MMsxbQbvDS8y0q4jw0+fBv0zHbUVhzyM83meOoCBrt7w4aRt2Y4xgu4M2w84xLIPy1+
oi57BnfzNQGDx8JHZHorQ1D5RIU1EOPlMLONM3qFrqKOiC/SYslYWFBa3IOeRSFFkgcygpjpzqJm
WYesBMSIZYQkMIV5luMwn7+XIXRuuj+dzdvoMUinmwd4qKjAiL94vTZCIWgBUAqTImwG1cDArfhq
TyCHDxd3f4cWpbVEVDdkI8Gnd5LrTL8VhCnLM2fOaO9vh1eINX8NksTM2sx6RehLg8g38dM92ONQ
sWJIhKjI7mhfuZae6xY8x7JJcSSLvg9svvC6yjmE56gDbvm8SSFQ/+5onJROGzop+8M09YTXcSoW
SLz3InryTfp71qUH+aYPYBNYD46clYti7hk0qWVb9TcBkuWQG+PbIkOOQ7LvRPPTvsX/OkL+h2PV
c9+w954Z/sSAkTq8Nb03YvvGgDydM/OBdFs46CiW7snWOQ8W2rc6UcP4rpkV78aBhm7Jk6NSd/NI
wplSQFHHKkTEQmmx/c39jXbytHGZzU1bCPR2OCUKHS46bdK3LaAVLkGzVvyrWqGgONcbfpdFiAOk
Nu0E7qF/ULp8d2tTlcW7fhTwU30CGKKNXXCbwuj0aPNRPt3tTGx0PSVm9MC39PUhGszGxOamZABm
DlwvFBDcsixiSpZ6BLbMj7Pi0YmFbPOrAKN9hCAgwCbkBJGvBwFnc/Gz8T2mdFL58xdcl5SItbe1
ucQKeBVBtFhYheUV9Q0qp6NfpDr8gJDarKcrvbblq26Mhy3a8WLDEi/VQnP8V6WxatcCyUvjxqFu
sxd7RrHysC6SMKAfNAfe4hWxn6XWZdVzn46M3ES8yQFoaBHmx8VMJkq8Lf1qs6DycXCFx7Tatx+m
QTQe+Xxy9qns4+td4o3NYkOCC+w5Qd+KmJXJKZAqSEdKp5reQIv8tD+HCSbdf+K0WHakn9B3vmvK
u9ZcoJSnxeC28u6ajJVfCF3LPAdfv4Af4PgWtp0GTMijYn2ZwBZt8jAFW5IrZFyYMnfw70Lp3+Kt
GiirlKz3LwIzat1utJN6sZGpo7vIQ1RBZjEyVMMSGXjzrBsDW0x6krnTQiUbcb/gg1eHTZmaZl6t
FpKZeo4zSOEQdtM3uE4TrF66mYRiCnIoySAtb7LUlZAJ7lhGLkwQBU+iUWi3pCj9+LQOSbzl4eZV
5Fd1mBvCvuEtbKECt84LwlY+G24zG7ySlk1Q6ucg2kw9XN3eakBJVi/wMgNuUvc499WbxDPTyeab
RYfFmnIltUHUSZUOLrPZAww6sdLdI+PckhEYJ+n9wzG4gBy7vqPjK+7SXKw93ecAL/GmOcNSVZwc
JDaPhV3e3yfhehpwtpdnsytB89mZe1UfaRNFO//v4p4CRbMQEwNat7yTJeUSv5Iornb2i81/XlSm
YogLb6c9f47nucBA5H0q/Jpw/dZf7EZYPqY0PsGrpxMcpE2NJG76QB++QqZxU5oC7BPNFuY1WT41
s5ixWaygtbnQJICkB0666aAOhNzbGPfRzHBAUAEgf88tO6WjbZvxnmFaDlRL8gKH/vJpympEMfhz
lfEuKzbGPUIpfa4Ndg9HCe6o2eEergMvqbDE1gItwQjHY0LMc8n1LoZ5USkojtzoPNRsoKXCh2hI
gBeiXxQfLB2ki47x7hOQvPL6d5aDEOM3A+3Uixhss3Q6O+MxWFdeURLG0MKGQmtIOmfxN07JKKsD
/dOLz9TatApmbkxBmF0rvc9VaU1xqLvZyw2yYsOSQopTPUDmnGnTqv/uDap6/kf+/Vpivcq8BEav
l5mL1cAfFLRl2Oixqv0ggTMuCMiR/6eZTTA5EbeQAO/XPYEq29NvuX4XWys/n84CDShqy5cHk+IL
APwnFe8HgKoTKST0decnkt25T0uD3fbutkx4qrbaS+K/G1KYi0PlE+c4S0lU933H3DQMJOmqvCiE
JdnrqiNZPC6Oykz4IXFpViZl2pI+5DVugHCv6mXGWYP1EbYhnrcMEUvkEJReb9T4bssWdiZYLmlE
e1HvIebSBIkbopIHyh1Ez0p2eHu79YACZqyBadr0ZH3y+IfCFKnAydiwcYOfjwc6UTLCEZZ86V18
WQdc42mDYGslZxB3yho76ROUDsM8tZY7oSL+xxqGq5WcMgYMCsyhqTLS/h72blBCQ3hGB1PQwMMu
O1g+ZeXHpSDvniBgmGD21Nhnix0elcpq5eXzmkhI+rAqwhPrFV0foTfZoJebG/oOpBtl8tqUWxdK
udNVuLM/TuyH4zLdKNpDfhZLEozYHwFTcwjdt7vfTVz3QxMbQn0VFNa0XlMYqCTAtYtNXYgdIjdf
8Wz4i4zbQnc0mVhxm9d3i+xndyDwK3PHl4ek0f6AcBQ0n68r8COUDXCutum2/eZ5P8YYknjQk35q
7UBuWTMaJ9wyByqpqFrTWfnZ35DRv7Ro5Bz/YvZ3koRzGeuQMMDriRnisvoncUsTioxZIGat4ErF
aLzXsbPN3PUvNep05mzTxRNgWijoXYcjBehGqJKTnTNZlhvvnUfn6mdpqqqLHUoBXVFjMnIeeKj8
YYc/j4OzYILLCkj1pBS/e5DlXhpWnVUJZ0zYJh4hbZTX3DK84IF/IQ9UKBbGJXTHbfWAVLISNsOI
ZfBF8c9QAGEKegXUk7AGA/yJBhv2dZXgURfPLZ0QvKJATpYGFhcRU3iQmn9Gmv7F3lXyKgmm2OwH
sr9JCAcaRC5+8yrOzAyRm/9RQDgxsuJ6GWluvENnxkS/HndvUZOxuVc34DmkT5lscGZCfK9/4pQ8
d0pBCCYS+zFhaKDauJhxdWGL3X81o1/je5ScaAKY0g31BKFoRWoKfY4qOJ7B+eERgf2NnUqIQquX
wWmBvjTqaZHXymUkuVRWdwkAFVyQLMi1InkTmi+jT0/rSCv5+ZGIl9edJDsMXYrUpsZKqvHejdWq
8kRrcHKekaRvaKeY9cXG01iJzW/PB+vqdQjzaPRZHzHF2SKMj2bh0Z3uNKIZFcfG81K63gUtxz25
knsz0k7ic9LypUm0TCLM3feoYga8YpWm2sNT3CvFG+BneMKrQjeMJTTpON2oI0caXNzOoEZxvL85
TEsZncd8/qbEk0K+/u3QbF0Tk9CmZ+uO8fMXE3CeDljLkZ3KpfD7UMSwyfCDhQxh1oS0suhWFYFd
ygH0OanD6QIdCNj9WS6rNPbuSdQ+uqf9WKP6K1QoL1sUGZia8Eww0hWf57n5r5vL3JTRZ8cx+Jdq
i6QxXSa2JawVmNj3H4Q59lI4gvfycMshH70PvBJh/e3NmgznePY1h5nrnCa3zQfUxU9EUm2Kj4Ti
3AcEHLp8RbcDRuZBjcfYTJ3qF42Hxba/fyBk38OFv0zlhLz/Z6v+qeRMJXplpLYMcx2PFIXb/IBG
mIXe12h/c5ZPqVMaOeZn62a6+hObrlam4e9U13s2TubH1OvBUCJDzOfIYgGhsx167tA8bNUMSJTI
nHPyR6CL4qf42gtwS/P+bQ7Ds3UzWBwak0QpiANnDn1JMprH6F6+kVHnJZ9AQvy5dEPjNxLtp1+y
IGCY5onvLJahPgvUnFrICfA4ay2ZXVF+PfYaFoQYbILKVN6/oUPE04YlCxfcFw75sikEJFUh8o4U
dHjAhOt8CljjhqSoHKjlPuFGaacvlPLOI+nzL4scltNwctBaxAGrlUjsPh+Ali8GVrMNT7uqp0HZ
mLt0mcxdUzUxEl/YjW1UQZrrHKr23V1eH9hBTUBtywq3PEb4awdxkHWiwdprfckShJNg6bUcy2Jd
jN7FT9j2/QkwbHYqlE+FyNrZHS7ZV0Xwh1WyMOQmx/Y6EZ225UurckvO/Q9w+hV8wn6k7mUGXopL
Eii2GLPohGRrUbpVaoOKTRFBGjJTKJQQNtECNYtt3znv0Sq/+HhWZQELqGDG2ucOgabR5t+6I3+P
cDInrZ/vZd5+zA+TsJxaPsQ+b+Uk2vza+jCvyF2+mc5OB5rlxEfO+8sViRuMUf/7vxon0GNN9/Ri
DGslyuDVD5mTSxAk3he+wogQX3XQabK19zRlC55yFixkfC4ZC/yJhCgrU4cVPuFLVqJvBiwSnuI2
eRBW4phro3lESZ5sKln5RcoHIRVlrlMOl7RqhUngteSivJMU6sgbJSzO/TysnWIEEuDksx31gVBr
tNT2uwKCNA8f/IUoImNQfJvke+42JmKCCtDTOt5r8WJWzV/ebS5g05jwfEmo/1L+yVApxHCi+I7Y
I+oVcwFz5z94Ig9XgKwrS7vs8RFbr58t+GSPWxUkDBG5dfsHJzjfaXwX3q3L0IpyZ5HtG42mzAHC
xzdXru/vL/VaMt9h61GWILr/6+1Z7Nl4oPzXQzqJaA0wJf2ZWcQQDmgYTHFqy4aADxLvamXHv6My
01Km7TXI2zZke06ivqF6eZnMNh0GF5OGSCCi6uvz8/ASfTdP71p25Qri4dTfT/86u6FDuSFfbPAS
BgxW9nHM+ACwqMOs/MTuhyLQz0j/tlUH1C1r7rBepzifc/ZXyhymgLECgHHwcs6kPG3Q0RzZylmf
VICdEusfLam0xojbAtB6e8DC4b2sCfsFAHMhJek0I9TtUi4LBXncyNWnUePBT/okj80LDWUcGx9r
EM7FCLS5xiD4TxjudjrL7ns2qwXCfxAcIhp0E8RlsOzvQ9gJzC0qD7mRK9xhXnBTVQ0fNxx+eAe1
ZkK22Z2vpV0azg9NmqYFhYeIFcDt8zYg7Ue83aGDtpacpHe/7q0ZlE2OcNpMa9RSqVE2ZruqOvs5
5q3UK2KOXsmntEJVo+IkAXITNG237CMuffNywNK8vbcbbsflLnhC0y4b9KTisJOZCZf3faY2zD9F
GreBQ+E4YiA1kGWVXPVq5T+/0lmMtc4ovb4e8xIrpknfBdjsDtJP4yRDiU+5O7khk/r911wwKv1C
Oh7ryptLqLQXj/ddy0Lmb0YCrmzdWNmK2JkLO10CzZrzUrf4jbvbPBAvFUfcLyXfmx7+F/VizSn2
a+cs2xL14NWfSn9eRXz/xMiNuNDCvXgMWkZeJE8cGUasL9VvycHZi/LaJRUvusD8DaMG8/HGfgSX
o2JFxGYi5VK1CK1vMAp2mTnI1dOK4BE0WnGTRaBKWslTcmPLkJQMGXWwDrDixgAXbX13xaFXBS3k
OEoluDIRqzeBhM1km1ub2svR1BXQ7gXAGUetM8dqMCBieqwRJOZcwVRy6TkquSsDFFJ71acneHhb
E/Ae8OPoNBZEMZna369Q1LBWCDgXGuIq73uBAFvkaMgu9HjRZg595F73AL8xJcFsH2feBdp+xbXI
Idya1YK6JpSWngkix2CZsYBl4QPT2A2qINjxj0S8kCf/bSdFKoMzYbKl/H0VwQ1XR0lBhilOUabF
m5mO8LcqP5ivuVNKcAy9LObvqH5EyC7Oqlz3+nW1spXL84gDgWhQc24aWmCYOuS362NwaRF/Bfa7
kbbnSoap0r1MV6QHuTeEK6+bUajGJDQVv2CTd3tbI5+mGHT7vyyN1Rvs3gVCWmiAJlFnyQqI2IYK
NFMUEsbg04Hw2UP+/L182hq6HcdagMjkoK3sXYxJLlfL5UTboe1xu0thOoGM/IdxnxGZQeragr85
zpuWqq826HTzVFwhlf/rgOtTrpXLAfR4XURK6Sop1BvyW9PbPMttpA/WASgig5QC5AeTQTPfTd/1
eRTukVzrYzjr5Ji0eaPGJkQWNVoOjYI6f9exoOGN8J05KARzlfEWkG0jHEA7Su4zE+/l7mx5ohJh
Xhkr8uVrk7OFWzleceYtPszK7T7xlFNCt0fEIfYUQUlqKR/RR9Krgmu1coXGyHX45vhILZ+aD+r8
4aHecs2wPgTDrnCRNKC6EfhUNo6+0m2bWWS0S53sQ/QzXaoKvZHvGtzpJkfj7+vEoyjWosy2kDJR
dbdDybPzgPXN/jhb07BPg7KpmRnyR+9hud48Im5bCi6wTD02QihKZlJa73o2E8G89HqqLyFs6blP
4f09E6Fb4mk6Zr0J62JwaCU7/D5kxAT81WHRFquZstt7DGjaZuIS+2lhjClOnjEpk6gXN2r8FxSC
0pSAYd5f9uAacOl5ZErpWFqxbfNsOEDmJfE+YZo17YhA3629SKt0uihJxxqOJXjvmGDVgkrPNvhZ
TEsEuAcsYah5n6cuVMWBXUiUoB3jD2S7IBqQwKdWbKUxZNaBHYrNtYpJ2/amjZQHnMFdwMzlfZIn
jgZao6Ek5wmu+OZtcGSlr6SmiZgmjZr7BmaMBysV4jVSRqgW+Lb/TvNIAr3OWrLymxRFCNb15JgF
220KZZ4tN0SL2MO1lwNcYwwCzFb9Z0Gi/yeYgr0hsH9TuIVFFwIO0y4sFwbC2fjFlXnSYK4oL8IF
XoyOtQS1gqdI+HhU4MSHihZ5QEaG9G2JxTb6K/eUKsTbk+CyXqceDLwUgOEH2P3PWDWJoWcY0+Ia
IAooy4CHT4Oa8MUWfO2lyRXFYIhSLeIhrnAiWEh6u+7g8CZcnbgbEKnJPB1Fo4UW2uh2juCN8WEX
v8JoFpLvce4hQrqaWAEMSoc7nd1gn/8U4vZMpb8acOL3xCeoubNac//Yei74AwhSCHsKrs1Qdqep
XkcMN8d5tyRMu6AIkBPoE7nO8j7fmU95dBHtLak21npH4TKnh9aYBHrYjlf1HSXFATYjJqimoYJ8
de+CUWHKIc3h04hbrcWXnylWMX1yioLcPkMbsoScgaAqvzSJ6sy54gfhGw+838ETb1a2d/SQZ+5O
OeJA7ReGnMLGTtK9ZL92symMuYyMJcIFp+MeqezzgnGavdgs0lk00TCRsdu1RjSnf8yWa8JkxG3+
U0CkTVTOl/Df4bGXEwz7Y37s1XgGK8QcbcsqXTeNR5CIHrpFOz/KXiLXfDbmi+C1GlnVXFjZ+GOt
yBR3siL9ykY9bQKcegyT2azj/cWXUv9znfTOn//HDjLjliSVLmnn+e/1wXT6PBhadZXpynyybiyl
Y7+ADbh1nNyGhhUb+cr0MZm3KaWCdabTBIEVNCvt2PaxCrttkJ3TidovHj9HM2Ti1km297bcDvjF
drhPfISWcB6RowyYpYFwhhnJGPvYOiC+VsChNMcMvNQ7sgtVBqEzTdOxgF+m8bpu9YZ7FuOYopP6
YjaVuAVeoAOK8A8DdFGCGEooZxI36agFk8XaIJY71QWpFG9fwkJ/WwC/XLb3OtAsqlIM3tKBZ56a
1sQHQKDgshP4HX3Ke8g8AhaexxzVg6eIWXyek/7g6dXwiPje2T/CwaV18o7Nt1G4gHrmxjgH1knT
D3jUfSHjsO1wEcC7ROfKPRyVHzoSjvmBUQc6nBVWM42IUbixzywZA3GQn9ggLtnEMj4QtguGVJMS
sOIV699r8IHE9+1YC14yuo3lHrF6qicwIuexOUfUeBwznFNIT5HYkkPtCd4DmDbY2IR3Rgz1rWsV
Px05wdUApsTPB9cYGWNWw7qFGutJEWhNuSCIgvREmL98zMFMChU3m7VVvfqM3+Pma0X1ZbGxqFG0
0H5WPtRGRdDMCLznWz2A6me+laeObX7XAiDQtyod3ys5FHGDEQSauqKWApM/amDsB2k8ugT2axXI
a4pIdNpRrLIfDkYLIw8pYcYuUuF6E+JfBy/HSppdtvC7Z9v7wYfdEyI8tiNuqdouhxvdgXcheKq1
yd85q3CpT7T9BF+kEZEE+ZGjAYZ/CtTEaVmz5aan+l7a8ahbT5OcrbAAMCexqk6B6X5kqRAJAzpW
iOJEJI8Ept/HeI8W/Lp4iKioFj+UMiTRM6g5byrMB9iPOllKqYCpz2eprXcPAjR8grxjJ0uIdNb9
Jr4iWY3iemz8kvKbqT5JVEw/PmAPyuXYScuy+hxBLUs+XIa/uX87zwN/M3vfEbvC7bjxQSY0xghN
mIMOlUOMyibkjM6OJ6N63YV84j6E6kbT+RFiuTu8HJHyK37dPMONy9/hkNeyS/r63kas/RyFSJwb
Fw4igi0yJxludVrhOwY5bpMqU8vYSpIKZ1X+PKicWkchSU5q2uze46vrVMPRqMeiZn2ZoteKqqFA
HzCrSM4hRTcIFJdHfd4DZjX2I2zqh6BF8Ijbx7JhstSKycq9VZ87yTK0+uExy/0ImRv9iT65owUC
d9hOGdH7kd0S6bU9mGSNXCJP1A+5ICWZ/z2fgpRWA53g2r2zSjMrPY/8+CroqKlq1zDYo0c+i6T7
36u+h01jPqw5zu+bvS6RF6Dy0TPUC96elQD1+G3gjxuIzDpu1AoP6WM2ONvK06obP2yaHWNP8yXl
kd5HDGWibBW/PPZjxjF9cuKxcr92DnFbfNPrUGTO/arcLiFUYqE/K4Tjf+nMv32AWAIWJo+icx3K
amZg6EllW6Or2cwjVgaB4/EAnX/YdLDwRE8Esih2X6F/flBAdEJeLCeNBOmEAGJRH/0GgIOJi0mR
WHM3mF9VxGW7D1O0JCPM0YLVh8HuFM+Dhgx3Bp5AwBlNTWbdpFa20WkONJlIf3zg1YpEUebALMHQ
GqO4dNv4t+kpcuWzmWbqYSCoVOlWD+1fVPI/qV2Ai0W0FfOkD1y6zpl/N+3OUxxxzLOgMkUScaLx
ifmJ7gaYiPRKQNuddcGClGVtZs3FOG5/tomHQLzBGA9+ublFkBpKMvXAV+XaY3HzHhJPLsdva7Iq
zsLXQTh+R6UUYSEk2KAxl1jUYk4cf0/TiZaoegYlkGs25WXHeaX6bs/H7k7cThn2fEWIQXCZVGNe
PVfqOkWOgwgSWNZovIgZVxrFgZwfWcM7dUmJ1CC98NlLNsZy6rQpRkUsn6HbUXuQS+3w06SIk0d8
LmTWz5zPV1E9XwaSEBvuwj8NU04Cu2a6ADcvy0b8srT8OhjMI3kBm2AUoXHK8LmUvgJaYGjGHdVj
ssG8DNuAMa2wrvcLVtYiVzSX1oW3lpTXMFeFMj1H4KPIYfvyGLMSb15PxjX0YM1PNwvtn0cFfoQa
w01bPdY95KIhUR0lE13pg3P9U3ujwgFdF26J4A017zFjNdeKQRstVRRfEyG0IgHZ5/VkhA+ZledV
HVHMbmIQz6qqyuUi/MxOlk3yBQ6zJKbNyQYUKop9eEScUFS8KVtUfG7EACffTIM/WVUfjb2z0BSF
uFzIBAR2L9nf4NTCY7Rk0kY6tQSNRg/fBcRZWwC0za1xVXig/zHB0PEXh+Z/fMGcDWoXq308wOLW
vRvmue0clOGm9yG9Oc46IkbZQ6xcHpymBJKnvzTzzVyjUNLu2AtZWkOp7tL6qZ9nmyAbs9gfHRNv
VGPQjg8xsbmu4qiKuUGBSGk69/Z0r6yrtW6wBjp2hp2CEEephHut5Q3YJ8KhQ+U+cBs/74AavwE8
TLateJjFWmB2Gty28lFOQ7Xl6A2SXqBF/1MWB+1NJJM7SPeyUqV5jG3nauHCjCnEoFp1b9Fcgr9L
ClJ1P4v21oJ7nRbdGJG53A+rMHdVI6EyLt22ZGCAZoXHcAWQvPM0uRwYdsG3qzJ0jTWIdl1PCqjw
8GnVL8pQ0WLJu/LaSr1fesN60sfQ1Z74mae1PfAcTc7UwYK2gbRAaesQv5uGEUoqUL6Wbb8gj01Y
HorvVDYnx31E18FAU1toziwMd7Cq1u6sMB4yQJlaOo8G7e3NymI3VzQitqfnt3t3bQYcF20JGofn
/hUkKv2ACV5DH07VA5eL+19NJk5gC9VXEBzQNZp0hGvFkX7ymbjN/KqKtBa7EWIi7/japRgIS6zs
OTgOuQ79On/l1WUu45+BHzwBWa389o34jMs2SCu/VGDyNQW29DAgPRt3sMZmZujxFFeH5YplNTC2
3ALAD5URXkljLkmiIxdtVVyPiKWGpMc2vfTRXMkZkYE6ueoBnBvWEBTNaYah5uHvLc8goFR8Bs+y
VUf1CUVtID78lE8JuuxZJLvOc9Q7R/Lph3aZcmvGcynQUOUARKabbwoUbFxLzgLAeIejQ4LoZfVA
ljOtJJre1yffzMppzdyVkceGW0aPCxOo9vWENaljL5Px9YBrsW9hVuAoTLiiKc7jRwwAlj+En10u
0lMwbT0s2vRuHfXOmjBlB11abN2D19n2xhjFn5aw1nhPMblecsqXGlrcIHfWuYq1weXt2l4o8vp0
jQ1EO6S2q5/qEwV+eAD+pHeOXelc45wJeJZS+K++WDLUCJw27m84l575oYcOa0C1wbnkl21TN5gq
G3cPech6A5G60NI/d6DYRG92lFt6pIGZ1W0yvBWPFInG+HB3bGi8uWcYLGqp3Abgkl6UMY3LmQtK
eqd3g7bQ+dZRsVvotV9ZVqzzEcnHGDBoa4ue5mt6T0PRM/cJR9MY1UIXEtGPSNz94TrjyhxgJfom
o2gWR1J1KJZdksy17velyLe9yZwM1thoZXvYbXXfwrSb0hXlDMAKThXHoRFxnp6az5osUr7K4aVI
u1Z2bixIwdyBRT4pN25uCGtnr42k7CllDQk5CAvRUeI3EGG6m7G4GpuIyfhHt0blU173sa3ZHfH+
JArb672tqok5E457P6jfd0/aAQ8xUyTDUEly+QLlQLJuoQScCaBrJKuoBJGILQ6Xeg5ZjdlWe7u3
O9dW/xbCo5kzKpOv4G9enupaJ4LTfhsMobRvCkg0tjbDBwFXuK+1wy0lG+NZvaFuXk+1Ytprv2+0
XA49f5CBq7h1bl1gg8Ch5goDt4Ru742nkdPuqlHZgR10XGAdwzrFms91aOoSTZBvItp+3i3PrhQG
u+hN3t8M5HdnSKoYm0ME8lBwp7PKcEglMe6YxHIY701IU/QkQl26VHjJuR1OZcB9jdV3APLpoXaX
okyqWpqvt1VhJf2HeLm8CgKCGD7WGWsvn5QeHuzxWh9IQltw9JdDCirBbJTYLCqrzfnO0WsqFphn
2O7JXvtp3LagcQcwGdCsvaFZsGdoADldlBOBXRO9dfJ82Zueq87zHqjZob1DyR7zBkqSmyN22zUP
HrHixNtT80G7q5JgaeOutACb0oU0sv1ASd4dysNf9H6hueSzLUIUxQ87aQbJlghA5P6e2yw8EpHo
oYRisRCOp+p+ItC4e+WLfxA6UwsFjlq3QI36YiPdDA95ZCyb+iK/+XpoZ2jR79cPabyPhzc2BWry
MSJrVdJq5emoHRu/scqw6CCeIGJlGG3E9sk91LyLr9ClitSlLx7l5ysRHDBRByh8YPKQkbhyqc0v
u8xpc+UqPambMGj5AmUtua/BFvzRbbvBvQyzhqKklpCmABnFB/F1L7NebanGl05L6jyNm/lTZo6o
g+ummCozkD86zJ/9cufDBWBDmlrNu+dPuNusAw7/mAz86LXL2sCFhYU4Fj+zIWsfUZDxDZmoJP2m
/Vg0kfwrq3geH4oml1/mL3Ho7rZyFKj2RQTieYNCWnhpScpSePZxKGDLhsnAp5cSt/Cxjo9fQ9bn
mOFZ2b4Ex6dQSl1tHDaMCBkrlau+mSjbbaxI260BkeiJsML+v2MCIF3+i2YPTiUn185xIAg1X5pB
+6oQz7TtFcNTY54zuziqfFSf8ylcFeCKwWx7GnYCti9jv3kSE7wkh+ObkqXGGZOoGh8nZ3YWa4Fd
sJHPeLn39rbO+owZ3FD11mLA4Wgeo5oCHc05EIHGFvbAAm1X8mxJVVu+Lg+WIXz7JPtac8JxSjdw
VEKa61zPzjOI4gB6Hfe1DXYH04HipVVpONAP/D0vbVqylHNCYq77kXl+XmNJg68o1iFyQC9Y6SS3
z0B8Y9nfro/FnNjUmuoFlj4DE7pEVmGLNox8HNOsuWeWTACv1YG/hUk4Hsbf0gfpx70AD94RfSJf
rgW2QTrHGVofbZGON44+YYpBM3CwNL8k0nEiLIK/73BmZgZvmrzySvGQBLP2h0GYZRaJGiIp7/IH
o+snOE4Z1mJlOKQy6/FbWm/FbhXDboRqzp7lQNGv5Hjvg+nx3oxm9Xv951K1SpYBNLsvjNLkAYa/
KvGFjqA8y6wze/j6RnIvUCxfMLDLrLuLzrESpQ7pQJ7g07VQRmiFlX/vfFVFGGXDGNkZ0DiD5DFW
tdMOH3WODzHnz4adHjakLOa33Ix+UqxZKodtS/xH+uvbz9IuACCJKdYUD7wy09nzhXn3ATjTMd7z
m4aYeAcZ1syyJxTaVM/rTaJoh43mYm5Ljtm5V7Pqu8cWciK/xzs0INU67Nxt9lqmDeDMBjm4jWOd
aEUG7PCvoaKaXAv9nxLPFTUlSe9r9Hnn93+fqDlbjwHc8FBxY4NfcqsM0gmVdY5q79omP2XWt4xa
+FjqN3zuE2Q6d1S1OiebQPaSBZmyDknyuT9DYzNfpiPuU1/D8eCgb3nnvz/3NEv2or9mGBlPwA6W
j2/StA2BA+OHZjmzX86trC2TNHbBMOveFg36sPUO9j4X5k5jqgNE0FnojM2zN8TkoaEw1vPDAbib
2J77YHdNRKV7uYKRXXAo0ndsYEv15P9ied0wz8BxlGcUyDNS5VMnL/WHncBbCTRTx9POfA+b72z/
9jpLE1tbRTxS4Bm7OMBP1mM3slaXKlJRRgWda15CYb440ic9ooEVdcuZFbO1eG5IEfwxrJHqZa3x
KB/nRYDbevTHOCzey75AU23SrQJDpZ0kSaqEL1JS2njmYMt/3Qgj9HdwWBKivtp/di0K1itRtqZc
VjSCW44GY56aaGhsosE4gBrfcJqxnEwdTgXLpySpb++efbPQaBgliXAew5LlQznoj9KTZIlU4fiH
daA8Gc04p7ystbLXwHaV3mpJxuL0t0F/iEQkWhHKs7r9cs8qD9q0+UpnVanXNJda6uxV4cTzlINW
L8ckMtTg5o5+iT9+FvVk7Po7UuroqDjk+3MYbU3+ig3qabPseJeAfqFVjzRe4btqDcJIlneTEl9T
PMWDirdvFMdd91YSsAb8Y6aV8Z3iEkjaVmW/0rLThzfJcKOL18AH8WTORyK7xTURdwcZBuSKOI+P
rVpUA2mglNOoZc0G5aNqTBm32MdHWZ/AxSvcEaWEEbo0WRCggS1lAy1RdFifTyrCHUAvQQVFMW6e
TUVcLgkt9duZ/H/Tb+lIFqe38VATAxPArM57zGl0AwMGn0iJk8hVGMhf6AuAq9zDvoxduibco3tB
0cUqteqVXjTxEfvHER/oElQPx1a1GWX0hp8hgaUpTZlz8TldKHl++XuA0rJ1fa7ZOTgtp+hC3mmv
MFS4WDQN9++maAfJIInLEU8hOXOKAGO8UJXQyXDoEEZfMX2htLY6FAUjHfmi65uMLPjbI8GhCPLk
FskAsSqH46mtdqbH6/pibxVKq0oF+rIJcAQGzSpIbhfL1DO1rRT+WYkaINHl72qe3NExhl+jirpE
9XYflQkIqqGBqo2wpVGajSmFdPOvJVP/8Q3nY6yjtIfIlDtx+OvjrSbB4CLdo4tJODmZo+6EWIeX
C7Fvb0D/KwiC8Ci49wZ2sLoJwN7yCgqbonR72wjaboM8QZqBGYkSoOVry5WiiiEQuQ0iFp9JSypy
W1IEHJz+uR+ywWG5lzGY4HIqEt4hQenBkss7MotScQU7Mo470IvlalI+hTHs/91MRXUyLKVOW6jH
5bgB4g2IGtByGdDvpYmV0LBM/v3nrxLGWmlff6pIjFLNAg1+rdbINivoF01LIoZ8OTcFhEsJlhHS
G6RIuAelYwR3vdWISOwJOVLR9+5yDaQD7UEhnQvuGUM3N+71OxpwSpFqSc/NHtiP+KTd5C45r1OU
klDOvHHOXIHQaxO8XOF7ZFt/+RNnWD1WagmQXawlIsW0FZGi3nK+ggN4IYtTYgE3mT3PxLISErDZ
wGecTirI6l2xPmmDzSuFr5LMWfULT/Y2D9hAYYiq0pkk0bdTtnaSKYSkFQ/fJ4iuYoda+sogwOZx
Kfscem8Y1XtiNof1Bo+OX97TmU7t1EKixPtOjDv3u6svecifnoIH0ZdtgxmVLN05rTlg7O+F5j2H
2r05ie96Fc3+pEe2/y4xEXxH25JUiN+udW8e/HOSqOQtYMPnUbQ/weZTyVayNdMMb55ay3iu/v58
D3eEjVMe/AXR7Fa9aUs1YBBnyHbID9sBILqCRn1hAFbDwxurzPBUqDPV7kjwZ9ESBVzi1bHIdQNk
F4ehejJZ1+ULovTlTrbOg62aQORAzmZrq8Sa8w7J0Ln69HxnFLeWED4+Zt/j3AnvsdjF7F8U/wZK
81TkjbdAnT45O3S6IN22DJvaZg7qQweMRBcaXpLoj9I83eKBGf8jk0+C3UfYuYHUdhIlCgHOwAmQ
QozR0sGGTZL+8V+XqzY4aI2A7obYSe5APUSv7oFaHRF+hAsnnv3+YJvEChVkGiR494c9xpdgoLcB
uOjuZeoEiecwGu5KFaUZijyZDztTUQeAQcMVB0bviNAxSImKU/HQyp/krrPDq05cHEstfG+5MXvB
9itMGvD9g1dBwAJFvYeu+kY2mkFaLfLxJeey4wDEGDny/qh/I1XmDMdKOXd9a1ozOS0Tl9Oiarsm
gzvzQigsqYpX0iKKUNeGtpOt0Jeg+yDKQVenNflo39fC5ukl2GECf8N8X2f4RMa7mOlpLfcY2oBv
O53kpxyJC4ud7kM3Dx+MQB4K8bAdcrbrws9aeWgkrbtpoKkienjDEfKGQ0Fja61ziogovTvIodVX
K1LEB9EsQpvVNWb0KrbL0af3EXD8P12Zs6k4olK1zxtJ6Y0Zv0fKdjd4ca6IeS7zzQxadvdLJOzl
3KyB9MJI2NMUXR7RhF7TN8R+db+IEeYgiu22zVHP1FD2zib7F5ztak9Cdspw+G69F6NFbsxqeJRi
yMR3tPJwrfMt/U2PAQhWgl4kirhjXGt+vV0Zx5j9lYq5HswONMIdZ6H/B7D7NM+OG1+r7oXNuaG1
dwD6R7sle/e8+5Mxqrd7kiGwQctYj7XD7t5ZTXnTh88QR/LXS5YQtU/xnkOdVN3vqLcBTrWBNSQ3
PpFVchEaYb8lW4KdTk35CvngJL4WpX2pOOu11lgwh9VrrZQG8xcvpsyJT4DkReRtjUV34DLwJkSE
wgevGkL8K13UOeCqLBv5u3J1YLfdMRR2jQO6Bj1yg5iQNAmh934DFhpKgie5D4MTYUqmPx1l+2ME
GeL10VnXpA41ilaumjjws6xWCH0hBn9FhhXkJCeavv85oJUboTggbzfZ3psKTxqus713wWoIiBQg
svPkVBde6EyaYOJSUFzPtfKRQaeL5Tq47dJrCaaCK/49HmJILSnFrkQvGmt2QGCu+dJCBm80UAp6
9zqWvgvYdmQXsc+aVVAB2s/zgw6CNUEOyJAnI3t86VQfkQj7pLoIw19wKic9UIg+AqHD2n7dTcfw
2APrAIURBTwKv6+7OjsN6Bl89M9U0DsRSBE7gkjuZslEpDd0HTZSf3J0dMo3A3638EW2glnFbsvz
lnkHVtzCsO2K1yriRYhrULbfzPdwu8aaQXHhHfM1jNtpQpbL3TDD19w/yYxcsrE74kdRQ8CkvVfL
3jBv0rmrMsXXM9aAJx5+dwFiNu7mXcf/SZzTirD+zAYpRtze77Bk4SFNauOEKX52IXw4KSb7x1yL
1EoMru/k9acj1CASMQl1ElO8cq7VxIwDsLrAH7p4gNtVWCEceqEVFT3tkK9RuHomcRKbnF9r6ozX
ecNKO6q49p0cgrQRtlWX8eglTJ5Dsyzf1/1//X02ohogsCV7/FHlyYBtvLYmhfzJtliaqvrF8P+m
nCIyB6L4cRVzme5Fr4VhV+ZHPnoqg+dJm4iSXuHdA+GIuLgSTpXkjbo083eS+Ksj9DGXoNi0XtZc
JXSmXh3mwDBOSbTxMITkI8PyMvODajEGlPM6nTi5Zp+D1XDsbdlK2/lrHfv96m7vu8HiB2J3m1Va
q6HJLH0UAj38xhgiNqld47gY+wDgeK32IKpYdw2frDLoRGpnDu1PI+qlXCbFgpROZUE0SqgMzUmu
UYNnlgQ9eqE73acypmp2WGTqcA2FX+D0SHw6YA+bO8+CNNyF9sLeDQ7zjK7yQSy4H6diaAgiKJG3
Q3sWKowhyw8eMqTsisxS4+2BUWnSn/BcvbRkVyHb17ypEm2NhmUHgBi5sXqQJq1Kj+JlnrXtofpE
VaEPle3INvfpWsB54ztDXRRiTqm9Y05ecnCHtalx/poQHgWNPoBLVwVtVybuCM7UT9uCH14Favuj
oVqYbYQi4Q96UrNswvxxPPPZ8ryXcgWz25PH5XsW3vYIprs40V3mpRdx5bLBVcF8YU97Rx3YMci/
GSak70mvu1wqjStdHWsm5tTnpb87QKIypgw9KS9Pq+iphEa85L2Wh3mz64DWt5WM04Kj6UPYcgoD
QZHTHXbvOHr0kMwzrp8OR620qlMtggTeUoUz+hCAkLX9t++Xer1/olxPxfztTxt0yAZQu8e0VnFH
dK43QjbapJyba5LkXsUGmJjDLMIIGcrNEBOHKHez7Xh22khaKatA4+TiNL2NkBT5GCaYd0La3Ak4
gMcmcAJfZMERBAC9b6p0HhhajxJd0OPkwo2tjdWLhnKd5b7/pnOHaQhH36gV0Y2QP1PZ3I5ogbfD
3DAEdKfQ7Axw7bI1vexYdbKo3f+uOORAYSGfvIr9NNlQulLhWicArtp2KAkRnr6Xyx9631LV1Ui1
zVqcG0vridDqIVO4tmbbZd5XjngGsPOkKwNGESsiRHSoXRw2xqhqM+Tluictv8k+S6l2Hk/AnPKz
FSeOgWtOEOjml5yHteJIAkLpbIMKHibQdzYKDvv4D/LFlJvRwvw3zDJj2YRJ2+vZ2KoyIJw/zPcW
rHwuZy6S/Y/kbRuETYqkTx9CluMPzdLAWkrVkB4emi4qwANSlIvvyt/Yzr2Bh/hXjUhSOXouB1j4
BjApwig9jSIxl5TEm5Jb2s5G5OcI9wcMjqXiIsT+qmoDTM/gl2rkk22ntH/Jm4cYEg7EGKu/ULRl
FCJasOb8nHkTV8ln935h3A4tjSGYtVgt77jMByEzKKKmamVtwAnSmIJjtPucsO75dKiwnVl0DcoT
LMXx7SRdneG8+7ZkufdghNqXSNd5Aeq0eWbRZg4JOjOi7vfzl05heOF1MspSyA3I5lDC2SP3BN4P
bWIg9y2LJqM9qpuxCQeYFDQmUi1vY4aqvY9fA/xiWCRIlVX2UUdETPfxCXniIS9gADoH+Ci15k6P
h/NveQFv0JF3C/jkw+sxMeltOnYp6QTpCRkgPFoQRsTPgE85/GrtfXmhlIfw0FYvzSkQ73p12Nlg
0sEdUxwtVHwE/IMO+U79jOF/38h2VBOYCxwWMKSXLLq44KH5TAv8WIBhu1kzv1n5/eERIt2FGo6v
yW7Aj8EwDsu/m74vvyvG8ehyga7DFrgrYK+FrnAF8lr+IP0oGXpJM8TM78a+bUjv+ILIyD4Iiwcj
tsbHvyK60qDdIkkoIj/r2cdbjyVSN50pLJB4onaGHd8cpymimGfdERk0Lhxe7L7oR32CaCGUCvrK
sDtPfvKH8l14OkvqDoQVhWftDwr6Ti0xbnWtqJc/Xcn7wAZ4/UasayP/VX4Tn8pePMkOgQSDGjLz
EkuRcVB1QuFRyjOFELxh6qHWCyakSZOqs//2fMN3p8MFsx50TiUt1oI21AXXTfcKhnhhFnLyDbCz
j2hpslWvI1vSKQyve6mpLQGeS8wyBWiwC+c/kzJszVU64fdcBcVCaHmi4Os4kclrvkv3M1xKASx+
BdDJrd/MFpoj9+k8iZF0QH9WSFU8nQi+wYD2GBICIoQVWcnFuru7urXxHReYA1NuTAyM/y4EwKa8
2xVdfKRVhFD5dn5fch/u9w0PhTcpyU9FbSCKdi9rJMqtcfeDcwB90Py+OG2tMZvoqjV78uEdeWXB
WAj96k0Z4+bBBhVR6xhfqj9cPMvbbux1p9lMZrjGC8wzpGguObvIGXeW+mvLTGMI6tcJZ+w+E3z1
0GvWC5R0Lq/FLHEpIgKCekyO8D2Lzpwezo2C1wbD/mCkQkBPBG+pOCDNeD0NZsZHx6gC7uUPSD6I
7G3YOz5mnx/HfdCVn0XFvcwX0zyZ/TOLbE4XV5fhxcjQxaVLnUugN98qoK7tiwjMPn7m495gZclW
lljHa1pHIB6KhqahPRFlK3ca2pTLh431F9IswFIXXL9Jc7PLEelYLg2XUtw2OeWQIW4tA+JUgngV
U1bT56aIaxn0jIOQitueK6DoHU6YVYQP4O1F+neMseg0zXymH0/R+QE4EnFKyTnhluEJe+Cbu7zr
sbkU2J1VtZiEzEFqumFYyjwkFvadld+s+exfm8S86RK11BX3+erOb8beOqi+ncQI7eUeeeh0kLTx
Jl3rIM5yue8eQ+lyoG95kBeuzw5+ZR73MEyOPWOeVgV9z40Brg1d+2mzpw4rJw2hA0kyc0cTLWg0
mi+zyfMlEhFBW/JySrrpMOnL2Wdt5I+S2syJrikzQhCT88KMuPIUyZJhBwVA2gDp/G+RNd/J0gqA
HFbIKlCmr1FGqaWsmDWdaZVUl5y/Z4cOEhe0gO5K97ETcMyO5Ejbjo5jGAavbQVJBFcz21JYOQxT
0ukI3zAtoW3fAO1U6ffs705kW1oKa2BRdjU5N4uBNe+ZAXt9sN5/annMlloosL5STtUYnv2xwUPf
cDo6Jp4v61WIjV+ZZvSHDf6sMCkR2DnTYd7+BihgN9VrP8FdfWRmEHyRVX2U90LDx0quZQ59KDK4
a1JdbSkkgnYiSyOXjGsXZatdcheogazY32BZXDKvr6EIXMgCA3XH52vGIoFahWJoGp0uB5sKFD13
GGBI6cBOP//iM/N9hZ3ORUDzqBcI2Zwk3zDVdHmQRW2o+PWImMQ578lQRcWh6moA/PhK5RKhpo1P
H4jjRUGWJ4KK9eYbx+1QShAoLrmwsk32l1qO5pWfbk+i9wjAhUTVocGDcP4WMygqKmJigu2sjs1L
62/FPUkRMU2YjMXARvRin2LXyQ5bIHmqD3QAB8cjaRNlATvisGnlqbZxYHQou64lDKtNeHpQ9l9J
Q2Y29KE2qYJzTEQo8ZFvnMiLJZG70qjq4vFGEZ8mKVS+USV+VRQ+rmH6iKROMQFyaiN/3ZBhCk9E
5YgSzQwHMq/muI25omKZW1zhfABZ0Wq9Gd7sNRpMhbWuy1ft8QUF76TVJ7y5OVCwe/LibtNNgFR5
Rx1Df+D742HJEO/4yC2DOndLxdbhLgMmHzmOMzES4LfP9Dcep5CRIMKbRQejy4jZ0EVeSir2+xuk
3Ky9zb6AOHFshPdLjv5OdDY8LK6lW0N9d0DpDLsZjWyYFTFEsw/GjU5dF2FjzUZuGs8643IfsRnt
3CAaXatc5el5Bmi9+A+AhjjpxsiMtE+LurauWxjYAV29Kjw+FMtZx0gQxLjT8npLvJXqVBLQ0L4+
PGNTIxBCkVRn4v/U4bSaNCbYlXXisaSAsXW+RBcGnC9Hmry3Jct0PcwcqZB+T14Dvu+f6ZCODpBq
PP3lMeT8r1gOHWGsBtLnI9ZlGfqsrqnPdGWop+UWOg5IMgmZ3wIP/0Xn1KmyVP5ed5mXmX5RlHnL
5A5LAJujFwMRnStGj9XIh8weJFW5I4XeRpSI91OHeJyqIbTIX0aqd+722MKr9QGcUgxPsg+6d1h8
ka1VfS0Vdxv1Hg+IsR8Y0p2k0AGrYj/JPlGtkvr0qQiGabGkL+OQXoePYjLpsqyKLBp2f8y/2MuN
XqJ2V/nxUja4vQRqTyl0hxXtcXdS2TFm1yFqiBAPpkIkNBQ4/Q0g4uLaoHBnqXoNPLbglowJ5+1t
EO64hSHdhoVg7hahPo79kSlheXPFLIDPnCogk3wNnfOljA+Vq3FLQ5GfrdOxdUhBR+nfrZb2E/te
pbV3XS9Tvts969hz58eeDflQf/7w+HViZvRpLt6DRe/vA+0a6gJZgkRcs3IqpuNXMFAzAFH52mZk
E0UyaahjKRezmHojFhbZazJJJJ81If8Gr+V51OCzoC2GA3ETzt019sQF8O09oCzMe0gbB1ZQrdoT
u52EDTXXH1SMfe9lEUano1aEjUtkXiyLWCkqK2/si/GzzANLfx0GxmPNSUIdQx8SQyw8ZpdnRL4A
79PbsaXD/IUqrO74xkfMx5YUtFWFdQ8Jyio9kxV2c/SUqJ4b/dr/wM0EbQPCVydeDOuamSDxU1tL
6KR5xhR/IpD0dkdLKU1cK3AN0pv2LCb1k+B0WOpNZuFxDIty1Hn+YV3+Q9ulaGnXtWkBHvPZRTMs
rP2NISdTYnpC7E521a6ebBWBCeUgeMCMLoiS3b31vWdpKKzm4bqpfrDzKDpPHEjjS8a/N/VN8P3M
QCFIZ17PLExF5XAvQQoGFw/JC+BxZdiTnHaMCiCrKbLiOpCF/WqZsejMDNrZ7eed/DoRWp45+dzV
LOQggvz3iWLt0hUBd2uFzdB30Pg9/94FUgA4w9PPDf1BQJgFyqwnKUzbEEEoYKXkvrI0fXvfjlfX
VdEDj8ODrtpF8AMNKTOZP82JfZc/xL/oJ26aCyQHu0Y/RQ00B13e4ubsxx9QOJhoeqGCXyJyEN0x
k2O6YP6AQc2gvYfE7l6JF+6Q7ssX7H32NwKCaM6OA0e2omxwrevyT7J6NkJrnTWtLjZHVC/arb/v
mEaTbF3+KPGpoLZ65R+ylHENwN/p4oCbhZV8FIYEPmHs0ZxFJZhTihlaUlI2p9Y9Oy7QCL+ccl9/
kcHlzduc6HnCdrXgEwypw1VzIen67kfeC2FmhOjOCqBO9iLtNUE+Jqx2C+WCrlxBxX+mbtrA3xiQ
/UdJsG2i+GMAQu4RMCoa3gSgKn62+XweusT5hw3o53o02wrqVCU2iCMj29d6XTC9jZsJBmAmF6Uf
P950eEMmYS1mVpFeZNozpQbtvmxl1TaETtiba8vhwTntOqKkhROexrL7No/h52cabxGeo1DZwQgw
c/ez8Xvb3qc/gWiHUABXT3ZZALm+QK4jyj3jIacvHuwPdb68J2S/MGOmEjj4ybMFKaS7uPuGWSy/
a66fCvKUr5tO3rW+WkB5rV1zwadq2LBnduZN6ZWi922EFcAG2zUyQYq0QURVSeMCkc8EeHmOpLsl
rUXCA7t8SBn4iKNop9DfufEy962gqdxgaL5q+c51/x9Ke6jMT08h/C7HK+xlavEo3HHAECZ5TydT
IMF25ve1K24aT22XtR0YzYxhvneAwk4gndVrFjsqtPQxluVkFvvLnNASlcQO41YeodHIihWCtmDe
fOL5nYCQaX/7AYj4nsoab0LVxYlG3BT6viDLevCvsIzoFi9wRtgiyJKmgJCa8YQJrOABPuHFAA7z
3ClVOJMCgmxa8ftwGCxc9nN3+cZJDA4rPCa5gqMTdAYYwsF2dakbhE14XOf4UaAcISVSLMbDATlo
ETMYL1kgLHDfgzDyfL45foQRn81UVdGCfdyZWVSWuJCgkBuLWRpEl7RtfNMh8bH3POch0b+7lt53
xJJNjXMbM80CZyz3vGSRcpBhloqlxW6uwxmfo4ePxHYIY3gHOA+fnvtL4ovhzHUtXs/JpRNlUGDL
3gcgcnPeARLXFc6H3kPtx8tt+/k57ES/RKS7Nnx4hcV6+Y6fEj6sKCWEj6peVLQ0QBdnhqKTKAJ+
LltmXG1MfQEvGTFteVnH6Gm4rV2PfZhwF0MO6Xe1WCqObj95gKR3ZrHwWdhEUgrosyPiHGCCttXE
EImZm/dnwiu+qtCr97vcyoQYAP4r4UI+6a0uDt827VW7pB1V3Awogh9uUZa0/XuTmHA2wgbubk9W
PKWcvalQ2b9spAY4iYT0igTlXuG8eR6HXDSG4RM++0AohJJtRIW8GfbjopHufhdkoOORa/o6I7tY
ktBrjAwsXEEBGX8s3lzfj5hd/eiGJYG5aHrK+oEVVaS6Y9KSte35Gu8QAWe3eZpx3NQyTzzv0yYI
dMdL1wTZZT3zv+Pc6Hbsv+peAL8/iu94UcolE6u7mClTGLtG9RYQni7KWVuEk1hPdqxqCgc7M7Ze
cPr9dCCB63cw2JpJ01KzvDTJLhOUPqkojI8s5aJqZu3/tkIyCpsgU8DIr7y2zTPpS1z7999yzGDT
RgGJyLyjT5Yt9jk60nX4ZPMsXhmZJiFIU8POFdJbBMUQdZn29blBgxz3JpxnhiAaT5/yn00w5hAM
OfUEgIAa5SAeEQHqARTZJGxAKmkc2BiW15lCPO9w3G5rdov9Fp39w+diVZZrroUk57X54pderlEp
OfwdkHYk6YYI5UK+btnYNfJ+xD+1srSEQB54Guh6l6nhip++1E9V2tgW0aBfon27H6AmBDoccQYi
dugDidU+euz5/oiBT8Dr8tVSCV0aEaATYwM0TptcvY9Po6fULk5/fyoJPtSZsn41iiRiZ/qj3nxg
2ONvBQnLjce3VtCmK+6XHxfKWvJQmTb4Jznfi3UR1wXcuhp3ryl1NQz06WfI70LRaaLX6cyPSsNN
zA8SV4l+2UuKsb5CEuTaN1I3HWXShCH6ESelTjqQmElqIHjZjr1R3iNhyiTKWiaEbHq2KeId8Sw0
IDyoGdMHmd7UxQpkzIAslgj3gsE9K6UrQ3k7i4WJii2hUgilTb49dAJrPCwy/v4dfveEaFfED4qY
L8XZD6P7P21MKktWM7jESWcKHpNWrRoCaJF9h/lXCiqbf40mfy7tqC1/C2BxTNcJRHIFMxyIgO/o
gutv3Z2ist3ZWDYCEd8+ratBShmCNPd4XG0nMa+XoF+28v6NApX34WKw3/Uk8Lv+GPf7f1Kug35y
NZm6Q5yYOcI4gxQBAkukAT+FOtPAwPZ2vKZowBBMXG5762Pb60aBSv1iK7/wgRkKjVTaBRmTXRdr
aDRw8xZb0dFc8YZghelw0y/1RUUR5Ub0Zag/LLm8CwBGUfpJfHZ2VPdrxFsLzy1zRvXRLKfeHyza
LdezU0cqIZMd20SeEIZOiKsACFY5g0oEJO5Ici0NdHP3HtNPBna5LZqEIrxYexsl0QCu7FvBrL5u
MVVWlDXfM7eyf+knKH9CFYWFZby3W6vDusqoc46InCfh6RHvQlaxyb4NFYta8Sqj8Y+4Kx4TDnEV
ru90ybvoPPlOm3fLUes9qqaWVvPeL5rpOWc6YBGksazu9hFA7DqZXj1gZj0fYQT/NgOfbumGc/bo
CWfmN5fq+0r8HruVvPwofI375vk42/n6xR9+XGdBfBxbO/fDGvH0ntNtg4FJT+y5A+FhRSVgxkCS
5mOISb78N9BINb8CTXFF+cNZDSg5Z7TqXBT1evSHM7GSaIhEGu/l4T9L4C+poswodnjFBuTsMX8y
RiQwAFBx7Wntlna+0aLg+U5UIp6SWpbgYxympKZeMjHiZLsWnNqKTbGJY/IS7wJjo+nRHtR7M2Yg
CEyYzF6x9QuUR2O5SVvaydHvsJtFFIXBbmy/GdHessemwIR1wt041YwFt1N59AcpQ7gIum//S+tx
+vUj1QSUWlUEKjQAX+JElq0oQ687qa7bGCxv0s+YRsnTABtox6GGpUBeaZdfX161jD+9drntCoIu
J/LZ2h8r+XyMgNCJi362nfeXDLWIaMN6etYNs7Tvq0PdupJt0hEP+0DKz3PrAgMyNO9kgSNgbuCB
d2qppFCyqCKiGXM6BV2g1X1xO+7xGO2BLg53xDTYEgyzPxJlgJoUYpTrM8HNwNTd4yLQYmIOGEZS
vRp0rpgTn7PXjkYsVXXLsYop24RUB4UzQvEkF6w4UugHcjAL8DZKZMFU3zQJpx9fviuXFxZzMND5
2F7hboX/ytVGfENYfnKX7af61Dhn1NEjDDtVMwkYz9J+2mmjz8t8KoNNr62jG0Bd0vyZWpxZI0XP
CpQGx4CUv0OJC4RUQWeZYfOX5g6QZnbpvMTc/g7IEmpoif8jPweb5f8AlKmvmNjK6PLHnNnOojgJ
PEZ+PTz0/SSlC9XWJdc099PXihyKb+TpGCmB24WocjoGwIJhTecBrsI9fGxDY2iSYxQkXW0eWu/j
1e1/xXfkoFgg4jUa4lPD3VzPFDrg+AZAVI2ldq3XIKy3lJQzT62X0XkiLXqiQ4zdROKe+PBKIp/d
zVwUQhExFdEAg3cB2wUh5P8wsqnyKJbN6ZYp02xvKA7kmRNDqY2ngRzacAVteVKvPfN9xGhwrsnp
Rmtf13dfEEXR0Z0xL0hPAiuzE9paCyPV1g41LlL7K3dF3IiK3zqLu5aboOuWDAr+39FudBDCK9gm
wLn5zCp1BX9rWJ3u67TpmII0aK1UnRSwd9UwMOhL0vZatNjSkbg604L1MnzpCHHMjrSL/KJGlu0m
JZd2TckfL3AM0ioyQ38VMa4TRmzKggAwjMXtlsplQEZaXjnet3x3eiqTrbr8RrUs289SQgPxjlMF
QnPpnVJEK5BrIW9Zh9jdxtI0VAqN0gM+NSMt4WLKteKVlKRygV8dNTegDwPOgoO8yZRhv5Q09Wsw
dxDuuGEySmiCR/8unWugJx8HWp9tnIZXTEm4k7EHUW+RhAR0ovApUVCirw60KS4Di4O6yxyaEaC/
T6ZaJYHBCdqFgo80hiJIUg3AocsUGYx9sznmkVmFEdDtJikIFyi+xsuM0BbfzQaka1rFVmB7ZSug
w+VZ656/v2fNNNyF4jymGZHyPC8GRt5TgbOAMM6sR+RtLyY/qYi3nSeDRjimNB3LWkgRyLNhRqnB
ItvbuPLuaO3kf6Zu/eLU4sNAkbCVBn0PSIvbaf0h9HhlFkByDBejmfKoDMq7jPNVz47uzLMj8AFM
Q5tSmzp5zaIkkP8r2yUItb6TM/syLXRvpSaQkKk77ijxq8q4RmzOZOUByMPi+9q1EYiMiXdTp4Dj
QK9QJCT/wb4lOLVWohaUgBwNvrl7zDKkNvKApWCkSZ41OSFcYzJkY+p3O08+f1u8mN1zli8Nb+W9
o6OXwSopK4CP0umjq4bzUAml+2Vxz5/kaSLKb7HUlOK0PtNlXEDXOx9U5yP9pJlseYT2rO1Ak2sv
rYXi4RzlfiIsxx1PUqDOG/LO7cIgrAUNoZA9na5+SaswFXnkqZSvl3rRhoTHXkkvWwmxExhhyjMf
xlowtsy672ULoSMd+bYFjV9lwdvzWw9TS4ffl4C+GgsYy+IELgLSGYQ6B0Ad1kYizndzSMml+icC
tBSui0kWRgwrk1jwZgPPNv66Q9LtEnZ/7NnO60ekYLifpsy1eZIf5ArBNrKsjRL54Q1eBLSadHSN
OcOqAaV9eEKCEurqEYKV4grNwTmbSm3WzZ9gruiCpXgzVYot5GI8t9Nh51xNjJDN00LftUQ289N6
Y7UiO3mzh3vVdGNvYXXgtQakPoNBQyGZCD6c876ICsiTljKcbA5XtFwFoA/6HPxEiBqCH6i+RfvV
YzcpLa/8BIBjh581AzYVuJH3JsOxXZk/vHTvExOD4163ho8k2V8AHv8t+OWFVw4sKFfgt7M+2bRx
TVgTz8fBvef+1gz56ug1q/gYzRJ7TZiG6e+yM49LiZUFvBewZDfyZ4EMTUscZoyLaxbCrLr7nKf0
9eiR82969ZNOkV7ZLTDMzoVeOJfjoCTxrjGmoOqeWIWQe+r/TpVtMFZJcI5uR+AT3OqVv0r0QhyI
SkvdmncuWwxcwJz7WkRVn1Zms/Gk/Z5KUwrxgetHI5oPRbCV7WmwzWu8xQCAWTj9zYGk2GbYEDu0
Ty3Nz6964KrtVvfesghnz5uwaU9pOeQD5KpcM+YObXm9hqFeHR8J0jlBlFWpCwOXLlPOcWTRnXrE
TNsSq2yo6pw4I3616yn87E1+tDhT/yzL5+WJ94VxWPvU/WQBSEO7g539ie189Ucy1Asqwt2imJeR
ut8QickC6ZS/f7FjXb4opzAf0DwQ58vwyP5CisBKaoCk7ufAUdqKKK9yj80yjUpiWHb6G+uzU367
daxrT3VcPw5QZCF50GtMAA4JMhZMqTfVqVDvNY8YdNipgoNZfvWvP58KNgP52qOMmeW0hfIsg+Z4
QSxUYzSe3468CtighfzXbJeoVS0py9Nsvhh7O4QWpXWV73N/RMtF25622ve8Ab3pVBWGU/63gUpm
9nESNuk8meAMYDobhl4Y7XLJnTOk2w/b5ILdg7QB37UAWBkzYMdk4R76vmFbed0iZyXzm6J3ZkcX
rGsuMDfx2RZERSPSTxYz8Y3hMg73cAbFxW5TbtNrGyOcbwDBV1mTmeGEvtFR7phv9xGzl7C+1yox
tvkHug+1HDwWJY0kCJ2cwvduZmLk5aiKeFDpQmI3A+Xcw+BftMLNUY9METVaZoC2QnKu1CfsQlRt
WIfTqvzMfdvpA/lU5UbZvt/DC9Sj1K3QROlKSo7cq7kvOAGRGnYc6c7MvuA0EV/nyaXNcU8RWuxY
snpdfaZRUEE8ImGt/lwJ+g6ll+ZiZZs3ToFOHzekK24hzhEShOxJtpsVZmnwZNF+YTEmpvEcxMCW
4ztLjZn/ligiHtv9B/R+/Ln6o9SJl38/xCZYhbA1b56lBHkV03y2i1z2JJ7ZY8BczxTklhSnZMuc
RpAT8GVH54Nq9iZUmpKLKh45ALT3VUaAVzVoLeBFQzDANeN4Wr0MokSUwGkqh4a4Fy9JmQWXGtMQ
8/5iHn/hXLbFW0o0fe7NY5sDBvHR1TcZgC8lp4ySjrNuwBjqDwQYHnRrWgREFtm28bTXqO4k/a8N
ymDDRTFpbt1m0+johR6Xm7yQYY9CaWRZYbYP0M+qrO6OhyyU/ZPXNNHsyuMhyGTAqUKw9nvAx8sz
cZM3QIJ7FhzLLZFEHGGaJ1CB7u2eYnxY4k+CkwFcmSyRwkLkfh4djPX1Ax9dW+wPR3ZoYieUW5G3
FvwTpByZ1mplLE4+KFngRx2T8cPOBid+KDBSRUaYyPJNKoAU2BIejuaE16Bx65FifZq1us2xzDy1
0QFzS6VsroFQI+y8t0xhS0wW+0j04mIRZ1xXLRhLCuCGDCNvpRWbk8X7doFdlmc7/YCSTtWIi+rO
2QFXwD8I4Ik5kNMwnVgByrP6cd0QjX+3fwNz7JEQo8WfsMOpNxle1O5ueTZ2R+O5Ih1d55Qt+PpY
gaTstducbbdtqmKkGcgBsPtjIayr/oZ2MxaiEkLSZ49QfM7QRCnJSV5xUDwmPIC7VRwcoCFcNgYM
diDblwK66fOeIwd2AswUjJPGcOptVAOaQcKerek7My6Gsu411myNTUIb0CQlKuPegrCyJxsaoSxp
XQ/QEXT24DOc0xZwUAGYI43PCocQMiTjLAkcsf5/bDnnLMXQwLVJcSc6mrCyXUytGHjamq4tjQEu
B7TtyHZGGrzJrWjivkx08Q8+9A887w/0qVHhBsROsIJ2SdvGEXxvso6LNse+hk3wES8gtpqO+tpd
bmThrGTs8/HrSYqH163zsBxddcXkk/NFBd9uNV0c9iVTCyff1yhvPwQYgz4ihXhkZQh5mMMfKg4P
MCsQvd26+43nkisBy8C35IHoZFoINdFQ0W0UhYlOpokHLjGRicF+WILj7x1rES+uMEZrLJcsOoYC
eB9l8m5FdMBoZlg3Vmst04KavLuAfLD/hYJGKp7yIlp2SFZhqi4UOhMM20ArKNgxzJWfLMmxgHkg
O4EGtqT8cv0LibMF3wZI/inLc+ButjMGjXQcm/fviXS5DqEffIcosIZW1dioc7QU55xQpodPYp6D
ASm675Y17+USrxQXYdyX7btTefQpBusbXC5n+Cr3ZgBxMM5vlkKk8GtpG1aQTofS262diEX5yPbs
ZxGq9VaE0lfSGx/IZW1+2gsz+4RsxuUxKdr5cM7UQA5htG426ciSO1zQpMIAqxKBU6d/OBTdOaQo
NXgi8qj88BHe0SnNkPhSiDsBu8AQSfUytPlK+FlYiJb1wrZEYJqo2cpIjMk1BZpXAFxCAP+CzN5l
pgMVQa1fQx84ZuIy4ZrZ/Tms+4VS0AB6Yxa7acUFJCNFWzzAN8LPLma/4KJmEGSsdf4EghrsjTzY
B6i91EeVSi3jEsQtUEdxxNAB4+HhKEyq9BPcCdFpS8v3D6Ld29MD4F0pO2fn497lwXP7MzlPfe6c
7pzQMJQNLGNMpiQHoSz0W+87ZqB3Ff4YwFpfpxUNROxJ9x11wKiNYNQ4pWJs93pl2nA9wZlmyplu
VSPjJObgRGSB3ahHZlpYZ0omtwtLb5UMmBBzm3XT4jaixEA1UDAQrz7T8eOWWwhtns5mbmJ4GoDt
ZHk17ZjQPUzBrnVL5nA++Azzb5PqqRsgl1PcKxiLejPdVEAANDHSQB0gYO/X3QkoTP6psbrLTHx9
fAmlxCNGRdOta29ALxTWg316G1UCGkWydBhjRtn1r35f6NTO3zRqk0gkQy94DHjCXLDHP0mck03R
qC8us7+p6wrizDAy8e5+K3nHo4KAxLbIP6ooYKxDWzzrjuDMU8TGIDUzeA4EXZHNh+8G2RYXNGsc
ZDYbkPPq+xtIIQM2GYenRFKwXSbqRxOPUQIeyAqJV8paMBaERH95c8Kp89O8W1bHy9rmAA/RBYaK
jGoSMLmQU4qlzshtRhZWKGI8wpiOXyEYIUiNqAucEYgbSiekUj7/SPp4A1ZJykzXBYz9ccBth2nT
Ior/oa+JW99C+8jRwYjDev6EPAWM8C75Nuf6Ohl9vfY004WctZapbTujhA0WJTKPbUINWtRaMfcV
+FRdgbfoZ9OCoclyOdwtHn/RupH2uCmwnRD7vYHsSLKYlkmzM3ezdoIZKzEid2SNg/YT2yr+liXh
Kb1WLt/7o4VkthV0b/Rd4cPkBrF1YAciw/nDYNRaFDPdYZvL+YZpd9+OglcyY1oc9GztMY8gBGvd
49/bLY107k91lxbgLR7/DFzPTM9zEff7GdqM809vsN2EWFOYQY/qKTlSEDSqahi0aEkpmNNqUKoI
zELa7wMpOfKnvoAkl1WQ1hajG6U0NAK2TZ7E5R6P4pmBRN3xP9RDXqT66pXgD1v5xO3g2VChH5ab
C51yMt5cZJylI/6iHZb2B7dkxIK2I7yrJ3uThv/yBC8P/2zHUhfWazBpaxGipvBjZLH+ZrpZIoMQ
2SdHVDcCksLfJlU7fczU2GeOLp0gXenRk8TvPcCyvVvF1Gdzl0WDFJyBxYugTaKYv4uGEM3/QzIm
8nNqYoOqomb+uqkv6qFZVTw7AkGcJ+aLqFElD1JwiK/LdN86jRiWr7/40eGqf75AnnzBF2jZz8sP
1TXohk0R6sDx/9bps48+C22zznybB6lCK1J48hCweNSQMVDlVfN9FYVcd//rRJEQQBAq5sy+l6dV
ebif0tMfp5IkhD+eTSwTZgug7cmtwsEIXOWMXdYNtbFMVY69V+DQyhbx8yOA6e6yajeOZoPIs76U
5jlgMjKolHILtQBIAssTmcuFq0ieDefiIiKZO4d7Idz1MYRQs+v1WZk9Ptk1ItOoR3OVMzRaANDE
GoZoeHSF/zl+qEXqGLANAO2JEd0GP6jaucOIm/P73Y1mQBkSrDf1XAGtb9NlM9L60mTT6b8vKI16
C7UAgXa78D/Y47dv8cCTp2KCSmBrdXcJX8wj161qb0DIZeqxjS+zXE5PHfYT/qG6Xm3NbcgdmIg7
xVRAaHxGaN7kqaaqXGZnV5OqWDSZDwCtZMjNJk9CvBQsRgZ05UpQaPTVolKFhpIemRxzuTCFSVdh
DJW9A9WRWv17P6ZqpJZClqagn1ZgL7r/5tnrUboMVEMn0rxTZwj1yZpbI37hZTnfzdkLsiCI7IAq
JEoA40RxzgVLejJQYACtOod2OCJZNKkVoEwzicGbZri9ocSjINw7oJSJUFNRSl7NIySPOflNBJfl
RUMB+ar7PnDvAn131dhXcpX+CGJPQTjg5PP7yBfdueOi425IvJ36BQDylBGMp4GkH+MH3gHGqIzD
gHLZONljxHPO2uOK7sddoKnCBVxumZox5xeI5JkNuVmivDk0ozxgl5htKvpiZjocW85b6sA1IOGB
ZR6XUXI/pfc0uzTdKrWmiAPh0S89I8DRnpe04cRIwRGiMahO87yC9pLk60NN7wLZTaxX3OYycoJQ
MKywCMDbTw/0eua8HYrpztyQT0WOWhM1k6VdYCdlRT/QlveSqvB+AMVjPz3OSbMHpKzIcSU7SqYC
NW9E9DLQW1AH+VNXNIBGSJYLXRT0sxM5CmyMZxByBDMVQsF4PCmfjcOCeOG8pwzY0f8o7xjeZXHS
0BzI12biuEqNc09dNljG0mC1P+06PSsAruug/T3TyAGHCM4bqBBTPbBK61x9AWqPfTt8du9lQKJd
Ib1e7aWoVFEZZPNIvGKJ7WQOz9Iaz6gVkcGqcq64WIN5srxLCKCh6BjLFUhm2xD1zSYCUMLoGDde
YJRrv6Fd9qBK0+HGirzQhBu9g84VHWVoEUUCmoAxt8A7qy1bRW/wPAhfox6vNHsdWOnzCM1QDe4q
xi/XiqpayHfRouGCnP4NP3vwQBef7F7Y3PXyMkIrkHHQNR1+xg5cdGMze+2o2gb8gTguKurR6k1O
lDKFIZ7m+OVNs4XTe47ImjWXvlED+rP3yC9W72zfCJQ13c+AOMm94HmvzIPnKQganUt/JyCc9Y+6
pwVLvStXRC/LBnRzgsxp2hMtUoyqrITSHEyv27wYYR3y4qtacMqzxJrPTJirZz6wLCYOvgl1WpoF
/OpbcT75RBDK9XfLD7bZHWH+zAp67bELAsahrYW2Q0w8RZ97NI/Yz3ka5rijMWvgaZWeYvzEL8pk
HKa7XROfRAyLuMlSbP0GDkBel3AuFgV8X64LWnwY/+6FW48WuMDuV6lW6iSki2GkuvzqjfPWrLG4
SJBzjsTZUjJWpMBViAQtDyFwNlyLlPN3ud+XqyKzCaWbddAjh82YXMX86ok0aVR10p9Jw09N/f8d
DvBDJBrnte6R67KuX7FhmoJ5Ep2ibAEJd0w/Ggd1aNilohG+ZUOR2T22e7zZhy0dPuVGtE4BVgwa
WtwRJXySmjaKgIqosLP31URiPE6lEXBtwPtHF3pjfw7z5tGVAK6v8m/D7FfaLyvWSuystYTIrw6t
i0ZY7rmEodR91/p7/j8hC6ohiaIKMGS2aEDsIOOeLyMTbq4vxeyiNpCz1mUdmG/9wLS+uavO51F2
hEUczolLSkQO/YzO+eIgvP4k40fjxqTztswUUCqtJv9AXYTp0bidz9vs8r0xVu43aSBmjarqhm1Q
Nv9O7oIn5xAvhmNcO0THKvFYfYNqnpNI9ZyX82VgK76X7rKU3KrpO3UcD4ox6knMK68+05v7TQ6G
Qfxa1Dugo7fPeA6gqVgDYTQKnbNTQIIT2RRjLKpS/+7FfaptqT737KA8VhrHOT4n72pimjTEqRqW
MLzC0QUjf88f2EUZgVfzJH3mj+ev1E88QoMzjkHPD2DwZGMpk3Sv6ZZvj+VSUBg81Kedqut0+1Qc
s0ht/xFXHj61AOAq8eSJ4VAqXeEDIY45aZWub/QH3KvsVTSHum97ZgOfuF6p+WrCJQwcHp/BI/fF
JvKrTAeuNllQ8I8uohojJFo9rtVFURUPl3HsKpiI9ci5vUgeMAke8w8bjBeE3QhsowRaORPd4iya
t+Ek2L/9hhmslufTsEt7xrp9vIApP8ZQQv0Ury30mltyFtDOyau38vyutWEU5wFgLuqSvI60IwRs
LTd4F5p+tmvc+tVrqmEBM2qqOOyam06cymrlIBHznvHB/COrnyUmF2iTiFYIkvFloxsABkZg7ToC
BUCOvCx+mZCxLF2+br+eyYNTRD8pFb0C/wCUYz8Mu9xJ/JWDlZ4z34/OjCbraSvrYB8DZFTIKy5E
ui+qHSM9LPRgv5kVneryAQcnMIVveeWb7M+FiuFx9KHNDxa3GgMDzcBqbJk/4pctrhl0H08rkFx0
wbFy9eMrxD3ggDKlSzjcRIspU9up7cusU7YwnTX1YlzZYSosNL2iyazdOJBCSVXjBz5kKsAuAQsc
iodrkwhRoFYV9/wgRSV4U/6/vp9QCT3fMFtw4rWprBGwlwi7Ugyh3+Xch7DsXGBVg+H5D9IJeWJq
UhJySRi4MM2p+Jj0fKlSf0Rxq50SCh2kw2bkRy214ZlKOfm/Pj/1LOiKmEWlAmMupu4X5xr/1qN9
60txaMuKiMTS10bSe8xHwb74XRlEVYwuqVGPwfUrnf7SKqRyjxhpM8eyqTll/bRmKW1PAScvQe+i
WE3Edb/pVD+Jg8JwVuvsIyjfF98bEf6Y0xkJ6tt6oFd3AocScxbR8DDpWg2+JxtFRYx/5X2qPSpO
tZT+9bUEW/aKelHgVC9hZ/7sUFkN6jNUugphix5ugeLN4CUP3LeWwAJYnwRNclosdftNMkucOsfz
n7KfZJgjRFI1XgYmZ2NrWiGpJNHE+gyJth/nykbd/snuNImUI9hPDQExPu25NvDpTnZVF6/3IQtY
jKXWBw5R27SGl2vuFd+V6+cBChx+jA3LrBMq28D6zKDeWWPUvgHWKqklYA97Ed/ZEOZQiQFfvfxn
wXMAXfe/A86+lXdu7abbGZ0s9H0bOzv+nQKSIB8BsPM36i1JJL6J8lxADE71zW53AladXLWJEOIM
AHViiWjKxoJ4nfoTpLqF1baRr7OPJqCTCFarDPKlzUngSnS/o4L2MNwlyKixW3hPLZxYgxPwlY7P
UtKnv3lf/ML9w09ailUTQaBm4+J3PgLCGG4AOHS/B/YFegEOqR3ISOx2/URfAjYX3EecK2IBMkw9
1Z7spZcUQyFeZbbOdxDDtZAliNBvtShTNinlbgQze+pfLLrRw2aLAtAp3MMquwM1N5Cjiemq6G1m
sBR5o6IFMqK2qnYoSl5Cb69Nnauap3q9DAwsszoh3DNUToWPo5JGrcdfO5Xlq5c1LObMLbf8a7hZ
JlINPLcmGhOVYzKgDFaodpfwtXKZHMIkld8u6nOngxqGbYJKNR0UdbUHEh+HhZm1q5qiwP6Stw1M
KVtic7ZPYFSao7HFdfo9C4uOE+YL4LfRsk0034oqdgdA4u0DOY+qqm0D6Gaqcg7UHmtabu9YG2FJ
1+7+wZG4TbTmOXRTHukwbDrdhPWMYCr9/B8ut/bp1l0tEFvK1VDjIXfYk4Pl3JtdwkRXQn9Wk6nf
qMQubp7b49J+Aha35NcuDO1bPbMY5PfAs049eHuPj1ymF9CrLssGvDOM3P5VZ8H892s7sIjskX//
Zu89Nr8dd+rQcmjBZpNDNI3Ig8UggKOjOumz+aPq3/6hq3YPZjwMNQc+JEyBTGNrHfQ1+o+f/JOn
zooUQ2nHyH925nVL+VRME1RXs4GNs6gLZRQznn1UbNrKKb+khpmIthd6GH9o02+TY6uIdfERo1J8
17VajHdxEyJxXB4XskJNPZZg8cbhKBUHWN7zuxY+yYeEJu3vL+Ly2pTfPkZSsd8V5DIHLrDFqMBZ
7B1FtAEiYbNls6BbBhgpFteTbBvPsDHEIFT545nnsmLfx2j8ko4Km4Daouz/4Yfl9ovF9oFbeKJx
v398Aj6ZpBU7JP40i8wlTgwKgi1LtNBvD4FG8cyzue0cOJxDrnbMAB46Za0ORbq6L9c6bEMDoV5R
ulPD+7zSA/dDY0LAC/9H4NhhqvHPfSurP5AfaWKiMMybdDo3+FXrt1XDEt63bBtBI9Wabx3YT6ah
c3qCodopCfgikJOvjVHn5a0wRp6Xh6Y1sOfIHlvxrVFdsXHOZUhtGqxHkked7NjoGz/uVXPi0Xhu
4X2jEUpntCaDzneor7RLpzf/pBjOQ1wYGfzv2jJDUna6Jlrx1bFxnOiWDXoMzCAXvMEP2HUzN60k
dbocKlorTswYouBy7varaR1CDYj+Au0jzN+kJqxaceEIZ1GwHOFhCL/FV/QSlmgsz+bVh65pf5mQ
dlhAnb7I4F+iMu0kzbP26PdWF7q6KEENwZcG7H2axdTFoKQUgxRzU2JWnAYUiTPKTW2ICOUwRIUl
DT9DtlRZhjfs8HKcCzv6/AbP3ZkVqEn1Ivenab47XG/B7SGuJLx4PeyKmFFcoNui5orQOerPmq3d
4OGBRTGE6Zt1x+2UKeNVr9+VRLMKWdmCdWX5ek90TK8LD9CzZySgXWB1qzQpVMxN6/3iMcpvjvno
T4TQEbnLOD0rm73mzFtmkRsyBBiXQneI+CNsLsrZQtuuqnjqXkmufVnkzSkTEkaQpWWkaaeqpWsb
vvzrr6Z1lywKqgqaygBQ89VutIvN0tMFZJTPhrDSlHLcLpo928P6+LmNqutEikhO+ynoc/qXs5PU
LAqkyBZ+4rZbiPJ6BDOkavo2FeKEjXRMi4I43Qr60qH6fJFfymWDVzMeCiN1BjJqPHZ58d1VrELZ
tF/jtRDi2QVr1DLuxKY9OPsXLvaXIBxVOkm/+KkuD4RFDZc3O2xvIurvwM2INpmghTTvckcgYU4l
ecX5Sfj2eNfiXcNzul6JAnEuPF3LlxFPeguY2iU9cagPVv13zzYZyOAHPuNgpcRE6eVQwGBCPr+i
tDvc+JtZFw/gkJH2TQw6ZIAXTTV2CU7FWGsWgqVlkGA4ZftW0u5yqp8iSaItB7P/5CnK/iN6878S
7IO/xwtjpo/Q+tNEA7tdFJ7UONKLMUHN41F4lMfVBtH/VYdNiSScMt8mZE8YcId59Ts5xLkcqy/a
CHn0o376cDCNmXnjQB4Dc1IHjn2B3NatUe0Nv1uWp0p1mvT8Jnn7tLYd1bYzDgFDqPGobyTSr3VI
awNr+y5FGowkFJO4kMIq12bn+WPFq/KrEkJDe9wivckVH9H20iO+m6Iyw+qLPrsFt7/apcjVP0s2
ouBJFT4wGGc8pb0Slm8YLjzSo+kQXmUOkWNEDoBRiCErTpfGZfEgYqy1j0FcciP9qbpdkkrF+1NG
JptcFRr2/NCjr7Pgwrsdcgjf6rLoxkjsYkEj8YKqnPGo4Oh0PyPzz4g6Dcd7n/HRrdKOLMTTjO8K
3jPXUFC2qQkm5loqpHy2A80hw4ec7wdb7WaCddVTKqg57CQurhsynNN79ZFb/udT5vrXS/9gosQ2
xNTNDarbaJztlvFC8xQe+cV4/HszVUnd3H4j+QdXZmfOiZc+PPMW8BOASNrkQxdx6xSkZkFOE7Uc
uA9ArIKxq+rzqqGytoNP42Ae9LtrklChrwpm51KaWvGBTuigSve+Sv40lM8SRymDRXRom590XBWS
xPzd+PRp7XIm6oS+1Kn8s21zhhNI8A8TH8t1T7W5x27GbsZroUVUwx9bF6LTCxqPlCYJ6k9UYoKM
eBY63BEN2rX0bDOHmp6iYIfPnCNB8GmqpDv0WK8S/48U7MABAZpJhWxjXDX4ke/Y/NmNRQ53wwc6
85FV7SpbXrUBXYmqjb0NNa8O979gc01yAMGcyF1eeWiUoV6sJhzDj8O1CM83o8IcKjYlT79poS0f
EBYykZrw28sNx7nbddG2xJJC6sTRuFJzC+HD2MRJK8DyT0YtIQXNgy1cwhLixzfhxkqbKPvRVOUK
J/+ywPMUAZCM7QzHtZdBER1BfBwgEG8+l1iTYAV94tIJPaM8raBEUb5OUTlO8S87zuAfD1ONr/0x
IGg9ChXg4EjQKa83hBdKQLHy5hHbGONqQ2cKVAELRhiPJZuHNhxA+hBv7/x6DBmOnBSWi8YjSNRN
e7Vcen/WYWq14AePou3m76xuE3tcSSVhLcXN36D+6syvdY8Nu5tx3NcZgjwKhIUgODWcQeCI5wD+
1n7EGdmgvur/4u6+fUkOPY2c7BLY2WxekUxnZLM1snOsu2PlTpyANC4oeUNwQpACkrM2yj5YEwuA
d0FIsVsf9z6YgA2VwHDzu6LkHPBBpyLINpkh4kytQC8i561T0TQQpbgHTpkhTwgcOllyf+s+NZVD
ipgn+dEv0px+tayWWHzBdgbKj7xvmIuwHpJHap6JbIA5ThHLK5QJwAanWCVh5Jm/sl5GMXCNkZpD
hn7053LoLoewn5knrqkpUxsj06/hec9yXUjBGq5qCUlZS1nkpS4RM5UXDQQgG4A2eOubTuSjuLBx
+AkZ4rSn4DBi+iC6KRc6TeY3iwin2uj4WK1F0yCM+O/GXOMb9oXwlMw24CT/RjtbNftmvHOS6DPu
Op+QfeJqXfgVlTEyTjGBDMjYj/CudXhlihK1QZkA9wENHzJuo1v5tUb6VJfse/zCkJlhfKKqKf19
/peJv3wyQZ/Wjm7Kfau+lb865VltYthdLC1gjSM3ODhsDkhffFwnG5YGGTvj0wPChVCTFhEKI5rx
PMO9mf7cw7zEGWw6D18KgpfhE8YNfMAwObYD9boSA3PzbuAvHuEiGQ37M7cR/2VW4sTdNFB/2m7Q
A0tMoPkOrZLGFJ3rtJ/gBIGBM4OqpKRx6ny9Ux+EsYvOoE9VvVUwsb/Kzqnrn4728jDcc4Iw7Daz
rCEuM/rDSsEf5PZnwO2YLP+UWTN5LdkMQTiowSdALZw24Us1n/5F3/be2VXAwgL5873AyL6SPXCt
xXjlxcIbK/5KTMnlcpSiY8mfBRWc59J3iN9jyiyZaYUrOHznVqUDFlsFch1lHm7FWBkc0WhutUvR
vOnEa7Q6QdBjq2unl4K7bmqea4x9dJv7viD2oO49V8rJPulAtqG3LgHVd52OrCevmRuE+Lu2aWpV
dGKgZJc7LCf+PXq0g94YNj7Kb386t9ZuzuOeBOZs0/TFP3py5tQORQQmOmIS2re7vqvJK/fFdHjF
nz5KidCMhmD+LDBxdCsWlumfYxsFShXlLirEsBGJhczoSP9AdDBYgzEGpYW+0MUl8VLt5fpYFGKO
241SqdoPTf5GR3ZTH4/m+XmDyIH4h/z+xvT8V9GproRFV+tY72RHkLY9wilMyEtEXOodwzl5dxZ9
x4BqD+hZPwFfVrEe769jjpQ6loDi8ofYiQjBXDa5kRFvQQhbbPXnColmPben4a9084hl3eIlb4PX
MHQCF+HuKmbwCrpZPsA+7W9wxSlmPGXSvxLfJ/LsWw2KIxzusWWh+bzGoBhAzCOHLfbwgzCfOxo/
SQhJb+Z9gO2emOnslzggESOWde0lxVC8BW2CFhN+HsEwh2NOm0Lm1GTetbOs/tP91m+eyV4zcg1u
D1/HTyTLzwxObElYJvJwe67+gik+BYUjDJOu1sU6LnxcYapZ+1/dpVuOo9+88ZBIT2JMXi+2Be3f
NDH6whBweoZoII7Xyz+2EKgeZXnSjw3W1t53O3x0Dj0m4pGw3XfrumT9ASvhb0EOFTcpdTdiChbS
RK6pGclg4mzjTfpX9xkOCIVVgWHE8ERSFD0Iwj3t/RoCklczfktKrfhbubjJpEt2wnzOjF75cMjY
LbKh12wbG3vI5F0MUMU6GmpB4k1KVszeP8Cw330xN767KDFVqAQuAXB9vRJ4nQe/lTARIUOj3JtA
tIza6XT6kjhQIZatuhs+UPm+ps79ncRWi1V3f6LbSy0HbpjFKLWsgn7TDfXs5AYzHnoQtCI55m9g
A2+xxdUM4yLEqZwrqS+ghrRrZIsHKXSbZD6A8Z2z/mLmf1HJYok6j4jr1zJfP6p6Latx4bqMlXxk
dMX+3HFgS83Zjsm4JlYjz43en4xJ2Y4MLPlN6dQDoecq9jnKyLQfuI5kaBUQWDqni14zVgQGtS9z
PCb37IjlA70umXYp/AP4HHq8Qw0cl+Uyq1Pt4BY96DMSL+ggMohJ8nj7GEBo0QVLGgk57Ec9sFZT
MXJXtNucDO70yzPWfwxgXePtzRjk2Gv3Nze54y3WJ0dNgFRGlJf2M3IZgR5yrj2uPf8gNlXQz56y
c3OuQEk/e69LdP1ie0maVZ5eFR7nTdb3B5rRloAKs8Ov1jZWAwvL5InFf2PXw1CTOAd16vEool5P
qzA9m3VTpTO9HXTA3mcrfJeKHa75RJAWJ6Zjt28y5vGm0hOwQ7EA86nPLz6enwLJbQymdgdMjEcV
mK9hVzsWNdpe7w65VhxyveU9OBSetoyQNxzxYRdWRN5iNmaF6U6QR0UFupjKl6/f9qaJpOEUHE2a
Ur8k5CiySkQvnAN4fzbAFHP7Rr2wpA/W19jywzESAo30huPRMl6th+7NODOshMUZOFflGzIEOHDD
o9IgO9N83G1BXgeOiS6hx6aqYyy6zZW8XkNFlMs3iarydAVm59Q5cNC6J/dHU3akAk/19mKqEuX/
lnfEZFW/Hqy5qSlylBZe+cmb3oj5EkzyPeBRfzSdHoblpTKckdhlEfjzeSywSO2t+kMtMN5Yv+YT
p5MlqQ/OwyhPHoUj7K8/6yv+ZQe/zMu5x6ZDdgbC2WqWP96t6Q1HG1N61wjD12z1jOlj8Pkwgh8g
g4d3A8taSHaYPJTa3n7OrgZkXAobv9S9scPFEEqnRMoAW5tCQb+ZtiaWyGgzTT72byOCQ3v0EQYY
jVH7OGeZZX0l6Opma7En9/wEfMmPpEXR6J56IUZRbijcs0oDUt1Ti7wArGVDGngRS1ykCCulZXum
nVWQDORyRVGRT4F/6XlNiE7jfgL/cuQjYLrhKZzVfz1PbpL4pLZ9iE/nsBNOgiLTuJQkDFlokeGo
EO25QSV2OO6y399oXecsoXyhqRdCwp/uH71Q+Sy20F7Jdl8+zshbq9v3/dYPxF8qy7SMuJu1SoJu
iZU7EhApp0TKVk+wiakk4EH1CuaWQap+96nOJwiqvzQPIJc+UKSjYRFHpTbmBZB3iWOLBa5BYrTC
3W+s4F20LpgJHT2gqJDzIgFwTMDQETxauX9X6SwrBS5/khnwq0j8Y9ap7voEYmcYvZaZLkJNRFXb
zFxzzFwSHjyYovCSTRlowXkIsoYSbUzx9UXuSXSZvbagMJRh9g6TMnrPY9q28avUeWpjhDtjqzEK
8AbcgYtfd4FoAeA0U7gTw/T4/hUXZ//0O2kgLY6HwgVjwh8AV1sIIvoKMjwhruEmMnNwu4wU7j/5
TQNHstg3ovDtL/JWHsgJOJrds319VozvmHQzJauGERTG/+EzQYwCu+pOj73UTm+EdX0+PDgCEir6
XUkgy0txK4b5xTAKBfRRYn4fMFnBu/wHYXENjoTLDGaE8ihOJ+TA6zQxR6CWUJT7NPySfrk3JnPS
wWEBoWTfd00XHLkELHdoq6dhlo+htA4c2H5n9Ti3cDHupYy0eOKj372e+TzcVioQDQNwoeD311Eg
o1w/hmqNr3z4wjH1iiwUK4+giJuI54pGnAEDoUx2Xg8cfDUVnfO27ueDGGUf/fP2vayjiVBtQgyi
yf02XsPEacfA6LzKCD8eACxay0iJB+WIPCM6cxENPXI2mscXo9XCaTtxdC2uEy/vIbdVDfzqbV7v
DciegDrAyDoRp+nix8/AU+sAYwIa2gUXgJGkGSJH4XcTLYR/sWQqvLpGX2IFNF7NSWiqWMu7l5Ci
JuTdoVQllTCrmo3Nb9VCWGRiXTxj82/2u0TQkDUsuAs2sJMWqONom4xHtQlvi//isMbTH6xjAVY6
KfG+sn70UByD2PHlXSyWB0aJXXFiuWgqI0z1z7i1Jg2MjAc4HVEa4YUqmb62//8KNCzZzvrygwNM
WXw9OHR6ztJxpQ3MvTO7d956sqgia8x2dBosJY1gVYxXgYD5No68bejaupCo4+RubqAWtRU8nt0M
4S9xOh2vtVLD7y1kBlesnFAVcgYSzGEMgveuOifsJiNJrUP4fuZxRRVe3KLbtyK75O/wMvGw6FKr
LDbVGoZMH/Rn7tK04/oErShgFr4QDx22Ivn92gaW67Bys3D4XGf7QmbKKo446bvoP5HvdF4zFIdL
JSii5L/tYip0ZNPyJsoEEeZBzh9gDflgeC2T41lMF/hWBx5y4X1Oh1Fw92vw7qmJRs2Wq0u5EDdZ
uRwtstIk3kao6QGwuMXabCIR3bWLgJaWqq79sApJ+p2f7vo2Tr0AmAhvkyPegrjsgguaaOTmMqWm
igU2KGv7pQafDx1u5emrwwFv9Ht79z97VTP5E09BapBsJaNmtrnsSjxb5LCLCkQNyuDJ+bs0XeUa
l17a9b4WcAvxIGDrXGY3RMlQT7O8hT6wQ6D/V079fhQpb8q3m42qU+I6NYwmGoGfY/9EqW/MbaBq
b87FzdvRR7SVLlVyZ7+sP2AJnrH1gT7CsNklPiIftpV79JCKJ/IReAEHo3Q/OFZkiIDZAUyuwTlB
+nCYdGaDIp+ZK2pwajVd4AqwgrhrAyJ1tSZhItI+eVTV3+YWgrQ+Kb5ilBgLIGbSIbO+dmkJd/00
uv+mBsR5rqQI3jiEXLmEaZN7RcemMLfutolRIiH1QzlV+D9qiqxJ0qI/rU7mLwLX1BsamcTJvlIL
EtZu4WPQG/Tg6mHZYf8oaVLeE82+h565syVmLv8AEj+qks3QMtqlbQ5jukOtWQBOshZ2PqayVT3B
Qozb/sCeIK8C3GhUwWtuGNcW0wzjoM4cMiPQskaBFDdzEiQuwqGihTOh8cJXzkpJZN7BLmkiCzQD
Qeg6hv5OXdCEFft5EEeEx7JCR52tOb7V6mhePnUAkVzqVlyBpLHLz7ztDGueF7P67reCgjF1M6Tg
QnEy/+nD0A7eFFtI0R9hNOu9d3o4Y5kxVt95/ggmFb5twt2Wv5O72kKkK52fvHGdf3IuWM3p8zv3
Nr0v0FOtw1vWNwnQ7QnAARN3jxKewDYo92eRgazRYdzRWyceYtpg+4DaewUsmDYIGBRDJqUHff4C
t74aqo6R00Ox7Mul3r76Z0GISVH7UTWOKAyFs5ACDuYJrrUaXG2CX4yuTRzJysPLewEa5f/2f8XL
LqQU2ZIrPF0BcMFRS2eNpBEMuKsHdESEOfk5qnMIiOjcBjx4a6eYuGRVy3wGkShvHEHWVnPc9R80
75hLuJBSS6Vd6S1BNuIl0x+TJQnttrCc+in0vIFVnyr/n/U619pC405h3dZ5TlXhcQkvI7GSoogZ
V1+DLagXQi5Czgs4OBuIMHa04CZga+TPs4S9dJp5LlcGXMgAuq+yUS8hMtl7b39PZtikYCWFTZqA
mM7XViOCEubsnGggfc5ZPqDLQCjULH6c4vpJQEBhsR547zJNmCYgKLnQglhB5MMa+XTWE1AanWb+
vnDg31UfptVvYIv2DpQ6789/ymtmeQDHJV/X/uJj8kjDCpaiIFIj3UkFd06YejjPeZR1uZP+miyu
EXfEynb4yIxbbb9WqZPCl6Yh2MAHUuQR6PR9olJ6PDOG69VpDxuOWUF83AsgF7i0Z6CRTIEMVoE3
fD5bwxJmGrpLWeoZ65DS91qXveyDI56AhIixovyEpxA5mz8Hpde4T883vBJ1LszkMYX9TI2H9CEa
m93a/G2im60QpxYRZx2TomCZ7mLPOlHHLspnXQi99AN7QNgh0/iMa9kegbqI9VaITNRYKL1Mhox5
XXcELjUFK86nLCOsmM+y+lqed4EOP+aHy6qloAQiNkkgQpiBcx/QRUIn0I/EcKksuddrmRmFzI4P
D9z923SMzU8rGwMqOBkGmmfi4nZTmEzG/xOQastmenitirWpsTaz8B9hkMyW2RtzxKzuhz8tBFR+
UkyT/ikSJyBoEp9SkCWscRCN93ZYba7aJdDxoEbCs0Fefl3PhpvMMkxCfYS6cCZhQVJ/DxTyuE+n
o4/0Ek8m3LhawmIaOAjnE3z35vKokaCtt4uao8ka2zvmd0iybyfN6WkSqz8Izyq1Tqf5xfXJ45PV
TNPzhQUxMnZ11Gx/++LXAS+/vs7f/sHkxMS069x9hzxrAHiZZNJUkIXlx/TE5Q5dUU65UtPbSHYB
Kf9eF0fdkJo2n5O7zdBY4JnuGE58hIELZ8P4dJPVoVMo0kmquhEHSo1QELzMJ4acKUkcq3Q074tM
c0Oe4BVgk0N0MS+L4aNjlm8E/Sarq05/yojHIaL6BHrMKLyG6+AaWFn5rT4Uo50FfUrP1CzB6Xcu
NhJMQs+uqzRireTE/7sT49IX4g2iW1UaGLCd76g2IEE7GHiaZrRtanw4Hv0kwDn9ItbsUd5LFfx9
E5xd6UeV8n+5ZEyk5Tv7havS+Ed1b83LThkrg4ItgRn4jt+uyiqfh0kMs0vZ6cLAFYmLAKXPANqy
DuV6QOBUVr0i1IO2sQmYMLZOhPXbmJMZtglx8OOx2TdZ3biAvHKtkcLOb9TptqFizXoHITF6A0aR
hWwQsGveNImWvgsFswRhGyQhtGrRmiGuzTDAb+CBVL4mr5ezo+Y/gLlNFEZrnpPu7NGe/Ue8nvLB
6ck9xF/4lzjjfopt+bIKjqo89sZpdlKLFg2JwHf3wcQfKyhnXfd9539wikT4SzOOkjE4CG02dh6B
AK1yFHFPWjKar8+kkzc7MFGgLHZ36pnKsTgcIB1y6vws8+NYwu5a9B/6cJWg0JWjMz8FGxoumdfL
Qj9TrE0J6Kv1uP2rU4rQOcXorvXY0dw9jvLs/xLicIF1ZCWGmzcTpun9N+nMDUMup8hvjnVFPjJ4
UJYLoJ/5azE+D4CP5CCToBJLigU+rh9FWO4QRI//Mo4/0ZazdnK9sacJI3qzp2bqvlJN3K0uujd6
ure3nsVT3oUWFjVOAX2B0+qA+RUjbvgOO/cyEoFOaGMfvz+j+zhtguSpszMX70JIbfbp5i0hSrTz
QHEptwXlZId3ng9A9IP9av4zJ9aOddPYDR2RXCatNfo+efAD0AwdIbGdYJze2f5/DazZLxOs57ZC
oRFgpzbvYtEPE5ulSkGH8hP9RT1cZH7avp0lVncpkx905OK6268YMuZYpvIb40SXLCD3C53/pv0P
icVCKj/7orG2/pGjPY0M8kAfWeZJLUm55uVLqGPaNoxiTXd/DvuK5iD2amZHs/dp30pRdDRBLkwV
BbHrXok2JX9dLN+MNxl3+2/UHbcblBRN/UV+6FgTMCARgqU/F0dOFDDe3kRPwajmcVxcuM+Dx/y5
25qa6ZPmILNUFamDP8g28b19pUz6TOl9FEY7/WB3CtK8cFWnb5O5BREu1xSLqy+FVhV9+B9/AEeL
ts9W3Pr7WRB1uPDdZ80D9IgsJmmFw5OvL5S3aBzEUi5daGJ1dmqMritb8JwG+9NMZzNOPABAwiFy
EK5Q2hVi8PCfMYr8IT2MaRja8k75SCab9zPbAI9abUoEUjQ7Zf8pIROnmgxH6Qi9KAinha4i7fDf
S/30IrZGiaAzOYoYm8bsvsDnqaCnlAeViuUF8SjLbo8JSduZuIv6RTKQy1p18LnVGQ/s56O0r8SW
LC3rVafO4E8f1S3vgo8ONfXLyEXICNDb1BNXcoWgMjA2j41nr6QUxKp9NzF2pMr5lsOajFT1LfyD
561kSU/8Hr/0NqHdJPBnfNRy1TKYLoKPbmEA57t10xPtdydHLBdGC2e6qmXdZZXbuJdNyDxT4rVq
XUEWomRONAj6FZDhsVOoHvLg8q39f+dWF6xHRAlPgXvDEZawhMdAhN89Tq4FzRdStjpSyjCHRboj
RlEpqfQWZnkfPuS33FgIAdyvxz1Tj3QfQVwQ5utolX1h31k+uvyJ5CNE5FFlAsiEPRNbtuqUvdFC
HcnIuIEghv4yWKbY5L8u2JeUdwTxvg/yrsF68PUjlC1E6NbGVwjLbUoGjGpie8MSWMyaCl70oqeS
WVGxInDqEB0ex8IPMWZU6dHkVGMMV3D5qC+fkfFuD5s8hoetEUVfGEXJ5wQ7Y9oQLFXNkzSfRqNE
HGgfqIqrr/6kFcA60Qgyhqp/2P0546BQQY+NjUopioF5v4mOQWbP/4bcCdw8UXxz5yTvhalKWMOS
CwoQUDVgoRvFF731uPxvTO0RH4aM0+flJCVvlelTicUBog7M1NZdWRVlGv3jFx1yUY412VqVlFCL
Q27dtRQws3mI6oroVmD4efVXrUxt94vCV8UP97duyJGalHV/NyBNSsEL0sEPH72/7Ursse8Ed1JI
phcU0LK4n5H7G9VsRXnKf46UnX9P0T3UMtp3spJHuiwwo+10Wg2Z/Bbxex4tpPguofoZVVJKTvVp
VSXYk6JaDPz5N0AR6EfS44YUHHVQTyBt1/210C0rDbYWI2PeF8C2ishqwX5Wru+YAmtDRQvonJ03
DFB0nfqFUbnoNhGG9tBJz01kk5vbXiC8yRSK2Vt9QJRDFydnu4wN8lUorDqVhuFVOR2RXiZHNPT5
xyP2mXcRW1GEQT/tMB6AxyDxmaeCvEpJnErT0utlRsUR/q+f1YtG03NWrvN8P/DhVH98/17BmoQ5
+J2k7EsyfB1FH/x69MB8GhrmuVp0wNkbjeHOisQWBNCYPndsPH8iiZt//cTUuwPfKWfGSTo7i4IJ
q4uFJdJCmnR25uwzHEvHV8d0dBeHWm1xvpeuWhPbCdB5xU+jrpOpvYulYMRcMWfodguWAIcCllIj
k7DVjKHiwXUCodwNnMkc5cNj6R5qq9IbvhcSAZd6p/Sro6QrTaMGgo3XklPusJ4qAts/YeMZKgeq
ZyOVRXs3fmtdMJKuodNr+YwHNE52Sl8dDSRxhZbDICyEiqnCLL7rJzWN+cCTvg7aXcuHZuftwwIq
zUgRe+RCvhhmX4+/jRMOCKTq36D0sBwNSvlf8lhXGKqgThGvpqRw5ktQ7sTjCtRvIl9fmwDfSMO4
zBph5u56QgvD4tkfpWtQjcsnUEPqH0sttrh97pZa+Q6X2tkOa4hUj/SNo6/jS0yitiJ/E1D/MfoQ
JOrhYP4+PdDgvKwDwsoVdjr1FPrgMYwZQult+w7y0UEiFN5PHc3YNKINoWkc8bPzLp6d1A1bqI5t
VgXxrSUF34VmiOOapGaH+b/NhshirKgadS1WBlJBpmVAEso2PXPo/F8qgM1Hz7vkzRWnobXxNZRG
x8Y8FTHMFWqrRMMkrXnDWHpfrYl9U58LK5bHA5eohPPOQp9AgeIDXtyZ73nH7A52ieoKRuBlTymd
aaFQjTG7uHshNYWDNWy6vAtHjWnnzYCh95jCxgE2fz8TaP8vlikv9QaCJzn9EPboyvLvsrJo9ato
r9piFi3cKKnMIYVKyxEfs4mZCg351DM98eFf3/RfCfvNKln9nZxsuNLHzOZ6h8c8FExx4q/hC0IT
+suN+38DzuxICraNGyaostlowuTDBxdM6DSE6hwpBVHyuKLb5udzm5HHvd1SMtaLL67AcYiklzI1
6cJiSOiCuYz7AJ8zJDw8Ka9JEiGFrKTi9YKORhOswTn4ubh3YKFBQOQn/3AVfph83NXcLm1AwKzP
OcHS7hWrbncyBP8oW4P9bDO3l8nWoDMqANZT3dqzZIJ+/63yF1ssGbVNKDDu1/RveNVK0ZNO/AWE
iHWeWVHWhaNLT11WY6Fs+Wx3J8MhPx5NUYtbu1ITEIkiMvcO2aOwg8MJLgN3hieklQEze/IfJQA6
y5EduPdO43V4lXzeJ03tD345kLzy31qnJBU4oHBfvoiWMppVLzVkuJECiOEcoFJe1i0tqLSZwmzh
f4thB04p1nJNZvS61/aa/yeSoLU7edjDzeNAEwwG8aVe2wFaJjEPuJfMwG28B1Q/zOySMVXHTLL2
kEJMiBiRqgoYL2PsrIROL/+9pwHMDsd46UUfoZuhoE0Fxv9LNywrA/vdrnWmGP4k1mhYhUI4fc2x
kr1tz4lYLqKCLRxwrZvWllznYCt7hBte6g/JT7IyxE2L4KPnVW+a++GTi+OCiK7ewcvOSSjGXk4a
JYntekxqHOWsuWgeHaZxH64q6LbU7livTcHG6wIldo4vGGtmFRkKzgKUtjsygyvG6phzumy76FNo
K+IO0omxhDWg1kcSJyq39jfo2Dbib90aHDkSnjwyBF7AR9pTPEDhodb+W9KvOUlQiBUonomjYDpN
bV3R3rpfTIGsFuNLcTtmbCXr70B18nLYIVeCqGViBqQ+rKiaA7H/LquglBVgbemaOO0xyvT/d75V
j1Tozxf0qTNJiHnHV4GSJAxAL7YxxFvzYCBPr3NdvFrnBDpiweKYsSXQTbc1xjmhmEeY1wqR9HKg
TMWClQpRNFo7wXjtRVlcS3Pki1YwTaVH/DYG12jwt0w1dd+p5aAtNDppVh5gUtc3bj/rICtj3N4y
7ofVK66myCjwhylilES/ldX+6XcsGhpTc4fbvNFqe6e8BAxLekcHUag2EiczvK5IVquRzYC6JTxt
McpoBOZwnot2nR7KvvFYgZbmXtptwNcD9ATBjsSDcIZ+S6lFxLzbtKgQxdzh7YXs5BZdZMlzN3vo
G1F/mrl1hkQCXMeV4wcdoK9OK5FPN3kA1E3L0qB2/s/OcYdLi5VzN6+PiqhG4v/rU73HLaEryHez
scYqxoPMONI0pnOYhPyxHrfrRTrn0323MSw4iBt7Sakrlgxw6nsGxRzUaMoXHoNwJVPix513vWzJ
jPbCvrfIcGf50BcS70h+Wy2xp00xMANP6NcLy6iSeZVMWc4OgfhZBNXGhC6UuPpJ5iZ0b6fwlwgp
AkFeDMwsQhBx4seyIU6GXuFdEV9KO0Aoq73HI78dHJA40ucTeJE1XNciK3FMxQJieKRIuJfr/d49
sP00oHON7X20kB0fM9ZrOWTQde/1ktFk1y1kQWOlpWunSlwBUokOZ/72KlOuPlHsaGkmHLGmbhfi
AZJ1Pw3UkzebiqCv6QcMrNV2NZB9ZqY96sJLM+ofkQ6oXNW+QcwB6HcRNlX+WynVcRBDKjWQqa3o
+YrSQJ5jUkx06DPDKVGfH7A3O3vqNpKfcN31u1awuSMZLVI3jzs0WUVTGKaCIU7hKIPlHFbErNBx
NvD8UywvNSkNoICuw545MhshF8CuumMiBoWELi9pMIT+pNSh2HOvNo8GGu5aXtfKiECh7wY6RrQi
vikV+scbuR84yE+u7wGyPOlqpfi0djbVcqUMI55AOEhFG2CF8iuInRW9ekdQIx+6ve+49PD1nmWB
SynJ51oj6UqeJ/TvYl8TWy+n9vlwI6kiuJnEJd3DStDMLtDwLcA5cJM19obLL7MitpYICUoMVCFx
mzVdEPH6AtgOSPIY+AsqDB6GLFQwB658T4YTJshkXh/e92xLO2xOKOUL17gSuRe5q5x7eBDsaLol
OtDjiKZeJJ/a5oy9DCE1H9YmRjDr8/VdoUdFxfyDi35KBGujJ9lFalXF5FXLGp3+kUpifDd3Q8j/
RA7AFg4CHAD8avHMLKNclrj9RMkU5kysxhjZ0c8c85k7rUY0/bR+pcB00krJa20fLajulxDoiuI/
XMDTAR/7A8EEaLSZsMy73cgj9+aKagA7C+qsYN5shqo5eE4yCQiBNtcjVM0jGw+nvApUZsDtJLQk
5ZMj01uVnUkNnrAzhTXjnVuK54rQDCu2qD4oekCIfvwk7+zWK3UCAalUuT1hYUr7Q2mnv53k7OQI
7Zf/SF5uZGArLKqhUIEQumITrYIfdOXh223Lds0xogY5YCXDG2WFL6jTrX3YwPBa4jlNj6rXlAiC
m9Qb7OnHyK/t8t5Udnt9HuiD3NmVucM6pKnGENyWxCP80LFvAEE8ny+8yw91b4Mfyvw9+7WhQmBL
TUNQhiBzXizmaAztc6ebV54KQd5VM9JIjxdAHdGy+sKyXHbV4BaAGmK7bxlnQZ2eEQElvQYUNCiH
B0AX922/4U6tsKjTkbumRXC4a47T7sFO1B/5i/aC2QLWMZB8gsyR0drenpS5epniYt31k1TsxX3M
6tzZqDrjlO3H5XS3WnU6/VKeEkKVFIBN39Vtq//s2UqUrm0Ru+gXRh/WOVQ5pgK2rSAxejsJh4CU
Wjse+kACnMB8IIkU+vRl+gP7DFmRFIaoAMsU6acWeSvkJU3JZdrnteqFnWQyRlZJS+ficHltcgRn
EuKHyvo6Jb+KHdZM34z/8IuT4os3+HHXfogkYLlK9f/3S+6y+GXhmwWCedZ3nMqLzZB0nPkAafEP
gBJxGLUe8RQttU5wXvKxIdWRfxZ+jCi1CWSvSdApchGRTOaEnxdJ6/c1WhBuHHzf03JZNeEsiClN
+5fJ/xNXeKE0idk5OXCVDuvgnkBfEwzsJV89sE+YTuMPjxfgZteYLDNckUD/4TL9CFgvK00E8UoN
ACusEvAVvq5DcP0JGqrBYtFq8LSZZ3irQaSRQV18g02jvTnTWSag2FG+bLrGWNLCSynRx/aAb6AG
Kbj1WlMIF99FJQtnyR4XifUJjwKBE8lhxejDt6OGAUvAF8X/z3o50Eqll6ZhN0QEEWwL64FLt0pO
ZSDBWPGSfbjtDfTNpweUUPXsNw/OPX0x2OoNI0TulXi7XsHlNctHNa6MIJYTjLZW6m9wZyPvV76V
Tkxw+bVoKm43hTJh0bp5ejSs67rhjg1KDFqInhvOn76DdUuMx8vWlXr26nb51b48jxEvk3ujRfhX
mAmoXZykro/qrE+HHqcjXSihiR2OpvvbNXPnyvFvUvdqtcwfdtS5rgt6Ze4hd0YRHzvyQwDzjxsM
8TWu50BEqMq9iVXz2aZsUpDfRkPOwYt47lPjcEhZO+uavXcDSMeE0JLYyKDu9/rC/0qN0d0k8ZJB
CJN1sBjEkkPVYahrnIqx0W4dxMSGNytFuUBObhp0djK3/DRVe29bFrnQI9w21pAO2GJkQF+YJGdt
PZ4GjPLfG6AVJ1uJAASkdYwyc9ECEQ/OABiAs0V1W24+zbukzkB3cp6Y4lFQ+1ibpf6TgPvwcjwU
l2klL7q53C/tTaC0Wpxq1jibz44Lg3wyWavYzPfE7bDM83aKc0XqDbzEb1UqbSZTX9+x7Fhb0AtI
exuZuv7C1/LLOZobtE25kqhFmuf0pVPNgJL6At0x+eyU5I9m7I2U6slwUD44td+/Q+WUiGI7sYm0
La+h/E7DOFWLBptablA1i8Nl/iKim4sSXpN43PDHqq4sbeFqEiGxZlqRzEtTTlGyQAXZ6x8QFyD2
DDcxm0eRim3UGEquOxJ2QSQ6LmOj+NlNgA3wijZp3eFDwgf4DOys1lLkwOJWSiH9HG65oYsoD+Vf
TiWhy8KlNMPvAgrBEcqtgJWpIl+UBDJW8vl3mKkkdmca3v4PMLWBLRxvfyNp/YBvqD35PSI9cysd
kNQu4OYCMbplPXi7zW6zHJqgedsUlbRQPq34hAF+pG4Xtwg/BfKzq5kjAGmNDnDPn5Md+CU8yp2C
gQhKTK+8Shx81iDPoUJZ7R3oWYHGGn1Ng+qPKgHAQgD0/MzY7GJE7jsWuLwzTqeZ7H4wH+Fyf6bk
EMSSwPeqj51eEDEAQZxvOB4sN4bR/IZZBpK5zG6POBwwmlNLrBmAMatlVVFFabNFx0Zrptmy1krD
4NkIc+R6a4E/liiboO+UmPs1k1BorttcJsVDI/a35nE+3bByA5Fv+Ho3gf5cJaV1ux/An/0vfvwG
1twJaGZRoUasmJcprpkmKAjMnwkpSM88F/ubRn/cWYlE6TuZ9MVB5LD8qDD9EqQNivFwEHMeATeZ
lMi8gTq+iXUwLFRPXBA/Kj3mR3XkOfJ4gSp9esB5n8WXNzbMBxP9b555mlBi/krRGttOiZ45uYVq
X1+pQS6hD1+8K85QTyH89wxT4YWXbBb5VejAeHtGdZihljoP/js7yFpKkB5hFy9UCc683YgPY8y7
IBQXM8XY3JboeUtuyZ3MzigEvqUqosIXy6GrCGHr1yQsjYYDLvfqmGAfjOjTcLeDmWg7iJqCaVSu
qQa2lqssDaKSMSf4AwBybYTmEEJnQZJIJL0ssW0UqcmUmcAjNUxXPCYcjzkwLJYjQfGHKKgg0gSt
YbLB8gQnGP+9ndkBVP3tZUBG2ZJSbqFTTBoDj9KWvEifSZSeQ95EzJYecUdYx+Ly500+wWQhA8lD
4Uo/sL9yGluShQsE7UXBaCQvQdqWEEL9m3Patu5ZSX+ABLVdzzXnnj8kAG+YIOt882YjbYw75iAJ
qXcll2wp2wUm4iiVM4BLkjWOW/Un/rP/xs4+Z824ziGyzYzSudB8Rn2jYMmov0O+vpv4L7whzTHe
oRJw+NVUNwlreDakXGqy5AIZhxiRlOsy7eIgwbPBk3LNU+ptz20DpPy4K29ClXC8y3tzK7MSRDSU
RlTuHt3nFHQhSFbOHB7V72DH7xLV/wFj9Y5tIqZHPHS0bzlX02vFTVz1SEP9EF3B1rcX4Piwd6HH
ld4pPxvqTuvG34Cb/5vm44/PMF+HhDSW7xnMqjZaACtSOWLE/sIKJji4oO6vIAfJp00xF2ZW+5qy
aA5eMVzb0LmutjINSRr58oTQ3KgqzMhIqeDx+SDsXSB66zQL0gkIh+8O4yN+8iOPjf1zqDKvCI9p
ywALcWdRQCF12denN4kcm1AoLPvcxtGF/e6RClS/X81AJ4i+CetqZtHcn2kk9JAsJg8HlJcIHMFz
aYowcR/RN+rs19Au3fGv4TlU8a6SElnvynikm4xpkeF8gs7OaQ2Dr8TwqvPQMb+9DgXHKr+Q0Z3k
7I+0wngPyeQcj7ptns32G6r7OZxo8YfbbPpkMLvHzYrpEviFMtO/yt/eZSt9WXvvo5T83iSvVHO+
uwgnFg0blhw8Cy+c7EfQItpc5BA14mhAsUbl1bQKhPMepJwByEl2fEIpW2yHrtcvbibcCxTmC4Jh
Pzp5mrDlwQRkIoVNf21SsPQlQ8W89+LW7gXVeDOEej/6Fyg1Yeme7Bg7qMBQY3KGGl2eOI01r6qD
H236F5KNfvt6Vi0oyWUyxqvqDqc4X9yZ0ZNpKUbBd0oUxSbZRdNw3ETVrkaIM47fWpFb/lEjsu02
nMBs10NvZUAFlZiiBVEQkNzxUBU22IYcgW5OjMER25SRYL8MLfhCG2C26+TbcHsIyvLKffnQTQx0
KTDvZRu90DuzDA4srubexg/W4WTyxsVBUYFZapXfbuziRhoQfBwjkpRemh9xXskIkz7Mowk42K38
chyUMlABC9kqD171x4nOVleyRv47R2YOavRqk2n1Qv8b2HFcJihuHgBPoe8/sO5X+ZuHXGlpjRtd
acDfhJojddOrJSmna4SimR/qo4Pfx0VaNwQwUHWWFmspZDbJxqXmbbtQm84Ei14o5S5lFrl1c8D/
QxHO+3JPk23jMsZMuGV65W1AbFazDvi8ud0VsXCu6mXQjx2TchyXoPq6bsk1Gaks8/IfZYavdS+M
oIJnX5Iv6NKevCst+gIDp29TRy3/eAzAW26hl1/NVTllKtMy8QlWBqH8puonVZ8ogLyli44ZSopl
gf+Xi2Yr9irBI1VraGRyNiVJ4/7rBzIQrphAYiLfB3iQN5JlY2xRApGsp3Kue6L7qxI5kdHuvodM
K6rgMe9AxO88EiAijLr/C7xqakMUMUSD/zpkApBjx/yYKZPe5M/qTHLK/mlWBnhGiKDworQDNrYD
/k533hhUKXCcEOeifpKckb1CoksTIQeQiuzyl+nWOfrUylo6UjKvZbntsNwSE+ais3v4+r2UVhxV
haPHYwzyT9qMy9P24ukvodnRiJDlfvgFVGdYKs3qMZC+ul1vvY6n5d+H3vyZ7F/6+f65vwhuSXBG
A8h7YDWwch5s8twDZv0Baao8NhFpF9Ki7lTrQQEA4lH0W1qhzVl5dwfwhKNv7zchlfidNx4b7Y8P
0EGJSq8i53chW1rb6f/yjsCv9qopiIZRhiNJOPnffyaH27uR8AnH/sPnGwpMfRUtp+RprR5/uEsQ
bo1xO9ih8r4UEVS3zbrf0SRsd3jMaWU5b9zv9oNMBwYgOWYQdO3b6+2i6LJldAqsXHyRQ+T3pGzq
iYIGJmOhBM/WFGu11d7HhsK/kn11XpGKFMDQamWGQzixZsOQ+JqiNJFFMdj7evjWUBUGImC4GeCu
nPxdrO8DzcrqvVgWJ+ZHbzlauqfG/lD0YCNKlnFPzLOZkt80NmYLWwjIVB6AhrwDkvgL5cjhd+S/
yyCy4UsSrH9GOEBMbbILmuyTzd6rkRaLPU4hNm4kQAZtyMkkFQrvpcteDgn3e5wcwB9mHhhIwUef
ygLRsJMQpNo/WAH1i2Ja0SK0IDpyJzVvm74dfYYzmppsTnnMK9l0YuwEI3FVPBY3cZ+cRZ9jsk/t
NOMhmtd+ni5+zjlLawv7kcDYsCNwsVz1VAvhnvXc+IfJRnyu4z9Jnr+2DHtFTzB5m5gAszfBifKh
a7p75jX9zYwIuJrI3YKuoAfU0vIGjv5B9rItCcXTJLc9G2znRCtPCPZm6mJeVcu1WncXzP/IkYuS
Xd5ZANQPGPbuwzAAg1mKtQwaSqrzpuX5XEAao5dDbWXYgQtf5pFaIc6dNbPerZf2EQA78pIO0pje
6Nd4C7RU8dhohA2QNctf6QT/Vwi6Y0g+1xvrPjyi/ApZiXDPbwhrNEBWoCa2InSlPWMsHdszmPt3
Ez3qmnZ7ZM8AgLL9cSQkSfIi1jHamGg5jH8WCLbrFwV7dX36zhSnG3oQ10+7xIFSTVEURN09Chsv
Eacu8Sgw5tCuaezFapzJktdxw4yfz0rgos/TckDEu0BURaIchsYlLsSjJKOqauimr+TTnaTPSGBV
RXw6i0GFIarVGyz7qp8VLTckbEPXd8yiyl99Z1SFrzz+TFoEx9SOr4+0iQSdhS7Zy2oudVa9YDsx
oxv2qtCtdbMuer7txc8lO/UhA3/v/MpMQakfPFWnhv3UpcpKqExVwyvjPjnSqQtikqeVUQ9nmM+n
ZzDz1EqzgbZvTfsTH4xi73EAvQWPXS/otvDYJR0Q7bTp9rsnGlQD88NBulUmf7jI0skiHPSKCHt7
BxneWOA/lQ/zODbo9ojWlxVQCmpMDDHIHaq2RTkgYZD8FSMCYZNjsmB0qjvJDZMKtEmRi+krOL/2
ZRdL3xJ9wozNJ7AE2zEU8OJdtzCFZa/6nWivy4rWYxLOqMLK6yKqUK0LgbrINh5/VsTypB6unuym
0362dqlesByW6pvrLXEos8aMz2gvCisG/BOKlXS9NcLDaUSAsSzOZYJgJ+lKUTD1QNc6zKWm38TM
cLIMQzBuvIHCgfWyMrbqUSaYPIC4qzNm29yQfkCMGB10SUSh1HAu1fuh2wh+qdj0/VmXyEFqYb/3
eCmMrfggnbzMQu/rw8YiOEkZ4Gldk6auM2bpGYDBAk/0oOATSIRdS6IUZb6NIt7oVU6Nxo/rVRh7
FWaqUYZBaOyQrQI5So04xrmCatbS0UGmCUatXutU5zqlLd5tR4B+VPjgcH47HSohIVaLEgpVjAZo
VEaUfbTLRKbKdDu/EySu4nGOy6W+zRsZ4x/u54ZXD6916rlkLMB7toulf5ZwekmT0qSfVgxBa1Bm
c96uNema8m8kwldQuY4iM4s8j39kSFMHTssEYUkL+1wvxUbrBUbpMWYHMpnZLkzrum8/NV3xQfqr
Th+Nv30vaMO7Wq7N2X7ITVU/gVjQpiGRNzOyz71sKciv/rZdTd/FaxyD7LXibnQGHtyUHzOa5r8H
FGe2JyEPl35KfX+hwNAIsKNZ73eVMFwYI9sWiCEsFLitIhyI/IPoAZFK0vsQW1zUiIIdBFFFYPGj
yYn0dX3tUbNMPAjrRSEQBiTVzQSJz2yKgP/azNl0fKkvwuCIhKLWZ01xwne6O577KyvvYA4MvHMo
QZktZzNRZclore24FqZJ6szR0CJW4UiVsJGO225OTgl/F3ZRC9NSjFI31ud5OEBEhXP3zsE6EBS/
YvTQJ5iKrdwtdnGnmU8hWW3D5Gj0TqsbrPQ2vDDHAog/vpsRyPuNLeLWtd55fWjV+D22zkNozpB4
y/VPlMb+yp84/UD6A8VUCPAXldFGJt2gqBGZ2sD0vf5jQu00seVh+cHUyc4+bz57XZi4i1UA6kEk
3XgsYDbe7VKCFl0G4SLza2CbLfyuoqdKYC4qMDe1HQsrd5SiFSQWxkIYCSH2qPvwCwQlQ5wBQbH9
lVtueCcA0CjmUrygx36dEYq+WdSa//Os8PNwqg3zsCaHlv4H6OYUKSRlx+XKmJHoCIs6jzIbOPEV
CfmKuGVgAVAKFz1m85qZsx+CZJa3nxsbvOm/70ybrxwOG24sxo13/rYhIM/eyb6zgdX4FkCF39eV
VhXmCYX6bXqpG29jWEt8DVK7hhyCIyBHUwqOi9echFOlkesOeJeABWhUqDNzx1938jhISJfJr8ui
Y0yq9LN8OsTOBfxXx0QmPFJkReT+1NQSus1CHD4rO9RmwLrlLwIXqajOFYdodohrGDYo+5Gz+Vkj
bJUZf647RAN2/xYhFQTK1IqdlzhddIcIrjt9H0vB1cFW0zHMyUOPB3qfzAPC3AcxHSlNe5PRDUvr
YVTF1utvmgOOc6GfbIWy1iM6xHk/Na8DgVm/h80NtgV6y98Sm+NCibR35au15dY73paN7oox+qiQ
HxkWAxxT4C4vTX9WcIcxppWS7sp1egHTfD/peuMcc8WVmHuuOTSeeok4fl6Wg+rx/SntoyPTExeR
X2Q6a8iTAFl5j4Ip3hGah9r/if04NR+j4W8BBoVwirZpfEU1PUwysX2z95oWZ7/gUpa8N8E34CWN
iyyRG0tHB5nDl+iVFhubYx1dBZjWues6l8FDd+kwWdUSTsBwVEMHoqYY5Am912cib1UvCdJ5otAa
gXxqHWlIjssAt7C3uPZbEuj7QZhRDjEB27ciyJRrbf93OTGOvTvFUBE9XeLEpi+jZXQyfTAUFHYZ
wKrgy8Ja1zdzhh07HM7eXUGnm/hq7aouodRqCZvpa9OADFDLbupFJX/FPX3W/y0pLRKf7eS1HzT2
RCHNaRQh6qMp22CkANZDDxbc0zfrcwTklC61rO9+e8ShWi5OmITXP6k95MpLKpfhOAr34dGb+lHe
8DYwBR1fKGeNpIbjK3YQ4BTFLhJT5CmmgN5qv+yNKIm7tK/6nePm3d0CL72RewNeOQuPPChU4ipA
1W+W2DCSgspN2t37D3SQ3THwh4oPo1GK0GbjYyH0Q641b6t/Ogwbj269ica3diMbL4lzecyLJcOL
vg/Rm4It7mghPcmUlLQTimh2J8yhROldl0BGD3aHkau2tVqWcHX0H/LF2OKGnAEHZexBNtqUBPhe
pCBCKU3dPO27Ex2WB7kt2w0drtsgRIBfRMkqYjBQF090H92b7279nIiQj9BkMPMTNV4AZ7DeNha9
Bsrua2HFa1PzshJhDw7kE+kswoFRxc6xuymlN3YD0flV5lkmzZGVFnspUtNgKSdzZURqFXjTAcon
wzHrgu4/hv9X/IV9YAPfK1mx5XL6wV+A36io71XAi6Xht9NmEsjwV5+kzGaFt00FxhRp/Tq2lx+r
eKVllvlUBKs8PoXqEt2o/ssORBOl4weeiWj1e5Y0nulTmvGi28riZQpcdPVbnjySFmnEtshJhqY6
k76vjJeYmlG0at1mrN9k6cVGsjzss3SohOeWnEF5c2wiSTgdxDEV9grvfNonrTNIZ2Aero2rxx7z
3P2xhzVazD5zzOm1y0J/h9UicUCurVFCRSTwpx8DwBAj0EUCPR9I4u/CXU27LUzXQr3ZErayCUy8
Jrsrc+J2Rmo/DRROmwrm0aC18x9GXtx7x2qCvfkOW+Of+2WfjZNlxuyvpdInXGEGL2jx69Viy2P8
m1H4+2TCrTom0C8zEX1wHP/7CJQpRJ7QGWIugRBtlJdxAec2BxaeYQdtMTRxUpIRK7rkN2H9PJao
fTvV15NxzaTJhpobtAMyFM6mCpqY3dqy84cChwmuoArQwqoDDqT5vGJLSyfeYOwF07MLUvGahYCL
DeQR9nfAGAJ2xtWciqY30PqWYYOjILzAISoCo7vlEXicpR5tc8L/3rYS+pxQG2wB0Y6m85j5DozD
gWNEnWH6Kv4lwTaJywTmDm946BV0nkxYSpZbLJiDRkLN0i+YS4zBV3bb+u61bn4LW2GKcOms/9No
Pfaptknny/pLmT+9jcpK1eCIrgIsqu1/zHz+CfNswi87jA2FsQDyDamimJf7fezPF5M8tUr+LTdg
EJiKjkO/9wOGNNlTuYyxoiDalxHgKL2719qB+5VFtG/YhiXLOzP26//lck8LZJAxg9rav2OsgjMZ
QgLdq6EqMAdJGTSPBGg2nNETXcKb7mDf6+7NZMlcF6kbglJR1jIopiCFcNrO6rORbKSxnjug7iQQ
ZvUoJ0JY0gxcevOyb9my2toSx43bQ73sgkh0ZGTH339xuLC2bBYMmSIBDWjc/9JyYJoAP0pTk5Oh
+yBOycPUmjlK0W2UtiP2u8iScSanhlMnTaLWVgWVZl8idQ9RwNa1awTD4NP2IAqfGvgcQEzjDzn3
DcI+fiwRD7di3jdyQXMlqAVvRcGLt7zWrzmM3hnuCHomMfOY9TUCDzugf15waW94cibh/Rk8hFbK
9eoWYqEgdQIIe14nL0N9Gx9A2hlShN6Pzrs3amBOQJFANtGAYAVTYchZUUM5gDiFFYpZrntEnMTA
Se2ebmsE0pOMXqEbjSU+kN7d7Oz9HhQnD8dhMMRObBMnvz0Ih8Kbo7RP8JA2h/K9w74sPOW/t42H
65Bp2lhWz84yqhLu0bdiblhFjHPp0a6a2J8mccHMXArthnwiMF4gk6MRvTYYET0ZIJm0UHvu/D4R
xVoSuAhrECABP+13FzVqV+cPlavBPwA2aKpdeReQFVcP57FFj2rNxwMGQFFNtH59PPDaRpVLTtdL
mlVuSjOqDFTeVYOFg2g7hkE03tXwBVG0dIki8GJjfDKzZYFeBfFaPMUbLuIG8YAPUhyX3ZHUm9/K
+43e0XHboTnfsKa9U5iWpIueph0f/f94oMwgsFGuo3w2I7Nm0a6Sb0Qr3AVv+vmR+kaZ6b3nWZ0e
ba+Z04L5WKhHBGl9q/KULYgGV05nd3mvp7DvQqCxDg6Kt0JXF+U3LaESj8589A6UK7lIcFYl1ao4
H9/X6ixWMeawvtDd2hynkrwJ2rtTNMrMOfYnETJYoOKw7Oh7jx9IfGQ7Dl4N1bmBMkW82SqNHloV
oyGwh9I3wbWGNyguHaBVfjKenjbHIlv8uO0QGBGfDmwaI7N1AdnUVC/2LqOdj0bwc4yi2IsipzSA
GizNgtG+lgvvS0w2ERi0L93yh9sjp6/NMFkX8VGdO11e+Qp0oS5ndp00RjeJgZey5rxMxqEpUEGW
ndNO2sXCD0W9IaTCEw7a07kwpJXjbRLfDEKxMrMRoY0NfmHxBqq7++bPvvoDaEbYReOpzYSGL/N8
7e+Gfg+3FW8p0gHO5OIKe/YvjnEQmHYIWUfJrlbkjs23Hu1KvW99Au2JWNutTumODPl6r3S/P8uu
Jdwnd/ELB/mLMidP3a1VaT8KR9YGm8h9lmg5Nx5ldGWcN7teljlp8keu1VZq+Jx13MrHsKP74cZh
Mj4ma8uMGCPF0X0wtkeP7NUGV+efpP9Oem9TKDj2yujt31IXLyG5qL6FNCLtlgxybapSskGst98T
FkiSDQwdU93hZAn91WRpC110pXb5JsIgX42iQGR+rtMXDV7gGoN/NlFBuvlGQitqo6fHvRXEluxS
CjdElE1QqrRKJmslXL0HMw7Op0cY7UCyKxy5l26qMyzbfQpht+xC8JogNRaM3XyKUfw5KwrsqFOY
WGFENDJEw6Zjw7Fstmp1prwj27WlixNnvAmihgPC2NZlrVS6ixjIK9TeWBYZyIXNmRI6I1SwEgo1
k1mh4DBcCFG9FmjOOnKDI7kE3Lc1thXc4MEgwq++/TX9mVA0COpg4792uyTCnSBav1oPLmNcsgpv
Uph4GNBaSPmX6P/acpf0Xue8M4Kq+Zh6eOx03E04c+UYC2d1bxgGqAsS6ANFcMWl9vMM6RzXWC92
deu30BjbTEYj7m2CalKv3DkQGhUFjTmLaYfjY5x/D94EKSVLZHAp9/qnhobPGC35HOi+ouyTKuKy
Zqlk8Wv1E2yhGKEIbYPyoFYH8YClC4dieR43SeyoLhhVdrNfGMzUwWNPfnQFT+9CC4/22i2BSoho
jhADDEVo8UiRFWGNVeNesmAaA1wkO3EkKWmNoDDCUCTMOD8NUAAmqUhVFYRcMIztJUnErjE21u2F
CB/z2U0v+qM+VvcEwXCJIx1bhRpjiFiz4zE4936tHdno/xmzT8AK3Qwo3f09HZFQHj1u88rX0H5b
B0IqNc8UOvN28hsDJPsyBduUiH++a4criRQZT6XCkNy5ENVRIu5g7dyYNiAS0s/pEL4PEzFlOqo2
3HFEXSkVgX/vALeLrXMRq4GSYeScluKYv8nkOqtfunI8mnIvcKEsEI6wgEj+yFFB6cPwTpjE/8cU
uuyfwViKnWcA6+6Eprt13NgQLw3gb0Ni3Je2g2Fpb8bBEzaK/lKYleIURZrQPNvQFy3A4OOAPLb+
TvdfV/f6TmJP/gN/DfLwzjGvqcAhUhOuW4GVNDRA7oi+kizZEuXvtI0WblSCqFiQJPVGo7pLb2yW
BAZF6aQv+tu1FxhbGkerfZULuWCtbCezpYRSmLPmxPizSdvRisANELClOkLuA1Pn2XEdseM7R8IP
03KCv+eLo9LxEGywIyCgGlN+xxTyFLFT4s7TiqQIgw5t8F7SJKkE/L46cm6HRgcxM7VoHge2x8iB
O6NkJk5BjgpKKeMTLyCrceTHM1a8ywjo/t1h9FCJL/d53JIedU3V0+CGBCYN/YzWsupDwsJCGE4k
B2ISKITSzuvCpbtwVrdAJ3kzpJSuP8LNl9HfQm8LnNLUyjJg8zWucQn7o1Ki/tiE9EiZmSv6SRQh
K+f1DH1YW9E+m9LJmLNWNBdh6Qr6Ty47ebCerYUHnnhSuOSXslWev+vG9g9BQN5TxUN0HLeSDImU
Ke8w9beoX6Ba4eYKOY5zuuMy2RdNBJVkI5aXyp/3GZpbDH44izcydH8l4jAKDgLO7kZ+MwHkupAR
ivj2wv86Tq4egULbobEnd3MpPQaKea06FdApoaTGbDVp9nm+MRXMBHsOLBA8Bx7MRc5vwbmHygjp
b7moWmG8uRvvI89ECh4zX4k8jbPfOGNEambmC2ZTsDv33xp0MGBpqiWjQuKXxiShqME3jlzLNddz
j1ADpdgFHHU1Iba1QuOE0TTTmMSy0huYCzNnhHuVHwPp4by+CVRbodFajrvRVguyde17wXVp2bLO
UvpHdqSpNZHXYwtbc/ddKer7DELJEmOdcab0R3lKeDd/DGgHh2ZgEWIM9TIRTcqtbGwofxBnyPOo
/eDeOszbl1IxLJ2Il15uv9dY9NPUbSx6M9Sb9pNGdCJrfdmwIGyWafurbl9dI6bT9OqEGiuyRZ1W
rNYXPz3GPw49XBGvUg033ozP3ycapdztX0H0ZgoRlRYVKN6RHZKfhj6HIpST1HefhtnAs3MvlEar
F8tkRZdyAztXLKzI6w6+0EWT5705Oe0rloB7+S8FwUDVnpxUj4FR5Godc4Cmpptfynqmji/wROkI
Erq2ibTl6/gMPv/jLJ3clZ1jq8zwa481IMrNtfuYNvOtDsAVOsIyqbhVhJL4tc5tzAPchUWZwt8r
aeQaBUiJ8ucWvbTGyCE/3SpYMrjPfPCQkyVgpzyQJujy/zHIzzY1QDJ5oNb8gBQJYNKY3PvXK//G
Vsc/yOTnbgyBq/jTyfxuKrpoBMWaqYch+gIFvOYdn0ldtbKprQYigeqT9lpn6MTjh6M7rvAPt5dR
I2o55hF1wLhCi/p0r/0+jYNN2kKZMBblAF3wZ2Ns1kwz22XNpsGER1YT0qFWlmWbgFBqXiz75W/q
YuPLrzqQmoOu0+pif7KDN1mDfW460jrXQdf/K71dnhKyKTWeqDwtGGuv6sdjwGFbQh+vHELqJYNs
7LTty2f/88cA1wdrnuTpwkM48qWV7mM2q/79FAzekEDY9uOo6bAonfTa/uxnX9wAwcvqrytzIH5H
mInGyxtyzpiywmWL+ToH8CP5YyWLNlF9YhKXJC0KrErhNRuUs9yD+3/aqShhGTeEY2nr+j4r5j4g
mo3DjIym3RJ/fyBOoR2rYHnFi2/xo3daQVpjnnnWvzceuNMWxFKI/HOSdJ5TZDhff9fWx1uOq1Me
BDWHxD8g789P96Vc5UE3kyyrgqUJX/gyCnE8/2Epgk+aA9itoNhXL/LFUA/90RCZodZbhZzVtewq
m7BcixDJdJq28/ihoWC66GiwSxh9sJbFtSqFRpTVUhvsXwsvx2K01PAMGACj089lNkIWr/VzRmBD
on3PKMMldQOW1MeN+syU/8Fj3rMPRPFRR12HJul9tPstxQR46m9w0I7ioU/njZqyxVwwPqUAkp9i
vo0T5gKLtKKj9zzdgAhG5iruMGckrpUVZmU5zDb1acRk9+NsiKQfCL0F9kNKP48tO9BG9PAyW4wx
N9G+pB8vapyN6qQkoD0DriC98rr5ct6ozxsMOWSxZrnF2RMyKRXVdUO/3aAbziF7FRJ+x+qEPryo
CpxEWkAujFWzJL5n6KmExlcFdy5fuAmFoLxmAHItEIjqAx8ewRoRTuG4SIBgujXbq55aG6X/lB+N
khS7nI8Vw7INBLzW1AKojaRtpnXd5LeT0MN+AM2IINRPLMMYbUjWJR4RiV+PbqOfzukKHETuJF9m
zKE6nRcozzT3wXl1QMy7dkOhyexKmJNy39ZLvgMSxWh0MK8HhlMJC+Jrgc38/10ungkA3Drd8cBP
xsl/BD7RJ2uW4Sqdhc0cOxvnKeZgSt+tnfHtx7cfcB15TQnf4ht7hwT3ytgnuEAZkjJdQlzxaZBm
moLXdHjAYrzZhj6C/iTVeVDzWrqDlfCLG9v8QDjO6rkOJ4Vo/WNHWPPi+3MHqNCnGnxPwwcKh8j2
9YXGTNSB1Aj1PUSx3Tc2U/E+f6/B/10XjzwmRIRiGQlvJ2WqKn7Q5CQpDMU+jG1st0x5LaIeUj3I
zOzFq6KtXbybHMtyr1DblRIe3odx/bWeJ8fDRQEYHO7A8BvYqcCDDzUpjNSCdennHw1eT9zBdQmo
WMFonVim/62iyewHcDFUUratUKRYmmPkvBnRQX9+DLymZRkuuIJiPFh0nCMR9lrNtg93AIvZHo93
DgSvJiJGVQ5sxySLlvARfbc6ha4+GmGz01SMS6h0xSGAYVLSP7NFdgUd5Dnf/B241thGGKkX6shD
8hRu4C1k9Mt2fai3gNIXrJYbL26PUNzGx8txcl6sU5mgX7QORvYYAC+IGwTYR9REilqMhTSChTNf
Qz0hTH/YbQgQkhARHjoVvXCcToyEoJsBM2k0SFkaUEdwxOL/GESrHkSn4mhxY88qyCoE/7BhcSNl
OEiJ8G+wfFMPtMvNC4CxHSv4Aaf7EkA6nl5jXYSFwH0t3FTcwdW3Sh6w9h1BGgmh9fHrSsEwyEN/
bXCCamnAxQoMWiUAWWdrPtiN3i1Z9ct59Ro5UFNS/gXoCX6SJWBftWMVDGfuqNJ2FrWiKOllqT+o
gQf8EPuWpB++plwR9jKb/ZlWMUW8KDwkhmX7vvGsDl9gTyLEzUUbGygFuGon3OBTCsG1i8cMuS1f
3dtO8cmpY5ycwNzC6QtoDixgnKCdePEW49N/D4AacpK0bNQ0ytfKO68I6Mz/oFFmV/nP/cYuEEs8
ZHWihIT4kuwiaVFUv7RXoerStzY+kO9ghTpj8PnPFBVN8SCjMnwweJh9KcW/NRdh86RErRt4/WDE
pmqV8gpvKkw/D4wO7wEpHtLbBDljhMcBBJ7KpZlBluv6w8UPNbK9ZBsqY5mWSapWJMIKF2cKX+yv
8Y0/mEJ3Fe8TxXC0xHA2/eP4JKNkXJWwtUxX8CX9/rCg56CYY93UcGFJYqtpM8u0yqONxJsGH226
3pbmUzxPu93VfGiDAksKFHnmrydA9tniGIO5cZ0RTYa5xPUAnhEkkB5sRrKfMoufcGKqeazsrtDS
S/3fLs0Jw0NMxTzxI3IjBqj3evxzE/OK/lWH/FJQIIv4VTL4CVW4rQ1m5KwOmEGMY0s9iFFqBxmm
4JgJ1Jt2fXe7EHXUo041WGGeKnxOATlajSTX+brXetajqkUwkOsLX1hGi9wF7YJtUs/I2D0mxaG7
KW/2RNbMI+bZhu6KumRrKIW0bP383zlEb2zjJIRe0j4VHTcpsLV9LZnlZY/SQU6g93aFlxrsO/ZQ
bOuTCl5XcgtDtnoEj4SyXIucL2UKEuTC0iHwzqwAa/QkCq/fzIgjQJE28rDGTCOawhJVxNdQZvgu
K1xaCUyEricqAFuwoIQO5zM45PUsYJFKnHg77xxeHjzI+8qQyrUAhzlmB9ylrO1CxRhlZXKmR1JJ
XatVsxKhxx6rlh7i4YGTq/iOpN06vb2IW57oOvt+NEnfwVKoH/90+u38dMEETDDWTlbtNCPzNGCk
4QbWdNCUY9cnCvNpTrmzdVCjI5uzXWgdQM6QgBZe2RhRvZJOtBZ0W33pK/potImQWeLrjRexvS0S
1JiGMJUT77oXDygx9YWsP3DRbylWNvmdct+/Y701Vk7WyuBynTsyKO0flWj92waV1EKgCkC9Ztv6
ovl55t/bWTPx/wVHm+65sDjRDOP07l7AvQj2G+Bx+3L4EM1ilwNoaNYn3ODE7Vezf9VgTMIEeJzv
PXaDUp1Hh8nglTa6cyeQjseUavfdwCAXB/CNx5v+xp6DQpbCHouQz3vTHkTvMO10dJ8YWYNhjgmx
72rUuwXJwCC54x6odonj6TMKDBIBhF2vQpM5ASLspSp9zq8FDqNRiKk4TY7XO5Nh5syPBpJ0S629
64hulGjK3CTo65Lu3jfoK9nPemGhGVidO/FymAyA9VZyC8eckjsw6nBftzLD9MMg8qRM1QZDMUWE
G9ZQku2NZjEjZjxViev4mBNFrTB5Y2rvCMwLolMBpXNXottF6zbjCUJiWFk7i0x3xvqjB9I1G1Pr
ZgQZ3Nois9xQIevk9B406wakn0HkMYVDw7AL/A8LkzSoRN9qrWt3kT1FTz7GMRNFTMcmhnnoshs+
GvOYmtV8y8gJLgkr823SH5aqlfS1JHOw8dIFpTgIyD1zESzA6veaCMnBvy3Jg/pXauSFHdmUpz8X
WBVrkwcaRq5doxDuZurAiuvFCWSREaJrWCY6N7KX35SWOlbmOBrtRG26+0X/x4ohWZsgm760rVDv
DiejM2GctiRKahW8heK6yq5+ZjRRedzCw3Ef5y7C4t6wFF4Tn9Dc1FvLkGG6zIAyZ83/J7rwinFH
lAB3aLoC6IPRgjUSLBtI34FyoOAlYkmOmdjIDLxac8ChACP9QEb1AAKSIaqPqmGYQ8O+IUYNbus3
DB7eeKPJgU2q9SdIfcuYNh+66kB7bCp6JbwqcVlLQgAoKKRDCIvPioEak/vYUIMffqtjxY0DVR9C
p1+NIFkhUpr7BSM5vqggUuOf7py2QZX6rS43QAnqxv7imkOt6pf8phLAumv8O70sG+EE1Qh+En7N
5lYJvyUMGbWnj+m77Wl5okIw96ipPzSe4jr+0EYIHj8dytnKRqWf5nbpdTsLNaac12Xh+iF9MW5h
vCHeaEmP0iML7mti9Fcp8SDWCEJRi4DlvxzJ07bQzb3GO09MNoCq4sGahfd90dLYXnQazWOKHkQM
XdtKFaxGGrlLdv8VzZfbZ+KnGePSJZPxW/6B+4Mzbf38M+hNyltMcOfbU0FIzbd4P8kePy2ATv3o
tfzQbSS5Msut0LwE0+qr+r2T7Flceea18bfATGRkW0wTKKDfmYZkCCi81eysCsFY4Q4Ebx/E2upk
zPUQUGwuttwvCQp8saVNoXJCg7Du/JnVeMqaLQjRXDtLNtJS4p9vESiKR0eRT3Vxk0LNZ/xbfcE/
9526EdzOINTU2EtPvrAjb12bX167F8kTTKyPFe4F+A5qZkKQsMHLkbRL552jaz4JK1rHca08ajVX
q23y8O/IJY5f/yGCoJOzeFkYGq9lbKLMDmtNtNgl2XtKhM4PZMZKsOYRdygsXwWmt0D1T08GskCW
MhJm8SosNltLihxe0lQ5fWwuTz9GREkgZ7oVpQpqGXezpi/9Y3l+/SwqvhIxFz1dtRe1KH7+WC3j
rYIN+nXykVzU1WsIv1YIwYDI0ntQ8IFBIVT8PFMGAR+G9SAZ6L2Z74XGu04tSJ9JhsxGj1udPIy/
fMTXXo0/qlcA13IkYsN1TmdHm5CwdsZvjzlqMKttcsHPLUP7XUf2H2nBzo8kq7DZ6OQvpNwlA8+4
Hkf9WPv40WxpBuFKa6vi1RSMlD8TOhWvXWQc9QmOViG3446UltEbGSNlhiqWChAjVDI5LVCXOR3w
lbUaG/17LwqNBMqSivdWreAQwnghX2Aq5n+o3UwI4G98epeTpwwBCITLToIRRdiHGdooonipMGLh
Q0aKLfePbQhFIKZUhkhYE/5/Y81aE+FSuK8lfXQbdAqBF2q8ZUt0lBZosV/J3LVvLE5keSy3lE84
QCqvTNzV1TbonyvdXkyzL0lKXvRp+uG5MXF61nPm0ig/W+woZ5NT6U9nw6bC68Tej7Uggp3yuyrK
1r8glYQa03utEmorJaefDB5CeR+pXTfA8L2rQXgSd016mUuOKOeaO3++Z4MIpGEEWYW6ng0lHNiG
D+hWPR1WGXjwvFv4knrrSoXGDoF9a8HVByXS2ygcrHKFYxA0i4GouZhoi9Gpx6WLFgdGCxfpyI/d
ToIecvTBbqBlazNdGUn9jp+ShDTdKKz37Pkox+SZQsiEMcB/yFuKBfYunXlxNdAd6pAfo0T+az5v
2V3LciGMRMNQG8PI9jAGztaJHy7T8liWo/uFpZBZVvx0pbabjvBDGtnI1+Dw39u1JWfRqxKz/rGo
ozkGWOxtDRVcRvNBmOatJc4EMkIXgOf1Eit2/pw+fFV1p1AsoJOIhwNDhNCEzuveurMozX676Yva
dkmRL24GG/CM8OMrwycUv25hzNpNCh7mRvpvcyQAvvSgA177XS11AJsBLGXQmeKA6IMYl4FAuOkF
VARC+glCRgMWEp+S4gcJkSGLu34nmIG5+8/IWLNs39vejmhPgBNCgl7o1LKXUoCDvJSs+4tl8wH0
bxdDx/bs9ZsDdahQ++nzksV9vDXfjEctHtzxYb5f48keCoqyFRUDFWgg4JGt6wq72jsIDICHi/WV
xrE8ZytzLyQyMGaSge9Tmk2XB9N7z5A1gMKYVC0Ixq4WLJCcjhSdySD1LQSkhYaoLg76AAG3w6xh
tcNoA3GfCVKExFLLRIoKjG1medAJJtneViVyVh9bnU9we0kPiiaqmCtOxMfUzVOaRiBvjHI1ZGdP
DmlzsU7OY5kcVrl9CXhtkRejyjCR9Qh0bJ3UmSdVMSWj+lqVgEWqk4isK5eQcVtVsDSG0Z/XguZ4
BGC9SkNMT+az24TBAKv9V8+GAewEbU5D91Yoiav3lTD8+appOUSQzEexswyK24A7wA8pf9R+PUYt
Grxwlg3BqoOKCrTGt+cZyjFNg9Aupcw1Emd4SzHFPrDmwgaMzVkOVcUCmGQdeCDweMf5nImYCLaW
YVRKpmR09wa4Cjlh/XZA2TZvGQl+bQEjluzZFhZ/3aGEjFsILJZbW3vyQbCLmPHeb6GjYXZqip2x
Qy9qwVLaK7E0OWvDjpKDtH8oZXp5nzMBHxSfUPh9LqjcSfA52+xjtg/8boV9riBNwi1jQMGSVBlk
afHTEgB+XReVhskStYg6kKE9mgQL8wiR5eb/ZlLpCsljlVoBjq+8lMti6UsOKkcGMLZcXfe/O6sk
Pmds/FrsJwKZOQH+LkaTqrpNXYgIbMVaSw96em/2a2AWcEoLKuecjkoaqsMtKCr4i315cq//uqXy
DLLfsYXcs5hG4tgfwB1y/HVxFwlttMqonvJtAIz4m2H4TrCy6xo9+qHKE35w1QU1DZdZEaXTGGsP
hxGBH4Anpbt1C0/QKqhjtoOIuC9bPQyUe8EBZLTCENFTxpUTK5bpuU5fP7pdOvDIVfG04B9aCLgv
SLUk2GxdmMNbp/gXHoXz0FXaTskUQ5wI8SXoqaDdZnl8JJ2ocT4hYElDnQpZLMK8J+3Yx+LYWoxh
I+vvKNEjOJley5BNQgYbUm4zCsSze5IE+Qs/XIYh5Se19Yz8QlvhmjaBqc8LwdzNR2Iu4VJR1Tes
Df/nb76s0fxTSJwoYwON7ufRvz+76A2ZOy1yRuSKWS4kME0sUCRCKTsLNlwEVcmLJ2gULkyrKHKP
H3uRk3OmnL8HdSw6grUMq59PEJwHj/Zd/xvf7fRpWhwRl325XdEJGd+WudrfAa+L/MDMVDulKW/m
yx1Z8tWOl7IpaLasnm7zmtzGMgy2OwnL0Vhpp4QGwl4o3Ucr17kwllhxYI0vIk2zRWKjILO1ySd2
XiRgkNk0yaPFUEDqP8v3Yjl59l8dFM47KhmzdsC1eIuv7G6yX+uGxe3D9K3ZCsjnZNra+dDmzFJj
cUqNI+Xc0xjOeIT7YbcQb5g3Sn28+Scbqv4U++7K6VcC/d4KJYy3ivyInG7XXTyrzX5asTXF9b/z
la0jQBHuTP4G15XBb0VCebtjZ6hkheDWhcDU49qtAaQog+KZc4i1yJLlX2YFOw24332Eki9UOGPd
/wH/gbjyHnl3ilqw+VuAP80/OEEkFb8Cmpg5xuT62LLCmgl0ixIe01Ofj+L9Scn5Xwwj5nuwJOxZ
ZZcdM91cV667uz0TZaUmI35h5uD0drM1lczTvpYAwUFqhQxna2vWeEZz2Hhc0zvrkM+dsZz2DC7w
IvnvSE8pxi38fN+B2tXasHVzeRd4RuZHp+urIPaTNW6rkqjEaiKgGXQX7p0PQC4YCkNOKyqKtjsa
fjyCNxyPvwlXoKr9lyxTW5KfO56M1L4qCfylt71Hg0M0vpJBPh3ICm/c5tc3/p5SK1nzxlIH3pB7
aisyZL3NCdAYEVcmDCPpnxEdb3nipQz9Q4ig5zsni3pAqpoXSq6/8xRov30tLt4WA1ECRIVom7HE
2KJOHZ/fgB9HlcrTnk8l4SUMfZR5o+1XFjna5kmLLant4Yazj696G4YWy04waE4UqBFjQubVxFr4
XX2JuHf9QmUMon6EWBWdmsm2/HD8wVWUp9nCjwh4qpGs4bIJjEfk/Vviw6uaYHU+0bQj9LfJo2dd
6RF6VhwAPpfh2GKoFDzJDuUss5Ooym2LX+mVOJEHAO1C+GvAba5Syt588mMVwJeb5JguKc6wTI7n
eQY306wBEJFY4waBxYhvSY/JoKURNWu+LzYZCFcUCBVmE+MK5Cn9rB1hRN7FxSN60joyVAzicp2w
FqnnlzJgmiiYuldhM2agYfhvLp7j4Zip82BwessAL7V839kaygVYLQkALNYU8ADRzyzJ0tWCegnY
xuYV8H2Zj/ZmfC7T1RlW/371JIUCU8QVXcfpFKsLmL2K9/+8wbolUxuEYfK2spBOLCwic4fhG3H7
qBX5guswhUIiIY8DYeoNEv1DALUXHBlfsa2FHlbptzyDWOHdMBUnKUdEpGdlWWjNN1Fx1o4aKhE9
0dx18Ud3qNXUuhF7Ix9OKpNpoKjJD5dLd/ElH5dzbe1hK3B/aW129jeTt9ypkPhazJcvqC65MzqH
CbWKXHCK69HY2YQGCGl/1tqt6Apc3vdrwFbAAItNdTKVH7qn5SiFwu0s+dG60dDQwBECXIUIhxeL
ZbnkYQRP3yzAIfoam7Zn1XUHqX3192z05fANS2IXDbAxnTziOrbww9eYAn+zFL8KxO8SIX6QBlpk
mtxPFTCEGur0K0xAVbhnyU10pmB9GWrwwmvV1B6UxnYC4nveiEul8k7dt1oz+3pSKO1IGDkj4bKZ
Hkfp3mL5OTbJngkDkH9Hq+ICsc8NJl3/NHBmc5/xB8HfQGcC90hYIWLDC6UzYOQa+/nBpJ5WESnt
ijzjCpcAeYYIM1l9mjXb7kTZs6n0pUrNIAWgvpPyTO0MbcHXq8G+fyXEpClX7lUV9oynvUzxxtzW
377XZ+tOK6PxAkDlCpH5/oAfP5Zb0B01yTUlg0FAA9b6PfEulGsJSLA2x96CESGhB2RSUWLU5ryk
DRcyeBYN4AZMxkc+HVnHuAU6DNwG35+oKU7Dl4jHgDCXJAQmEehYRMo2X93TOv7+rHszPWyVghrH
tVXvikSXqmnYXmVmqp7FuvrB5ZTmpM3sGXCDH+G0C1lxGKsHjEeTWnFjv5N4Ul/IcTKQMvu+W2oy
llbVkzz3V5y8pm4j6eek5O11xH4pWhrnL906g0bh8rcV/lyIQ0HBqgxZsOPzEmE1WGTZBuKaR692
s34MtZEqKMucUixI1hn+zokwehkPONRpr9AD0TBd+NpP3yLjVNqNovxZY48QEU7aM4+Sn0ujT6+H
CX7kVSOwG69waYNCL4pY08NmVxX4AYc5JzamZvWBPUMsdc0/pP1th3EnDccpikx2fN8cZz2iVvkM
DRuOU4hIQRTDkxE04oQOuMfpqP0BmYyp03NdcdaSU4qc/mxzAxBMbXWbCKePLK3NRp+Zf5+qiodg
1eeMXe2WoaEg2K8VPBTHcoqdEX7NQB3Jb0bampqTL9VkkgqIcgCAt4C4mxRR//ICTnVhYX/awsoM
Bf6Hehb2O/xasaracGRERy2Eir/1o860Rbrd92KNKRGOZK2V1QrxLXJyrLDqdcOx8BMllcWHxvvt
8qCBkuHQ/k4wW/NrtVMUAOBJruURfwfEAi2RmDuRkf3o/5RxKPy67lEbM011YUWhULvg1Ce8sch/
09JTV+fceSPRxPjd1vwl3uwWXKmmd6AngjhvMqIlpsld3I3xx3gEZ+JX3QBXz67eTCMYFmsntVP1
fP9s7aWCFaEamB9M381J7Vn9v80WTPjIdWrYjFBu6Bu94d35sitqwDBIwowvJYIss6CJCW3gmJdx
I5+ryWwfNvxO2l94gy1jjp09vbB7tnJWq/tTC9idaHPJt0tYnuCOR/7bovXMEkTscZS5JS+t32yl
Y6mUVC02NYk0y2ClVCSArppygIZKp5Dkt6z1fMkXkMMKpbWVZfIa/+jUOcSOZsgY1bXAx8oCFeck
3XqYAl/5Sb9a0yWRTp/4IUR9I+NNqqFaCbg/beF8ET3dRluhlhSiEiBnXnMlJqHE8+kPxO2CDl/L
Rpe69GKrxVo0a8uH7pZT/wg/dbMmmqCmxwOGNWppSln/cDHc7YnR59n41iw8gMFo06oZLtB4WCmt
HXCvS1GNKk4xdikfxiuS3CE30OBKViC1ZaFwlmrqzE+gk35HvEdHOoOEeD9/4BcLng9IerGYxVtF
4l4dZxWpdW0Fy4SwpPgwxv3MBREu9/IKVgTwbVwxQtnl38GqXp7gv8h6oFTYhL58b0a0FWjtWIKv
9MgNI+XnzEhllg+tOKkVOqBTdbcsMq0H82cmps8MSt+TK2odYPxWNVpxE10aW3dnQhIW4oM86vHH
S2j35xxXAXeDQoEGT0EnNPDOPX8AEqQmFLZ+I3gBLpAcjP5/uH2vR7oWQlr3Y8u4PP7QgU7KbkMf
pFd+6Gkjz23LElFHgwjN4ORNuoQqPCDKUHDTCSUpfeP0557Y37ZC44VpvJfXMbGeSQ+dJ3QJWZi/
SwXPfhnlt1xP52RF+KGA7a/qT1OgU29TeFxhgqLXfJhT+WzQ1SmOW0/Ile3uoPkHZlTvOSAICjz/
phsow5iT0ZIMdclYt7S4ydukX5R+MenK6gacvF4Woc5V4HJ9xUSDIIa3Fl8Q1niiYD69Scv1EVVo
vrwSx/ia540DxB0GhWfY8CTYpUv9dzyBFmAzmS65EnU0NfyYJi0vmjhCRgFfT8UlTB1sJ1ZSdRP2
KcpwJkp0bmlmyuaMMDprXzMPD1Jnw5u8m1FT6xxoKRHxZ2x5NbU82b5YfKbgcs4Jfg626N3gJvKx
Vu/X4yMjz27bJ8FQFfera2SBcrzGUKKfJkrFgI7uxkqzMrqcYCUvMUSvbWo8NZj9TAGSoOtVdLru
ES+8gI2uK83i0AclsZ7xOGD7gvsnWcKtJPKooOJPVCnNr9nPgehuP2ihT+1FRkDfZw36gbTCS62y
JgEWIcd1SpMwUpgWDrTNH6f8aTnsn8cvFiXiSGOwndcomM/C1HDEpfk7Up4M203+N7LWFDcp2xTA
lpQ5ILtMgbH7L0o7dj+KpSxESihR0H+wfwyJhp7Dkr1dT+V2F5nNaQrNfBlPK7cWSxGWqueTPHaw
CtKjomsPtmT7vYnNWlR5M7TgDFkjsfI5KZT94wbqQcoOEvFHlSXR9WX0bQ3WemASZLEm1QsZgqXQ
3rRtlGp0RpVj8ygWDoerlEY9NxkgMNDZMi+FBnizFyyfCaM5RmlkVqKGB7l2du1e/i/XghpzWR5J
KHQ55ftMNUn6hnYtoJWgRA300RYbnRC9FK5hRdM5ptICbWKWEuz7czJ7Hc0sVtGNhN4GkJlNlJ7y
DiYAoMFUSH5KB/p5e88by3mMA/OHByNB7opcphMCxGStw1YBh0sDVFgBI5Zi4iFjGD9WnV+U7ypd
0keqOF7RaWFJBJqNyf4Er+4wqKS3f1sUVXsNjxjm6eBshJPDesf8PuWc2xZU2DO/ptBsoJoBCpOl
XqjW5lhUpeYUTnjPMXp96ATlyB03FkmX/OvNXuvSJLsSwrHTtNpSetCmJdjoQZL7x+rXyaHyET9H
d5O3FiSuL6joBy16dKvFfeuGKKrOl8VUn3GvVL3HxzTG1k2nEaBsxnKWp1qO7E8ibsuSyuC7RSQW
zDQIgKR8sawhdgntCKb9Fi9zz0YmSJGy0QncchcfXDT7QZq+y4W0bYg0ybGakScr0z7vsxKZsh88
23b+bgxLu52YavRRjayrdVtNeS+48PYRWUjvySfCwp8oS7i2TeuogM5nZO+lzqgrGb6eS4iPrjDq
dcgRSpA+ZvuPvr4WGBG685CntCK2B2/o94YElavcsUH5ZPnxxFmgKQs6Jvtux54gdVcBzDK8Zrwj
0ow8BfjsIZPvdW/eVOkvtk3RjMjmHezREAzZgK7N8YMPKtGvd8YfFctaGE+84NAkPUVhM1+vTsJ7
wXxqy+jdejbnEa2y+hcqvRUZDxMrR/k+xM2FYbtPs3HDQeC63IETWCyFV1fTvmatfLDwk09zyxaX
CHNpw4xfaYp026qjHzEU2ijb3th7n5xCEZQ9kYKzJnEqjmFLcEkVwx8SvbRORFvwD+XAbJGDpQU8
RLldNNAI8FhRTKj0DYyZ30TCh1jre6Rki3pEqw60wdmv+AvKFU0GXRCUqaafdpP31qt1rM/x6njp
KgAAyBnP9318kXLTayyxJNV6RxncRdTFGP3qwQne7mzGB5jMevgbwpRMoc3bUYy5RmWSm/IPwd9r
rBaIQBeBLmxTkub7eJ43ceaOGpVtbpDPI94t+JonRuQmX10ommG52SZ26Ng6vlq/YDUVUW0fVBrX
yQebmKjWS7Qcu5falPybv4v885l0YfMJasfZpTBAnq0N/pslj7BeyaRgOCFN8s1VX8DMJeWk38rK
kppDr1rcFx4tFqMFMTnrFXf+qYHduyv/6ZalnYu1K4Rd1zHADR5745hP1WM4ZZf0c1LaXbN+3t8p
NhXA6PnXXX59KM3Re3rSZeRtGs7DZt4BZ9XadbyxspYlFNXLfyXGFvGY01Vq9LIChSycGEVPldSq
NrI/fxF3K76dys2Nc7yILKGvmVW8XRQlSYBQYTo/SbzypZDLMYwFXt+aa4XKGyrVDIBoVQcfV283
3QNN2n9YKMVxRfTzE+3cQvBp3bQzXrBdd4Hw9iWk3hDV1R2w+OzAMFG8syMf1roDLCEXm9xTSM8M
o27g1+fOISo+8q/4ApKTnGUf0j4g8Vv36qXS9RbSJnp6xNWjxRQKq6+z44Of7AGGgLJBke0sCsjx
oPUThhqbizUFpdjUiKmnxDYPeskJpo0pknmpjrZaA9k89+OQLBhQ4h0ocM+qDZBCeIbHaW66asrF
HTLzJu0m4rfTr/4fpkpq5li13Cnvmd2ID+NM1TXeMpAghVXzM9QuUis6rBolxf/nR/gLZMIXPD9u
RJcyNg3cBmBQQjEUaDyC7uzXaSykLIvZ9Z3WSTjCcnAIzdXgTOp4iWfwrV2bs+fCeCJvo6hXoYO7
cJKkFuBfD8KtLAicguXjzoFd5Dv1VCd7Mc5/gwG8VRls62uEdpYte0VcQtyfEYZiN8Eza1oCnNg7
vzFVCFfFnfKyC2V9zkkyvhWHLCDAKPiVyM3bHE6K/Id7NPTAhz1js15myGNoCs62AomXA3WVWEin
xRpPvl0xNMqlQ0Z/2y/vtgbyy91gqG82Dop8+6IOrK9nPQH4ZBCnMe8hjAHWnaYQYuJ2czlv67C+
NkQULpEeE3QsaBB6WauWx2/hpEc8vz6heLHTc96j2iN21teXMDu55ZRTTRXPZY0lKortQcGIhjbu
pfpO5ddCSmaQ5kGcuLRxkgiHQpnFBa5jO0eL5hosxPU6q7SroGlftyckcO4BeZfzxYwFaJW6Xakj
cglHySDu6g1byPZQbwNALmZ1xKtwkr+oJH19MRAQlbqIHaJmImYvCZhekWg5FBS7OvZFsU8U/jNm
0x+12RIrIvC+X5mmv/MxXJcY24nOJqObOStb4qpod8w84yThV5wO6oEjtU3+gn90EJbSh9/Fv7lh
47t5bwgUlind5EReCBK2QKndQ1RG+zC3boS5D9YUnNB3bNeF9pv5KKdxCoPuiOf6JkABc+HHgWIw
llAIy3PfthgU2RCq2dR3J+rUUKSmiPVAZc2ZtknYOTo/jfxYQ8mfcb1/q46tfjsQ4V8ABWGlG1Mm
feRNRANKx18Nb/NjrmlAn8Zu+PBI0lQy01BoKrNWyvXNwl68JmEbV4AjADpG9hAs+/4Ym0/P1Prm
rj/TnRFI1OYuoB0bulsMUnkYRHUMn6gSANncc1d61n/P1XDHkrbDNjft1s65S0PxgJlQsZEl/4w/
9BVqNI/yhrzwfF+MGHlj1tx0/VzXnQsZUiTyESVhzJI/AB5Y1UrKbTX270SdPDO2kcznoDp78qQG
gnvGjt/Vev7qQQoFjMBYkxZtBQ+gsIiL7INa2nG+nlYEYT04231Kry+KzmVSG1Wf6FGOk+Y274jB
mY8q28XCmyZyKtyG4Tn9MxyNXja5zSbwGEuOcCqhWP6+dCgdLTdHQgF8kJScqrMO1KoFimAvyVZp
jRwx+vrEsfXJ09YsgpFXysVaOYnDx+Aezk9s67UBvsm2umZo/wgQltZFLF7ruIsNe4oe8cD3omVb
Zhnx/0h813qM7lkC1ZLNP83woXRc1XKV/eJPQAs97P4g7KxAhdJcGFvzAVpZ9Enrk42fsasFbmN5
H2IGwknGCymEVzNpWOAHF4gY3+c67MZyIlj+g0/k1fxvGLsgaky8yIwg4ZoXi78vz32RwCZbawhP
Ad4mYdOnUBqRUAX79uLQPI7p2kDea3D0yqY+WTsPJMwWOLZbGfiFDlqO//WDUlGFyAGp281YMhFi
tESXthffUaH9MZKfOXoGyqR5UgecxE3vmh1vCq6aueweJ50RNmLnNnnC8h6m02MZQ+CWLUdUlLDg
LqRep5iGFSyLyeJJrouAsqoKtdpuEXLIC+ck7hgFmk7Yc1hv/Vk8vPoKlQBWAk/aghu8zqtY3oUw
sorhGTBj7A5fqPwWLE5kaDsaBkoe91QJXP6pXNrOzWH5kxzJNOil03z9paVKpAdCu3AlN5osYz2s
9mvuKfSwYf9o3Y1obBcL2njnezbyKNV4I5mFzwUboOFy+4OTudXr6W7rSJxVEDVbyhFp+MbnhaNR
scZpX1oxk8kC875vAipYdjZ4NoH4Y5BMo283TWAT+HqZjyEY9Uhbz4tI/P3/K/5oidpbiGKkv9Co
PY0wlvtiLQFv3Gp7vIptUb8RhlptycrSsn3widRh82k4zZOyyabLDy6+QqDhJcF4lDiI1fKyissz
fddbI/MWGR9PC+reJtcO1FkoQR+BwBGbA3v088TgNbg0a6VZFEfL5E+kLv0rCXkLlr0kpTxk5PO9
+XRD+Ob2IDEVdjZsafBV7TuZAU+nPenyhtZ+IU9h3ip4xok0ZjmtFGmKukNhvFylnAr6p8jEjCVu
ph6fiEQ+3Lwxl6glLFwFRE9IRhB1pajfAnz7Q1+fGiFFazPc6W/wO01PI4Z9tf48eEgI3zye7/Xp
J9X5asUGw6REypliGpqA2wJRH7hWo3GOOzzXhXABs/6WXW0TAe6yLSRXu8kXhvDvDY98FCiV10dl
8fPDLlVt8zosFerLeXk8HiDIZJOnCKq6Y7gmZbpVpvLAK/Vyze4AddJ5Gr/gqY4J2UTIR7Qz5RKG
zRS+a27rcDDzWVH+Fus+EJNfm6qzui9i4k9bMYO0ukyK4oby2ifRG0sTdNcJQiHeMbQ2kHYK3RZQ
1nkpJCJVKDzuONTKGgi+nroLtWk8Q9ujQlFMnKaF9Q0rGb/FOIceFqcevDd2DA9TK33oGlmxoMdz
dH0mERbcWlUOp0dKWZ8IqIZ90vCwycQhL0GQw7UY9JLFTcuEVAabvZQ6AEfYc8re9M2Lb1nAC/C6
n+N36RUjM6vXyJ6Xw+BUzYkLIo1OhSEiI6L/WUtV4/o1EJIm/4VH1yfMLBPsRwd+HxPWiNb54KZi
+IxFKJEr9lFbXBaOZ8P8fmi995+BvDI/5PNLjVEoJExBXVgyBPS/SbNosOTK4lyNSReDx2CcMrRn
ex8FW1DlKnIWXoy5pMf76EC6noTGNSJirFSrifcc7bisGNXsffyl8LEDf2h87jECotJzqeQeqjFc
ceRnwT27K72W4z9wl4BMJZhMuSSsOdA4nznUsh+9wodgv0VGIxezeqrXYR3bepHyHFf4cmxHq+Ha
mPmY7h6Aq5/DWU1HvI/9BLJaRWOgso8yHmkccdq/rTOXK1N12Bk99l39Os2GVZOFzI+3vBfew+9r
qJj8DCXIDg0TeIZKNri9l4ZIrD4blY2mBzRqm08tXpaPYdlMIkWmVSL1eFNlB3KsJ0IypEPPeVbF
AYmacEvN7SjT8qOI1gauG/2JfhgDscGVcB0M+F6oQdsAbpvau0U5vMf2AuWOgCeaJdoEYX+/we2a
ro+eJ9wSLqPsBi8N9rMGRZzGOL+GnOmPgIua12JNhL7Bs2PVhQTyYEUUOhok8x4GAFtChb8tW7cp
IfEUmst9kqULuDWg/IqS/zawsUxMumAbsEu3OPv1S41R7mNV16nKPiFFi+KlsvdRzPlXCQBau6/j
8ReAP0O0MrJl58A4CEcnTXl5h1NR6DXuavGaV3Vy2A6JEyHxJjcUNT7UEv4PzJFdVJiWbFbIm1Em
yGXDLj/Tmn7A7iLtv6YzbxZMHgOTXCvI+PBqoEgU2opmcqCo0hpgGlQklMqVbl3vgl4oSaguJ4Ay
jRIcp1Aq4ViqbI4gvkGmv/A1KyjRiYNjbc/qgg1bpobTWokYmHXkP5LkHWNhaniTGVkdw2G7Zw2r
YSuhc4vxFm3Dtv/EyJXRMEfi1DQKQcs+o1QNOVmlDgbl+jAUHn6YWUevJsQ5wRSr3NsFbuaq47Q2
c/nRaMi0MFggXR7WfN/I7jg+a6z/xva19KrXWlO48isDR2KXHbJb8Lcg6FrTdu8fcVdromciqP1E
FhDM8e7bDQBsZQ9oI3+rh6PvJdV72esDCJnC+3i2vHlmf7ERvlXyeoG8mTCWq1NO913hy9emKSQ7
SIY12c0waxZ6v3tGPL9lBUzppFvZye9VRX9r/lVJjJdsW7R1FIoEXjzLTuWX5tJnJ35WxgWXN8FR
qlQuQ8jB7aiZRujBqtPZV21656T+QV32y0MZby/BSkRXx+oVuA/F3w9DkJgdEPHAZW/ilAGast4I
fbKAxV5jVdeJ4l4AytEP52L4F8DSRFw9pRoyZ8u2akAUQkeW0bn2zeDkv4gxL/LrQhnOWJI2shJO
1BNvSCEtkq8JjmdjxmS+I4CHTHXDEcoa6PhHXi+/vvSRfUsP3tViQlZnV5HCTLRYUcGVUaP8d5/q
i04J1HWNQ5ImU9Pw44aQa3gC23tyBRjfsCUKS/ZdzdclYi/eyBOqXiRL4r4mIfUp0gCV+iSppCDU
f8Om+ad2qLQ6k2/8+ktl1myfmAuVo4zdy5mVWijyFxZX90vZJ3xNwz9lmMnvEpR/hw5+zugUOBUG
GdKCay8MQ4X/gkbBehBBMuw29Y+PxyTD9z9lH0EofrgG3QHsiDDvCqhGqx4G6Ycfdfe8kvA9+/Sz
WpSqOEALA0GmDTd4tE5XBYOGKnOkKZhmZbb6pR5F+rSWyhu9Nt/tGGN4izrfppOf/WAF2M2GXejk
hTnXfUFt8cyLeKrGmoWf1PgyGuPGd+b6hmuc1gZVXhzL3zb0iM7M+djARTtmu7B3neM5mOMgIpbA
EQx2/Ihj52KQcZbvi/7UHpuRSVvmuRZd+Fn+CYjcHj8wDSfUgJpxZcEEjtYHQbyG1rUptfNPeS9H
PNjp+Rg6Jt6pqCMuEwqLa00Bz6ZGIPXUhmTBgo+1l79076OGCGQyUhdbYtFw4A+SSGrFTlJBJ00G
wPx/c3PI+UJJ4eiTZKPla24VJSRNWOPsC/4cF36h8bcFGiX/xcb0erOlK0gdflEdQRCqq78c1w/E
FHKOsKFVye6CxMPF9ni4yEdUXIcSHKPEJhj5I8WVBxsngjyL+sFeuZm02/yoRgBeLeHFn+ZeWzIZ
O3vgsEMD01hSNNK5SJ32RdHn/qIy/VrgJsws+Nqb8OcHc/0QS48SINAbPT1qsTxGl03ufNf48Ac6
M66Bk9zumaOzw7kY9dbdVe6anMDwJ4Lf3LFJKwIcnd4Xgkm3uW47Js1t9PZPkshw9ijQznvg8VyI
D71l4MedRRE43ucyckqNLWI1bxdy0je0nWr6IEpmntRwDD1tTmLxR1kNUJVzb+YsbM4NGTBsgZpg
ZFxy9tNH5VNMDS1MtUZTp8j0NemlO65Bko+UsIGjSCK0DWxRcRfoN8ARP7PIiBusvRNhdWtVKgYr
W6cFLxrNxSUdmGu3GAyEnx7T87BCk4eGaWngDT0IoRsGnrh/lDT/dEMddnqZB+wtrxXbvmzuBnwB
dMWra3sSvyYukUZAcOhNK3rhsShftTQFgH/FmoUti1U/lm4EyRfZtYoexd39JtT8xWOMkfOPq0Jo
5fm4apLkkP8qkj9UG2LSufXL2LXVddrG5+TWoeS5L3rYquUy76t4YbWwwz/EC3BbIL2II9uMjJCr
JwF5ZeIl96DYb44pSWKPKfZLnt1IHyoTbslqx2fXHmbcHZKiymzGOflB9JHeZlSMJ0QSmJyGGCBF
S26j1+buvULjkK5IghyIKP6zkGLRy2H5Uz/H03FyvTW/IaOXuB397TiVXXxomjSeLM+6+VDNiFYu
vRNaEik1R5xaV/9BhCvqpqmKpaKUfesJd3GJf9GN0ZASZf8K6DNdCw8nsKVhT0KhgCyT5l7DVMHa
bGFNtK3GDTwk3Js8UzXDLGK2yh4H4ib/cDfeGu6lF/XX3ufRssGN9Rn9A+kII0K3ieDTJHZ3PUbM
dgoSP+oEoywLmMmix9Y/hQwjSwwWrU8yPWRiufOfJN0+daD6czj4BuvsVxIOi9fnEMG2rCvIJtEQ
HHFhkIyb9UExmCRXD82Ut9zxOKL1ayhzlljniQZtq10nZNOhmfGjvbkTvTKxL7qx540jwJVpKLzr
qdDmvOpQtwELdX53jCkpmjS0XSq4Z8wNO6G1F8uOIgye+updrWFi11KmYcDgDYBxRxNCt8k7flDt
Ln7BW5n/QY+5DjQwOunF4lCJKzy93TvA1zxR0CVYukYqaII9iYU0aOy+hAteAf87dWvU/4EHq1rW
G+417uaH3YWqZHcrMz2UZT9PcJETzcpWNOeeIImFtW4ymZ6GNjvIhiln+N8mjMOJD7K83rM79S33
qDFZJnfXcOH2GKQn0/d6mEODMwOfkiFklrErtm1Lnk10Py3/eTFem/SYnxh1f5ltHNp9tflZedYg
G3PPmglO3bTY686uLTTX4DLDzpP/5HYQIe1xYicjCzhdWHw6jtC4xdMwlWXnEDCrAqOlE2cpdkGX
yBQStM2/dXiTCDBNJG3VMX8cRoKy5T6CfxODgKhNL+WeC53P9dJrvleYFCUszNlA0n8Osxeu6kt2
NwHJpmbgSlspbwGRT22PcFZUvRoizQGzfuDRRwZ+h6yGJ14wRRHvpyNWGLQYK+NgMU3T0UxwdE9n
+LOOu5J2WRw7pXX1FhBuh6C8lhAGjEi33XylHu/IEPYOSLntIaGj7dtWLZCiOiFu2TpcLu9GApv0
YbnT/mJrbHf0V9j8ruBdVPWpulupCZiQPFsBVWNDjGwLES1KWz+KvMjEoV0KAXrTi1P56AC9jXCc
8nhkCN39JAX1VTsyhPpEnaKm+h/YhMpFfX30eEGZ7KRoA8er6vAYVLklsDuAhegYVtFwVcw+TSRk
zVZeo5UJn1KT8GI611yuCjl4aT3ObdPZsSi7xAanTLzDv8QwftrSU3KKGoqs0inB01+ZIcb7PUpo
Xo3WSLNpH+cOq5BKCrpRj3rSOAbMwx0IaNbhMrDTHADlKDb9jfnv9iFZzmYNhciJo5GRAaegfEHS
oppQzAOAGSZfHLfPt/J9g4Gee41S0bvEp50rBaM4HLv3k96+Lg4e2bF41ae/wWKbrxLIJEg1RsH+
IlRyoOnOqfL7G7KwmjGocq+oDwNn0FeTOnsbNy9Bthvq2WOs1D4mxByQD/HPfahSyOU49UpnoXy2
6wt0k9UlSbDcMze4dN6uusGyaeF9Fv584rQtkSiU78zYY1VMTKKMQz0EvkVKddmdhQF5+0K7SBeD
KmjJSZlrM8+ScgNcgrJOoLAuBStuWQESXku+nvAPVqzNQnPFSg3wMeliogcNF20+7xXSsVvsFWH5
2lsnt2JQyrZIBmIfyR2IXYieIaGBtXq9R8wsRrD6nKS1qZcevWXPKaaff/5KFUDSIlMi++4VIsUi
Y20bAr27jl0WRH0X1iQE8K+ue8Kx4vKjkIHMbagvH/KUzpQFpGvlR5LtpjQfLXf2BsDq1JFB39As
jNlmqmF1OaW1hIPEJEunZr+4y+72/iZKritilKmNRzKQ4OOSqJ9iYbE8KHhcIlxDa9cbHi2EsFvn
NXiTCgVmfy8FxPr6x+/Yq7EEWOTHTKDtMHoiGpXh7wlEOnEOFb8O7YXYTxnsGC0fvEE0ZpQUApB+
mEHyoNrgUYRG4H7w/UEdz1SDsThJ8VuNQ13uKxgDEyQHw8XttIsrSF/Z7oN5rY8Y55Wt4aZKp48Z
aky7uIyCc/WTzRZN90M5Bo61frIk6dluiewe706MujKesO86o33bEE6j6q89RHAiypzdD/LLUAgh
cGvQ1Zp1st5VLZYi8CC/GOTMY5nmBRCXKJXGCZH1XEZ6xqSphDWF54Ydlm5HLPCwfN45rBbDjfjx
qMgSUUqrQycFSAKaO7YoUNNqULEITQAbs759ZpRAusUkG8r0XYpICU96CoPXbmqlkx2VAc9wYzRj
/TiKFeUROKu0m1uKrB2FHwDHym0C57TsCucHxW1XEsgN4jzNxzF7hlYOgUrFjYw+p/K0JNBr4TOA
JUdEwmjghkmyDgBwuGXhed0DcPgtBuB2jGyEK/PDSIwZo+oOZq3tLET0ZXZI3Z+1vbaQNehKn5/8
+z864fTc6oYFuitImRfbtL8Q9Frd/snswx0XF0vhu52r46m5bXv3daqnebo32wN/aRWog0yUeq9U
UXVurC8blhiuoXKTgm9aphvohK6koQq5OcbI2GLgVRLLYLiENxP4CDDCPhQWclvj4Q86U1GMbTME
+wFhjjxMYQEk/BXlNSlNyFRj8KMqw6Cj5dmwnxl6iBVhNCrtHaRAeTMkqWT6YSxHjx8RPMBq1J2W
XG7Haz0P5wBjKu2D9SAyMWEtvgHRsC8tjsZmFkMpwljVJEGpoSNbDDA8tx+Qjls8Gw0E6EbCXfoS
0TWXjHofpd9xdI4nvKj2AlQXYvAoVgpPdIjiXL1tMTTCF3UtRfMn1HqK/q1mJfxFRAj2bjv+clDW
6YCDHMpsXR7/EQL9fxrEhXTScyrWPbSwjp4Z+NJEjOXxfpZU2ls+wuBS9KuLU8jHvIkirzNl7tIh
YUazfH0z+1tWmEpxTD2NUNUpS6wZdULd1UBLTvHJKefpmu/E1pRovYKq9XOQb/9JRwnXn7LDhZm5
qas72BPW8sewFjd/jiQPiaswnfMCccXNAA7N7Xj1J8UH12XHP830J3kg7eogFH7qpMz3/dQM5azJ
Qsz5nbj8xKqLK4+xcjm5krnnT+b3ta6WLI5ghzg4UPk7sl4rr7OujGQ5UzeDhg6LD79ujABYOihs
mybkA1j9hcIrTXYH3zYsjKlhuFY9WjlhTqleAJozT8L0b2k7kLn9nTd0hYOhNJqy9C2mnsMfXb0G
2bH92RQ7nXRaoMOkvvJZViI7VHm7xYvG8I+twDxEBVsK2uQeJgpZAqoU4ib4Gf2yuBCAAwCxGVog
zevIjApDgRwLYt+WBnFOmV5LDwN9DcJpz1sjmG1w+1GHxEoalwE+9AAbZZs1nvyCbAu5HZxU3KG2
M8Hpeb8R1U+mldEMndwDAeu72qxwTVdZ4v+7MHoY+jqV0EItWx82HMyv4FXUHPehwMheFp0Sm5jq
yrvB4p/FubNPyEhj2TJWEjmlhdK1tR6KhiYum6aa4UVimMc1sF4uYbpNwiJ7+eiMYTl0mpJUWJVL
hI6g+8lz+TzRPpy3HD970vEJuIagfSvywIWOWiAz9JJqavF1lzbGdGUnLoU5mKlAfuEv788F/iaj
bA6H14vcltD9XqGS3tkQU7GKQJ5t0ad5zCfyTzuTpFTQW3GQppQx+Di+31B9021fAb6pyNjbHv5K
ONb4AcoNsFv39I6eYth+hb3bP4F+mR3lA8H71ZfVho5eVIWyvByoyQNTg4WFg+n1rwQkE8byC47P
iugxxilEzsKuUCqvp5G0rPT7eijJlRxyTBn5/Vt1klT/ZpyLZBfLOnJ/YdxJxeH/siQJHDScG0X+
ZwLunAQ7qj4dPkrPRUFyewKIe1CUPCH46RMTZ/oYinA+fTVxOdTSm6u+MFEVE7D96QJVYpo01Ek/
doh88mc/6oeWX1fl0nP43GW8pU1hxJZgRSg9bxiVsYNFwPXBw+KJ4oFu2FLJypH6hHQ++iQPD48n
RXrOnb4EerZxRzg6K0Ks43Z5GNUy79BIm4w1Lqu0mz7Drxll/vrT5F+Y8cyQoCt8u/YxXgtUBWhm
Z4ti6tnGq0uhberu1q46iCPRaXFOSpef0IOXStijVHh6tMQmYx/FBL2ZYlhK6Pots8yv1jhESJ16
rdL/pTSqZeY2gzpiMZcEyfSqNJwPpeavXqa1Tfa7jLiNExFjwbXg+BSl0a0wwPq7r142Ei/rQmjE
6eJ1bBZ0WgXhrTXhw+m+adas8bHF+k9gRT8s5qA9ByNKtuw4w3Pz6CfsPnh29Wh3TfsHrB0PMBZx
XA4ooq5jdwfjODsAUJ5wtxVYALL0PdrCzQzvR865fnswPSMNrAZSmnxWXu3PPNEQGyN82fPC5Z5p
5T0QLWz3hSKTD8dNRzdN/07sqjN4Ko8YjLnK8WAOY+7DJBxG4l4G5A9zqnA5jyASHj7puOcTB/de
4dDEWTZNZ9SLBtmAM/AfgxLInl2ffTQqj/esDXeKX77onQImsmkbq4IaSEBCZB+hqyGfbGcL3VBf
bW7E2Is1EgOYzsHXqUet+66ZNBtjIAvh5waXbb8H4g3xxRo4TarmPq822EVYP8i6JdGfKy/5H2ob
WlA7Bd3sOvucfYR7kyyPKpX8jJfMn2hBE4awqBvr6ldF1Cuj36Eaj1FiSagheJhT51+hYKlXxEel
2Jn1qBJIymbVe8J1fAyJqlha11WZpfShE/ZxK5IyzcC1+Nlmh7GwchU12tbBDCw5HfD8bpBVv/Rv
xSyAfFFIqJA843Naa/sNPONkUDESRscVRpPzTZY2qPuZ8evMUu2cu6KO0Vt4FKsx9PLLtwt2Rs97
LXFkegycUlRl22D1OgF8aERxGgm0dVIGWMXUidSaSUezSHHe7lYbJBFBjrIG4yUFcdyRe7xNN7Oh
bZ4jY0R98fiwR5USCCtOGfrlBJl+taQJy1SXl1cgnvAA25D3CfSIcp4UaoC5HdWlKoLpHuwNd7+J
MwdDaUuKk49nmzIuWPsQc5/w3Q1lZI6sJwspxTf2aCO9DVyM0KUPTFVr++Xd1+jLnxG3xboxnpPS
65LKvvgl7ymXrijAwrmDSdzUIl4DzA5LcrvThoYbhATUzwmxDjOVey71dfhghxYnXsOY9zAusu9J
LwnN70g29mlkvnqyty/TGdApRl7i1dtWE6AastiOeklLq2lLtoQgjFh4uiTdmKEuFtidI2grqafi
c0TSeYVU02nl3ashlZBaOAvcEV3FzmuXyvSjFw22fyHUBmd+9abB42uZDW4JHilzhuR4i9biCxDC
WfLlrNsCkRm/SSpDJVUyzaDIf/uXd23JEueJVBLdn5dAINAc5dU+RdBZxm+riZ8JEb+A45taVe0u
rpxqUaj2PeSvBTX/hXXYZ+/ScQoJpxWqi211w1fLw8y/pN1YVRkVxZOSsT9SVgFtuh70zPhvi3a7
g2B2yFzDeiClGDNpPMBmdNKRr5X+UH/Y0BqX1JnR4pGjTCvUcz0trctlIg+UI0wfPNDTbHHC4hNN
8wgsN6h6BWWprw+q7X+G2MVj0eimH9mskxqpN0hwjais0PHqgd4m8XxqEFxBbcESYjcKV982FPnv
k0PENt7P5Ld5bd8TzJvIL/7QKnFDYYyxFlcgl8zLe1zvax36dclq4jxh0JSaV5BZVelr7Tad+MM4
VpVbMX9v5RZKg6JLeldUeMiOBPU4G5w9KLtyeyGjhzIs8LiodPxyPnemrj0WaAfCdrUkyY+L7BPX
kcQogeqeV0VlbQy/hldEnN1uusFM5QxsJy9fm5h1rTEiATCMfNit1tZBYTFPIUqOVqGl2mE+i6e0
5aumWebRIC9Ycs+cXkaV/P62leiOmR/TEUBH40GnlABMV2KC0f7g0tEYkkh7QAGDk/jPDRm2+xen
bL3afywL079qnz0A6+6mzRWJIHJn6dDTtJcEGAkCs7jHD3Zp03rnW8vRJpgxQ5Rb6dJIjg5UoN1Z
pkcbshAzE8ezcmc6cfBXAw1h5D9sH3O+nWOXteuwPZgtAaoKhAyVeOxBomloU9IqKZP5QqgHGAsw
2qc2I/AmgCRRhHxPlNan6r7GrNf449nzaEhr8qv605gLh+gniR3GF7jfCfWxNFWnCVctsg2YwWJO
Qo2U8yisnBmsKzw6Q1Nm7VTdEm/auZ0S1IHtIfDiqQi5IfyIxHFMWtck9kg3gRWX1TsnEAW6dRmY
yj9nNj7uc9BE7DJ3j1C7R42f1Pnaqduo6cOVj8i973WuFVRGx9xAZvbLkT2/HGRv5H2Jfy26S0/b
dL0iPyL8wy1vneOhqCB5EjXlua3EJdPbYRlmPqXhCa9UnzCrXvcU9aHAe1fTUsOL5JpWr7nQpYvw
9CS9rXgDTGyz0+anf4lwqCRveXuhCPemvrp0ZByGj4pc7SSV4Dn7R3eyjU4cwN7/hrqfHOIqY3ZD
bVhtUBG1Lyaa5vwHBin4EhUw+b5+viGNi45Axp/mL78/Pn0HCYvZ0kiyIFJUn5LnhGnUpRkoc+5A
fQMC5yiGGNAHqP75cfTNWRu85W0t1nRaJPzYfKnq41f2bMEKZ9brP0AI/GBpOXJYmdLE1hpfLqEL
FkKdJah6ik0kzu16O9cR+mDgikpfomCOXOt58RLomRhgZjQbV0I35HE8LxrAf1vosm1AYvQKDBSa
N3tiY0f6aSL+xKbsGMbEjMakg78/Mywk9BuvnFyc5hjHGVGyywUHM4gBKnLX7qhWAweIrYqXSb/0
CVuJQvmJyE9X5/hJT5VYoMpmpB/mjksNVm1pGiTVSeW+/cvVzaHlyAmN/saxjuITq4XjX5pT29++
I8BQmA8fY6AjAXL/l07AdR27zC3PrW4ljbYJ7dGFbs4b9MCyBBxfROmlWPK8BiWMIYsJ40Jsw3fV
6syXD0MWPU+eUclJwhmDl+o/str2ZL43MpJ/dsCojdcVGyhQkBYl1ltYYAPnY6TqGTNrHt09/rU3
dBTUC8aybYP7II+1ruHAhsTd1BSZGIV4uJTDVTPARkNOPvdW05HVX8Er5PoXIYbKlsJnkqReM5/X
RrcsSOU2VfCAnj3kio/ZmNPpF5zIIXgBebmCHNtUy3qjrt7bq9qm9xCfAT34U58eN+1fkGJNukf4
XM3NY9DiyEO5jlKusQbo//m49P7xMOIZXgFWyG7IwRgA/K9/2we5Au2qfZnxVcyPYO8GwBfyyjlF
//5LKyHROtv4qv+sS7sFFxpAK5t/lmh6eDcNY8pwwH+GaPkyk4xN6PxIpm8lwoNGfZYeYE84icTY
yAc5mEjmk+Z8JMwoTH6HZU9NtgbfQuGsH3QzI3oM5QE0jKJ5BCscqE1MdFOVWCOWY6jEI7rV2hly
kaH1wADAwTtN+I+FA7uyM2pu1nWrKfdkH4Rr1vHefIeyEFmfx/weqWz7mrYpihzg/sabKanYLu0y
kgSWhOFGjb4mZpw7KCvYj8MXGuk+5V1sZ3yQbffHRwVdNN8hNsOXMRAKycoZQD9RH217DUyqztlq
aLVSG34tcKtzue3Z9QyK7aTrIWNK43D7CxoqB7LY+Dl86ABc5QgYRXIpXvpogoQHEibuRTC9V+8F
39JMzyXpkBl0yTy4csUpjYxeOn2FuhDDxiuCMvB7ZW5RKJGwO0nfAQ5OxwpWyMJxjUelWKx0Aynb
gU7mo1rIqmLlWlc/waU5WHGtPOC/DzB8HesDMCt26rgs7WwMFMIszAUDp5yVBPHpZrpAltkcrskH
GUmq0Z9ikYyACzpmlP76y4NjlkO8yDKnWDN6vw4VOs302joyhTdW98JXBRtNCas2jpYPmXqpFAYQ
jPD7z5lmdseiIJO8dNgEuK1u4PNKAzL1O24vJnrs0lLVGPdxmTpik90rYbX2dlRdIKjloZo7R85E
qnwcXyA8QYRDQ5Dba5rHg2Biydkc+7D3me2p0g11QXsenlqotSUl7vNDhMZD/LntoIa5u79amKjv
MN/4pnrfM4rwcY1ZXcX7DKw35pESy16pT4rY7CNb9GrcKj1gkdFzqlPeTpuCApOuuEV1J7eovYlR
wa8JQo2d3mnmzD/Y66LARwiJ9mv3p7prjd7SNql5CgSTrZFsmLoyIjGzxojx4D1ZKbQiTQ8vptW7
Vpw/A8gQ1GfZpbvpO2emWrLq4uUcfS1XrnTOyTtmc3B5rF7bUaxqkxXslSjDTj46y1/7vQT6MAVK
0Ciko6cCpuVmfV2Anbbz+7wP1hvAQPpEJceqFmXg4W5NXli4fOZsWZiazl/bOWWd+oWP4sO7Qnxr
bVL6D04AlRlQ2LzKHQPbpFLQjWLyeLgTJqAhERyzXQckVhmNXfSwxayxWOTknKwZ5Zn9WKccFBOi
5yG+xeDZgtZzgRD9HCecCAi4LXcaVuQwrWXASGbA+1BKNe9T/43y4KKjsiYi+G+yL7aRbPcbgyJZ
/GSY6Ac2pVMoiXHmErxgBzcPOhfbXjGdUeGMlX9mCmO9XPXukbVELFkXXYq9t9Vnc1zjBPJP1ube
RlxWWwS8cwf+Xi0JIhPvrFsFmEf0tA81FnNGLltU7EaW44k94/Z4nohRO9WPaRK7RvKImCbBhOoP
4sdXH0CoDXIatECcZGdL34fO+oSZiMe7dT7JNW2+GX5aetMqBB3ZxX6mX24Xce6P+vSA/hCA8lhG
4Cla+rGzU/i69d/w22u7OG/jzAHfxlrKCpqb+3wMjUNB9r9V/2XtU76DxbexYGJ/uc3X5CN2H5H+
ONwk9uhZ3Et4IBaR9BR32yaFAm4Pjdu5iuPWCDvJ5gICLB/s42/K74LtQ/+4J0e6a9yYQ/AIV/x5
wITfDNqYcRhoH3FBMrNssIh7Q0/ilbM7yCiLwMm8Q+bcp+ZM7N3KIBAezhR/uQqH0pFgeb8qDWRQ
B6aEQlXgPW7eH/1w7zQjZyEMrNIZ3n2bmGaW3EHrILw0vgLeXCN2y4fivBnryzNdkW6myIDKBoLC
Yo/r7wj/UR+Tlhrw3M35w1dWj/cWqdlqU4KD6RM+oEa/XEnDv7M8w8HTPpZRr9F384osnAW0dwJ3
OV3kiUEcMwPxb5FT43RH71x40lyiY3BuceyuhvHBAdrA7MyAPsWbTHSp7pp+WioYJhpPvduCOfIU
vF4lbZbk1vazY/DRW1PiK1iSBXTQJ+Omqcj34rMcowlxgWobT7YqO7iJ/CBwTjAKEvTEwryNr+4Q
kZP2kqzunOJlYRGTpRjCbQnplcz/5eScWyUE8Gb9ackbdBpvNZ21wFEe4QStIAeG3aM3/YjPE8v1
9JeIaKqeB3TJs9R0jADrh8a7L6KWZvErE29+i9IhIZllVbgo7feUkDjQto9Sb6ymRZ2GKcu8T8rh
qKeCG5jt5zb+BISVcYLQauPSFHDVnJNfSh+CabIQxN72+fajxyqRA4+o5xf9leJzbkzrpe36xLm5
Khs7K5wBTlBqfL618yGbE30ZuaGi3YnMxDmvwYyQdOHuMdCEsO6Mag68+dV5ShKegePfFme+ymV/
/VVz9/BOO9GCSX3/DCAtWkz1BgtRXR11ERGxcPNqG9EG2b/vazldPQCLp6f/Qsui/EuQrzi+twc+
uewEYJVIaOfEhLbCtkzxdhPArKgS8eVhtA4icnZMKg90RCPwvPJAu1USYp9ucUaiuCmtp3ynop+d
6QjdCe/bB/+PZ1Ugx+vUq6m7aUj7h4MJ1STv1RMQj7VK89R9O3aWj2i7za1iSQiWi3ZrcLucJsFV
QCZC7rBt1dBnlTn8+lWeu6zg0XylOBmc4RsEF5pVZzA+MtOHSYIIMbFg5akpH17OZgflyZn7Lk+P
7+Ar5zYt9/A5Vp8dSJ7xjuKqzDFADnYoCfpkMGXuTCRtvJvAKogHhdUHuKeEgb4tG91AwMXyPrRM
SaTXWeJMif3bXTzl/VzM2kd6dLSawXoWoDiQIWHVYiMIGHg4Cc+3xKr/IBSOyAi+GzB5f9zS+qAi
H2QUjwt5hhP8h3mxtrBLSUTw5GS9MEtsGqsGvoD+qc196U800dGMQE07mzRFjeiVZHE60Gj5ER0q
kFCwiGmzoWzYKDY5IHAcFncFaHWvcOx6BVoGopR+z2Z7MgLbbYT2ptKQ78oSHNif7ILnuf5Gj8Pi
J9EX/kl6k4WOmA99u6if0V67TElQnmVkyrQv71uH6o2atokDEmLvUXfUSuFMRaUpe7rb3nt4r7WP
o50phORQ4KVJ75NI1CAWJD/sY8XcAdbRkzxpgSj3x71Iu1kii1bU3gAdg/zFkivtMl5Y3+pbSJYX
FDA8Lq4mMQN0EUOuVWIbjCJSuMiJbaPL4BGoivP+a2vuT2MHFqF+ZmZc4ftD/T9RfvWeYu1i0WRS
OCofkirOPnQIqaiH+02mJBDuA4vqLe6Dpn98siwS9C1SfYkaRKMBOGuiMK4ixRSY3sn4kV/nb1yn
9AKYcC3JCOnfyvV1Q1xn5iW6/o4lVR7HcvMtDSTCGHWoTMcdM57Kzb6UdqdckSwkp/ts2aeuRHzP
mvkhxnXSruqAk+T7MtEb1EyOXpnzjcuWxtAITFBQzUzE1hTqB7ktT05KfefJuVWihfBdymKkvkjP
sYJ3tzf6zOXjJpz3QkBERSj/Z3BeqeItcRKbMohF8MaoN12L8O3UPbUydf8D8zVTNM/BaOQidx3X
MtKJhtxWVxvteTZxJfcUUJTylQFwsy0C8iE1osUIEcxlzG+cdk+CLx4lntvIH/G4Yvi5Wy0Ct2kM
E/Mdj0aIBJtnoZ5jziR+sq3sJ7D9GXfbdcox5ntoM7RyDFYe0aWMAx29e4tqZzIVzrlWRTnvIll/
3ElgFj+lU/7WwCxFgQDgX1tPS61YdtHatXKWZdOV9plm6azL2BFki2qB+Rl4GKhYt+3gaZS3p21s
jcJK5Xn9aBGrcNW4KG1uTKCPqT5Pjy7KZdxgtIiABewTk9ni8RSHMvjRzkSvCIDLJuxhpa0WoyCy
1YoI5+Z70DwlAKNU1kWSHFMEq/Ap2D3x8hFljws4lr22pMosf9sx2i0Go4qt3Um1pi/ouB5/5biM
oZBWpGczG4fARc6SI88ZPUaFCAqkrkR+4ztC6iX9WsAIcPVrcutcfc72ICVzH1ToYSCYjBrUzXpT
9L4/S07AyXcaRhfWD1/wvp130zTDLwQpR36zITFw6WreeTehIpxGoUzz/zRpooLMBMpe71oUZhhy
KH4qnvy04/4+zRvcgkTgeRCxtgWDrHsvkyFsruzjtcIJLZjc6itAfcjwJtk6ppalKmnuiaSCPZeX
M1dTzzgxY6NKs7peFgi7vFogdLIxP6+HGQ2zBtYUaN6Vnlh5aNuwHlh1VQP6hn6L+CmP7kl8YmJf
SoRdbDhC9Y7fh3MIwAjAeHQe9l2vsdHgdzQhr8W8UZ4t/FN5Smj9h5WstAdxohEA+yJHe+o16zoO
zS5FBLuAZl2tO108nu3etIqa0Sn6j2x8eRNGZtgMfhmu8KyjYJaxLLVIbJB5gF3b1Q3qX+uqkamT
odPCxc6j+4wkPnoPC+9RQRP1ZXBW9U5uL9KzA2xbqOIQn5MTb3KsUSxPQDre+T4l7UjDDk42EHKA
OXElQAlUldIfRO8qw2XdYr2G0DTV2va0duQBJD41cZN/G3RpxAvj2ONL4pzvpRu304FsYZpguOPa
otQz7sfDGTi4nuQ0tR8Fz+AZcqGQB+3oPfy1MUqIrAW4BwRjiWX2W4jpDPe4gwbDQCf5DXoNgC93
q/HqBJbbixZzCHIDK+MuwkStueL+t4CL8lb7wlKaeJV9sPpQ7+y60m2Jk1jwZRHp+yVfj4GVn93E
aGf8SA675D7quodAaAFwZgrzGalpNhRCk5XP3yI6Rjzhw2aAtxsOrrqvh7QiE5SSOE2//KNSn2qw
IKo60n1VvqLuMvcwgm2CoxHz2s/ENjCDsxjk+pIf3xsvD7m/ej7x24/BnXXsg8XPNYO4Whh4QoVM
2NQvFEiHPkOLGKV+RR07phHsKqCKBCTiA/xwaXGPmCjS83AeKrzO465MJkx1PxN2YAgQW9p37e6E
EN0CORBLisr6M0ejEZLbDNbxofIiyGVwBb03xYhJE9PFz1Vhdh3oFc0wExjKwFBK1cE3f9+WeiNv
glxU/iL1rOM0nrj8mIkiTn9inOkB7d+Znit73DtLYq6t9WSNs77R2OkgturiynxewY3SsY9vfeBs
9FxHgtPg/XjSt4cA0H6+FwLKmwvu0ZB895dJ4ugq0q118nk0MoVgnPTt5p84GWweXO5Jq6z5CQSX
01PlwTvjYQIlDOsddxbHa+LkQDrLGA8sa01lx9QjkRH/7YpKaqUHzEVkRCgDT5qe5hFtXt+1eriN
MuSauWxLhYycqFsAWUKRXkBPKmQnFefDAxnuacOgz6JtMb86fXYzagg9truj2P3wUB2ht8InWGnp
8gyhhTReecDkV7W9/Ddp6gxAoFpVUk0xiTrIGJQDznrV9loR+W64c/1fEBTws4ocRbK8gpfQ9mSF
D6ayHTeStHEu8+3Nl5UuMW3AqbuT70QzhELmjIzjUQ/J+yBdi86xqjaCi2fAhwRGNep9HEb/W900
77Ziy2nvuTpkQc6bL5+scFipSxIRc3rng2rnaPhfpjsqMr6DY4z8+DmLY1lpWfAVn7WTYvVmSeTT
QoiDDhTSQLS8x/D0bF1cOplabkHBZDmcBo/jeEv/8zahuIe1cywIyqRwMpcXQqm87Jkil/kNU72Z
ZU+icJYEU5SuEsWT5KbwKyuduKZMyOGdRyI4vXL3keuw5cP+T/PMK6T5e/fz3dC4dW9NTss1omhN
d/alEspSrqH5qoOT9tth+v6xWioVaUMFP9Vs9g33zOmKUuU1PrB0+7Ir+ZbV9mOJU7U32gzbkZB2
QUK8Q55FcJWg3k+mlziV43EBIVWeZUFo3BByvUJuuAJQpPxrCIKLsPOU/GJ1lJlbCi8kvu4vLZ31
V03yxsS7JlKCYTWu4h579kKVzBU6owz0YuoBu3VTLdb+9GV3V/B58FPVGWkKlvzWpgB29i7viOI6
mKpmjPMKjgr310z2QyoKMudVDpo0ZXM1mzEsYlvrpP2T+ZktLC36/6VULu9DPiWK+olf9rvhiPk2
674LQuUkdoQWM6IinbqKpfK8lAedyk0wqB4WgKKaK2SuQ2kyynprl8sCgTDe0r3WTH4eicH27K0e
ejVPVxD7MdKqSJcXyVlnxTQpvN85xIiYCA+qlUo4O5K3kv4iApQgngraGYEP6ywUjWpdQ9GzSTZb
zUZjm2d7kRwPqswe8Kgdw+qrY3UnvdKWvwX+nOGvJDSSpKv5I0SFYk2wzaoK5fJs7cF2UtvkQDaY
SEHCAMHT86LsVqu8dTelsk/tv5IZxHbxDCh/hjV0OCleTfOIDYHJWJYfgUyYJSKuzf9d9uqnhleG
CV3ehARnaKohUch16Nsx3NQk69SDrb6aDuRzwPGDCGvqYaBdPQrMl4osUxfRpT5zgiuJydPXCvv1
xBoQsq1MFic67qaF2y/JY5lh8KPSKFmAdiMjVjcyNDEICOxPUfamWLjHr2fu7F3lc8IlhuDVu0qk
u2JnJrciT0oY0BZrXpez4ij46LcvEc/uBLNeHIRE9XPrFuxqv8q/NL4Kvi4Q8yukymH7+OsI9kk5
Q+Cf+Vz+hL0w2m697DEBccp4kqHFG/NKTCYz4o/QiZ4w+kC/I4CLjYbVxm1Y9R1jwZVlfhunsbhX
lv8aFot8aZ01c67GBTWqnWs5uWPZcrc88Q5sDL2THJTPvQu2bl+Ex0ovm7v0vbiRH5LvydtvxSCY
r221bvsEmdWrMVbPyoBwWOlj1vlStkF0SMNwfQ2XpSKkfUHm3BR9bnnoMgdP1AeesoLXM0lNmyrV
Q9YstGbzud5ieNi2ATPZYVlmN2XvmHnAvmcvZFARHzoEawIl6ACPi+dzQEFe7iexSlD93ZXxBobS
5tBc8uuLt1XVW7l/hX5lw340PoXgJsmvnoBpilxaIZ4Eh2UIH7cebf3AFjdITm/zfCVs00fBty7m
we0AdiWSi406MTo1vqDuueKQ+b3zN66WawK3KwFWjRkx8Ap4Bi7Tnt4NHvJyKjs4uddB3WxOVPcT
I0s5u9boDIDlIILlLWHRI7UwczxCysEm62++VBG2BSHiRpt9QqljSu0BEFrH7gqdLSc0cF0jHWW6
c2kooiLbT40ckD49zyhlN/yyZetG2lG86ASJkx2Jl0x5y2cdrPin2YDogNel2ToURGIYGYB/bLY/
RIg98NFNQ0LN2ybn1RoSJlCV58YVDBDg105k69s7dkWVSIcywSZfWCK6zzGdxuakp7NWvD3zKsoH
7eQkx6Im9kZJm0VznGm3GQtVoZWNJVGUupO6Q4SoC5a4g4EJC3fJGzcyy/lpkh8iu1MPyhzNrIZo
50l6iW6KH2sltdeKsohhs8+XSB99TFz4NaSuYRubO7ozBVy2iSS1XrZmeUSfbVXcb2UMaTRZIEAb
FMbVMK9ABJ4o4qcXRqP3J54MnKotbu0ZUbl8DGeiDFzE/XxBepZn6HYrUor7UPStclXPIuxSTRXA
wRMGueJzbI8oFa/nd/NYQDDnLSCAWcUdulLSJKlbji3eVjOaBJ+EYF9GtvQ8ecI7k9uBNqF2vKyx
5iRJi6XqIqp+ekNF4JPNSqQpayXtngfwUQw8IjwwxwLcMZ7yrlBO2j03hiOQcHB6nVz0bLiD1qiT
FFN6kTaeA/9NxcGHuoO2DShst7PlF5M+DrOl/vY1Elab94sxNBziza9ZcxtqbJEa9yoHMd2ArMBe
pBJMnpNa+22T7ksIUtpswzE9rFeHA0SXvrUKMwV27pfzKrrzdrzXCW6VzjzwlPJb6eWf6KNbqRP4
TFDyCn1aHRludmY0IOWg2cuSVH3lWsDp+P4avherrZK+ImNDuHaCl1YX+yxrlSKxiDtcdnryHlZr
t9hdUSRWMa1EWm2vo4n4ql6U4dUnzBJmzyPcb0gszSi1oSK6ouQFhpzvvtLDXywlc7i3RO/IWZ+A
Jsw6MlcCV+xQJVWv6jVB6LP/2r5GDDyH0anCxQeOhUUmASjo7F/FyqYqMh3VCGZAhl8l2zJJodz8
IsudwiBvX6e6l0CGjJgb8Za4jcRWnOOhduWcrO/u/4ZfWSp57uFwgeSkUua8AX8e2zQUgtJMviN2
nCka0UlGLL1kMPNdQhm3QC+QAlrtN7nIg51PYoZLfqUcLiIzzWpUaweFy0dczZI1asYQtg3zWs3o
YwhBYAPEfrT92Wzl+G57xPxd2auBX+nXfRhByrQl6PeNyzxsC1yWL0Mkwyta/5Q56I0yN/qtgUFj
Z4ohuRXRY9LKUiiz5GU1VXDYgELnECobR2rS+/+cDhVGMtLo4fasrkzzYv10WuwwKfQZP2m7ZuYI
zDmVYD9ilFXKMOBjTKN67854/BNva/BkyNh9sfSghTObzlhN1P+zOI8eOHd58khWvebGeIaDwNzN
JBzn5X6RRKphlKs46Gj6obrR7CCHSJHFAW1AabPQUnyV+04VM4HO3hyhgm45wEJgj9tFcGjwjLf4
WXwBI9KmrPXxzs3UFNq6g8g/zhSoDx3KkjlluO9vmmbaTtWhd0RBWVSxO0hjCCqfbXPLtW9L8lOF
5zlG/CUkwv6fANAA8YQknptbNlfu6QMu9PJNn/t/dYYBv2m1gK6Q7WV3Lk0SUZPDqG/WGspKLaXX
vji4w5G6b9NuVF2TfSnEw3E0J1XilY+4YvmkrGRFemhhjOI0taxBN1QZUDkIah3PCbhfteglJCTF
mD9vw93Ul7dIBCG3ir68uhwm65vhEE1WEJrWB1dK6pJsBolaAOOmbAkHQRtRyIMOzCl1SSysNNKz
muFRfGvF9wUTz2xEV9i0BUoxmFat2b/js1+KEhvVSy1y4oMPnxE7LAQv2iNVv8bEn+nPG/8pWdYw
X1KBneh5T4hRRmZfLNsmGZOCqJO5TwW9yrijbRMCzkY28yiD5JjTmI5EH/4qxzfy1DmCOG8/WA8J
xsofbaYni6fDc+EovAcGYPQm57/VMdbTiVZjLbvXbmC37GVVHPkUHcQ3tfkOCmJ1jMHX+iN+oeCP
iiJfHWaOpshwpJuWsT4F7wrmM37Z3DRq3tUPSbkUyIQ2lzcpEI1hRTXsVH7qWQP01Q3q1Fznw6YY
OvfCeVSMCKzsY9nXDtGUkVZCPaEWYH6t4Ls9DXy6VVQwiJPtiyVjYIwysv2xKSxL7DmLjXG+o453
8iBOoPIxMUOnzCRLkK2aI8bFsLDa0nO7Skn/eXNmezimAfPDp2joZkr7LlUMPYd5DuJdo7EJD6/7
LCGkJpO0O/L6+QmHJrgch9TDt9mbf7rii0N+fkEIbmZQ1dCJf9L+wBZHBAmO7R44Rwo4IkyLgVz3
R1aWlyj1nTZm7WlC+8U4oazVXtrSmDe/qQoBwMvVMPF4nN5ENQiOg5By1eh1trN62bsKJSO0HN7E
+4Xx937hvewx5945mVphjm7cpSSU50CLexLDhNFdSMWsm4oWXGgmqB37Fbt8f9gXGHaO1IRctHNG
HXjrxPngGhAa2K2hOF4fzWaSAqtmby0SkhW6rc3GzIim+WTEVlvdx+TLZB90KoMrN4H/7hor+Y2Q
yBPXvJKS4z2+rHWvA9A5tKdV7j9UHMtpBbKwqAlgsAEPl/+xXre0z4Qflu0qHBfFYrTXnVxdGoTw
tox3XVTtP5odsxhtQQkSsRyb+a54/dpfqWIe39p0IDzFr2W1feSCQwMhXWEzXwEHj0NjWCPcMFZA
NQmJAeAi39a6Cy8N1TmrZ/N9g/2g1P6hp2agZ3nG03ygnQywyOUcjSQR/8AJGwrVCFEoKo7N5lm2
6CvrJOUEyZxnGU7pCjGZh3f7pfqOm0Ur1cUEdYjYg/zshA20kvne5tI/2fUlOd6kWOkPB0mXk1IZ
/LdaZ42xBEpMmAMFkb3Ckd2khEtoG7ZanfGMEpjUhZPpWqshmFt+ZNXhO/GxIlhpBN6eub5pCkVy
e/eflLnHPlPNsr4IqfNdaTAAswmUqaVvC7xgqUbYZdCjOG0es1A9wTKDrLqBc9q/BfNCKdIHAuQT
Yd/sz5PCBMKyq+6qEMGeMqoGrbuXTAkEgedMiw/pmkNBd/jers6PXKfiBthCxbm2wH9Q3eYlgStM
Na8xY40AS9Wr4Oa6zSaHdDD6B86ZrEhrXfhMygC4ppACDPXb3ciDged+YHmpjgl+G2qcSmEX08mf
JjlHwLubpkuftgeX4VwNl8kbA1mqh1JXjrht2j5u2R/dpWF+EmWyWoueMIEn/qi9B8zIcbElOXqc
w9CSyPvNloSFbqsbMtQNhFBzqH6xYbM74D2+6d85tLJMMBZQhNOHBqlxBzx109Kf5cv4S4riztPF
fDpAw7HZmfezzEWl44vD4egaWst7lAgcLxpGj7bAPAe3ZVkCTG2LW7wrtElctaT34exO0wpQzNg3
N1KcrX1KRFiFvjMx+PVTTTQ/blIdWY3prs5cso4ClvOhOoeb8f38aFl4c5xAi8+U3FHkO7LfOfZ/
IxWpoQ0bqwZvbXw50ONfY2eL3cE4hXDyf4CMA0puwzuBW+oVfkGtk7Q7DyeEuQFFc3V4r/JpksWJ
/VbKNQbunjJ5+cbW5NoT3XFkDIudB0XcqfmLpSEE46jdEasFxHC2ovZ2nvKRRJQS+krOq+m6tvop
bVE1NTr9b2YQshVFl6JSiGVfCFaUS6QfLhhTPMrz6Uw398Iug/NY36YXFbzaWZ1qcNoAW4a3nU4t
GsPqg11wmIt8TqNXutTIdMJ7ecZJd15k3p7ZRT1Fm56JuFnk01eeQaoL2tUqPVeAjaDcCY/yGZ3Z
L5fBUCYKJIazsoOcd+3qvMOzmrA77ljG4vX6SQXNAjqAVddpUhGPYGPFI/YL3MaN2kRNcvtYiHYP
s/oSvxv3Z6bKIGEFnbWtjVWk+ZKII/EXIaKgoc2knUSqVPgqXuvsy87b4BIADdqzmTpqAqHDkzyq
7UK7QdzsiWZBrvtaHm7WQV8r/A3h89gao+QhT0r1xfV0IaB4XGXXar9spYlwVzS1PdPvNHBnnYgb
Sn7med3ThAVZedc1sRxUEeLfSpNAhBoPjQZwVpD4p5XbC1dkBnuzc4SCdXNGnLoCkzxWt+4XPEGb
uv3YGH9Jd74XWpGxX1hYQv/4lZDm0HcfHigP/DBatzAOFSGPf5x2KUnjv6FRgxdpCoLKmvYqqV0Q
W/ytPrf4DP97PXk8aJFt7uGpdWIaHA3QJkU5W34eW7ZY2u/hhyx8TeKuQmV1Fy1OzqumqptDYBZW
tDcx2bEvyHUzEDm9kongIKSneJh5qiLIOfrOYl/uFRATOPpnaaEgy2BSmf5Htfn/T2Nvm9MoLUbI
wZKyO8bFlzDGyO40VoS6nitE4sgmmuV1SMZnlQD3B97bZ2uU7Teqn0RHnWlp/R2yQd9kxQ+4KvGH
pOizDNmj390Xi4EcKbU+L96E20zzn7ZfT7J3uRcD2sEW2FsTwHRyBMbf+2HSEL2ug2twL06fUdop
HerbTLFsq6kl37zEjZ9XL8WJ4+nHc3CNSCdep0heQSW+EZuH1ObIkNGbeWgBbIIHskGbKuC67sjF
aImDPL6nHWqLBJCEV0kq8Ck+ytZzt5QqbwCdjI1K+CYjQKm0PYkt2sZv9T+LY84u7yk2eEZRguZk
FzWRjDA6yTC+sw1jGphY627Mm6RPWV9Vito+qFE+aRo98fIu3/Yxu1agbmdoYqZAg3S+GL5atptm
Np1q5u/n8JuzK6LS6/8vyMHo8S8Zj0oG06FZidk6Ao11DWhm5q/uyhUdtoQhiWNqosmGWskjWG8Y
2dhLuFFuEu1NFOk7cL4dSRYfupWpK97zGA3FQwAd432hvBRbmoaW9+fLxsVGmLS3i7eIM339xyex
2JK5c9m96QK2STgp1ybk0fyAxg64Aa5vUdvlQJEdP0jDeTiXf69yKuBNrxFVuwroZ5LSyI18UHp2
Y1z6ojAZ6pA83KFAKklcTp89xwu6W6a75jdDjPrIzcT4v2F9M1uG8iNUe7v2k/EUZqsl2iRtGcGD
E+pzZKpH/4gP+A3iKSuzHPEtAEE3H4pdoU/V3mFdHuswy11S+WMaGySEeddEGGc4mRXhQ3b4HKbh
3Xo9aSJc6kqiydY+breRkzridELicgVltOficN7ZVBQa0EWqW0WGlOzxKeOPd4TLD15tNfzvVAKa
HQ+XPdt0y5KsjhyNdpswIiGtrWEkVkyhfUNkrAOh8aMYMkFGV9Ysnm70V3JuJfkvwbN0nAD8MXwW
UzTODVMb9/N8uMz69BLObfZIwksPIoR0ZWYty7ShhEMNcLq3dMdVsw8pBl2IBkhdjwaShC106ioF
EQb6st2IkOpcM/HebZDUMG2sZmbnvv5YGGSKrHINpR7yNJfVTLM1Le8S2x3oqqdGnolYl8XJRyTg
fTeNLOI10byyUp4n4qI8EQTnB/VpBr8BToK/fDQFrzUcLS6Dpv9TLbhdzMpwofrxq6m4+R2DRbF0
PeBTb/10pUJVs1OmvYuG8fnD9rRuHBnwQID4hLwACI31MEwI0wROizeIi1goPPFeGW9A1EcgVpU7
44lXhR7um/tACgS37VqyaFZ4LF1EufeZiRabtT5K7YhqVvrGLEBS2noXfhqgo8mHsyXsiQxYhIuQ
yPbftJzxo9IBd1BX+hypOxRuqrbn1SvyOGxHoTYDwUPlwirDgId717TN2+elik6bZX/W0Td+Fluc
mgv7YqbQuQLTuwR3EnmRbefiHYwBZrfx86r2e/omG59He1vB7EmrVYjzAcOhzDFFb3sHbSjfGgPL
2EbI7QCT10jig1sjR6KuoD4Qm4g4+JuCqXHWoDxiuiEaNwuARI5O/uKOeChZdQFGLnd4No+SCR+U
ZUK34+UHN+3XmKsdrPxJ9MUa8Ws/IhAWx+dCM8OywIxvBqmHsQnAoi/2gwtI6qsB+wQPR8RK4hYL
z3RvvGWLNczurthXcHC4O5ifY3lODGS+YcGTBgYrqRed835wCOo/5v/FU173SBuTgETE+UWZiknQ
oLc08gBP3l70DW7HLy6ondh8nHahl0nLYPymH+5ahBouOtxALPAFCrMFjGuzP23uQQ+tD/lixU40
Rh+vNdkt8GgnU+2F56f53RRt8BmWk0t1KwaLTHAiDY8mwIgjemzhiVfJ9jC0EWdiW2lf+9XVn/Qr
7SYeo3j8BQ4twYYSReaa5UAWbQw6SokL1arwxd8lXIuzKpFKPx/FG9nQ7Q2/LtTFUug+EMJTxEEm
E3MnaWiGv9Z3alR+fhEiDeMDQ+hPzw7xGrNtYohHAtRIr8gZq9BKcI4j2lKgijkojg3eBtOUckyU
QgTFx1BMAyna5ddJAAWTZOeZinYkicfen3JzCt53DUOarxLGkjBGFSoyKGpdhPVwMgwyMC7Uclej
pGhpVQ/w6QEaWmnVGjIBX3vMLFSIc/ZetTTwTey4AFoAeBZ6mMdfoJRTGGdoXxwiKXbUPKyJUU+W
6XBUiiaXaMyRteQU5b1k86NltXhfc3LbptvE2jCXlKvMc3yg5/CEWTWJ5CpsaDwObvnZa1swbTO1
IIT8fdjwBDp17q4SVmuRXryWKmv0Uy0HoPTK9epDEo+Mup35XNqshWOQPNCRPyApV80eG8HdqJwt
Ydrl4FtLue03retqZ/kwpexMOTqm3Fza64aug/+qyzkAM65oHWlQZFc9H1GYrffu44yaRWOrisb8
lEeCzmKqJiId1/lWH9X9GrcMEs5UMR3GcHgbhQUc3tzTu2PURrXrGOW96GVuDN+3CBCw8hIIkI7W
+iO3e1q5q6bU1k65wpRhUROd11LFED2UOW8ACmbZgm+qLN/47JWwlMq3yBgjGFvxenw6mRqSBdNj
eqRAIYcAmJGMctIqA6ndkZObvRFmr9oN04tprGa3KK4rzDVNFdOzLnveRhJJ197DvmVHYO/6DDN7
DuCfTMUkNY9IjUmePCCMtHrrKIAI8P2tV+CkL2yOpBWN8IBDQOoPACN/EswygEkCSCxNGhoyMtgY
0csMA7NQcM/41Kk7LkBfLTN4Ow6AElLD8iE73hokblyO4/urbmVLAzXETKNRw55uN9OrTxFzJXWI
6tOA48oNx9u2EtoqCC2RH3uji0Bx5SUFvk15YFwt3VrdrPsVaS5VcetaU+kXhIFAzjasy8PaNrjk
+sHpOdeC9v3VlkhXDIMuctfAOjZ/xU5Pf3HzNiHN20Jjp0MNIXOddlu2dPvC9SNrvsD50HcLS3UE
gyhu0+GFXVnp9FxYA99E1LDV4wBC3bHZQiyaIg5deqc6TL7CtYvxtvm1VGQ7XhX9RBTDOLA3niWC
hJd6qwpAl+qXCJm1gdOYecAIRajmf0Gjt6+wSrOuBp+H/zr3e2NrFkCs9v4FauMv3CMkJDKGRJGy
aaBEflzIZtv50cN6NVZmpvDppgnFcazUiZuIyEfmjMPEIGdAG/1jIcFt+SbJ/p/6zsg3EdF1Zd5w
7Bl7mzB+C1qvy5QYZ+wByUJRSCkzbKkVvMZ9QkISKB4L5FYhV5EQqNyp0QYzPo5zn9OS7UWhV9vF
srg7zq66HXT5pEfJ7EoruKEduYJtmZG0PZD1WVGOMRFDJLr1F5V35R2E2bXtayPISoaW9zLRoXje
Ef5VZYZBv7ka8WGxcJoeTGcKY//duDHGIH0iLr40E7Zkeb7m6reFw4OU0TxjZ51SqNLwg5/1JZL3
l2d1ssxPcWCFCewOn++bkG5iu5jpj3NE9vlULbWViFJ8L1s/9ea1XG1roNtSmXhOLcvYBNkwLWpy
4qboJYBTQLoCVIvY5gS3b0T8aZ9hg7YLYI6yZFy9xceYyIlFrpTi5YB47oVv9t/0Yt+ucdFLvJfn
lv7kmXBjK9PvawNH7iUht8Hz9vCkz59uulcBDqIdk5aQxZU09xU85cphYGgSEaWTowD+GyNpbPen
oPEeRr5XLv8bSnj2g+ulV1PACA9GmCur727UwpwBlfxDavF7gmL2f6qOMWfWhGQ3mzQpC4C2E9xf
KM7bvI+Iv16ZUvWVo7Vi9qTZUCz9Z6Jjai/LlCn0skFEGGmCRzUjs7a0QV7lZOdRJWqs8avuG975
dTu00hMPgfLXkIxVfFkXJvjr4cd2xF8INGFFOqGapOdhV9Zi73uFQG7W+cUDW+DyAAzwWTB6g2Kh
baHlc32ug3C+syr8XTXrEFX2Kcs84Skav1TT3UkyFgE9BcryJezZbWBnjv64+uZgKrw2dk5VvO8w
msUeahqp+bi8RyQ5bBf3hr9lDLT0fG9zN0YQJFW13QVNJxK8ud+uuthFsqqS0xZ1GqI9Cb4Z6wQ3
8rX4I+XCl4v2cocEbEHhFhA4Z7Y5qdhuvw3Z9zuIpZbu76lhv3uGGzWEnxtv8s/4gzwuZdqUJH/Z
s31DvB/YBBG9WZ/G4YmJXznEVvTuHjmuZdBh/cZo2dwI7YCVXmmVl/TIJJVzgssAeZKRK0RzDclh
nzvJbgz/fSj4vvYH+QoUZ5tgcLliCqSKP4HBf44NFE9SyLTPtpVX7JudikNPP7JMuevTIf8uBXX7
xFHPJxcoMW1aXccaW4uEGKNaJpwrwBVB2H0uIuBJGf2ptnQaabP1365w7snFR7rG7dAz1x43Vvbk
FxB1XdnCY2BUohmIC9mCc5+Jsmf2nOfJ1a7CqRD3nUm8HfacXDpyQTmGkVDXH3MXN7QgfTkkidN1
gqNIF42HOauTHm4aZ3Q+a9VdZ3NGnFL7nWJ9CwjZa2jxF6eOvhAPRxcbgdMAB2ZwL4JgimK9sF5F
jWs5lpdp4uX4wIgzGvVDyUfLFv8qUJngfVHXZRgywjIQdmLTCl1OSZ2nXXPM1RUJFYJCzX2Dy9Jr
JHDTbZCOwocg5i//lNz3R+f5idQeF0XtcwbD3Kk8wNb6ZIF9H5C9rriRuHFlM3BdtDzK9VCy4tfk
qKPXRxV2Cq+jkgpVQPVsqEo5BxPIgmxdoXfqjDxYUqecGqLLSvYNUoCwvKeQis3gj1cy2EvcmDTW
pZjQhM61I7N7mVRkeJUn2g+Vj57nIUvm8vp+Z/WHXkrYgPua14WKpWYSqepleayc6YPmWz/cfke/
OfiOJifeVshKDf20/MdD+99GAawmoK/7iKdK7dAB8lLtjIBPNxLx2+rr/JMSBBA2pH1kMlECSAKc
2+WbvoI8yjLA8Ykud23ruqBn7JNKergfNbXCKBx22O6kQU5hYn9ytUnRCqBXaEzgDAtuRlC6hLy7
8owgS7IhyG4n6Dvsw+fnbelLn7s3VMVJzQgqE4n9AD723Ca9LW+2cRFpPl0D1lV6m8WFvQ1U5G08
AbjHatgVdhxMtNJWuuBOdVTd6pdgK/PN5RXVCfoPiiJHUfraPuskIFNTTXmHnlSLQiy8vemGD9Pm
MGP2qGE4d7Xc+0VLfRsGviHyyof0yLHuYNJWfhaFksd3O30F8iyRawvTDgaXkpC5G0ZX9rXB17ab
GZlmOWMUIN12XMmlmyjUXTiskhNq0DE4UcEkNTSqnebfG9F4Elrug8hAttyQqL2R7NPrYsO/Wrl3
KC/Fi+GOvU0teDCmH13AWa4kbZhH+eIF1oOAkQjFrJNpSepz40E7KWO+RT0WMLgdvHp/RzFi79hs
j3dYL+jBeGaGwgn80ZRsS8sVI2uBZ2oqqkxdt9vxiRflkRug7N4f/mIpw34llzo5fcoFc1mkOHVL
4YA3ncYLGYHfGQigfrMufsvXVESFVbSfI5A/Osc+a5dcLaH5n5z7P5Up0vDNEbBX/WcaGEeijAS+
FQwVkVjN8uxQKsOQv971SiXDpRSt8FRo6v5stzpsWaKfkNJ6yAmgrWXTY+RQlhBJQB5Hj2nAX+Q3
v6gzz1KUNyYgPJoXhRJbmiUlF7wHQYA0ao9p7PGcQDEn7Ms0pefnqNuSAooWQG0qtvCndHpSRbC8
STw19oV8/2u0QTLqkFNjDSb8CnRM8o7/y8S999rD2auXGxlHle2HWRq43oTYcoEQaWKgAaulp+S4
R9f9i7Pf3yEoGZ3CX5KkbCCNen6VDl7Qxj3IM6Iia72OXXCmX/mKYLeinQitv61sKf++1SBKMfWX
ZganhAeaR3caQ2iivhxVz68sM5c0to5m5niorokVt2Q9HUy1pWMejtypgDevuSUMOoYb5u+f5PrT
4zG4Og4B+yVSpx8ZPIkBVajVkwpXLLm7amHwraQkcAfBG2Kwef208oYHB1iAmGggUHURfoYStAOF
xRNTIC2IK/gcgn8BmRL0352XBdEEkYAGL6HO/MkKfsJYgU9S+0UT0GLxdf5hFX+MoN3TocHUGVTv
GDyhX8w8+4Zywmn+IgfAI1eS8g9xzTefSQsfGUTNghQ+Ez1IDa5t6YTozi55TR0LprT5+B+T28CD
b3vT0klDlXNIBjdHy4OqL4w1j4AEwIc2VrUw5L72jpa11VasxGENlljdfT4UgYqFVeeJlWINtfqg
37El4lKN0o4hcd2VyrTZ2uT+sXROoGetzDoNfrnP44Y+r0Ph85fvTz6w7twuNQNiaZ+wCCCTRlwe
f89f/ZDK5oP9QQ+Z9QrOHSb0MrPtzwmkt0Vt+ZSWzfnFQrDygAWC39GAyJZDY5Rq9rJicPkE4Dbv
gU6afM165mRcOMKat32sbtWED+/4tlmrsJkenLR7BeTpfnFLHgRBq/Hfdl+0f1fwaOdfRY2OQ0P6
x2jqonBcCtoYp4cbHI41U2EfatK5xlwsRT9zQYnhpwET2ExiL2edPF4OgwirtPPwAOG3f5mflPYX
aIxoloegULu7u5WL1yXkrwHA1GnSE8Y29qTL6sEpwpjJagbDKTeZzVH5Zr4YdadiFR7pWuxAQx5k
7VCCEQYmDxEJAYjbtuXLXpvPBYOLeOmO/2msX7n4gWbkyv0o+aAMjoM0+wNiejMeAZ15C1wq1cMi
t6S3jdH/1pegESisnCvmWElam6BuBkenq42f92u1TqYL3uxKlT12LH8sPn17FS3FP82qM/eTWDhe
B20BSjmtkLzpVl6BcZcGzsq2LxyrRCGDOS5CHhRmeMekVRFBs3RGtcEOl3CAKKYpxqX+p3yLIQDx
KJTWrRt1uhRHCEdjoPVw9nnzvFfY0ls+19WQoRm3Qg1p9KTQZDSFYVy+v9g7mJElSVCLELkVVtmj
UuYQmeT1mbYoANZxarb/UIWjdyMU0RBDQMdkAc/z7nNKkZrZ47IEllbdvJj5nS0/8j7Y6Okfm/q1
6+8gX85DZ63cwuYub/xTl/IUm6swKUYwny+k53NTPhuOoJxgm9nDepQ3nRB2StqhUn1/GAaesxvS
Thn0fJIbGKW7Fb8c3MN562JsB7omWM7x8PTN6lywsISI6gEb+ODv+pViN34zaza3ySiWe0x8arpM
ieQrMDM3fdxloJ4eGJ0OGqUQzlrUKxqgDxADpXg7UK1YOQZlAHMxIjp6mU3DsLdBgW02unQW7vWG
3QhJkFHBHOp7IUP1FdQmYSn3qwHlzGiKV66bqCZ1wNN24RIheQdcrl2hA8iZbsB5U4kal2NDPvaE
/mjqtPiwJu66rt6xlu5CYQZI+2Cpsn0pNo/yCSKYIvpg/apKHJ8BUnADbr9/T7Fz7vTmWTE2Bkec
YYf+htLdcvumWCSLsO8335rct5GBj3FK8IvhZfJ4v6gA7stgHTcF2SIEDdmbe4vJYEF0YkO6zeSD
d2jiz/9vtyxM8VKzArmy+lOt/U+xDgGXiQ3SSca8JuQoy1A32QwO87HRFuiPVg==

`protect end_protected
